magic
tech scmos
magscale 1 2
timestamp 1711438170
<< metal1 >>
rect -63 5738 -3 5998
rect 5970 5982 6063 5998
rect 5827 5917 5853 5923
rect 2487 5837 2533 5843
rect -63 5722 30 5738
rect -63 5218 -3 5722
rect 3927 5617 3993 5623
rect 5407 5617 5453 5623
rect 5527 5617 5673 5623
rect 5747 5597 5783 5603
rect 5777 5567 5783 5597
rect 5887 5597 5913 5603
rect 5777 5557 5793 5567
rect 5780 5553 5793 5557
rect 4727 5537 4773 5543
rect 6003 5478 6063 5982
rect 5970 5462 6063 5478
rect 627 5397 693 5403
rect 5327 5397 5413 5403
rect 527 5377 573 5383
rect 5727 5383 5740 5387
rect 5727 5373 5743 5383
rect 1927 5337 1953 5343
rect 5567 5337 5613 5343
rect 5737 5343 5743 5373
rect 5737 5337 5773 5343
rect 327 5317 473 5323
rect 2947 5317 3033 5323
rect 3367 5317 3433 5323
rect 4387 5317 4453 5323
rect 5407 5317 5493 5323
rect -63 5202 30 5218
rect -63 4698 -3 5202
rect 3727 5157 3753 5163
rect 1627 5137 1693 5143
rect 1347 5097 1373 5103
rect 1607 5097 1633 5103
rect 1787 5097 1913 5103
rect 3107 5097 3173 5103
rect 4167 5097 4273 5103
rect 4487 5097 4513 5103
rect 4907 5097 5033 5103
rect 5707 5097 5833 5103
rect 727 5077 753 5083
rect 2267 5077 2313 5083
rect 4807 4997 4853 5003
rect 6003 4958 6063 5462
rect 5970 4942 6063 4958
rect 2987 4877 3073 4883
rect 3907 4877 3973 4883
rect 5347 4877 5383 4883
rect 3027 4857 3053 4863
rect 3500 4863 3513 4867
rect 3497 4853 3513 4863
rect 4580 4863 4593 4867
rect 4577 4853 4593 4863
rect 4920 4863 4933 4867
rect 4917 4853 4933 4863
rect 5213 4863 5227 4873
rect 5377 4863 5383 4877
rect 5580 4863 5593 4867
rect 5213 4860 5243 4863
rect 5217 4857 5243 4860
rect 5377 4857 5403 4863
rect 3497 4827 3503 4853
rect 4577 4827 4583 4853
rect 4917 4827 4923 4853
rect 5237 4827 5243 4857
rect 2727 4817 2753 4823
rect 3497 4817 3513 4827
rect 3500 4813 3513 4817
rect 4577 4817 4593 4827
rect 4580 4813 4593 4817
rect 4917 4817 4933 4827
rect 4920 4813 4933 4817
rect 5227 4817 5243 4827
rect 5397 4823 5403 4857
rect 5577 4853 5593 4863
rect 5397 4817 5433 4823
rect 5227 4813 5240 4817
rect 5577 4823 5583 4853
rect 5537 4817 5583 4823
rect 567 4797 673 4803
rect 1527 4797 1573 4803
rect 2307 4797 2433 4803
rect 3747 4797 3813 4803
rect 4507 4797 4573 4803
rect 4687 4797 4713 4803
rect 4987 4797 5133 4803
rect 5537 4803 5543 4817
rect 5487 4797 5543 4803
rect 5807 4797 5853 4803
rect 2327 4777 2393 4783
rect 5487 4777 5513 4783
rect -63 4682 30 4698
rect -63 4178 -3 4682
rect 947 4657 973 4663
rect 27 4577 133 4583
rect 867 4577 1013 4583
rect 4547 4577 4613 4583
rect 4887 4577 4973 4583
rect 5867 4577 5913 4583
rect 3807 4557 3833 4563
rect 4647 4557 4673 4563
rect 1257 4537 1293 4543
rect 1257 4527 1263 4537
rect 1247 4517 1263 4527
rect 1247 4513 1260 4517
rect 4647 4517 4673 4523
rect 5117 4520 5173 4523
rect 5113 4517 5173 4520
rect 5113 4507 5127 4517
rect 5427 4497 5533 4503
rect 187 4457 213 4463
rect 3807 4457 3833 4463
rect 6003 4438 6063 4942
rect 5970 4422 6063 4438
rect 627 4337 653 4343
rect 1287 4337 1313 4343
rect 5760 4343 5773 4347
rect 5757 4333 5773 4343
rect 5757 4323 5763 4333
rect 5727 4317 5763 4323
rect 4647 4297 4673 4303
rect 5547 4297 5573 4303
rect 587 4277 713 4283
rect 867 4277 993 4283
rect 2827 4277 2873 4283
rect 4627 4277 4653 4283
rect 5487 4277 5513 4283
rect 5527 4277 5613 4283
rect 1107 4197 1153 4203
rect -63 4162 30 4178
rect -63 3658 -3 4162
rect 1127 4097 1193 4103
rect 3627 4077 3653 4083
rect 927 4057 1033 4063
rect 1087 4057 1153 4063
rect 1827 4057 1883 4063
rect 1877 4043 1883 4057
rect 2647 4057 2713 4063
rect 3427 4057 3573 4063
rect 4467 4057 4553 4063
rect 5267 4057 5313 4063
rect 5327 4057 5353 4063
rect 1877 4037 1903 4043
rect 1897 3987 1903 4037
rect 2227 4043 2240 4047
rect 3053 4043 3067 4053
rect 2227 4033 2243 4043
rect 3053 4040 3083 4043
rect 3057 4037 3083 4040
rect 2237 4003 2243 4033
rect 3077 4007 3083 4037
rect 2237 3997 2273 4003
rect 3067 3997 3083 4007
rect 4157 4007 4163 4053
rect 4157 3997 4173 4007
rect 3067 3993 3080 3997
rect 4160 3993 4173 3997
rect 1897 3986 1920 3987
rect 1897 3977 1913 3986
rect 1900 3973 1913 3977
rect 6003 3918 6063 4422
rect 5970 3902 6063 3918
rect 1447 3837 1473 3843
rect 5167 3837 5273 3843
rect 3807 3817 3833 3823
rect 5600 3823 5613 3827
rect 5597 3813 5613 3823
rect 5747 3817 5773 3823
rect 5597 3787 5603 3813
rect 5597 3777 5613 3787
rect 5600 3773 5613 3777
rect 3847 3757 3913 3763
rect 3987 3757 4053 3763
rect 4427 3757 4533 3763
rect 5427 3757 5493 3763
rect -63 3642 30 3658
rect -63 3138 -3 3642
rect 3007 3537 3133 3543
rect 3187 3537 3293 3543
rect 3627 3537 3733 3543
rect 5667 3537 5693 3543
rect 5707 3537 5793 3543
rect 3540 3523 3553 3527
rect 3537 3513 3553 3523
rect 3647 3517 3673 3523
rect 5047 3517 5093 3523
rect 5207 3517 5233 3523
rect 3537 3487 3543 3513
rect 5560 3523 5573 3527
rect 5557 3513 5573 3523
rect 5880 3523 5893 3527
rect 5877 3513 5893 3523
rect 5557 3487 5563 3513
rect 3537 3477 3553 3487
rect 3540 3473 3553 3477
rect 5557 3477 5573 3487
rect 5560 3473 5573 3477
rect 5877 3483 5883 3513
rect 5847 3477 5883 3483
rect 3507 3457 3533 3463
rect 5687 3457 5773 3463
rect 3627 3417 3673 3423
rect 6003 3398 6063 3902
rect 5970 3382 6063 3398
rect 4687 3317 4813 3323
rect 2467 3297 2513 3303
rect 3520 3303 3533 3307
rect 3517 3293 3533 3303
rect 4320 3303 4333 3307
rect 4317 3293 4333 3303
rect 4607 3297 4633 3303
rect 3517 3267 3523 3293
rect 4317 3267 4323 3293
rect 3517 3257 3533 3267
rect 3520 3253 3533 3257
rect 4317 3257 4333 3267
rect 4320 3253 4333 3257
rect 527 3237 693 3243
rect 3667 3237 3733 3243
rect 4007 3237 4033 3243
rect 4687 3237 4813 3243
rect 5347 3237 5393 3243
rect 4607 3217 4633 3223
rect -63 3122 30 3138
rect -63 2618 -3 3122
rect 2687 3037 2713 3043
rect 1807 3017 1873 3023
rect 2487 3017 2573 3023
rect 2677 3017 2733 3023
rect 2677 3003 2683 3017
rect 3127 3017 3213 3023
rect 3267 3017 3373 3023
rect 3907 3017 3953 3023
rect 4367 3017 4433 3023
rect 4487 3017 4543 3023
rect 2657 2997 2683 3003
rect 3277 3000 3313 3003
rect 3273 2997 3313 3000
rect 2657 2967 2663 2997
rect 3273 2986 3287 2997
rect 3740 3003 3753 3007
rect 3737 2993 3753 3003
rect 4537 3003 4543 3017
rect 4847 3017 4893 3023
rect 5587 3017 5673 3023
rect 5787 3017 5933 3023
rect 4537 2997 4563 3003
rect 967 2957 993 2963
rect 2657 2957 2673 2967
rect 2660 2953 2673 2957
rect 3737 2963 3743 2993
rect 3707 2957 3743 2963
rect 4557 2963 4563 2997
rect 4557 2957 4593 2963
rect 5853 2963 5867 2973
rect 5853 2960 5883 2963
rect 5857 2957 5883 2960
rect 5877 2943 5883 2957
rect 5877 2937 5933 2943
rect 6003 2878 6063 3382
rect 5970 2862 6063 2878
rect 3767 2797 3833 2803
rect 4567 2797 4593 2803
rect 4713 2783 4727 2793
rect 4713 2780 4743 2783
rect 4717 2777 4743 2780
rect 4737 2747 4743 2777
rect 4727 2737 4743 2747
rect 4727 2733 4740 2737
rect 1827 2717 1853 2723
rect 2607 2717 2713 2723
rect 3767 2717 3853 2723
rect 4527 2717 4653 2723
rect 4987 2717 5113 2723
rect 5687 2697 5753 2703
rect 2947 2637 2993 2643
rect -63 2602 30 2618
rect -63 2098 -3 2602
rect 1507 2517 1573 2523
rect 767 2497 793 2503
rect 2047 2497 2073 2503
rect 2127 2497 2153 2503
rect 2167 2497 2213 2503
rect 2327 2497 2353 2503
rect 3007 2497 3093 2503
rect 3387 2497 3473 2503
rect 3867 2497 3973 2503
rect 3907 2437 3933 2443
rect 4767 2417 4793 2423
rect 5147 2417 5193 2423
rect 5287 2417 5333 2423
rect 5607 2377 5653 2383
rect 6003 2358 6063 2862
rect 5970 2342 6063 2358
rect 2607 2297 2633 2303
rect 2247 2277 2313 2283
rect 5727 2277 5803 2283
rect 1907 2257 1933 2263
rect 3800 2263 3813 2267
rect 3797 2253 3813 2263
rect 5167 2263 5180 2267
rect 5167 2253 5183 2263
rect 1273 2227 1287 2233
rect 3797 2227 3803 2253
rect 1267 2220 1287 2227
rect 1267 2217 1283 2220
rect 1267 2213 1280 2217
rect 3247 2217 3293 2223
rect 3797 2217 3813 2227
rect 3800 2213 3813 2217
rect 5177 2223 5183 2253
rect 5177 2217 5213 2223
rect 5797 2223 5803 2277
rect 5820 2263 5833 2267
rect 5777 2217 5803 2223
rect 5817 2253 5833 2263
rect 1147 2197 1193 2203
rect 4987 2197 5033 2203
rect 5777 2203 5783 2217
rect 5817 2207 5823 2253
rect 5727 2197 5783 2203
rect 5807 2197 5823 2207
rect 5807 2193 5820 2197
rect -63 2082 30 2098
rect -63 1578 -3 2082
rect 3147 1997 3173 2003
rect 3707 1997 3793 2003
rect 5887 1997 5953 2003
rect 3777 1977 3833 1983
rect 3777 1963 3783 1977
rect 5567 1977 5713 1983
rect 5927 1977 5953 1983
rect 5000 1963 5013 1967
rect 3757 1957 3783 1963
rect 1087 1917 1113 1923
rect 3757 1923 3763 1957
rect 4997 1953 5013 1963
rect 5617 1957 5673 1963
rect 4997 1927 5003 1953
rect 5617 1927 5623 1957
rect 3717 1920 3763 1923
rect 3713 1917 3763 1920
rect 3713 1907 3727 1917
rect 4187 1920 4243 1923
rect 4187 1917 4247 1920
rect 4997 1917 5013 1927
rect 1047 1897 1093 1903
rect 4233 1907 4247 1917
rect 5000 1913 5013 1917
rect 5607 1917 5623 1927
rect 5607 1913 5620 1917
rect 5597 1903 5603 1913
rect 5597 1897 5693 1903
rect 1807 1877 1853 1883
rect 3607 1877 3633 1883
rect 3727 1857 3753 1863
rect 4807 1857 4853 1863
rect 6003 1838 6063 2342
rect 5970 1822 6063 1838
rect 1927 1777 1973 1783
rect 3287 1777 3313 1783
rect 207 1743 220 1747
rect 207 1733 223 1743
rect 2307 1743 2320 1747
rect 2307 1733 2323 1743
rect 217 1686 223 1733
rect 2317 1707 2323 1733
rect 507 1697 553 1703
rect 2307 1697 2323 1707
rect 3117 1737 3153 1743
rect 3117 1703 3123 1737
rect 3267 1743 3280 1747
rect 3267 1733 3283 1743
rect 3547 1737 3573 1743
rect 5787 1737 5813 1743
rect 3277 1707 3283 1733
rect 3097 1697 3123 1703
rect 2307 1693 2320 1697
rect 2907 1677 2953 1683
rect 3097 1683 3103 1697
rect 3267 1697 3283 1707
rect 3267 1693 3280 1697
rect 5607 1697 5633 1703
rect 3067 1677 3103 1683
rect 3307 1677 3353 1683
rect 4127 1677 4213 1683
rect 4907 1677 5013 1683
rect 5887 1677 5933 1683
rect 4287 1657 4353 1663
rect -63 1562 30 1578
rect -63 1058 -3 1562
rect 2327 1497 2353 1503
rect 5407 1477 5433 1483
rect 557 1386 563 1453
rect 1207 1457 1333 1463
rect 1527 1457 1573 1463
rect 1647 1457 1733 1463
rect 2487 1457 2523 1463
rect 2517 1407 2523 1457
rect 3067 1457 3113 1463
rect 4427 1457 4463 1463
rect 4457 1443 4463 1457
rect 5307 1457 5333 1463
rect 5467 1457 5493 1463
rect 5587 1457 5653 1463
rect 5787 1457 5813 1463
rect 4457 1437 4483 1443
rect 1867 1397 1913 1403
rect 2207 1397 2233 1403
rect 2507 1397 2523 1407
rect 4477 1403 4483 1437
rect 5107 1437 5133 1443
rect 5587 1437 5613 1443
rect 4477 1397 4513 1403
rect 2507 1393 2520 1397
rect 5077 1400 5133 1403
rect 5073 1397 5133 1400
rect 5073 1387 5087 1397
rect 5707 1377 5773 1383
rect 4747 1357 4793 1363
rect 6003 1318 6063 1822
rect 5970 1302 6063 1318
rect 4567 1257 4613 1263
rect 4507 1237 4633 1243
rect 5547 1237 5593 1243
rect 2967 1223 2980 1227
rect 2967 1213 2983 1223
rect 3827 1217 3853 1223
rect 4787 1217 4833 1223
rect 4980 1223 4993 1227
rect 4977 1213 4993 1223
rect 5460 1223 5473 1227
rect 5457 1213 5473 1223
rect 5567 1223 5580 1227
rect 5567 1213 5583 1223
rect 2977 1187 2983 1213
rect 567 1177 593 1183
rect 2967 1177 2983 1187
rect 4977 1187 4983 1213
rect 5457 1187 5463 1213
rect 4977 1177 4993 1187
rect 2967 1173 2980 1177
rect 4980 1173 4993 1177
rect 5457 1177 5473 1187
rect 5460 1173 5473 1177
rect 5577 1183 5583 1213
rect 5717 1187 5723 1213
rect 5577 1177 5613 1183
rect 5707 1177 5723 1187
rect 5707 1173 5720 1177
rect 307 1157 353 1163
rect 1687 1157 1753 1163
rect 2507 1157 2613 1163
rect 3007 1157 3033 1163
rect 3087 1157 3113 1163
rect 3247 1157 3333 1163
rect 4607 1157 4673 1163
rect 5067 1157 5113 1163
rect 5367 1157 5433 1163
rect 5447 1157 5493 1163
rect -63 1042 30 1058
rect -63 538 -3 1042
rect 1847 957 1893 963
rect 2227 957 2273 963
rect 367 937 433 943
rect 1267 937 1293 943
rect 3567 937 3653 943
rect 4667 937 4753 943
rect 5227 937 5273 943
rect 5487 937 5543 943
rect 1407 917 1433 923
rect 2367 917 2393 923
rect 1867 877 1893 883
rect 5537 883 5543 937
rect 5627 937 5693 943
rect 5887 937 5913 943
rect 5517 877 5543 883
rect 827 857 853 863
rect 1367 857 1413 863
rect 3087 857 3173 863
rect 5517 863 5523 877
rect 5487 857 5523 863
rect 6003 798 6063 1302
rect 5970 782 6063 798
rect 3467 717 3493 723
rect 4187 717 4213 723
rect 5227 717 5293 723
rect 397 667 403 713
rect 5753 667 5767 673
rect 397 657 413 667
rect 400 653 413 657
rect 5747 660 5767 667
rect 5747 657 5763 660
rect 5747 653 5760 657
rect 147 637 233 643
rect 247 637 313 643
rect 927 637 953 643
rect 3467 637 3513 643
rect 4307 637 4413 643
rect 427 617 473 623
rect 3267 617 3313 623
rect -63 522 30 538
rect -63 18 -3 522
rect 4367 437 4393 443
rect 1207 417 1333 423
rect 3707 417 3773 423
rect 2047 397 2073 403
rect 4487 337 4533 343
rect 6003 278 6063 782
rect 5970 262 6063 278
rect 487 197 533 203
rect 1507 177 1533 183
rect 1307 117 1413 123
rect 2727 117 2773 123
rect 3967 117 4033 123
rect 5427 97 5453 103
rect 2627 57 2653 63
rect -63 2 30 18
rect 6003 2 6063 262
<< m2contact >>
rect 5813 5913 5827 5927
rect 5853 5913 5867 5927
rect 2473 5833 2487 5847
rect 2533 5833 2547 5847
rect 3913 5613 3927 5627
rect 3993 5613 4007 5627
rect 5393 5614 5407 5628
rect 5453 5613 5467 5627
rect 5513 5613 5527 5627
rect 5673 5613 5687 5627
rect 5733 5593 5747 5607
rect 5873 5593 5887 5607
rect 5913 5593 5927 5607
rect 5793 5553 5807 5567
rect 4713 5533 4727 5547
rect 4773 5533 4787 5547
rect 613 5393 627 5407
rect 693 5393 707 5407
rect 5313 5393 5327 5407
rect 5413 5393 5427 5407
rect 513 5373 527 5387
rect 573 5372 587 5386
rect 5713 5373 5727 5387
rect 1913 5333 1927 5347
rect 1953 5333 1967 5347
rect 5553 5333 5567 5347
rect 5613 5333 5627 5347
rect 5773 5333 5787 5347
rect 313 5313 327 5327
rect 473 5313 487 5327
rect 2933 5313 2947 5327
rect 3033 5313 3047 5327
rect 3353 5313 3367 5327
rect 3433 5313 3447 5327
rect 4373 5313 4387 5327
rect 4453 5313 4467 5327
rect 5393 5313 5407 5327
rect 5493 5313 5507 5327
rect 3713 5153 3727 5167
rect 3753 5153 3767 5167
rect 1613 5133 1627 5147
rect 1693 5133 1707 5147
rect 1333 5093 1347 5107
rect 1373 5094 1387 5108
rect 1593 5093 1607 5107
rect 1633 5093 1647 5107
rect 1773 5093 1787 5107
rect 1913 5093 1927 5107
rect 3093 5093 3107 5107
rect 3173 5093 3187 5107
rect 4153 5093 4167 5107
rect 4273 5093 4287 5107
rect 4473 5093 4487 5107
rect 4513 5093 4527 5107
rect 4893 5093 4907 5107
rect 5033 5093 5047 5107
rect 5693 5093 5707 5107
rect 5833 5093 5847 5107
rect 713 5073 727 5087
rect 753 5073 767 5087
rect 2253 5073 2267 5087
rect 2313 5073 2327 5087
rect 4793 4993 4807 5007
rect 4853 4993 4867 5007
rect 2973 4874 2987 4888
rect 3073 4873 3087 4887
rect 3893 4873 3907 4887
rect 3973 4873 3987 4887
rect 5213 4873 5227 4887
rect 5333 4873 5347 4887
rect 3013 4853 3027 4867
rect 3053 4852 3067 4866
rect 3513 4853 3527 4867
rect 4593 4853 4607 4867
rect 4933 4853 4947 4867
rect 2713 4813 2727 4827
rect 2753 4813 2767 4827
rect 3513 4813 3527 4827
rect 4593 4813 4607 4827
rect 4933 4813 4947 4827
rect 5213 4813 5227 4827
rect 5593 4853 5607 4867
rect 5433 4813 5447 4827
rect 553 4793 567 4807
rect 673 4793 687 4807
rect 1513 4793 1527 4807
rect 1573 4793 1587 4807
rect 2293 4793 2307 4807
rect 2433 4793 2447 4807
rect 3733 4793 3747 4807
rect 3813 4793 3827 4807
rect 4493 4793 4507 4807
rect 4573 4793 4587 4807
rect 4673 4793 4687 4807
rect 4713 4793 4727 4807
rect 4973 4793 4987 4807
rect 5133 4793 5147 4807
rect 5473 4793 5487 4807
rect 5793 4793 5807 4807
rect 5853 4793 5867 4807
rect 2313 4773 2327 4787
rect 2393 4773 2407 4787
rect 5473 4772 5487 4786
rect 5513 4773 5527 4787
rect 933 4653 947 4667
rect 973 4653 987 4667
rect 13 4573 27 4587
rect 133 4573 147 4587
rect 853 4573 867 4587
rect 1013 4573 1027 4587
rect 4533 4573 4547 4587
rect 4613 4573 4627 4587
rect 4873 4573 4887 4587
rect 4973 4573 4987 4587
rect 5853 4573 5867 4587
rect 5913 4573 5927 4587
rect 3793 4553 3807 4567
rect 3833 4553 3847 4567
rect 4633 4553 4647 4567
rect 4673 4553 4687 4567
rect 1293 4533 1307 4547
rect 1233 4513 1247 4527
rect 4633 4513 4647 4527
rect 4673 4513 4687 4527
rect 5173 4513 5187 4527
rect 5113 4493 5127 4507
rect 5413 4493 5427 4507
rect 5533 4493 5547 4507
rect 173 4453 187 4467
rect 213 4453 227 4467
rect 3793 4453 3807 4467
rect 3833 4453 3847 4467
rect 613 4333 627 4347
rect 653 4333 667 4347
rect 1273 4333 1287 4347
rect 1313 4333 1327 4347
rect 5773 4333 5787 4347
rect 5713 4312 5727 4326
rect 4633 4293 4647 4307
rect 4673 4293 4687 4307
rect 5533 4293 5547 4307
rect 5573 4293 5587 4307
rect 573 4273 587 4287
rect 713 4273 727 4287
rect 853 4273 867 4287
rect 993 4273 1007 4287
rect 2813 4273 2827 4287
rect 2873 4273 2887 4287
rect 4613 4273 4627 4287
rect 4653 4273 4667 4287
rect 5473 4273 5487 4287
rect 5513 4273 5527 4287
rect 5613 4273 5627 4287
rect 1093 4193 1107 4207
rect 1153 4193 1167 4207
rect 1113 4093 1127 4107
rect 1193 4093 1207 4107
rect 3613 4072 3627 4086
rect 3653 4073 3667 4087
rect 913 4053 927 4067
rect 1033 4053 1047 4067
rect 1073 4053 1087 4067
rect 1153 4053 1167 4067
rect 1813 4053 1827 4067
rect 2633 4053 2647 4067
rect 2713 4053 2727 4067
rect 3053 4053 3067 4067
rect 3413 4053 3427 4067
rect 3573 4054 3587 4068
rect 4153 4053 4167 4067
rect 4453 4053 4467 4067
rect 4553 4053 4567 4067
rect 5253 4053 5267 4067
rect 5313 4053 5327 4067
rect 5353 4053 5367 4067
rect 2213 4033 2227 4047
rect 2273 3993 2287 4007
rect 3053 3993 3067 4007
rect 4173 3993 4187 4007
rect 1913 3972 1927 3986
rect 1433 3833 1447 3847
rect 1473 3833 1487 3847
rect 5153 3833 5167 3847
rect 5273 3833 5287 3847
rect 3793 3813 3807 3827
rect 3833 3812 3847 3826
rect 5613 3813 5627 3827
rect 5733 3813 5747 3827
rect 5773 3813 5787 3827
rect 5613 3773 5627 3787
rect 3833 3753 3847 3767
rect 3913 3753 3927 3767
rect 3973 3753 3987 3767
rect 4053 3753 4067 3767
rect 4413 3753 4427 3767
rect 4533 3753 4547 3767
rect 5413 3753 5427 3767
rect 5493 3751 5507 3765
rect 2993 3533 3007 3547
rect 3133 3534 3147 3548
rect 3173 3533 3187 3547
rect 3293 3533 3307 3547
rect 3613 3533 3627 3547
rect 3733 3533 3747 3547
rect 5653 3533 5667 3547
rect 5693 3533 5707 3547
rect 5793 3533 5807 3547
rect 3553 3513 3567 3527
rect 3633 3513 3647 3527
rect 3673 3513 3687 3527
rect 5033 3513 5047 3527
rect 5093 3513 5107 3527
rect 5193 3513 5207 3527
rect 5233 3512 5247 3526
rect 5573 3513 5587 3527
rect 5893 3513 5907 3527
rect 3553 3473 3567 3487
rect 5573 3473 5587 3487
rect 5833 3473 5847 3487
rect 3493 3453 3507 3467
rect 3533 3453 3547 3467
rect 5673 3453 5687 3467
rect 5773 3453 5787 3467
rect 3613 3413 3627 3427
rect 3673 3412 3687 3426
rect 4673 3313 4687 3327
rect 4813 3313 4827 3327
rect 2453 3293 2467 3307
rect 2513 3293 2527 3307
rect 3533 3293 3547 3307
rect 4333 3293 4347 3307
rect 4593 3293 4607 3307
rect 4633 3293 4647 3307
rect 3533 3253 3547 3267
rect 4333 3253 4347 3267
rect 513 3233 527 3247
rect 693 3233 707 3247
rect 3653 3233 3667 3247
rect 3733 3233 3747 3247
rect 3993 3233 4007 3247
rect 4033 3233 4047 3247
rect 4673 3233 4687 3247
rect 4813 3233 4827 3247
rect 5333 3233 5347 3247
rect 5393 3233 5407 3247
rect 4593 3213 4607 3227
rect 4633 3213 4647 3227
rect 2673 3033 2687 3047
rect 2713 3033 2727 3047
rect 1793 3013 1807 3027
rect 1873 3013 1887 3027
rect 2473 3013 2487 3027
rect 2573 3013 2587 3027
rect 2733 3012 2747 3026
rect 3113 3013 3127 3027
rect 3213 3014 3227 3028
rect 3253 3013 3267 3027
rect 3373 3013 3387 3027
rect 3893 3013 3907 3027
rect 3953 3014 3967 3028
rect 4353 3013 4367 3027
rect 4433 3013 4447 3027
rect 4473 3013 4487 3027
rect 3313 2993 3327 3007
rect 3753 2993 3767 3007
rect 4833 3013 4847 3027
rect 4893 3013 4907 3027
rect 5573 3013 5587 3027
rect 5673 3013 5687 3027
rect 5773 3013 5787 3027
rect 5933 3013 5947 3027
rect 3273 2972 3287 2986
rect 953 2953 967 2967
rect 993 2953 1007 2967
rect 2673 2953 2687 2967
rect 3693 2953 3707 2967
rect 5853 2973 5867 2987
rect 4593 2953 4607 2967
rect 5933 2933 5947 2947
rect 3753 2793 3767 2807
rect 3833 2793 3847 2807
rect 4553 2793 4567 2807
rect 4593 2793 4607 2807
rect 4713 2793 4727 2807
rect 4713 2733 4727 2747
rect 1813 2713 1827 2727
rect 1853 2713 1867 2727
rect 2593 2713 2607 2727
rect 2713 2713 2727 2727
rect 3753 2713 3767 2727
rect 3853 2713 3867 2727
rect 4513 2713 4527 2727
rect 4653 2713 4667 2727
rect 4973 2713 4987 2727
rect 5113 2713 5127 2727
rect 5673 2692 5687 2706
rect 5753 2693 5767 2707
rect 2933 2633 2947 2647
rect 2993 2633 3007 2647
rect 1493 2513 1507 2527
rect 1573 2513 1587 2527
rect 753 2493 767 2507
rect 793 2493 807 2507
rect 2033 2493 2047 2507
rect 2073 2493 2087 2507
rect 2113 2493 2127 2507
rect 2153 2493 2167 2507
rect 2213 2494 2227 2508
rect 2313 2493 2327 2507
rect 2353 2493 2367 2507
rect 2993 2493 3007 2507
rect 3093 2493 3107 2507
rect 3373 2493 3387 2507
rect 3473 2493 3487 2507
rect 3853 2493 3867 2507
rect 3973 2492 3987 2506
rect 3893 2433 3907 2447
rect 3933 2433 3947 2447
rect 4753 2413 4767 2427
rect 4793 2413 4807 2427
rect 5133 2413 5147 2427
rect 5193 2411 5207 2425
rect 5273 2413 5287 2427
rect 5333 2413 5347 2427
rect 5593 2373 5607 2387
rect 5653 2373 5667 2387
rect 2593 2293 2607 2307
rect 2633 2293 2647 2307
rect 2233 2272 2247 2286
rect 2313 2274 2327 2288
rect 5713 2273 5727 2287
rect 1893 2253 1907 2267
rect 1933 2253 1947 2267
rect 3813 2253 3827 2267
rect 5153 2253 5167 2267
rect 1273 2233 1287 2247
rect 1253 2213 1267 2227
rect 3233 2213 3247 2227
rect 3293 2213 3307 2227
rect 3813 2213 3827 2227
rect 5213 2213 5227 2227
rect 5833 2253 5847 2267
rect 1133 2193 1147 2207
rect 1193 2193 1207 2207
rect 4973 2193 4987 2207
rect 5033 2193 5047 2207
rect 5713 2191 5727 2205
rect 5793 2193 5807 2207
rect 3133 1993 3147 2007
rect 3173 1993 3187 2007
rect 3693 1993 3707 2007
rect 3793 1993 3807 2007
rect 5873 1993 5887 2007
rect 5953 1993 5967 2007
rect 3833 1973 3847 1987
rect 5553 1973 5567 1987
rect 5713 1973 5727 1987
rect 5913 1974 5927 1988
rect 5953 1972 5967 1986
rect 1073 1913 1087 1927
rect 1113 1913 1127 1927
rect 5013 1953 5027 1967
rect 5673 1953 5687 1967
rect 4173 1913 4187 1927
rect 1033 1893 1047 1907
rect 1093 1893 1107 1907
rect 3713 1893 3727 1907
rect 5013 1913 5027 1927
rect 5593 1913 5607 1927
rect 4233 1893 4247 1907
rect 5693 1893 5707 1907
rect 1793 1873 1807 1887
rect 1853 1873 1867 1887
rect 3593 1872 3607 1886
rect 3633 1873 3647 1887
rect 3713 1853 3727 1867
rect 3753 1853 3767 1867
rect 4793 1853 4807 1867
rect 4853 1853 4867 1867
rect 1913 1773 1927 1787
rect 1973 1773 1987 1787
rect 3273 1773 3287 1787
rect 3313 1772 3327 1786
rect 193 1733 207 1747
rect 2293 1733 2307 1747
rect 493 1693 507 1707
rect 553 1693 567 1707
rect 2293 1693 2307 1707
rect 3153 1733 3167 1747
rect 3253 1733 3267 1747
rect 3533 1733 3547 1747
rect 3573 1733 3587 1747
rect 5773 1733 5787 1747
rect 5813 1733 5827 1747
rect 213 1672 227 1686
rect 2893 1673 2907 1687
rect 2953 1673 2967 1687
rect 3053 1673 3067 1687
rect 3253 1693 3267 1707
rect 5593 1693 5607 1707
rect 5633 1693 5647 1707
rect 3293 1673 3307 1687
rect 3353 1673 3367 1687
rect 4113 1673 4127 1687
rect 4213 1673 4227 1687
rect 4893 1673 4907 1687
rect 5013 1673 5027 1687
rect 5873 1673 5887 1687
rect 5933 1673 5947 1687
rect 4273 1653 4287 1667
rect 4353 1653 4367 1667
rect 2313 1493 2327 1507
rect 2353 1493 2367 1507
rect 5393 1473 5407 1487
rect 5433 1473 5447 1487
rect 553 1453 567 1467
rect 1193 1452 1207 1466
rect 1333 1453 1347 1467
rect 1513 1453 1527 1467
rect 1573 1453 1587 1467
rect 1633 1453 1647 1467
rect 1733 1453 1747 1467
rect 2473 1454 2487 1468
rect 3053 1453 3067 1467
rect 3113 1452 3127 1466
rect 4413 1453 4427 1467
rect 5293 1453 5307 1467
rect 5333 1453 5347 1467
rect 5453 1452 5467 1466
rect 5493 1453 5507 1467
rect 5573 1453 5587 1467
rect 5653 1453 5667 1467
rect 5773 1453 5787 1467
rect 5813 1453 5827 1467
rect 1853 1393 1867 1407
rect 1913 1393 1927 1407
rect 2193 1393 2207 1407
rect 2233 1393 2247 1407
rect 2493 1393 2507 1407
rect 5093 1433 5107 1447
rect 5133 1433 5147 1447
rect 5573 1432 5587 1446
rect 5613 1433 5627 1447
rect 4513 1393 4527 1407
rect 5133 1393 5147 1407
rect 553 1372 567 1386
rect 5073 1373 5087 1387
rect 5693 1373 5707 1387
rect 5773 1373 5787 1387
rect 4733 1353 4747 1367
rect 4793 1353 4807 1367
rect 4553 1253 4567 1267
rect 4613 1253 4627 1267
rect 4493 1233 4507 1247
rect 4633 1233 4647 1247
rect 5533 1233 5547 1247
rect 5593 1233 5607 1247
rect 2953 1213 2967 1227
rect 3813 1213 3827 1227
rect 3853 1213 3867 1227
rect 4773 1213 4787 1227
rect 4833 1213 4847 1227
rect 4993 1213 5007 1227
rect 5473 1213 5487 1227
rect 5553 1213 5567 1227
rect 5713 1213 5727 1227
rect 553 1173 567 1187
rect 593 1173 607 1187
rect 2953 1173 2967 1187
rect 4993 1173 5007 1187
rect 5473 1173 5487 1187
rect 5613 1173 5627 1187
rect 5693 1173 5707 1187
rect 293 1153 307 1167
rect 353 1153 367 1167
rect 1673 1153 1687 1167
rect 1753 1153 1767 1167
rect 2493 1153 2507 1167
rect 2613 1153 2627 1167
rect 2993 1153 3007 1167
rect 3033 1153 3047 1167
rect 3073 1153 3087 1167
rect 3113 1153 3127 1167
rect 3233 1153 3247 1167
rect 3333 1153 3347 1167
rect 4593 1153 4607 1167
rect 4673 1153 4687 1167
rect 5053 1153 5067 1167
rect 5113 1153 5127 1167
rect 5353 1153 5367 1167
rect 5433 1153 5447 1167
rect 5493 1153 5507 1167
rect 1833 953 1847 967
rect 1893 953 1907 967
rect 2213 953 2227 967
rect 2273 953 2287 967
rect 353 933 367 947
rect 433 933 447 947
rect 1253 933 1267 947
rect 1293 934 1307 948
rect 3553 933 3567 947
rect 3653 934 3667 948
rect 4653 933 4667 947
rect 4753 933 4767 947
rect 5213 933 5227 947
rect 5273 933 5287 947
rect 5473 933 5487 947
rect 1393 913 1407 927
rect 1433 913 1447 927
rect 2353 913 2367 927
rect 2393 913 2407 927
rect 1853 873 1867 887
rect 1893 873 1907 887
rect 5613 933 5627 947
rect 5693 933 5707 947
rect 5873 933 5887 947
rect 5913 933 5927 947
rect 813 853 827 867
rect 853 853 867 867
rect 1353 853 1367 867
rect 1413 853 1427 867
rect 3073 853 3087 867
rect 3173 853 3187 867
rect 5473 851 5487 865
rect 393 713 407 727
rect 3453 713 3467 727
rect 3493 713 3507 727
rect 4173 714 4187 728
rect 4213 713 4227 727
rect 5213 713 5227 727
rect 5293 713 5307 727
rect 5753 673 5767 687
rect 413 653 427 667
rect 5733 653 5747 667
rect 133 633 147 647
rect 233 633 247 647
rect 313 633 327 647
rect 913 633 927 647
rect 953 633 967 647
rect 3453 633 3467 647
rect 3513 631 3527 645
rect 4293 633 4307 647
rect 4413 633 4427 647
rect 413 613 427 627
rect 473 612 487 626
rect 3253 613 3267 627
rect 3313 613 3327 627
rect 4353 433 4367 447
rect 4393 433 4407 447
rect 1193 413 1207 427
rect 1333 413 1347 427
rect 3693 413 3707 427
rect 3773 413 3787 427
rect 2033 393 2047 407
rect 2073 393 2087 407
rect 4473 333 4487 347
rect 4533 333 4547 347
rect 473 193 487 207
rect 533 193 547 207
rect 1493 173 1507 187
rect 1533 173 1547 187
rect 1293 113 1307 127
rect 1413 113 1427 127
rect 2713 113 2727 127
rect 2773 113 2787 127
rect 3953 113 3967 127
rect 4033 113 4047 127
rect 5413 93 5427 107
rect 5453 92 5467 106
rect 2613 53 2627 67
rect 2653 53 2667 67
<< metal2 >>
rect 136 6036 163 6043
rect 156 5947 163 6036
rect 416 6007 423 6043
rect 876 6007 883 6043
rect 156 5896 163 5933
rect 16 5547 23 5573
rect 96 5560 103 5563
rect 93 5547 107 5560
rect 176 5527 183 5853
rect 296 5667 303 5863
rect 356 5608 363 5893
rect 376 5863 383 5993
rect 876 5866 883 5993
rect 1056 5987 1063 6043
rect 376 5856 403 5863
rect 596 5860 603 5863
rect 593 5847 607 5860
rect 1016 5863 1023 5973
rect 1016 5856 1043 5863
rect 796 5687 803 5852
rect 367 5596 383 5603
rect 516 5596 523 5653
rect 676 5596 683 5653
rect 176 5427 183 5513
rect 136 5376 143 5413
rect 196 5346 203 5593
rect 256 5467 263 5563
rect 116 4947 123 5043
rect 133 4860 147 4873
rect 156 4867 163 5343
rect 216 5307 223 5373
rect 276 5340 283 5343
rect 236 5127 243 5333
rect 273 5327 287 5340
rect 316 5327 323 5343
rect 296 5316 313 5323
rect 296 5303 303 5316
rect 267 5296 303 5303
rect 276 5076 283 5113
rect 356 5046 363 5413
rect 396 5388 403 5563
rect 456 5547 463 5593
rect 536 5527 543 5552
rect 516 5387 523 5413
rect 576 5407 583 5563
rect 736 5527 743 5563
rect 616 5407 623 5453
rect 636 5407 643 5433
rect 696 5407 703 5493
rect 796 5487 803 5594
rect 580 5386 600 5387
rect 436 5340 443 5343
rect 476 5340 483 5343
rect 433 5327 447 5340
rect 473 5327 487 5340
rect 516 5076 523 5253
rect 256 4987 263 5043
rect 136 4856 143 4860
rect 173 4860 187 4873
rect 176 4856 183 4860
rect 396 4826 403 4933
rect 296 4820 303 4823
rect 156 4667 163 4813
rect 293 4807 307 4820
rect 13 4567 27 4573
rect 96 4568 103 4653
rect 133 4560 147 4573
rect 136 4556 143 4560
rect 16 4307 23 4553
rect 113 4507 127 4512
rect 116 4336 123 4493
rect 156 4427 163 4523
rect 176 4467 183 4513
rect 16 4107 23 4253
rect 96 4227 103 4303
rect 196 4267 203 4593
rect 216 4223 223 4453
rect 236 4343 243 4513
rect 276 4487 283 4523
rect 356 4523 363 4823
rect 336 4516 363 4523
rect 256 4348 263 4373
rect 236 4336 253 4343
rect 336 4303 343 4516
rect 376 4427 383 4533
rect 396 4487 403 4812
rect 416 4787 423 5043
rect 536 5027 543 5313
rect 496 4856 503 4893
rect 556 4887 563 5373
rect 587 5383 600 5386
rect 587 5376 603 5383
rect 633 5380 647 5393
rect 636 5376 643 5380
rect 587 5373 600 5376
rect 696 5346 703 5393
rect 796 5388 803 5473
rect 836 5383 843 5433
rect 856 5427 863 5513
rect 876 5507 883 5563
rect 956 5527 963 5813
rect 1196 5707 1203 5993
rect 1216 5856 1243 5863
rect 1216 5807 1223 5856
rect 1416 5860 1423 5863
rect 1356 5827 1363 5852
rect 1413 5847 1427 5860
rect 976 5567 983 5633
rect 1256 5596 1263 5673
rect 836 5376 863 5383
rect 576 5047 583 5293
rect 716 5087 723 5373
rect 856 5346 863 5376
rect 876 5327 883 5374
rect 976 5347 983 5473
rect 1036 5447 1043 5563
rect 1076 5527 1083 5563
rect 996 5346 1003 5413
rect 1136 5343 1143 5433
rect 1096 5336 1143 5343
rect 1156 5307 1163 5473
rect 1176 5387 1183 5433
rect 1196 5407 1203 5533
rect 1216 5376 1223 5473
rect 1256 5307 1263 5343
rect 1176 5247 1183 5273
rect 596 4927 603 5074
rect 636 4927 643 5043
rect 536 4856 583 4863
rect 476 4767 483 4812
rect 556 4767 563 4793
rect 576 4767 583 4856
rect 596 4826 603 4873
rect 656 4856 663 4893
rect 676 4820 683 4823
rect 673 4807 687 4820
rect 736 4787 743 5074
rect 756 4907 763 5073
rect 876 5046 883 5153
rect 836 5036 863 5043
rect 836 4856 843 5013
rect 856 4967 863 5036
rect 436 4556 443 4593
rect 476 4556 483 4613
rect 376 4336 383 4413
rect 456 4343 463 4512
rect 516 4343 523 4613
rect 456 4336 483 4343
rect 476 4306 483 4336
rect 496 4336 523 4343
rect 536 4336 543 4413
rect 336 4296 363 4303
rect 216 4216 233 4223
rect 16 3347 23 4093
rect 136 3996 183 4003
rect 136 3816 143 3853
rect 176 3816 183 3913
rect 236 3387 243 4213
rect 356 4087 363 4296
rect 496 4107 503 4336
rect 616 4306 623 4333
rect 556 4287 563 4303
rect 556 4276 573 4287
rect 560 4273 573 4276
rect 356 4036 363 4073
rect 256 3927 263 4033
rect 76 3263 83 3293
rect 256 3267 263 3873
rect 396 3787 403 4073
rect 436 3847 443 4033
rect 516 3907 523 4003
rect 556 3947 563 4093
rect 636 4087 643 4773
rect 656 4347 663 4553
rect 676 4526 683 4753
rect 756 4667 763 4853
rect 896 4826 903 5233
rect 936 5076 943 5153
rect 1116 5076 1123 5113
rect 816 4820 823 4823
rect 813 4807 827 4820
rect 776 4507 783 4793
rect 856 4627 863 4812
rect 853 4568 867 4573
rect 896 4556 903 4593
rect 916 4567 923 4993
rect 956 4947 963 5043
rect 976 4856 983 4993
rect 996 4987 1003 5073
rect 956 4767 963 4823
rect 956 4687 963 4753
rect 976 4667 983 4693
rect 696 4336 703 4373
rect 736 4336 743 4373
rect 716 4300 723 4303
rect 713 4287 727 4300
rect 776 4187 783 4493
rect 836 4487 843 4523
rect 936 4487 943 4653
rect 956 4526 963 4652
rect 996 4607 1003 4823
rect 1056 4767 1063 5043
rect 1076 4827 1083 4933
rect 1013 4560 1027 4573
rect 1016 4556 1023 4560
rect 1036 4427 1043 4523
rect 1076 4467 1083 4513
rect 876 4336 883 4373
rect 1016 4336 1023 4373
rect 796 4287 803 4333
rect 856 4300 863 4303
rect 816 4247 823 4293
rect 853 4287 867 4300
rect 996 4300 1003 4303
rect 993 4287 1007 4300
rect 1036 4283 1043 4292
rect 1016 4276 1043 4283
rect 576 4006 583 4033
rect 636 4000 643 4003
rect 633 3987 647 4000
rect 473 3820 487 3833
rect 513 3820 527 3833
rect 476 3816 483 3820
rect 516 3816 523 3820
rect 556 3816 563 3873
rect 296 3763 303 3783
rect 276 3756 303 3763
rect 276 3727 283 3756
rect 356 3528 363 3772
rect 496 3727 503 3783
rect 533 3520 547 3533
rect 596 3528 603 3653
rect 536 3516 543 3520
rect 636 3387 643 3933
rect 696 3907 703 4034
rect 736 3847 743 4013
rect 776 4000 783 4003
rect 773 3987 787 4000
rect 856 3967 863 4073
rect 876 4047 883 4133
rect 913 4067 927 4073
rect 916 4036 923 4053
rect 736 3667 743 3783
rect 756 3516 763 3553
rect 796 3543 803 3953
rect 896 3887 903 4003
rect 936 3947 943 3992
rect 996 3987 1003 4053
rect 816 3587 823 3833
rect 856 3816 863 3873
rect 996 3816 1003 3973
rect 1016 3927 1023 4276
rect 1096 4207 1103 4873
rect 1136 4856 1143 4913
rect 1156 4887 1163 5193
rect 1216 5076 1223 5113
rect 1276 5103 1283 5413
rect 1296 5207 1303 5793
rect 1256 5096 1283 5103
rect 1256 5088 1263 5096
rect 1236 5007 1243 5043
rect 1116 4507 1123 4812
rect 1196 4667 1203 4693
rect 1136 4567 1143 4653
rect 1216 4556 1223 4673
rect 1196 4487 1203 4523
rect 1116 4347 1123 4373
rect 1216 4336 1223 4493
rect 1236 4487 1243 4513
rect 1256 4507 1263 4933
rect 1276 4907 1283 5043
rect 1316 4947 1323 5693
rect 1356 5687 1363 5813
rect 1396 5596 1403 5633
rect 1376 5427 1383 5563
rect 1416 5487 1423 5563
rect 1336 5167 1343 5333
rect 1376 5108 1383 5343
rect 1416 5307 1423 5332
rect 1456 5227 1463 5373
rect 1476 5247 1483 5933
rect 1676 5927 1683 6043
rect 2296 5967 2303 6043
rect 2336 6036 2363 6043
rect 1816 5896 1863 5903
rect 1576 5596 1583 5633
rect 1496 5487 1503 5594
rect 1656 5587 1663 5833
rect 1756 5596 1763 5633
rect 1796 5608 1803 5863
rect 1856 5707 1863 5896
rect 1876 5787 1883 5894
rect 2356 5863 2363 6036
rect 2576 6036 2603 6043
rect 2636 6036 2663 6043
rect 1936 5860 1943 5863
rect 1933 5847 1947 5860
rect 1976 5827 1983 5863
rect 2036 5843 2043 5863
rect 2336 5856 2363 5863
rect 2036 5836 2063 5843
rect 1936 5647 1943 5773
rect 1936 5596 1943 5633
rect 1556 5307 1563 5333
rect 1336 4967 1343 5093
rect 1413 5080 1427 5093
rect 1416 5076 1423 5080
rect 1496 5047 1503 5173
rect 1516 5167 1523 5273
rect 1556 5267 1563 5293
rect 1556 5076 1563 5193
rect 1576 5127 1583 5373
rect 1596 5107 1603 5563
rect 1736 5467 1743 5563
rect 1676 5376 1683 5413
rect 1736 5346 1743 5432
rect 1616 5207 1623 5313
rect 1656 5287 1663 5343
rect 1756 5327 1763 5373
rect 1776 5346 1783 5433
rect 1853 5403 1867 5413
rect 1876 5403 1883 5563
rect 1916 5543 1923 5563
rect 1916 5536 1943 5543
rect 1853 5400 1883 5403
rect 1856 5396 1883 5400
rect 1856 5376 1863 5396
rect 1916 5347 1923 5453
rect 1936 5447 1943 5536
rect 1976 5447 1983 5594
rect 1996 5566 2003 5693
rect 2056 5687 2063 5836
rect 2076 5608 2083 5833
rect 2316 5647 2323 5813
rect 2336 5667 2343 5833
rect 2376 5747 2383 5953
rect 2493 5900 2507 5913
rect 2496 5896 2503 5900
rect 2416 5787 2423 5893
rect 2476 5860 2483 5863
rect 2516 5860 2523 5863
rect 2473 5847 2487 5860
rect 2513 5847 2527 5860
rect 2533 5847 2547 5852
rect 2316 5596 2323 5633
rect 1996 5427 2003 5552
rect 2056 5487 2063 5563
rect 2196 5507 2203 5593
rect 2216 5547 2223 5594
rect 2436 5566 2443 5673
rect 2036 5376 2043 5413
rect 1936 5346 1943 5373
rect 1967 5343 1980 5347
rect 2076 5346 2083 5493
rect 2096 5347 2103 5433
rect 2136 5388 2143 5453
rect 2316 5416 2323 5533
rect 2456 5487 2463 5733
rect 2556 5707 2563 5893
rect 2576 5867 2583 6036
rect 2656 5908 2663 6036
rect 2796 5987 2803 6043
rect 2676 5860 2683 5863
rect 2673 5847 2687 5860
rect 2716 5747 2723 5894
rect 2756 5863 2763 5973
rect 2756 5856 2783 5863
rect 2976 5843 2983 5863
rect 2956 5836 2983 5843
rect 2736 5767 2743 5793
rect 2556 5667 2563 5693
rect 2556 5596 2563 5632
rect 2716 5596 2723 5653
rect 2756 5596 2763 5773
rect 2956 5667 2963 5836
rect 3036 5807 3043 5863
rect 2976 5596 3003 5603
rect 3096 5596 3103 5993
rect 2356 5376 2383 5383
rect 1967 5336 1983 5343
rect 1967 5333 1980 5336
rect 2376 5346 2383 5376
rect 2236 5336 2263 5343
rect 1876 5287 1883 5332
rect 1616 5147 1623 5193
rect 1616 5083 1623 5112
rect 1596 5076 1623 5083
rect 1336 4883 1343 4953
rect 1316 4876 1343 4883
rect 1316 4856 1323 4876
rect 1376 4826 1383 4853
rect 1287 4816 1303 4823
rect 1276 4427 1283 4812
rect 1396 4747 1403 5032
rect 1536 5023 1543 5043
rect 1536 5020 1563 5023
rect 1533 5016 1563 5020
rect 1533 5007 1547 5016
rect 1496 4907 1503 4953
rect 1496 4856 1503 4893
rect 1436 4687 1443 4823
rect 1296 4547 1303 4573
rect 1316 4556 1323 4593
rect 1456 4526 1463 4753
rect 1476 4727 1483 4823
rect 1516 4820 1523 4823
rect 1513 4807 1527 4820
rect 1493 4560 1507 4573
rect 1536 4568 1543 4813
rect 1556 4787 1563 5016
rect 1576 4807 1583 4913
rect 1636 4887 1643 5093
rect 1656 4947 1663 5233
rect 1676 5047 1683 5193
rect 1616 4876 1633 4883
rect 1616 4856 1623 4876
rect 1696 4883 1703 5133
rect 1716 5076 1723 5233
rect 1956 5167 1963 5273
rect 1773 5080 1787 5093
rect 1913 5088 1927 5093
rect 1776 5076 1783 5080
rect 2053 5080 2067 5093
rect 2056 5076 2063 5080
rect 2156 5076 2163 5233
rect 2236 5227 2243 5336
rect 2376 5247 2383 5332
rect 2416 5227 2423 5473
rect 2476 5376 2483 5413
rect 2616 5388 2623 5552
rect 2716 5427 2723 5533
rect 2716 5383 2723 5413
rect 2736 5407 2743 5563
rect 2856 5527 2863 5593
rect 2996 5487 3003 5596
rect 2716 5376 2743 5383
rect 2916 5376 2923 5473
rect 2496 5307 2503 5343
rect 2596 5340 2603 5343
rect 2593 5327 2607 5340
rect 2636 5336 2663 5343
rect 2216 5167 2223 5193
rect 2196 5076 2203 5133
rect 2436 5127 2443 5273
rect 2240 5083 2253 5087
rect 2236 5076 2253 5083
rect 1736 5040 1743 5043
rect 1733 5027 1747 5040
rect 1836 5027 1843 5074
rect 1896 5027 1903 5043
rect 1696 4876 1723 4883
rect 1716 4826 1723 4876
rect 1676 4787 1683 4823
rect 1656 4683 1663 4713
rect 1676 4707 1683 4773
rect 1656 4676 1693 4683
rect 1496 4556 1503 4560
rect 1693 4560 1707 4573
rect 1736 4563 1743 4933
rect 1773 4860 1787 4873
rect 1816 4868 1823 4913
rect 1856 4887 1863 4953
rect 1876 4947 1883 5013
rect 1896 4987 1903 5013
rect 1776 4856 1783 4860
rect 1836 4747 1843 4823
rect 1756 4667 1763 4713
rect 1696 4556 1703 4560
rect 1736 4556 1763 4563
rect 1296 4487 1303 4512
rect 1336 4467 1343 4523
rect 1556 4447 1563 4523
rect 1756 4507 1763 4556
rect 1796 4527 1803 4653
rect 1836 4647 1843 4733
rect 1876 4687 1883 4893
rect 1936 4856 1943 4893
rect 1976 4856 1983 5074
rect 2240 5073 2253 5076
rect 2396 5076 2403 5113
rect 2176 5040 2183 5043
rect 2173 5027 2187 5040
rect 2316 5007 2323 5073
rect 2456 5047 2463 5253
rect 2376 4987 2383 5032
rect 2476 4967 2483 5213
rect 2516 5076 2523 5233
rect 2056 4826 2063 4853
rect 1856 4556 1863 4593
rect 1896 4547 1903 4793
rect 1956 4667 1963 4823
rect 1996 4820 2003 4823
rect 1993 4807 2007 4820
rect 1816 4520 1823 4523
rect 1813 4507 1827 4520
rect 1896 4507 1903 4533
rect 1536 4348 1543 4373
rect 1116 4306 1123 4333
rect 1136 4207 1143 4334
rect 1327 4343 1340 4347
rect 1327 4336 1343 4343
rect 1327 4333 1340 4336
rect 1236 4247 1243 4303
rect 1276 4247 1283 4333
rect 1356 4300 1363 4303
rect 1353 4287 1367 4300
rect 1116 4107 1123 4173
rect 1156 4167 1163 4193
rect 1033 4067 1047 4073
rect 1073 4048 1087 4053
rect 1116 4036 1123 4072
rect 1156 4007 1163 4053
rect 1056 4000 1063 4003
rect 1053 3987 1067 4000
rect 1096 3947 1103 4003
rect 1176 3967 1183 4233
rect 1207 4093 1213 4107
rect 1236 4036 1243 4073
rect 1256 3967 1263 4003
rect 1056 3816 1063 3853
rect 936 3787 943 3814
rect 796 3536 813 3543
rect 816 3486 823 3533
rect 896 3516 903 3573
rect 1076 3516 1083 3573
rect 736 3447 743 3483
rect 876 3447 883 3483
rect 76 3256 103 3263
rect 16 3227 23 3253
rect 296 3067 303 3153
rect 356 3083 363 3263
rect 356 3076 373 3083
rect 296 3003 303 3053
rect 296 2996 323 3003
rect 376 2996 383 3073
rect 436 3027 443 3333
rect 536 3296 543 3333
rect 596 3266 603 3373
rect 976 3367 983 3514
rect 1136 3483 1143 3913
rect 1156 3776 1183 3783
rect 1156 3707 1163 3776
rect 1236 3667 1243 3783
rect 1276 3767 1283 3893
rect 1193 3520 1207 3533
rect 1196 3516 1203 3520
rect 1116 3476 1143 3483
rect 676 3296 683 3333
rect 936 3296 943 3353
rect 516 3260 523 3263
rect 513 3247 527 3260
rect 513 3227 527 3233
rect 616 3127 623 3293
rect 696 3260 703 3263
rect 693 3247 707 3260
rect 16 2867 23 2953
rect 436 2847 443 2963
rect 16 2747 23 2813
rect 276 2776 283 2833
rect 413 2780 427 2793
rect 416 2776 423 2780
rect 76 2743 83 2773
rect 76 2736 103 2743
rect 236 2740 243 2743
rect 233 2727 247 2740
rect 516 2527 523 3073
rect 553 3000 567 3013
rect 556 2996 563 3000
rect 616 2996 623 3073
rect 716 2966 723 3113
rect 776 3047 783 3293
rect 836 2966 843 3033
rect 916 2927 923 2963
rect 693 2780 707 2793
rect 696 2776 703 2780
rect 956 2747 963 2953
rect 976 2927 983 3233
rect 996 2967 1003 3263
rect 1036 3127 1043 3273
rect 1056 3247 1063 3472
rect 1036 2996 1043 3113
rect 1116 3063 1123 3476
rect 1136 3087 1143 3263
rect 1116 3056 1143 3063
rect 1076 2996 1083 3033
rect 996 2776 1003 2932
rect 1056 2927 1063 2963
rect 1096 2960 1103 2963
rect 1093 2947 1107 2960
rect 1136 2927 1143 3056
rect 1196 2996 1203 3373
rect 1296 3266 1303 3533
rect 1316 3363 1323 4153
rect 1336 3823 1343 4213
rect 1376 4207 1383 4233
rect 1376 4036 1383 4193
rect 1396 4087 1403 4173
rect 1416 4147 1423 4333
rect 1476 4247 1483 4303
rect 1516 4300 1523 4303
rect 1513 4287 1527 4300
rect 1436 4006 1443 4033
rect 1496 4000 1503 4003
rect 1396 3823 1403 3992
rect 1493 3987 1507 4000
rect 1336 3816 1363 3823
rect 1396 3820 1423 3823
rect 1396 3816 1427 3820
rect 1413 3807 1427 3816
rect 1436 3787 1443 3833
rect 1473 3820 1487 3833
rect 1476 3816 1483 3820
rect 1536 3827 1543 3992
rect 1496 3780 1503 3783
rect 1493 3767 1507 3780
rect 1336 3516 1343 3653
rect 1556 3627 1563 3814
rect 1453 3520 1467 3533
rect 1456 3516 1463 3520
rect 1316 3356 1343 3363
rect 1216 2960 1223 2963
rect 1213 2947 1227 2960
rect 576 2740 583 2743
rect 573 2727 587 2740
rect 636 2687 643 2743
rect 816 2740 823 2743
rect 813 2727 827 2740
rect 596 2527 603 2613
rect 96 2476 103 2513
rect 356 2476 363 2513
rect 596 2476 603 2513
rect 716 2507 723 2533
rect 756 2507 763 2713
rect 876 2627 883 2743
rect 1296 2746 1303 3252
rect 1316 3247 1323 3333
rect 1336 3147 1343 3356
rect 1356 3047 1363 3353
rect 1476 3263 1483 3453
rect 1496 3267 1503 3294
rect 1396 3260 1403 3263
rect 1393 3247 1407 3260
rect 1456 3256 1483 3263
rect 1356 2996 1363 3033
rect 1396 2966 1403 3073
rect 1336 2907 1343 2963
rect 1336 2867 1343 2893
rect 1396 2788 1403 2952
rect 1416 2783 1423 3033
rect 1456 3008 1463 3153
rect 1496 3087 1503 3253
rect 1516 3063 1523 3593
rect 1576 3547 1583 4493
rect 1616 4087 1623 4493
rect 1796 4336 1803 4473
rect 1676 4187 1683 4303
rect 1716 4043 1723 4333
rect 1876 4307 1883 4453
rect 1816 4247 1823 4303
rect 1696 4036 1723 4043
rect 1596 3987 1603 4034
rect 1636 3927 1643 4003
rect 1676 3947 1683 4003
rect 1636 3816 1643 3873
rect 1696 3828 1703 3913
rect 1696 3783 1703 3814
rect 1616 3516 1623 3693
rect 1636 3486 1643 3753
rect 1656 3747 1663 3783
rect 1676 3776 1703 3783
rect 1596 3260 1603 3263
rect 1593 3247 1607 3260
rect 1536 3107 1543 3233
rect 1636 3227 1643 3293
rect 1656 3167 1663 3433
rect 1676 3307 1683 3776
rect 1736 3767 1743 4073
rect 1756 4027 1763 4193
rect 1813 4040 1827 4053
rect 1816 4036 1823 4040
rect 1856 4036 1863 4113
rect 1876 4047 1883 4272
rect 1836 3967 1843 4003
rect 1836 3747 1843 3772
rect 1876 3767 1883 3973
rect 1896 3887 1903 4493
rect 1916 4427 1923 4554
rect 1936 4523 1943 4633
rect 2016 4556 2023 4653
rect 2076 4567 2083 4913
rect 2133 4860 2147 4873
rect 2136 4856 2143 4860
rect 2276 4856 2283 4933
rect 2316 4856 2323 4913
rect 2236 4826 2243 4853
rect 2156 4727 2163 4823
rect 2336 4820 2343 4823
rect 2293 4807 2307 4812
rect 2333 4807 2347 4820
rect 2376 4807 2383 4854
rect 1936 4516 1963 4523
rect 1956 4336 1963 4516
rect 1996 4447 2003 4523
rect 2036 4520 2043 4523
rect 2033 4507 2047 4520
rect 2116 4387 2123 4593
rect 2176 4556 2183 4793
rect 2396 4787 2403 4953
rect 2536 4947 2543 5043
rect 2576 5040 2583 5043
rect 2573 5027 2587 5040
rect 2436 4820 2443 4823
rect 2433 4807 2447 4820
rect 2476 4787 2483 4823
rect 2216 4687 2223 4773
rect 2156 4520 2163 4523
rect 2153 4507 2167 4520
rect 2216 4487 2223 4554
rect 2093 4340 2107 4353
rect 2096 4336 2103 4340
rect 1916 4296 1943 4303
rect 1976 4300 1983 4303
rect 1916 4007 1923 4296
rect 1973 4287 1987 4300
rect 2076 4267 2083 4303
rect 2116 4300 2123 4303
rect 2113 4287 2127 4300
rect 2096 4276 2113 4283
rect 1916 3827 1923 3972
rect 1936 3947 1943 4073
rect 2033 4040 2047 4053
rect 2036 4036 2043 4040
rect 2076 4003 2083 4253
rect 1956 3847 1963 3953
rect 2016 3947 2023 4003
rect 2056 3996 2083 4003
rect 1976 3816 1983 3873
rect 1936 3727 1943 3783
rect 2036 3767 2043 3813
rect 2056 3727 2063 3996
rect 2096 3887 2103 4276
rect 2156 4207 2163 4353
rect 2176 4267 2183 4473
rect 2236 4336 2243 4693
rect 2316 4587 2323 4773
rect 2313 4560 2327 4573
rect 2316 4556 2323 4560
rect 2296 4348 2303 4523
rect 2356 4343 2363 4633
rect 2376 4447 2383 4713
rect 2396 4527 2403 4593
rect 2336 4336 2363 4343
rect 2373 4340 2387 4353
rect 2376 4336 2383 4340
rect 2416 4336 2423 4453
rect 2296 4306 2303 4334
rect 2216 4267 2223 4303
rect 2176 4187 2183 4253
rect 2216 4083 2223 4253
rect 2216 4076 2243 4083
rect 2136 4036 2143 4073
rect 2213 4047 2227 4053
rect 2116 3816 2123 3993
rect 2196 4000 2203 4003
rect 2193 3987 2207 4000
rect 2236 3987 2243 4076
rect 2136 3907 2143 3973
rect 2256 3967 2263 4303
rect 2336 4227 2343 4336
rect 2296 4048 2303 4113
rect 2273 3987 2287 3993
rect 2256 3816 2263 3853
rect 2296 3816 2303 3953
rect 2316 3847 2323 3992
rect 2327 3836 2343 3843
rect 2336 3807 2343 3836
rect 2136 3747 2143 3783
rect 2276 3780 2283 3783
rect 2273 3767 2287 3780
rect 2356 3767 2363 4073
rect 2396 4043 2403 4303
rect 2416 4147 2423 4273
rect 2476 4183 2483 4512
rect 2496 4207 2503 4573
rect 2516 4526 2523 4553
rect 2536 4387 2543 4912
rect 2616 4856 2623 4973
rect 2636 4927 2643 5313
rect 2656 5307 2663 5336
rect 2656 5127 2663 5293
rect 2716 5076 2723 5233
rect 2736 5127 2743 5153
rect 2756 5147 2763 5343
rect 2776 5167 2783 5293
rect 2796 5267 2803 5343
rect 2856 5307 2863 5374
rect 2856 5187 2863 5272
rect 2896 5267 2903 5343
rect 2936 5340 2943 5343
rect 2933 5327 2947 5340
rect 2856 5076 2863 5173
rect 2656 4856 2663 5013
rect 2696 4947 2703 5032
rect 2556 4826 2563 4853
rect 2716 4827 2723 4913
rect 2736 4868 2743 5043
rect 2776 4967 2783 4993
rect 2796 4987 2803 5074
rect 2956 5007 2963 5333
rect 2976 5147 2983 5374
rect 3056 5327 3063 5343
rect 3047 5316 3063 5327
rect 3047 5313 3060 5316
rect 3096 5247 3103 5373
rect 3136 5347 3143 6043
rect 3336 6007 3343 6043
rect 3976 6007 3983 6043
rect 3196 5896 3203 5973
rect 3156 5860 3163 5863
rect 3153 5847 3167 5860
rect 3156 5787 3163 5833
rect 2996 5088 3003 5193
rect 3036 5076 3043 5113
rect 2776 4856 2783 4953
rect 2796 4927 2803 4973
rect 2967 4874 2973 4887
rect 2967 4873 2980 4874
rect 2636 4787 2643 4823
rect 2876 4826 2883 4873
rect 3016 4867 3023 4993
rect 2656 4556 2673 4563
rect 2596 4447 2603 4483
rect 2676 4467 2683 4554
rect 2736 4526 2743 4593
rect 2676 4367 2683 4453
rect 2756 4447 2763 4813
rect 2796 4727 2803 4823
rect 2896 4787 2903 4853
rect 2956 4707 2963 4823
rect 2896 4487 2903 4693
rect 3036 4647 3043 4913
rect 3056 4887 3063 5043
rect 3096 4927 3103 5093
rect 3116 5046 3123 5193
rect 3156 5167 3163 5613
rect 3176 5566 3183 5653
rect 3216 5627 3223 5793
rect 3213 5600 3227 5613
rect 3216 5596 3223 5600
rect 3236 5383 3243 5973
rect 3296 5863 3303 5993
rect 3296 5856 3323 5863
rect 3516 5843 3523 5863
rect 3696 5860 3703 5863
rect 3496 5836 3523 5843
rect 3453 5600 3467 5613
rect 3456 5596 3463 5600
rect 3496 5527 3503 5836
rect 3576 5627 3583 5852
rect 3693 5847 3707 5860
rect 3793 5600 3807 5613
rect 3796 5596 3803 5600
rect 3576 5507 3583 5563
rect 3216 5376 3243 5383
rect 3176 5107 3183 5343
rect 3196 5076 3203 5113
rect 3087 4883 3100 4887
rect 3087 4873 3103 4883
rect 3096 4856 3103 4873
rect 3136 4868 3143 4913
rect 3056 4767 3063 4852
rect 3016 4556 3023 4593
rect 2916 4467 2923 4554
rect 3076 4526 3083 4773
rect 3116 4556 3123 4753
rect 3156 4707 3163 4823
rect 3196 4647 3203 4993
rect 3216 4963 3223 5043
rect 3256 5027 3263 5153
rect 3276 5047 3283 5493
rect 3316 5127 3323 5343
rect 3356 5340 3363 5343
rect 3353 5327 3367 5340
rect 3416 5327 3423 5374
rect 3436 5346 3443 5473
rect 3496 5407 3503 5453
rect 3616 5427 3623 5563
rect 3656 5447 3663 5594
rect 3433 5327 3447 5332
rect 3336 5107 3343 5293
rect 3536 5287 3543 5343
rect 3333 5080 3347 5093
rect 3336 5076 3343 5080
rect 3376 5076 3383 5133
rect 3473 5080 3487 5093
rect 3476 5076 3483 5080
rect 3516 5076 3523 5133
rect 3576 5043 3583 5374
rect 3596 5346 3603 5393
rect 3656 5376 3663 5433
rect 3356 5040 3363 5043
rect 3353 5027 3367 5040
rect 3496 5027 3503 5043
rect 3216 4956 3243 4963
rect 3216 4826 3223 4933
rect 3236 4867 3243 4956
rect 3256 4856 3263 4973
rect 3293 4860 3307 4873
rect 3336 4867 3343 4933
rect 3296 4856 3303 4860
rect 3356 4826 3363 4913
rect 3376 4767 3383 4933
rect 3436 4856 3443 4913
rect 3156 4520 3163 4523
rect 3196 4520 3203 4523
rect 3153 4507 3167 4520
rect 3193 4507 3207 4520
rect 3256 4447 3263 4753
rect 3476 4667 3483 4873
rect 3376 4556 3383 4633
rect 3416 4607 3423 4633
rect 3496 4627 3503 5013
rect 3516 4867 3523 4993
rect 3536 4907 3543 5043
rect 3556 5036 3583 5043
rect 3556 4868 3563 5036
rect 3596 4947 3603 5332
rect 3676 5307 3683 5343
rect 3636 5083 3643 5293
rect 3716 5167 3723 5513
rect 3736 5487 3743 5563
rect 3776 5507 3783 5563
rect 3836 5447 3843 5594
rect 3616 5076 3643 5083
rect 3616 5007 3623 5076
rect 3676 5023 3683 5043
rect 3656 5016 3683 5023
rect 3656 4947 3663 5016
rect 3676 4967 3683 4993
rect 3616 4863 3623 4893
rect 3616 4856 3643 4863
rect 3276 4507 3283 4553
rect 3436 4520 3443 4523
rect 3433 4507 3447 4520
rect 3516 4487 3523 4813
rect 3536 4707 3543 4823
rect 3616 4667 3623 4813
rect 3616 4556 3623 4593
rect 3636 4587 3643 4856
rect 3656 4767 3663 4893
rect 3716 4856 3723 5132
rect 3736 4907 3743 5413
rect 3856 5407 3863 5913
rect 4016 5863 4023 5993
rect 3996 5856 4023 5863
rect 4056 5767 4063 5993
rect 4096 5927 4103 6043
rect 4596 6036 4623 6043
rect 4133 5908 4147 5913
rect 4616 5908 4623 6036
rect 5236 6007 5243 6043
rect 4096 5860 4103 5863
rect 4093 5847 4107 5860
rect 4296 5747 4303 5863
rect 4376 5847 4383 5894
rect 4736 5896 4743 5933
rect 4356 5836 4373 5843
rect 3913 5600 3927 5613
rect 3916 5596 3923 5600
rect 3793 5380 3807 5393
rect 3796 5376 3803 5380
rect 3776 5307 3783 5343
rect 3816 5340 3823 5343
rect 3813 5327 3827 5340
rect 3856 5323 3863 5343
rect 3836 5316 3863 5323
rect 3836 5287 3843 5316
rect 3876 5303 3883 5333
rect 3867 5296 3883 5303
rect 3756 4967 3763 5153
rect 3856 5076 3863 5293
rect 3896 5207 3903 5563
rect 3936 5507 3943 5563
rect 3996 5527 4003 5613
rect 4116 5596 4123 5633
rect 4036 5467 4043 5594
rect 4176 5566 4183 5673
rect 4096 5527 4103 5563
rect 4176 5467 4183 5513
rect 3756 4856 3763 4913
rect 3776 4867 3783 4993
rect 3736 4820 3743 4823
rect 3733 4807 3747 4820
rect 3756 4556 3763 4753
rect 3796 4567 3803 4953
rect 3916 4887 3923 5393
rect 3956 5376 3963 5433
rect 3993 5380 4007 5393
rect 3996 5376 4003 5380
rect 4016 5307 4023 5343
rect 4056 5227 4063 5393
rect 4096 5307 4103 5374
rect 3973 5080 3987 5093
rect 3976 5076 3983 5080
rect 3956 5007 3963 5043
rect 4036 4927 4043 5113
rect 4096 5076 4103 5113
rect 4156 5107 4163 5343
rect 4196 5327 4203 5733
rect 4256 5596 4263 5633
rect 4336 5567 4343 5633
rect 4276 5427 4283 5563
rect 4216 5287 4223 5413
rect 4296 5376 4303 5433
rect 4133 5080 4147 5093
rect 4216 5083 4223 5273
rect 4356 5103 4363 5836
rect 4416 5787 4423 5863
rect 4456 5827 4463 5863
rect 4456 5647 4463 5673
rect 4556 5667 4563 5893
rect 4596 5860 4603 5863
rect 4716 5860 4723 5863
rect 4593 5847 4607 5860
rect 4713 5847 4727 5860
rect 4796 5827 4803 5894
rect 4896 5827 4903 5863
rect 4420 5623 4433 5627
rect 4416 5613 4433 5623
rect 4416 5608 4423 5613
rect 4533 5600 4547 5613
rect 4536 5596 4543 5600
rect 4736 5596 4743 5653
rect 4396 5527 4403 5563
rect 4376 5346 4383 5473
rect 4396 5387 4403 5513
rect 4516 5507 4523 5563
rect 4556 5487 4563 5563
rect 4436 5376 4443 5433
rect 4596 5376 4603 5453
rect 4616 5447 4623 5594
rect 4636 5467 4643 5594
rect 4716 5560 4723 5563
rect 4713 5547 4727 5560
rect 4756 5487 4763 5553
rect 4776 5547 4783 5693
rect 4896 5667 4903 5813
rect 4936 5707 4943 5893
rect 4956 5866 4963 5893
rect 4996 5767 5003 5863
rect 4856 5596 4863 5653
rect 4936 5566 4943 5693
rect 4716 5376 4723 5433
rect 4456 5340 4463 5343
rect 4373 5327 4387 5332
rect 4453 5327 4467 5340
rect 4816 5346 4823 5413
rect 4836 5388 4843 5433
rect 4896 5376 4903 5453
rect 4836 5347 4843 5374
rect 4576 5340 4583 5343
rect 4496 5307 4503 5333
rect 4573 5327 4587 5340
rect 4136 5076 4143 5080
rect 4196 5076 4223 5083
rect 4196 5046 4203 5076
rect 4273 5080 4287 5093
rect 4336 5096 4363 5103
rect 4276 5076 4283 5080
rect 4076 4887 4083 5043
rect 4116 5007 4123 5043
rect 4336 4987 4343 5096
rect 4473 5080 4487 5093
rect 4513 5088 4527 5093
rect 4476 5076 4483 5080
rect 3893 4860 3907 4873
rect 3896 4856 3903 4860
rect 3816 4807 3823 4853
rect 3876 4787 3883 4812
rect 3916 4727 3923 4823
rect 2573 4340 2587 4353
rect 2576 4336 2583 4340
rect 2736 4336 2743 4373
rect 2556 4247 2563 4303
rect 2596 4267 2603 4303
rect 2716 4267 2723 4303
rect 2476 4176 2503 4183
rect 2376 4036 2403 4043
rect 2416 4036 2423 4133
rect 2456 4036 2463 4073
rect 1736 3528 1743 3613
rect 1796 3486 1803 3513
rect 1696 3296 1703 3473
rect 1716 3447 1723 3483
rect 1876 3367 1883 3483
rect 1916 3447 1923 3553
rect 1496 3056 1523 3063
rect 1496 2996 1503 3056
rect 1536 2996 1543 3093
rect 1516 2907 1523 2963
rect 1416 2776 1443 2783
rect 1136 2687 1143 2743
rect 716 2476 723 2493
rect 753 2480 767 2493
rect 756 2476 763 2480
rect 636 2367 643 2474
rect 796 2347 803 2493
rect 816 2447 823 2474
rect 153 2260 167 2273
rect 156 2256 163 2260
rect 656 2256 663 2313
rect 693 2260 707 2273
rect 696 2256 703 2260
rect 16 2187 23 2253
rect 256 2187 263 2223
rect 456 2203 463 2223
rect 516 2220 523 2223
rect 436 2196 463 2203
rect 513 2207 527 2220
rect 436 2063 443 2196
rect 436 2056 463 2063
rect 76 1923 83 2033
rect 316 1956 323 2033
rect 356 1968 363 1993
rect 456 1926 463 2056
rect 576 1956 583 2193
rect 636 1968 643 2223
rect 756 2147 763 2313
rect 816 2287 823 2433
rect 856 2387 863 2443
rect 896 2263 903 2443
rect 896 2256 923 2263
rect 816 2203 823 2223
rect 876 2220 883 2223
rect 796 2196 823 2203
rect 873 2207 887 2220
rect 767 2136 783 2143
rect 76 1916 103 1923
rect 56 1707 63 1793
rect 116 1736 123 1793
rect 136 1787 143 1883
rect 156 1736 163 1813
rect 196 1747 203 1773
rect 216 1707 223 1753
rect 136 1667 143 1703
rect 116 1216 123 1313
rect 216 1223 223 1672
rect 236 1448 243 1813
rect 273 1740 287 1753
rect 276 1736 283 1740
rect 336 1436 343 1923
rect 476 1923 483 1954
rect 476 1916 503 1923
rect 356 1667 363 1773
rect 396 1736 403 1773
rect 496 1707 503 1916
rect 596 1748 603 1793
rect 636 1787 643 1954
rect 656 1767 663 1933
rect 776 1807 783 2136
rect 636 1707 643 1734
rect 656 1727 663 1753
rect 716 1736 723 1793
rect 796 1736 803 2196
rect 916 2047 923 2256
rect 816 1956 843 1963
rect 896 1956 903 1993
rect 816 1927 823 1956
rect 876 1867 883 1923
rect 936 1847 943 2333
rect 976 2207 983 2673
rect 1376 2667 1383 2743
rect 1076 2507 1083 2553
rect 1376 2527 1383 2653
rect 1073 2480 1087 2493
rect 1076 2476 1083 2480
rect 996 2307 1003 2453
rect 996 2223 1003 2293
rect 1056 2283 1063 2432
rect 1116 2427 1123 2453
rect 1136 2347 1143 2493
rect 1316 2476 1323 2513
rect 1436 2483 1443 2776
rect 1456 2567 1463 2893
rect 1416 2476 1443 2483
rect 1456 2476 1463 2553
rect 1536 2547 1543 2773
rect 1496 2476 1503 2513
rect 1236 2446 1243 2473
rect 1176 2440 1183 2443
rect 1173 2427 1187 2440
rect 1256 2387 1263 2474
rect 1276 2436 1293 2443
rect 1036 2276 1063 2283
rect 1036 2256 1043 2276
rect 996 2216 1023 2223
rect 956 2196 973 2203
rect 956 1827 963 2196
rect 1016 2007 1023 2216
rect 1076 1927 1083 2223
rect 1136 2207 1143 2273
rect 1176 2256 1183 2373
rect 1216 2256 1223 2293
rect 1276 2247 1283 2436
rect 1196 2220 1203 2223
rect 1193 2207 1207 2220
rect 1196 2027 1203 2193
rect 1196 1956 1203 1992
rect 996 1903 1003 1923
rect 1036 1920 1043 1923
rect 1033 1907 1047 1920
rect 1096 1907 1103 1933
rect 1256 1926 1263 2213
rect 1276 2147 1283 2212
rect 996 1896 1023 1903
rect 1016 1887 1023 1896
rect 460 1703 473 1707
rect 456 1696 473 1703
rect 460 1693 473 1696
rect 456 1507 463 1673
rect 556 1467 563 1693
rect 916 1700 923 1703
rect 536 1436 563 1443
rect 256 1327 263 1434
rect 556 1407 563 1436
rect 316 1400 323 1403
rect 313 1387 327 1400
rect 416 1396 443 1403
rect 416 1367 423 1396
rect 596 1387 603 1434
rect 553 1367 567 1372
rect 196 1216 223 1223
rect 253 1220 267 1233
rect 256 1216 263 1220
rect 196 1186 203 1216
rect 96 1143 103 1183
rect 76 1136 103 1143
rect 76 927 83 1136
rect 196 983 203 1172
rect 296 1167 303 1233
rect 316 1187 323 1273
rect 476 1247 483 1363
rect 516 1216 523 1353
rect 676 1347 683 1403
rect 736 1347 743 1493
rect 776 1448 783 1693
rect 913 1687 927 1700
rect 1016 1587 1023 1873
rect 1116 1847 1123 1913
rect 1036 1706 1043 1813
rect 1076 1748 1083 1833
rect 1156 1743 1163 1833
rect 1176 1763 1183 1923
rect 1276 1827 1283 2133
rect 1296 2087 1303 2333
rect 1336 2307 1343 2443
rect 1396 2427 1403 2453
rect 1416 2256 1423 2476
rect 1476 2387 1483 2443
rect 1536 2387 1543 2533
rect 1576 2527 1583 3133
rect 1653 3000 1667 3013
rect 1676 3003 1683 3293
rect 1796 3267 1803 3353
rect 1736 3067 1743 3263
rect 1856 3187 1863 3252
rect 1896 3227 1903 3263
rect 1936 3107 1943 3713
rect 2016 3516 2023 3593
rect 2076 3486 2083 3613
rect 1996 3480 2003 3483
rect 1993 3467 2007 3480
rect 2016 3296 2023 3413
rect 1996 3227 2003 3263
rect 1796 3027 1803 3053
rect 1656 2996 1663 3000
rect 1676 2996 1703 3003
rect 1696 2966 1703 2996
rect 1796 2996 1803 3013
rect 1696 2788 1703 2952
rect 1776 2827 1783 2963
rect 1753 2788 1767 2793
rect 1796 2776 1803 2833
rect 1636 2607 1643 2743
rect 1556 2516 1573 2523
rect 1556 2307 1563 2516
rect 1656 2483 1663 2553
rect 1636 2476 1663 2483
rect 1396 2203 1403 2223
rect 1396 2196 1423 2203
rect 1416 2127 1423 2196
rect 1316 1956 1323 2013
rect 1396 1968 1403 1993
rect 1336 1867 1343 1923
rect 1176 1756 1203 1763
rect 1156 1736 1183 1743
rect 787 1436 803 1443
rect 836 1436 843 1493
rect 876 1367 883 1434
rect 996 1287 1003 1363
rect 1056 1327 1063 1653
rect 1076 1627 1083 1734
rect 456 1186 463 1213
rect 576 1207 583 1233
rect 696 1216 703 1273
rect 596 1187 603 1213
rect 356 1180 363 1183
rect 353 1167 367 1180
rect 540 1183 553 1187
rect 536 1176 553 1183
rect 540 1173 553 1176
rect 676 1043 683 1183
rect 656 1036 683 1043
rect 196 976 223 983
rect 216 923 223 976
rect 340 943 353 947
rect 196 916 223 923
rect 336 933 353 943
rect 336 916 343 933
rect 433 920 447 933
rect 436 916 443 920
rect 76 883 83 913
rect 76 876 103 883
rect 316 847 323 883
rect 153 700 167 713
rect 156 696 163 700
rect 76 627 83 693
rect 136 660 143 663
rect 133 647 147 660
rect 176 367 183 652
rect 236 647 243 833
rect 293 700 307 713
rect 296 696 303 700
rect 336 696 343 753
rect 396 727 403 914
rect 456 787 463 883
rect 496 747 503 872
rect 656 847 663 1036
rect 756 967 763 1273
rect 1016 1256 1023 1313
rect 833 1220 847 1233
rect 836 1216 843 1220
rect 967 1216 983 1223
rect 807 1176 823 1183
rect 756 916 763 953
rect 796 887 803 1172
rect 856 1147 863 1183
rect 316 660 323 663
rect 313 647 327 660
rect 376 587 383 713
rect 496 696 503 733
rect 396 627 403 692
rect 416 627 423 653
rect 276 396 283 453
rect 136 307 143 363
rect 176 147 183 174
rect 216 143 223 353
rect 216 136 233 143
rect 316 143 323 493
rect 336 408 343 573
rect 396 396 403 493
rect 436 467 443 663
rect 476 660 483 663
rect 473 647 487 660
rect 536 647 543 773
rect 696 767 703 883
rect 816 867 823 913
rect 856 880 863 883
rect 716 696 723 753
rect 816 666 823 793
rect 426 453 427 460
rect 413 443 427 453
rect 413 440 463 443
rect 416 436 467 440
rect 453 427 467 436
rect 336 367 343 394
rect 476 367 483 612
rect 296 136 323 143
rect 316 107 323 136
rect 336 127 343 353
rect 376 187 383 363
rect 496 363 503 453
rect 553 400 567 413
rect 716 408 723 453
rect 556 396 563 400
rect 496 356 543 363
rect 576 356 613 363
rect 636 307 643 394
rect 416 176 423 293
rect 696 247 703 363
rect 776 347 783 652
rect 836 467 843 873
rect 853 867 867 880
rect 896 767 903 883
rect 936 807 943 1073
rect 956 1047 963 1214
rect 956 747 963 953
rect 1016 916 1023 1033
rect 873 723 887 733
rect 873 720 913 723
rect 876 716 913 720
rect 916 660 923 663
rect 913 647 927 660
rect 956 647 963 712
rect 976 666 983 913
rect 1076 883 1083 914
rect 1036 876 1083 883
rect 1056 736 1063 876
rect 1096 767 1103 1693
rect 1116 1587 1123 1703
rect 1176 1463 1183 1736
rect 1196 1487 1203 1756
rect 1256 1736 1263 1773
rect 1336 1706 1343 1813
rect 1376 1807 1383 1923
rect 1416 1887 1423 2113
rect 1456 1963 1463 2293
rect 1476 2187 1483 2293
rect 1496 2226 1503 2253
rect 1576 2187 1583 2223
rect 1436 1956 1463 1963
rect 1476 1956 1483 2093
rect 1516 2087 1523 2133
rect 1516 1968 1523 2073
rect 1436 1867 1443 1956
rect 1236 1700 1243 1703
rect 1233 1687 1247 1700
rect 1356 1667 1363 1773
rect 1396 1748 1403 1773
rect 1436 1736 1443 1813
rect 1476 1687 1483 1853
rect 1356 1487 1363 1653
rect 1496 1527 1503 1923
rect 1556 1787 1563 2033
rect 1576 1767 1583 2173
rect 1616 2047 1623 2443
rect 1696 2407 1703 2553
rect 1736 2507 1743 2693
rect 1776 2667 1783 2743
rect 1816 2740 1823 2743
rect 1813 2727 1827 2740
rect 1856 2727 1863 2813
rect 1876 2747 1883 3013
rect 1916 2996 1923 3073
rect 1973 3008 1987 3013
rect 1896 2967 1903 2994
rect 1936 2907 1943 2952
rect 1936 2827 1943 2893
rect 1913 2780 1927 2793
rect 1916 2776 1923 2780
rect 1956 2776 1963 2853
rect 1867 2716 1883 2723
rect 1733 2480 1747 2493
rect 1736 2476 1743 2480
rect 1776 2476 1783 2513
rect 1756 2387 1763 2443
rect 1796 2407 1803 2443
rect 1767 2376 1783 2383
rect 1776 2226 1783 2376
rect 1876 2256 1883 2716
rect 1936 2667 1943 2743
rect 1976 2667 1983 2743
rect 2016 2523 2023 3133
rect 2036 3087 2043 3252
rect 2076 3227 2083 3273
rect 2096 3008 2103 3673
rect 2156 3528 2163 3713
rect 2356 3687 2363 3753
rect 2376 3687 2383 4036
rect 2433 3820 2447 3833
rect 2436 3816 2443 3820
rect 2416 3743 2423 3783
rect 2396 3736 2423 3743
rect 2396 3567 2403 3736
rect 2496 3727 2503 4176
rect 2556 4087 2563 4233
rect 2716 4207 2723 4253
rect 2756 4247 2763 4292
rect 2836 4287 2843 4373
rect 2936 4336 2943 4433
rect 2976 4306 2983 4333
rect 2876 4300 2883 4303
rect 2873 4287 2887 4300
rect 2516 4007 2523 4073
rect 2616 4036 2623 4073
rect 2636 4067 2643 4173
rect 2556 3907 2563 4003
rect 2596 3947 2603 4003
rect 2576 3816 2583 3853
rect 2656 3786 2663 4073
rect 2713 4048 2727 4053
rect 2756 4036 2763 4073
rect 2556 3727 2563 3783
rect 2576 3627 2583 3733
rect 2596 3687 2603 3783
rect 2676 3783 2683 4034
rect 2716 3816 2723 3973
rect 2776 3787 2783 3814
rect 2676 3776 2703 3783
rect 2596 3647 2603 3673
rect 2696 3667 2703 3776
rect 2796 3747 2803 4153
rect 2816 4007 2823 4273
rect 2916 3828 2923 4253
rect 3053 4048 3067 4053
rect 3076 4007 3083 4213
rect 3096 4048 3103 4303
rect 3136 4187 3143 4334
rect 3276 4306 3283 4333
rect 3196 4300 3203 4303
rect 3193 4287 3207 4300
rect 3236 4247 3243 4303
rect 3296 4247 3303 4353
rect 3373 4340 3387 4353
rect 3376 4336 3383 4340
rect 3436 4307 3443 4472
rect 3676 4376 3683 4554
rect 3816 4526 3823 4573
rect 3873 4560 3887 4573
rect 3916 4568 3923 4613
rect 3876 4556 3883 4560
rect 3496 4300 3503 4303
rect 3396 4227 3403 4292
rect 3493 4287 3507 4300
rect 3536 4187 3543 4303
rect 3136 4147 3143 4173
rect 3176 4048 3183 4073
rect 2996 3947 3003 4003
rect 3053 3983 3067 3993
rect 3036 3980 3067 3983
rect 3036 3976 3063 3980
rect 2976 3828 2983 3893
rect 3036 3816 3043 3976
rect 2816 3780 2843 3783
rect 2813 3776 2843 3780
rect 2813 3767 2827 3776
rect 2836 3747 2843 3776
rect 2896 3727 2903 3772
rect 2916 3767 2923 3814
rect 2196 3516 2233 3523
rect 2176 3407 2183 3483
rect 2236 3467 2243 3514
rect 2316 3447 2323 3483
rect 2153 3300 2167 3313
rect 2156 3296 2163 3300
rect 2136 3227 2143 3263
rect 2056 2687 2063 2993
rect 2116 2927 2123 2963
rect 2176 2827 2183 2994
rect 2136 2776 2143 2813
rect 1996 2516 2023 2523
rect 1896 2267 1903 2513
rect 1956 2407 1963 2443
rect 1696 2220 1703 2223
rect 1693 2207 1707 2220
rect 1696 2107 1703 2193
rect 1796 2043 1803 2253
rect 1916 2227 1923 2313
rect 1956 2307 1963 2393
rect 1996 2347 2003 2516
rect 2076 2507 2083 2733
rect 2156 2667 2163 2743
rect 2116 2547 2123 2593
rect 2036 2263 2043 2493
rect 2076 2476 2083 2493
rect 2113 2480 2127 2493
rect 2116 2476 2123 2480
rect 2096 2440 2103 2443
rect 2093 2427 2107 2440
rect 2156 2383 2163 2493
rect 2176 2427 2183 2593
rect 2196 2507 2203 3213
rect 2216 3147 2223 3313
rect 2236 3307 2243 3373
rect 2273 3300 2287 3313
rect 2276 3296 2283 3300
rect 2336 3266 2343 3453
rect 2356 3227 2363 3353
rect 2376 3347 2383 3514
rect 2396 3367 2403 3553
rect 2433 3528 2447 3533
rect 2633 3520 2647 3533
rect 2636 3516 2643 3520
rect 2536 3486 2543 3514
rect 2416 3367 2423 3473
rect 2456 3447 2463 3483
rect 2416 3296 2423 3353
rect 2496 3347 2503 3483
rect 2536 3427 2543 3472
rect 2556 3447 2563 3514
rect 2696 3383 2703 3653
rect 2816 3516 2823 3673
rect 2976 3627 2983 3814
rect 3096 3747 3103 4034
rect 3156 3947 3163 4003
rect 3136 3747 3143 3772
rect 3176 3767 3183 3783
rect 3116 3647 3123 3713
rect 3176 3647 3183 3753
rect 3216 3687 3223 3973
rect 2716 3487 2723 3514
rect 2676 3376 2703 3383
rect 2456 3307 2463 3333
rect 2396 3227 2403 3263
rect 2236 2996 2243 3093
rect 2276 2996 2283 3093
rect 2316 2967 2323 3033
rect 2416 2996 2423 3173
rect 2436 3107 2443 3252
rect 2476 3247 2483 3313
rect 2616 3308 2623 3373
rect 2496 3267 2503 3294
rect 2256 2827 2263 2963
rect 2216 2508 2223 2774
rect 2256 2687 2263 2743
rect 2316 2740 2323 2743
rect 2313 2727 2327 2740
rect 2336 2723 2343 2994
rect 2436 2887 2443 2963
rect 2476 2827 2483 3013
rect 2416 2740 2423 2743
rect 2327 2716 2343 2723
rect 2413 2727 2427 2740
rect 2256 2567 2263 2673
rect 2456 2667 2463 2743
rect 2496 2627 2503 3253
rect 2516 3243 2523 3293
rect 2516 3236 2543 3243
rect 2536 3127 2543 3236
rect 2556 3227 2563 3263
rect 2596 3187 2603 3263
rect 2636 3227 2643 3252
rect 2676 3083 2683 3376
rect 2696 3187 2703 3313
rect 2736 3296 2743 3353
rect 2756 3327 2763 3472
rect 2796 3447 2803 3483
rect 2856 3407 2863 3453
rect 2876 3427 2883 3613
rect 2976 3516 2983 3592
rect 2993 3527 3007 3533
rect 2800 3343 2813 3347
rect 2796 3333 2813 3343
rect 2796 3267 2803 3333
rect 2876 3296 2883 3333
rect 2896 3327 2903 3353
rect 2916 3296 2923 3333
rect 2816 3266 2823 3293
rect 2956 3287 2963 3353
rect 2896 3227 2903 3263
rect 2756 3127 2763 3193
rect 2656 3076 2683 3083
rect 2536 2996 2543 3033
rect 2573 3000 2587 3013
rect 2576 2996 2583 3000
rect 2636 2966 2643 3053
rect 2556 2867 2563 2963
rect 2556 2776 2563 2813
rect 2516 2727 2523 2773
rect 2576 2727 2583 2743
rect 2576 2716 2593 2727
rect 2580 2713 2593 2716
rect 2356 2507 2363 2613
rect 2536 2587 2543 2613
rect 2147 2376 2163 2383
rect 2036 2256 2063 2263
rect 1796 2036 1823 2043
rect 1616 1956 1623 1993
rect 1676 1926 1683 2033
rect 1696 1847 1703 1973
rect 1753 1960 1767 1973
rect 1756 1956 1763 1960
rect 1816 1926 1823 2036
rect 1936 2027 1943 2253
rect 2056 2226 2063 2256
rect 2136 2256 2143 2373
rect 2236 2307 2243 2443
rect 2176 2256 2183 2293
rect 1976 2147 1983 2223
rect 1936 1956 1943 1992
rect 1856 1887 1863 1954
rect 1616 1707 1623 1793
rect 1693 1740 1707 1753
rect 1696 1736 1703 1740
rect 1156 1456 1183 1463
rect 1156 1448 1163 1456
rect 1193 1440 1207 1452
rect 1196 1436 1203 1440
rect 1236 1406 1243 1473
rect 1333 1448 1347 1453
rect 1136 1087 1143 1403
rect 1193 1220 1207 1233
rect 1196 1216 1203 1220
rect 1276 1187 1283 1273
rect 1296 948 1303 1253
rect 1336 1228 1343 1353
rect 1356 1267 1363 1403
rect 1396 1247 1403 1473
rect 1416 1367 1423 1513
rect 1476 1436 1483 1473
rect 1513 1440 1527 1453
rect 1516 1436 1523 1440
rect 1456 1367 1463 1403
rect 1556 1367 1563 1673
rect 1576 1467 1583 1703
rect 1796 1667 1803 1873
rect 1836 1767 1843 1813
rect 1856 1736 1863 1833
rect 1916 1787 1923 1923
rect 1956 1920 1963 1923
rect 1953 1907 1967 1920
rect 1996 1907 2003 2033
rect 2036 1926 2043 2013
rect 2076 2007 2083 2253
rect 2156 2167 2163 2223
rect 2196 2220 2203 2223
rect 2193 2207 2207 2220
rect 2236 2147 2243 2272
rect 2256 2167 2263 2253
rect 2276 2047 2283 2333
rect 2316 2288 2323 2493
rect 2356 2476 2363 2493
rect 2396 2476 2403 2553
rect 2476 2547 2483 2573
rect 2376 2268 2383 2443
rect 2336 2187 2343 2223
rect 2376 2127 2383 2254
rect 2296 2087 2303 2113
rect 2396 2027 2403 2293
rect 2436 2263 2443 2493
rect 2496 2488 2503 2513
rect 2556 2507 2563 2553
rect 2556 2476 2563 2493
rect 2456 2427 2463 2453
rect 2516 2387 2523 2443
rect 2576 2427 2583 2473
rect 2616 2446 2623 2913
rect 2656 2887 2663 3076
rect 2727 3033 2733 3047
rect 2676 3007 2683 3033
rect 2693 3000 2707 3013
rect 2733 3000 2747 3012
rect 2696 2996 2703 3000
rect 2736 2996 2743 3000
rect 2676 2867 2683 2953
rect 2796 2963 2803 3153
rect 2756 2887 2763 2963
rect 2776 2956 2803 2963
rect 2696 2776 2703 2833
rect 2733 2780 2747 2793
rect 2736 2776 2743 2780
rect 2676 2740 2683 2743
rect 2673 2727 2687 2740
rect 2713 2727 2727 2732
rect 2676 2687 2683 2713
rect 2656 2476 2663 2533
rect 2696 2476 2703 2653
rect 2676 2327 2683 2443
rect 2736 2367 2743 2553
rect 2776 2423 2783 2956
rect 2816 2867 2823 3113
rect 2836 3007 2843 3193
rect 2876 3008 2883 3033
rect 2916 2996 2923 3033
rect 2836 2927 2843 2953
rect 2796 2746 2803 2833
rect 2816 2507 2823 2853
rect 2856 2807 2863 2952
rect 2896 2807 2903 2963
rect 2916 2776 2923 2853
rect 2896 2687 2903 2743
rect 2956 2707 2963 3053
rect 2976 2667 2983 3293
rect 2996 3167 3003 3413
rect 3016 3347 3023 3493
rect 3036 3447 3043 3613
rect 3216 3563 3223 3673
rect 3196 3556 3223 3563
rect 3056 3467 3063 3553
rect 3147 3536 3173 3543
rect 3196 3527 3203 3556
rect 3236 3547 3243 4034
rect 3276 3947 3283 4003
rect 3276 3907 3283 3933
rect 3336 3843 3343 4173
rect 3576 4147 3583 4373
rect 3596 4147 3603 4334
rect 3756 4303 3763 4453
rect 3776 4306 3783 4512
rect 3836 4467 3843 4553
rect 3896 4467 3903 4523
rect 3736 4296 3763 4303
rect 3796 4143 3803 4453
rect 3836 4348 3843 4413
rect 3876 4336 3883 4373
rect 3896 4300 3903 4303
rect 3893 4287 3907 4300
rect 3796 4136 3823 4143
rect 3413 4040 3427 4053
rect 3416 4036 3423 4040
rect 3476 4043 3483 4073
rect 3467 4036 3483 4043
rect 3496 4007 3503 4113
rect 3396 4000 3403 4003
rect 3393 3987 3407 4000
rect 3316 3836 3343 3843
rect 3316 3816 3323 3836
rect 3356 3827 3363 3953
rect 3276 3707 3283 3783
rect 3336 3747 3343 3783
rect 3376 3747 3383 3913
rect 3396 3707 3403 3814
rect 3456 3667 3463 3772
rect 3496 3747 3503 3893
rect 3216 3536 3233 3543
rect 3036 3296 3043 3353
rect 3116 3327 3123 3483
rect 3196 3347 3203 3373
rect 3216 3347 3223 3536
rect 3256 3516 3263 3553
rect 3293 3520 3307 3533
rect 3296 3516 3303 3520
rect 3316 3407 3323 3483
rect 3336 3387 3343 3473
rect 3356 3467 3363 3553
rect 3376 3443 3383 3633
rect 3447 3616 3483 3623
rect 3456 3567 3463 3593
rect 3476 3587 3483 3616
rect 3456 3516 3463 3553
rect 3436 3463 3443 3483
rect 3356 3436 3383 3443
rect 3416 3456 3443 3463
rect 3136 3266 3143 3333
rect 3056 3207 3063 3263
rect 3176 3227 3183 3294
rect 3196 3263 3203 3333
rect 3196 3256 3223 3263
rect 3156 3147 3163 3193
rect 3076 2996 3083 3053
rect 3116 2967 3123 3013
rect 3116 2887 3123 2913
rect 3013 2780 3027 2793
rect 3016 2776 3023 2780
rect 3056 2776 3063 2813
rect 3116 2767 3123 2873
rect 2933 2627 2947 2633
rect 2993 2627 3007 2633
rect 2956 2476 2963 2593
rect 2993 2480 3007 2493
rect 2996 2476 3003 2480
rect 2776 2420 2803 2423
rect 2776 2416 2807 2420
rect 2793 2407 2807 2416
rect 2836 2387 2843 2443
rect 2416 2256 2443 2263
rect 2416 2207 2423 2256
rect 2516 2256 2523 2313
rect 2496 2167 2503 2223
rect 2556 2147 2563 2223
rect 2596 2187 2603 2293
rect 2616 2226 2623 2313
rect 2647 2293 2653 2307
rect 2636 2167 2643 2254
rect 2796 2226 2803 2313
rect 2856 2256 2863 2293
rect 2896 2256 2903 2333
rect 2156 1926 2163 1993
rect 2213 1960 2227 1973
rect 2216 1956 2223 1960
rect 1913 1740 1927 1752
rect 1916 1736 1923 1740
rect 1956 1706 1963 1733
rect 1816 1547 1823 1703
rect 1976 1527 1983 1773
rect 2016 1706 2023 1833
rect 2056 1748 2063 1913
rect 2156 1767 2163 1912
rect 2196 1803 2203 1912
rect 2276 1907 2283 1953
rect 2196 1796 2223 1803
rect 2156 1706 2163 1753
rect 2216 1736 2223 1796
rect 2296 1747 2303 2013
rect 2336 1956 2343 2013
rect 2373 1960 2387 1973
rect 2493 1960 2507 1973
rect 2376 1956 2383 1960
rect 2496 1956 2503 1960
rect 2536 1956 2543 2013
rect 2636 1926 2643 2113
rect 2696 1956 2703 2153
rect 2736 2127 2743 2223
rect 2796 1968 2803 2212
rect 2876 2207 2883 2223
rect 2856 2196 2873 2203
rect 2856 1956 2863 2196
rect 2936 2167 2943 2253
rect 2356 1920 2363 1923
rect 2353 1907 2367 1920
rect 2396 1867 2403 1923
rect 2436 1847 2443 1893
rect 2176 1547 2183 1713
rect 2280 1703 2293 1707
rect 2236 1700 2243 1703
rect 2233 1687 2247 1700
rect 2276 1696 2293 1703
rect 2280 1693 2293 1696
rect 1633 1440 1647 1453
rect 1673 1440 1687 1453
rect 1733 1448 1747 1453
rect 1636 1436 1643 1440
rect 1676 1436 1683 1440
rect 1816 1436 1823 1473
rect 1993 1448 2007 1453
rect 1916 1436 1963 1443
rect 1416 1223 1423 1313
rect 1396 1216 1423 1223
rect 1456 1216 1463 1273
rect 1396 1187 1403 1216
rect 1476 1180 1483 1183
rect 1473 1167 1487 1180
rect 1156 847 1163 883
rect 996 703 1003 733
rect 996 696 1023 703
rect 1176 647 1183 753
rect 1196 663 1203 883
rect 1236 863 1243 914
rect 1256 887 1263 933
rect 1336 916 1343 1133
rect 1516 1127 1523 1183
rect 1556 1107 1563 1213
rect 1576 1186 1583 1233
rect 1596 1223 1603 1273
rect 1616 1247 1623 1403
rect 1656 1367 1663 1403
rect 1736 1327 1743 1434
rect 1896 1407 1903 1434
rect 1916 1407 1923 1436
rect 1796 1367 1803 1403
rect 2076 1406 2083 1513
rect 2316 1507 2323 1733
rect 2336 1607 2343 1813
rect 2396 1736 2403 1813
rect 2436 1736 2443 1833
rect 2376 1667 2383 1703
rect 2133 1440 2147 1453
rect 2136 1436 2143 1440
rect 1596 1216 1623 1223
rect 1676 1180 1683 1183
rect 1673 1167 1687 1180
rect 1380 923 1393 927
rect 1376 916 1393 923
rect 1380 913 1393 916
rect 1656 916 1663 953
rect 1236 860 1263 863
rect 1236 856 1267 860
rect 1253 847 1267 856
rect 1316 823 1323 883
rect 1356 880 1363 883
rect 1353 867 1367 880
rect 1316 816 1343 823
rect 1196 656 1223 663
rect 796 366 803 453
rect 1316 443 1323 793
rect 1336 767 1343 816
rect 1336 666 1343 753
rect 1396 708 1403 873
rect 1416 867 1423 913
rect 1436 883 1443 913
rect 1436 876 1463 883
rect 1376 627 1383 663
rect 1416 656 1433 663
rect 1296 436 1323 443
rect 1180 423 1193 427
rect 1176 413 1193 423
rect 1016 396 1063 403
rect 856 360 863 363
rect 853 347 867 360
rect 547 203 560 207
rect 547 193 563 203
rect 476 146 483 193
rect 556 176 563 193
rect 496 146 503 173
rect 756 146 763 233
rect 816 188 823 253
rect 856 176 863 293
rect 896 267 903 394
rect 996 183 1003 352
rect 1056 307 1063 396
rect 1176 396 1183 413
rect 1296 408 1303 436
rect 1333 400 1347 413
rect 1336 396 1343 400
rect 1136 307 1143 363
rect 976 176 1003 183
rect 1116 176 1123 233
rect 1256 188 1263 393
rect 1356 327 1363 363
rect 1436 363 1443 653
rect 1456 547 1463 876
rect 1496 827 1503 883
rect 1556 827 1563 914
rect 1696 886 1703 1033
rect 1716 947 1723 1213
rect 1736 1127 1743 1233
rect 1793 1220 1807 1233
rect 1796 1216 1803 1220
rect 1776 1167 1783 1172
rect 1767 1156 1783 1167
rect 1767 1153 1780 1156
rect 1776 916 1783 1053
rect 1836 1007 1843 1213
rect 1856 1187 1863 1393
rect 1976 1347 1983 1403
rect 1916 1107 1923 1183
rect 1996 1067 2003 1253
rect 2016 1228 2023 1403
rect 2076 1347 2083 1392
rect 2116 1267 2123 1403
rect 2156 1207 2163 1233
rect 2056 1107 2063 1183
rect 1827 953 1833 967
rect 1856 928 1863 973
rect 1856 887 1863 914
rect 1596 847 1603 883
rect 1576 696 1583 753
rect 1696 696 1703 813
rect 1796 807 1803 883
rect 1876 886 1883 1053
rect 1907 953 1913 967
rect 1933 920 1947 933
rect 1936 916 1943 920
rect 1907 883 1920 887
rect 1907 876 1923 883
rect 1907 873 1920 876
rect 2056 847 2063 993
rect 2093 920 2107 933
rect 2136 928 2143 993
rect 2096 916 2103 920
rect 2176 923 2183 1213
rect 2196 1127 2203 1393
rect 2216 1183 2223 1473
rect 2236 1407 2243 1434
rect 2256 1247 2263 1393
rect 2336 1228 2343 1593
rect 2416 1567 2423 1703
rect 2356 1406 2363 1493
rect 2436 1436 2443 1513
rect 2456 1487 2463 1692
rect 2476 1468 2483 1553
rect 2496 1443 2503 1853
rect 2556 1787 2563 1923
rect 2516 1547 2523 1734
rect 2556 1667 2563 1703
rect 2596 1647 2603 1703
rect 2656 1667 2663 1773
rect 2716 1748 2723 1923
rect 2596 1567 2603 1633
rect 2676 1607 2683 1733
rect 2496 1436 2523 1443
rect 2416 1400 2423 1403
rect 2216 1176 2243 1183
rect 2207 953 2213 967
rect 2236 947 2243 1176
rect 2356 1007 2363 1392
rect 2413 1387 2427 1400
rect 2456 1347 2463 1403
rect 2516 1406 2523 1436
rect 2396 1187 2403 1214
rect 2176 916 2203 923
rect 2256 916 2263 973
rect 2287 953 2293 967
rect 2156 787 2163 883
rect 1496 667 1503 694
rect 1556 627 1563 663
rect 1596 627 1603 663
rect 1556 463 1563 613
rect 1556 456 1583 463
rect 1576 403 1583 456
rect 1556 396 1583 403
rect 1436 356 1463 363
rect 916 147 923 174
rect 1396 176 1403 353
rect 1436 176 1443 356
rect 1496 287 1503 323
rect 1616 287 1623 652
rect 1656 627 1663 694
rect 1656 396 1663 613
rect 1756 366 1763 533
rect 1796 403 1803 693
rect 1936 666 1943 753
rect 2196 747 2203 916
rect 2276 847 2283 883
rect 1856 643 1863 663
rect 1856 640 1883 643
rect 1853 636 1883 640
rect 1853 627 1867 636
rect 1776 396 1803 403
rect 1496 187 1503 273
rect 1676 187 1683 363
rect 1716 360 1723 363
rect 1713 347 1727 360
rect 1776 347 1783 396
rect 1876 367 1883 636
rect 1976 627 1983 733
rect 2236 687 2243 793
rect 2316 787 2323 883
rect 2356 867 2363 913
rect 2107 656 2123 663
rect 2136 660 2143 663
rect 2196 660 2203 663
rect 2116 547 2123 656
rect 2133 647 2147 660
rect 2193 647 2207 660
rect 1916 247 1923 433
rect 1976 396 1983 433
rect 2020 403 2033 407
rect 2016 396 2033 403
rect 2020 393 2033 396
rect 2116 396 2123 433
rect 2136 427 2143 633
rect 2256 627 2263 773
rect 2313 700 2327 713
rect 2316 696 2323 700
rect 2356 567 2363 713
rect 2276 423 2283 553
rect 2193 400 2207 413
rect 2256 416 2283 423
rect 2196 396 2203 400
rect 2256 396 2263 416
rect 1996 327 2003 363
rect 2056 327 2063 373
rect 2076 327 2083 393
rect 2296 347 2303 493
rect 2376 427 2383 933
rect 2396 927 2403 1173
rect 2416 1127 2423 1183
rect 2476 1147 2483 1183
rect 2496 1167 2503 1393
rect 2536 1347 2543 1493
rect 2556 1447 2563 1553
rect 2596 1436 2603 1513
rect 2636 1436 2673 1443
rect 2616 1267 2623 1403
rect 2676 1307 2683 1434
rect 2696 1367 2703 1653
rect 2736 1567 2743 1703
rect 2776 1687 2783 1933
rect 2916 1827 2923 2013
rect 2916 1748 2923 1813
rect 2796 1623 2803 1733
rect 2936 1706 2943 2073
rect 2956 1767 2963 2393
rect 2976 2367 2983 2443
rect 3036 2407 3043 2553
rect 3056 2446 3063 2673
rect 3076 2667 3083 2743
rect 3136 2547 3143 3073
rect 3156 3007 3163 3033
rect 3176 2996 3183 3113
rect 3227 3016 3253 3023
rect 3276 3007 3283 3263
rect 3196 2776 3203 2873
rect 3276 2843 3283 2972
rect 3296 2887 3303 3113
rect 3316 3007 3323 3333
rect 3336 3127 3343 3294
rect 3356 3187 3363 3436
rect 3336 3087 3343 3113
rect 3376 3067 3383 3413
rect 3416 3327 3423 3456
rect 3396 3187 3403 3263
rect 3373 3000 3387 3013
rect 3376 2996 3383 3000
rect 3476 3003 3483 3293
rect 3496 3267 3503 3453
rect 3516 3307 3523 4133
rect 3576 4096 3613 4103
rect 3576 4068 3583 4096
rect 3600 4086 3620 4087
rect 3607 4073 3613 4086
rect 3667 4073 3673 4087
rect 3696 4067 3703 4133
rect 3613 4040 3627 4052
rect 3676 4056 3693 4063
rect 3616 4036 3623 4040
rect 3556 3967 3563 4003
rect 3596 4000 3603 4003
rect 3593 3987 3607 4000
rect 3676 4006 3683 4056
rect 3736 4036 3743 4093
rect 3556 3847 3563 3953
rect 3547 3823 3560 3827
rect 3547 3816 3563 3823
rect 3547 3813 3560 3816
rect 3536 3467 3543 3772
rect 3576 3763 3583 3783
rect 3556 3756 3583 3763
rect 3556 3727 3563 3756
rect 3656 3747 3663 3993
rect 3756 3947 3763 4003
rect 3796 3987 3803 4113
rect 3816 3943 3823 4136
rect 3836 4006 3843 4073
rect 3896 4067 3903 4113
rect 3853 4040 3867 4053
rect 3856 4036 3863 4040
rect 3896 3947 3903 4003
rect 3796 3936 3823 3943
rect 3796 3887 3803 3936
rect 3556 3527 3563 3713
rect 3616 3587 3623 3693
rect 3596 3547 3603 3573
rect 3636 3567 3643 3593
rect 3596 3536 3613 3547
rect 3600 3533 3613 3536
rect 3553 3467 3567 3473
rect 3576 3447 3583 3483
rect 3616 3427 3623 3453
rect 3636 3347 3643 3513
rect 3536 3307 3543 3333
rect 3613 3300 3627 3313
rect 3656 3303 3663 3613
rect 3676 3527 3683 3873
rect 3696 3856 3783 3863
rect 3696 3827 3703 3856
rect 3713 3820 3727 3833
rect 3776 3843 3783 3856
rect 3776 3840 3803 3843
rect 3776 3836 3807 3840
rect 3753 3820 3767 3833
rect 3793 3827 3807 3836
rect 3716 3816 3723 3820
rect 3756 3816 3763 3820
rect 3816 3786 3823 3913
rect 3836 3876 3883 3883
rect 3836 3847 3843 3876
rect 3856 3827 3863 3853
rect 3876 3843 3883 3876
rect 3876 3836 3903 3843
rect 3896 3816 3903 3836
rect 3936 3816 3943 4113
rect 3956 3827 3963 4873
rect 3973 4868 3987 4873
rect 4096 4863 4103 4913
rect 4076 4856 4103 4863
rect 3976 4787 3983 4854
rect 4056 4727 4063 4823
rect 4116 4568 4123 4873
rect 4136 4827 4143 4854
rect 4147 4816 4163 4823
rect 3996 4556 4023 4563
rect 4076 4556 4103 4563
rect 3976 4526 3983 4553
rect 3996 4287 4003 4556
rect 4056 4336 4063 4373
rect 4096 4307 4103 4556
rect 4136 4343 4143 4613
rect 4156 4523 4163 4816
rect 4236 4627 4243 4973
rect 4376 4963 4383 5074
rect 4416 5007 4423 5043
rect 4376 4956 4393 4963
rect 4256 4587 4263 4953
rect 4276 4867 4283 4913
rect 4296 4856 4303 4933
rect 4316 4883 4323 4953
rect 4333 4883 4347 4893
rect 4316 4880 4347 4883
rect 4316 4876 4343 4880
rect 4336 4856 4343 4876
rect 4396 4867 4403 4953
rect 4396 4826 4403 4853
rect 4416 4767 4423 4933
rect 4456 4907 4463 5043
rect 4516 4927 4523 5074
rect 4536 4947 4543 5313
rect 4616 5287 4623 5343
rect 4736 5340 4743 5343
rect 4733 5327 4747 5340
rect 4616 5207 4623 5273
rect 4956 5267 4963 5613
rect 4976 5567 4983 5633
rect 5076 5608 5083 5933
rect 5116 5903 5123 5973
rect 5116 5896 5143 5903
rect 5116 5627 5123 5896
rect 5236 5867 5243 5993
rect 5356 5866 5363 5893
rect 5176 5827 5183 5852
rect 4996 5376 5003 5453
rect 5016 5407 5023 5493
rect 5036 5447 5043 5533
rect 5056 5467 5063 5563
rect 5056 5427 5063 5453
rect 5096 5346 5103 5453
rect 5116 5327 5123 5592
rect 5136 5566 5143 5753
rect 5196 5596 5203 5653
rect 5236 5608 5243 5813
rect 5276 5763 5283 5852
rect 5316 5827 5323 5863
rect 5276 5756 5303 5763
rect 5176 5507 5183 5563
rect 5216 5527 5223 5552
rect 5227 5516 5243 5523
rect 5176 5388 5183 5413
rect 5236 5343 5243 5516
rect 5276 5383 5283 5673
rect 5296 5547 5303 5756
rect 5356 5596 5363 5653
rect 5396 5628 5403 5893
rect 5436 5727 5443 5852
rect 5476 5667 5483 5863
rect 5536 5827 5543 5894
rect 5596 5843 5603 5863
rect 5656 5847 5663 5894
rect 5576 5836 5603 5843
rect 5576 5687 5583 5836
rect 5336 5467 5343 5563
rect 5376 5527 5383 5563
rect 5300 5403 5313 5407
rect 5156 5287 5163 5343
rect 5196 5336 5243 5343
rect 5256 5376 5283 5383
rect 5296 5393 5313 5403
rect 5296 5376 5303 5393
rect 5376 5388 5383 5453
rect 4696 5043 4703 5253
rect 5136 5127 5143 5213
rect 4893 5088 4907 5093
rect 5033 5080 5047 5093
rect 5036 5076 5043 5080
rect 4556 4987 4563 5033
rect 4507 4916 4523 4927
rect 4507 4913 4520 4916
rect 4467 4896 4483 4903
rect 4476 4887 4483 4896
rect 4476 4876 4493 4887
rect 4480 4873 4493 4876
rect 4516 4856 4523 4893
rect 4253 4560 4267 4573
rect 4256 4556 4263 4560
rect 4296 4527 4303 4713
rect 4456 4667 4463 4823
rect 4496 4820 4503 4823
rect 4493 4807 4507 4820
rect 4536 4787 4543 4813
rect 4556 4807 4563 4893
rect 4576 4807 4583 4993
rect 4596 4967 4603 5043
rect 4636 4907 4643 5043
rect 4696 5036 4723 5043
rect 4596 4867 4603 4893
rect 4676 4856 4683 4993
rect 4696 4887 4703 4953
rect 4376 4556 4383 4653
rect 4416 4556 4423 4613
rect 4456 4547 4463 4573
rect 4156 4516 4203 4523
rect 4116 4336 4143 4343
rect 4176 4336 4183 4413
rect 3696 3707 3703 3773
rect 3736 3747 3743 3783
rect 3816 3747 3823 3772
rect 3836 3767 3843 3812
rect 3916 3780 3923 3783
rect 3913 3767 3927 3780
rect 3733 3520 3747 3533
rect 3776 3527 3783 3733
rect 3736 3516 3743 3520
rect 3856 3516 3863 3573
rect 3916 3567 3923 3613
rect 3893 3520 3907 3533
rect 3896 3516 3903 3520
rect 3793 3483 3807 3493
rect 3676 3447 3683 3473
rect 3676 3387 3683 3412
rect 3616 3296 3623 3300
rect 3656 3296 3683 3303
rect 3456 2996 3483 3003
rect 3516 2996 3523 3272
rect 3536 3007 3543 3253
rect 3396 2887 3403 2963
rect 3436 2863 3443 2993
rect 3416 2856 3443 2863
rect 3456 2863 3463 2996
rect 3576 2966 3583 3233
rect 3596 3047 3603 3263
rect 3636 3260 3663 3263
rect 3636 3256 3667 3260
rect 3653 3247 3667 3256
rect 3636 3207 3643 3233
rect 3636 2996 3643 3193
rect 3676 3187 3683 3296
rect 3696 3247 3703 3453
rect 3716 3447 3723 3483
rect 3756 3480 3807 3483
rect 3756 3476 3803 3480
rect 3816 3447 3823 3514
rect 3736 3308 3743 3373
rect 3876 3303 3883 3472
rect 3876 3296 3903 3303
rect 3756 3260 3763 3263
rect 3753 3247 3767 3260
rect 3733 3223 3747 3233
rect 3733 3220 3773 3223
rect 3736 3216 3773 3220
rect 3836 3207 3843 3252
rect 3456 2856 3483 2863
rect 3276 2836 3303 2843
rect 3236 2776 3243 2813
rect 3276 2746 3283 2813
rect 3156 2736 3183 2743
rect 3156 2707 3163 2736
rect 3296 2567 3303 2836
rect 3416 2776 3423 2856
rect 3376 2707 3383 2732
rect 3416 2627 3423 2713
rect 3093 2480 3107 2493
rect 3096 2476 3103 2480
rect 3373 2483 3387 2493
rect 3356 2480 3387 2483
rect 3356 2476 3383 2480
rect 3236 2436 3263 2443
rect 3016 2256 3023 2293
rect 2996 2220 3003 2223
rect 2993 2207 3007 2220
rect 3036 1956 3043 1993
rect 3016 1920 3023 1923
rect 3013 1907 3027 1920
rect 3056 1907 3063 2093
rect 3076 1827 3083 2033
rect 3096 1987 3103 2353
rect 3156 2287 3163 2333
rect 3236 2327 3243 2436
rect 3156 2256 3163 2273
rect 3116 2187 3123 2253
rect 3136 2007 3143 2213
rect 3176 2147 3183 2223
rect 3236 2023 3243 2213
rect 3256 2047 3263 2333
rect 3316 2263 3323 2413
rect 3296 2256 3323 2263
rect 3333 2260 3347 2273
rect 3336 2256 3343 2260
rect 3376 2256 3383 2453
rect 3396 2347 3403 2533
rect 3416 2427 3423 2573
rect 3476 2507 3483 2856
rect 3496 2647 3503 2963
rect 3616 2783 3623 2952
rect 3693 2947 3707 2953
rect 3616 2776 3643 2783
rect 3516 2736 3543 2743
rect 3596 2740 3603 2743
rect 3516 2607 3523 2736
rect 3593 2727 3607 2740
rect 3596 2667 3603 2713
rect 3500 2503 3513 2507
rect 3487 2496 3513 2503
rect 3500 2493 3513 2496
rect 3476 2423 3483 2443
rect 3476 2416 3503 2423
rect 3276 2226 3283 2254
rect 3296 2227 3303 2256
rect 3356 2220 3363 2223
rect 3276 2067 3283 2212
rect 3296 2147 3303 2192
rect 3316 2167 3323 2212
rect 3353 2207 3367 2220
rect 3216 2016 3243 2023
rect 3133 1960 3147 1972
rect 3136 1956 3143 1960
rect 3176 1956 3183 1993
rect 3216 1967 3223 2016
rect 2976 1743 2983 1813
rect 2956 1736 2983 1743
rect 2993 1740 3007 1753
rect 2996 1736 3003 1740
rect 3036 1736 3043 1773
rect 2816 1627 2823 1692
rect 2836 1667 2843 1703
rect 2896 1700 2903 1703
rect 2893 1687 2907 1700
rect 2956 1687 2963 1736
rect 3096 1743 3103 1952
rect 3156 1920 3163 1923
rect 3153 1907 3167 1920
rect 3087 1736 3103 1743
rect 3056 1700 3063 1703
rect 3053 1687 3067 1700
rect 2776 1616 2803 1623
rect 2736 1556 2753 1567
rect 2740 1553 2753 1556
rect 2736 1436 2743 1533
rect 2776 1487 2783 1616
rect 2896 1436 2903 1473
rect 2936 1436 2943 1513
rect 2756 1367 2763 1403
rect 2756 1267 2763 1332
rect 2773 1220 2787 1233
rect 2776 1216 2783 1220
rect 2507 1156 2523 1163
rect 2416 943 2423 1113
rect 2416 936 2443 943
rect 2436 916 2443 936
rect 2396 667 2403 873
rect 2416 847 2423 883
rect 2456 727 2463 883
rect 2460 703 2473 707
rect 2456 696 2473 703
rect 2460 693 2473 696
rect 1776 187 1783 213
rect 1547 183 1560 187
rect 1547 176 1563 183
rect 1547 173 1560 176
rect 576 107 583 143
rect 676 140 683 143
rect 673 127 687 140
rect 1296 127 1303 153
rect 1316 146 1323 173
rect 1416 140 1423 143
rect 1413 127 1427 140
rect 1696 140 1703 143
rect 1693 127 1707 140
rect 1816 87 1823 174
rect 1933 127 1947 132
rect 1996 123 2003 143
rect 1996 116 2023 123
rect 2016 87 2023 116
rect 2216 -24 2223 233
rect 2376 207 2383 363
rect 2416 247 2423 413
rect 2456 367 2463 553
rect 2496 427 2503 853
rect 2516 847 2523 1156
rect 2576 1147 2583 1183
rect 2616 1180 2623 1183
rect 2613 1167 2627 1180
rect 2676 923 2683 1213
rect 2696 1147 2703 1214
rect 2716 987 2723 1033
rect 2656 916 2683 923
rect 2716 916 2723 973
rect 2596 880 2603 883
rect 2593 867 2607 880
rect 2556 696 2563 733
rect 2600 723 2613 727
rect 2596 713 2613 723
rect 2596 696 2603 713
rect 2516 527 2523 693
rect 2576 627 2583 663
rect 2616 527 2623 663
rect 2496 396 2503 413
rect 2516 360 2523 363
rect 2513 347 2527 360
rect 2507 317 2533 324
rect 2413 180 2427 193
rect 2416 176 2423 180
rect 2456 147 2463 233
rect 2276 -17 2283 143
rect 2256 -24 2283 -17
rect 2376 -17 2383 143
rect 2496 143 2503 292
rect 2576 287 2583 513
rect 2656 467 2663 916
rect 2836 923 2843 1393
rect 2856 1347 2863 1433
rect 2876 1216 2883 1353
rect 2916 1216 2923 1273
rect 2956 1227 2963 1403
rect 2996 1247 3003 1653
rect 3036 1406 3043 1573
rect 3053 1447 3067 1453
rect 3076 1436 3083 1553
rect 3116 1487 3123 1773
rect 3136 1547 3143 1753
rect 3156 1747 3163 1793
rect 3176 1748 3183 1833
rect 3196 1827 3203 1923
rect 3236 1767 3243 1993
rect 3256 1907 3263 1973
rect 3356 1956 3363 2133
rect 3396 2107 3403 2223
rect 3436 2023 3443 2273
rect 3456 2147 3463 2353
rect 3496 2256 3503 2416
rect 3516 2287 3523 2443
rect 3556 2407 3563 2593
rect 3576 2367 3583 2633
rect 3596 2547 3603 2593
rect 3636 2587 3643 2776
rect 3656 2727 3663 2773
rect 3676 2746 3683 2873
rect 3716 2807 3723 3173
rect 3756 3007 3763 3153
rect 3736 2927 3743 2994
rect 3816 2996 3823 3173
rect 3956 3028 3963 3773
rect 3976 3767 3983 4033
rect 3996 3767 4003 4173
rect 4116 4107 4123 4336
rect 4156 4067 4163 4292
rect 4033 4040 4047 4053
rect 4073 4040 4087 4053
rect 4036 4036 4043 4040
rect 4076 4036 4083 4040
rect 4036 3816 4043 3853
rect 4136 3823 4143 4053
rect 4176 4043 4183 4193
rect 4156 4036 4183 4043
rect 4216 4036 4223 4133
rect 4236 4063 4243 4523
rect 4476 4523 4483 4753
rect 4536 4587 4543 4633
rect 4533 4560 4547 4573
rect 4536 4556 4543 4560
rect 4576 4556 4583 4593
rect 4596 4563 4603 4813
rect 4616 4587 4623 4823
rect 4656 4820 4663 4823
rect 4653 4807 4667 4820
rect 4716 4807 4723 5036
rect 4736 4967 4743 5043
rect 4787 4993 4793 5007
rect 4816 4856 4823 5013
rect 4836 5007 4843 5073
rect 4996 5046 5003 5073
rect 4876 5023 4883 5043
rect 4916 5040 4923 5043
rect 4913 5027 4927 5040
rect 4856 5020 4883 5023
rect 4853 5016 4883 5020
rect 4896 5016 4913 5023
rect 4853 5007 4867 5016
rect 4836 4887 4843 4913
rect 4876 4826 4883 4993
rect 4656 4647 4663 4793
rect 4676 4567 4683 4793
rect 4756 4607 4763 4813
rect 4596 4556 4623 4563
rect 4396 4467 4403 4523
rect 4476 4516 4503 4523
rect 4256 4306 4263 4373
rect 4376 4307 4383 4393
rect 4296 4187 4303 4303
rect 4336 4247 4343 4292
rect 4236 4056 4263 4063
rect 4256 4036 4263 4056
rect 4156 4007 4163 4036
rect 4187 4003 4200 4007
rect 4187 3996 4203 4003
rect 4187 3993 4200 3996
rect 4296 3867 4303 4093
rect 4136 3816 4153 3823
rect 4156 3787 4163 3814
rect 4056 3780 4063 3783
rect 4016 3607 4023 3773
rect 4053 3767 4067 3780
rect 4196 3707 4203 3783
rect 4236 3747 4243 3783
rect 3976 3247 3983 3453
rect 4016 3447 4023 3483
rect 4096 3467 4103 3514
rect 4096 3296 4103 3333
rect 4116 3303 4123 3573
rect 4196 3516 4203 3593
rect 4176 3427 4183 3483
rect 4216 3367 4223 3472
rect 4116 3296 4143 3303
rect 3996 3247 4003 3293
rect 4036 3260 4043 3263
rect 4033 3247 4047 3260
rect 4076 3247 4083 3263
rect 3993 3227 4007 3233
rect 3740 2803 3753 2807
rect 3736 2793 3753 2803
rect 3736 2776 3743 2793
rect 3756 2736 3773 2743
rect 3747 2713 3753 2727
rect 3776 2707 3783 2732
rect 3596 2436 3623 2443
rect 3556 2187 3563 2223
rect 3496 2087 3503 2113
rect 3416 2016 3443 2023
rect 3396 1927 3403 1954
rect 3256 1747 3263 1813
rect 3276 1787 3283 1913
rect 3296 1847 3303 1923
rect 3316 1803 3323 1893
rect 3307 1796 3323 1803
rect 3196 1700 3203 1703
rect 3156 1607 3163 1693
rect 3193 1687 3207 1700
rect 3276 1706 3283 1752
rect 3256 1587 3263 1693
rect 3113 1440 3127 1452
rect 3116 1436 3123 1440
rect 3136 1267 3143 1403
rect 3176 1367 3183 1413
rect 2976 1186 2983 1213
rect 2956 928 2963 1173
rect 2996 1167 3003 1233
rect 3036 1180 3043 1183
rect 3076 1180 3083 1183
rect 3033 1167 3047 1180
rect 3073 1167 3087 1180
rect 3116 1167 3123 1233
rect 3176 1216 3183 1353
rect 3196 1347 3203 1473
rect 3256 1436 3263 1473
rect 3276 1467 3283 1692
rect 3296 1687 3303 1793
rect 3320 1786 3340 1787
rect 3327 1773 3333 1786
rect 3373 1740 3387 1753
rect 3416 1743 3423 2016
rect 3436 1926 3443 1993
rect 3476 1968 3483 1993
rect 3516 1956 3523 2053
rect 3556 1956 3563 2033
rect 3596 2003 3603 2436
rect 3616 2163 3623 2273
rect 3713 2260 3727 2273
rect 3736 2267 3743 2553
rect 3756 2446 3763 2493
rect 3716 2256 3723 2260
rect 3756 2226 3763 2253
rect 3656 2187 3663 2223
rect 3616 2156 3643 2163
rect 3596 1996 3623 2003
rect 3496 1887 3503 1923
rect 3596 1907 3603 1973
rect 3587 1886 3600 1887
rect 3587 1873 3593 1886
rect 3616 1847 3623 1996
rect 3636 1987 3643 2156
rect 3676 2127 3683 2153
rect 3696 2107 3703 2212
rect 3716 2047 3723 2173
rect 3687 1993 3693 2007
rect 3716 1963 3723 2033
rect 3776 2003 3783 2653
rect 3796 2587 3803 2793
rect 3816 2687 3823 2913
rect 3836 2567 3843 2793
rect 3856 2727 3863 2833
rect 3896 2807 3903 3013
rect 3996 2996 4003 3053
rect 3936 2927 3943 2963
rect 3916 2776 3923 2873
rect 3840 2503 3853 2507
rect 3836 2493 3853 2503
rect 3836 2476 3843 2493
rect 3876 2447 3883 2474
rect 3896 2447 3903 2673
rect 3936 2547 3943 2743
rect 3956 2507 3963 2793
rect 3976 2527 3983 2963
rect 4036 2947 4043 2993
rect 4076 2967 4083 3233
rect 4136 3067 4143 3296
rect 4156 3266 4163 3353
rect 4276 3343 4283 3633
rect 4296 3528 4303 3853
rect 4316 3827 4323 4213
rect 4396 4087 4403 4333
rect 4456 4067 4463 4303
rect 4496 4227 4503 4516
rect 4556 4467 4563 4523
rect 4616 4427 4623 4556
rect 4713 4560 4727 4573
rect 4716 4556 4723 4560
rect 4756 4556 4763 4593
rect 4636 4527 4643 4553
rect 4516 4287 4523 4413
rect 4576 4336 4583 4373
rect 4556 4300 4563 4303
rect 4553 4287 4567 4300
rect 4596 4167 4603 4303
rect 4453 4047 4467 4053
rect 4467 4036 4483 4043
rect 4396 3907 4403 4003
rect 4456 3967 4463 4012
rect 4396 3816 4403 3853
rect 4336 3767 4343 3783
rect 4336 3667 4343 3753
rect 4376 3607 4383 3783
rect 4416 3780 4423 3783
rect 4413 3767 4427 3780
rect 4476 3767 4483 4036
rect 4553 4040 4567 4053
rect 4556 4036 4563 4040
rect 4616 4003 4623 4273
rect 4536 3907 4543 4003
rect 4576 3996 4623 4003
rect 4536 3867 4543 3893
rect 4556 3816 4563 3933
rect 4496 3787 4503 3814
rect 4536 3780 4543 3783
rect 4533 3767 4547 3780
rect 4416 3567 4423 3753
rect 4576 3707 4583 3772
rect 4316 3516 4323 3553
rect 4276 3336 4303 3343
rect 4216 3316 4273 3323
rect 4216 3296 4223 3316
rect 4236 3167 4243 3263
rect 4173 3000 4187 3013
rect 4176 2996 4183 3000
rect 4036 2776 4043 2912
rect 4116 2783 4123 2963
rect 4116 2776 4143 2783
rect 4056 2740 4063 2743
rect 4053 2727 4067 2740
rect 3816 2267 3823 2432
rect 3916 2387 3923 2493
rect 3973 2480 3987 2492
rect 3976 2476 3983 2480
rect 3916 2287 3923 2373
rect 3936 2303 3943 2433
rect 3956 2407 3963 2443
rect 3956 2327 3963 2393
rect 4056 2347 4063 2573
rect 4136 2503 4143 2776
rect 4196 2776 4203 2952
rect 4236 2867 4243 3053
rect 4256 2807 4263 3113
rect 4296 3027 4303 3336
rect 4316 3067 4323 3433
rect 4336 3307 4343 3483
rect 4416 3407 4423 3532
rect 4453 3520 4467 3533
rect 4456 3516 4463 3520
rect 4373 3300 4387 3313
rect 4376 3296 4383 3300
rect 4347 3263 4360 3267
rect 4347 3256 4363 3263
rect 4347 3253 4360 3256
rect 4336 3207 4343 3253
rect 4396 3187 4403 3263
rect 4436 3227 4443 3273
rect 4456 3127 4463 3293
rect 4476 3287 4483 3333
rect 4536 3323 4543 3693
rect 4636 3667 4643 4293
rect 4656 4287 4663 4334
rect 4676 4307 4683 4513
rect 4736 4503 4743 4523
rect 4736 4500 4763 4503
rect 4736 4496 4767 4500
rect 4736 4467 4743 4496
rect 4753 4487 4767 4496
rect 4696 4303 4703 4393
rect 4776 4376 4783 4513
rect 4796 4507 4803 4673
rect 4816 4523 4823 4633
rect 4836 4567 4843 4812
rect 4896 4607 4903 5016
rect 4916 4826 4923 4973
rect 5056 4927 5063 5032
rect 5096 5023 5103 5043
rect 5096 5016 5123 5023
rect 4947 4863 4960 4867
rect 4947 4856 4963 4863
rect 4947 4853 4960 4856
rect 5056 4827 5063 4854
rect 4873 4560 4887 4573
rect 4876 4556 4883 4560
rect 4936 4563 4943 4813
rect 4973 4807 4987 4812
rect 5016 4727 5023 4823
rect 5076 4687 5083 4973
rect 5096 4747 5103 4993
rect 5116 4907 5123 5016
rect 5136 5007 5143 5113
rect 5156 4987 5163 5273
rect 5216 5040 5223 5043
rect 5213 5027 5227 5040
rect 5256 4963 5263 5376
rect 5396 5346 5403 5493
rect 5456 5467 5463 5613
rect 5513 5600 5527 5613
rect 5516 5596 5523 5600
rect 5496 5507 5503 5563
rect 5533 5547 5547 5552
rect 5276 5307 5283 5333
rect 5393 5327 5407 5332
rect 5416 5127 5423 5393
rect 5436 5387 5443 5413
rect 5456 5403 5463 5453
rect 5456 5396 5483 5403
rect 5476 5376 5483 5396
rect 5556 5347 5563 5374
rect 5496 5340 5503 5343
rect 5493 5327 5507 5340
rect 5476 5187 5483 5293
rect 5576 5247 5583 5393
rect 5427 5116 5443 5123
rect 5376 5076 5383 5113
rect 5416 5043 5423 5074
rect 5316 5040 5323 5043
rect 5313 5027 5327 5040
rect 5236 4956 5263 4963
rect 5156 4856 5163 4913
rect 5213 4863 5227 4873
rect 5207 4860 5227 4863
rect 5207 4856 5223 4860
rect 5136 4820 5143 4823
rect 5133 4807 5147 4820
rect 5176 4647 5183 4823
rect 5196 4667 5203 4733
rect 4927 4556 4943 4563
rect 4816 4516 4863 4523
rect 4816 4336 4843 4343
rect 4696 4296 4713 4303
rect 4656 4007 4663 4153
rect 4716 4036 4723 4073
rect 4796 4007 4803 4133
rect 4716 3816 4723 3953
rect 4736 3947 4743 4003
rect 4576 3427 4583 3653
rect 4656 3587 4663 3813
rect 4696 3780 4703 3783
rect 4693 3767 4707 3780
rect 4653 3520 4667 3533
rect 4656 3516 4663 3520
rect 4516 3316 4543 3323
rect 4516 3308 4523 3316
rect 4576 3263 4583 3413
rect 4636 3407 4643 3483
rect 4676 3447 4683 3653
rect 4796 3647 4803 3813
rect 4816 3707 4823 4233
rect 4836 4187 4843 4336
rect 4856 4247 4863 4493
rect 4956 4407 4963 4593
rect 4976 4383 4983 4573
rect 5176 4567 5183 4633
rect 5196 4556 5203 4653
rect 5216 4583 5223 4813
rect 5236 4627 5243 4956
rect 5256 4587 5263 4893
rect 5356 4887 5363 5043
rect 5396 5036 5423 5043
rect 5333 4860 5347 4873
rect 5336 4856 5343 4860
rect 5216 4576 5243 4583
rect 5236 4556 5243 4576
rect 5276 4567 5283 4813
rect 5316 4767 5323 4823
rect 5396 4723 5403 5036
rect 5416 4826 5423 4913
rect 5436 4867 5443 5116
rect 5476 5076 5483 5173
rect 5516 5076 5523 5113
rect 5596 5047 5603 5813
rect 5676 5680 5723 5683
rect 5676 5676 5727 5680
rect 5676 5627 5683 5676
rect 5713 5667 5727 5676
rect 5696 5608 5703 5653
rect 5736 5607 5743 5863
rect 5676 5543 5683 5552
rect 5656 5536 5683 5543
rect 5656 5376 5663 5536
rect 5693 5380 5707 5393
rect 5716 5387 5723 5563
rect 5696 5376 5703 5380
rect 5736 5347 5743 5553
rect 5756 5527 5763 5833
rect 5796 5763 5803 5894
rect 5816 5847 5823 5913
rect 5853 5900 5867 5913
rect 5856 5896 5863 5900
rect 5776 5756 5803 5763
rect 5776 5423 5783 5756
rect 5816 5596 5823 5713
rect 5856 5608 5863 5653
rect 5876 5607 5883 5863
rect 5796 5467 5803 5553
rect 5836 5427 5843 5563
rect 5776 5416 5793 5423
rect 5796 5376 5803 5413
rect 5876 5387 5883 5453
rect 5636 5340 5643 5343
rect 5616 5167 5623 5333
rect 5633 5327 5647 5340
rect 5727 5336 5743 5347
rect 5727 5333 5740 5336
rect 5653 5080 5667 5093
rect 5693 5080 5707 5093
rect 5656 5076 5663 5080
rect 5696 5076 5703 5080
rect 5496 4927 5503 5043
rect 5536 5007 5543 5043
rect 5453 4860 5467 4873
rect 5456 4856 5463 4860
rect 5496 4856 5503 4913
rect 5433 4807 5447 4813
rect 5473 4807 5487 4812
rect 5516 4787 5523 4823
rect 5556 4787 5563 5033
rect 5636 5007 5643 5043
rect 5596 4867 5603 4913
rect 5636 4883 5643 4993
rect 5616 4876 5643 4883
rect 5576 4823 5583 4854
rect 5616 4856 5623 4876
rect 5576 4816 5603 4823
rect 5473 4767 5487 4772
rect 5396 4716 5413 4723
rect 5036 4487 5043 4523
rect 5113 4507 5127 4513
rect 4976 4376 4993 4383
rect 5036 4336 5063 4343
rect 5056 4187 5063 4336
rect 5096 4287 5103 4393
rect 5136 4367 5143 4553
rect 5160 4526 5173 4527
rect 5167 4513 5173 4526
rect 5136 4336 5143 4353
rect 5236 4327 5243 4453
rect 5296 4343 5303 4573
rect 5316 4367 5323 4613
rect 5376 4556 5383 4653
rect 5416 4568 5423 4713
rect 5356 4467 5363 4523
rect 5456 4523 5463 4573
rect 5436 4516 5463 4523
rect 5276 4336 5303 4343
rect 5336 4336 5343 4413
rect 5196 4300 5203 4303
rect 5193 4287 5207 4300
rect 4916 4036 4923 4073
rect 4956 4007 4963 4034
rect 4896 3947 4903 4003
rect 4876 3816 4883 3853
rect 4936 3786 4943 3853
rect 4976 3816 4983 4073
rect 5056 4036 5063 4073
rect 5196 4036 5203 4073
rect 5256 4067 5263 4333
rect 5276 4087 5283 4336
rect 5316 4207 5323 4292
rect 5356 4127 5363 4303
rect 5396 4147 5403 4353
rect 5416 4127 5423 4493
rect 5436 4347 5443 4516
rect 5456 4336 5463 4493
rect 5476 4427 5483 4753
rect 5513 4560 5527 4573
rect 5516 4556 5523 4560
rect 5556 4556 5563 4633
rect 5596 4568 5603 4816
rect 5536 4520 5543 4523
rect 5533 4507 5547 4520
rect 5520 4303 5533 4307
rect 5476 4300 5483 4303
rect 5473 4287 5487 4300
rect 5516 4296 5533 4303
rect 5520 4293 5533 4296
rect 5136 3907 5143 4034
rect 4996 3747 5003 3783
rect 5076 3723 5083 3893
rect 5153 3847 5167 3853
rect 5176 3828 5183 3992
rect 5216 3967 5223 4003
rect 5256 3967 5263 4003
rect 5296 3927 5303 4034
rect 5096 3747 5103 3813
rect 5156 3780 5163 3783
rect 5153 3767 5167 3780
rect 5196 3727 5203 3783
rect 5216 3747 5223 3773
rect 5067 3716 5083 3723
rect 4696 3387 4703 3533
rect 4776 3516 4783 3553
rect 4667 3313 4673 3327
rect 4496 3187 4503 3263
rect 4556 3256 4583 3263
rect 4313 3000 4327 3013
rect 4447 3013 4453 3027
rect 4353 3000 4367 3013
rect 4316 2996 4323 3000
rect 4356 2996 4363 3000
rect 4296 2960 4303 2963
rect 4293 2947 4307 2960
rect 4336 2927 4343 2963
rect 4396 2947 4403 2994
rect 4416 2987 4423 3013
rect 4473 3000 4487 3013
rect 4476 2996 4483 3000
rect 4156 2667 4163 2774
rect 4216 2627 4223 2732
rect 4253 2727 4267 2732
rect 4256 2687 4263 2713
rect 4116 2496 4143 2503
rect 4116 2488 4123 2496
rect 4156 2476 4163 2513
rect 3936 2296 3963 2303
rect 3816 2047 3823 2213
rect 3756 1996 3783 2003
rect 3696 1956 3723 1963
rect 3713 1907 3727 1913
rect 3647 1873 3653 1887
rect 3376 1736 3383 1740
rect 3416 1736 3443 1743
rect 3356 1700 3363 1703
rect 3353 1687 3367 1700
rect 3396 1667 3403 1703
rect 3216 1247 3223 1293
rect 3236 1167 3243 1213
rect 3256 1187 3263 1373
rect 3276 1347 3283 1403
rect 3336 1387 3343 1434
rect 3356 1407 3363 1633
rect 3436 1487 3443 1736
rect 3533 1747 3547 1753
rect 3467 1736 3503 1743
rect 3456 1607 3463 1734
rect 3556 1727 3563 1773
rect 3516 1700 3523 1703
rect 3513 1687 3527 1700
rect 3556 1687 3563 1713
rect 3316 1216 3323 1333
rect 3376 1307 3383 1453
rect 3396 1436 3403 1473
rect 3476 1406 3483 1653
rect 3516 1406 3523 1533
rect 3576 1487 3583 1733
rect 3536 1307 3543 1473
rect 3596 1463 3603 1733
rect 3636 1647 3643 1703
rect 3696 1587 3703 1653
rect 3576 1456 3603 1463
rect 3576 1448 3583 1456
rect 3616 1436 3623 1473
rect 3353 1220 3367 1233
rect 3356 1216 3363 1220
rect 3336 1180 3343 1183
rect 3333 1167 3347 1180
rect 3073 1147 3087 1153
rect 2836 916 2863 923
rect 2696 807 2703 883
rect 2796 827 2803 914
rect 2816 847 2823 872
rect 2876 787 2883 883
rect 2676 647 2683 773
rect 2956 767 2963 914
rect 2716 696 2723 753
rect 2696 467 2703 653
rect 2736 567 2743 663
rect 2496 136 2523 143
rect 2576 140 2583 143
rect 2573 127 2587 140
rect 2596 87 2603 453
rect 2613 403 2627 413
rect 2613 400 2643 403
rect 2616 396 2643 400
rect 2616 67 2623 353
rect 2676 203 2683 273
rect 2696 223 2703 323
rect 2696 220 2723 223
rect 2696 216 2727 220
rect 2713 207 2727 216
rect 2676 196 2703 203
rect 2696 176 2703 196
rect 2636 147 2643 174
rect 2716 140 2723 143
rect 2713 127 2727 140
rect 2756 127 2763 633
rect 2816 563 2823 694
rect 2836 666 2843 733
rect 2936 696 2943 733
rect 2876 660 2883 663
rect 2873 647 2887 660
rect 2916 607 2923 663
rect 2816 556 2833 563
rect 2836 396 2843 553
rect 2936 366 2943 473
rect 2976 403 2983 693
rect 2996 547 3003 853
rect 3016 847 3023 883
rect 3076 867 3083 914
rect 3196 916 3203 953
rect 3236 916 3243 993
rect 3376 987 3383 1173
rect 3396 1107 3403 1233
rect 3113 907 3127 913
rect 3107 900 3127 907
rect 3107 896 3123 900
rect 3107 893 3120 896
rect 3276 886 3283 953
rect 3176 867 3183 883
rect 3296 867 3303 914
rect 3173 847 3187 853
rect 3096 696 3103 793
rect 3256 767 3263 793
rect 3356 787 3363 883
rect 3036 660 3043 663
rect 3033 647 3047 660
rect 3076 643 3083 663
rect 3076 636 3103 643
rect 2976 396 3003 403
rect 3036 396 3043 633
rect 2856 327 2863 363
rect 2776 127 2783 233
rect 2873 180 2887 193
rect 2876 176 2883 180
rect 2956 146 2963 193
rect 3016 176 3023 213
rect 2896 140 2903 143
rect 2893 127 2907 140
rect 3033 127 3047 132
rect 2376 -24 2403 -17
rect 2656 -24 2663 53
rect 3076 27 3083 533
rect 3096 487 3103 636
rect 3136 627 3143 693
rect 3116 467 3123 593
rect 3136 567 3143 613
rect 3156 527 3163 753
rect 3236 708 3243 733
rect 3316 666 3323 773
rect 3416 727 3423 1253
rect 3493 1220 3507 1233
rect 3496 1216 3503 1220
rect 3556 1186 3563 1253
rect 3676 1247 3683 1533
rect 3716 1487 3723 1853
rect 3736 1706 3743 1993
rect 3756 1867 3763 1996
rect 3796 1956 3803 1993
rect 3836 1987 3843 2223
rect 3876 2127 3883 2223
rect 3936 2047 3943 2253
rect 3956 2187 3963 2296
rect 3833 1960 3847 1973
rect 3836 1956 3843 1960
rect 3816 1887 3823 1912
rect 3776 1736 3783 1833
rect 3816 1736 3823 1852
rect 3856 1807 3863 1923
rect 3476 1147 3483 1183
rect 3476 1007 3483 1133
rect 3516 967 3523 993
rect 3516 916 3523 953
rect 3553 920 3567 933
rect 3556 916 3563 920
rect 3456 727 3463 913
rect 3596 887 3603 1214
rect 3656 1047 3663 1183
rect 3656 948 3663 1033
rect 3696 947 3703 1433
rect 3736 1407 3743 1593
rect 3796 1467 3803 1703
rect 3856 1547 3863 1733
rect 3876 1706 3883 1893
rect 3896 1747 3903 2033
rect 3936 1963 3943 2033
rect 3916 1956 3943 1963
rect 3916 1926 3923 1956
rect 3996 1967 4003 2212
rect 4076 2163 4083 2473
rect 4136 2407 4143 2443
rect 4116 2396 4133 2403
rect 4096 2226 4103 2353
rect 4056 2156 4083 2163
rect 4016 1867 4023 2053
rect 3933 1740 3947 1753
rect 3936 1736 3943 1740
rect 3996 1727 4003 1773
rect 4036 1743 4043 1953
rect 4016 1736 4043 1743
rect 4056 1736 4063 2156
rect 4076 1956 4083 2133
rect 4116 2067 4123 2396
rect 4196 2367 4203 2493
rect 4216 2407 4223 2553
rect 4236 2487 4243 2653
rect 4276 2476 4283 2553
rect 4296 2507 4303 2793
rect 4236 2223 4243 2333
rect 4316 2303 4323 2833
rect 4356 2788 4363 2853
rect 4416 2747 4423 2973
rect 4456 2960 4463 2963
rect 4453 2947 4467 2960
rect 4496 2927 4503 2963
rect 4536 2776 4543 2813
rect 4556 2807 4563 2993
rect 4476 2740 4483 2743
rect 4516 2740 4523 2743
rect 4336 2446 4343 2613
rect 4376 2476 4383 2673
rect 4416 2587 4423 2733
rect 4473 2727 4487 2740
rect 4513 2727 4527 2740
rect 4556 2627 4563 2733
rect 4416 2476 4423 2552
rect 4296 2296 4323 2303
rect 4256 2227 4263 2254
rect 4156 2187 4163 2223
rect 4216 2216 4243 2223
rect 4136 1956 4143 2113
rect 4236 2067 4243 2216
rect 4236 1963 4243 2053
rect 4256 2007 4263 2213
rect 4296 2207 4303 2296
rect 4313 2260 4327 2273
rect 4316 2256 4323 2260
rect 4396 2226 4403 2273
rect 4296 2127 4303 2153
rect 4296 1968 4303 2113
rect 4236 1956 4263 1963
rect 4160 1926 4173 1927
rect 4167 1913 4173 1926
rect 4216 1907 4223 1953
rect 4233 1907 4247 1913
rect 3956 1667 3963 1703
rect 3896 1267 3903 1453
rect 3916 1287 3923 1653
rect 4016 1647 4023 1736
rect 4236 1736 4243 1833
rect 4076 1667 4083 1703
rect 4116 1700 4123 1703
rect 4113 1687 4127 1700
rect 4296 1706 4303 1734
rect 4016 1436 4023 1473
rect 4136 1327 4143 1693
rect 4213 1687 4227 1692
rect 4267 1653 4273 1667
rect 4256 1467 4263 1493
rect 4253 1440 4267 1453
rect 4256 1436 4263 1440
rect 3896 1243 3903 1253
rect 3896 1236 3923 1243
rect 3716 1167 3723 1233
rect 3800 1223 3813 1227
rect 3796 1216 3813 1223
rect 3800 1213 3813 1216
rect 3916 1216 3923 1236
rect 3776 1147 3783 1183
rect 3856 1087 3863 1213
rect 3896 1180 3903 1183
rect 3936 1180 3943 1183
rect 3893 1167 3907 1180
rect 3933 1167 3947 1180
rect 3936 1007 3943 1153
rect 3696 916 3743 923
rect 3496 827 3503 883
rect 3536 827 3543 883
rect 3736 867 3743 916
rect 3416 696 3463 703
rect 3216 643 3223 663
rect 3216 636 3233 643
rect 3196 396 3203 473
rect 3116 367 3123 394
rect 3236 367 3243 633
rect 3256 627 3263 663
rect 3356 660 3363 663
rect 3316 627 3323 652
rect 3353 647 3367 660
rect 3456 647 3463 696
rect 3336 467 3343 493
rect 3336 396 3343 453
rect 3376 267 3383 553
rect 3293 180 3307 193
rect 3296 176 3303 180
rect 3236 146 3243 173
rect 3136 87 3143 143
rect 3176 27 3183 143
rect 3376 107 3383 193
rect 3396 146 3403 433
rect 3436 367 3443 453
rect 3456 427 3463 513
rect 3476 447 3483 713
rect 3493 707 3507 713
rect 3536 696 3543 753
rect 3520 645 3533 647
rect 3527 633 3533 645
rect 3556 467 3563 652
rect 3616 567 3623 813
rect 3696 696 3703 753
rect 3756 703 3763 933
rect 3956 928 3963 973
rect 3996 916 4003 1213
rect 4016 1167 4023 1313
rect 4156 1303 4163 1434
rect 4296 1407 4303 1692
rect 4316 1523 4323 1753
rect 4336 1687 4343 2193
rect 4356 2187 4363 2212
rect 4396 1987 4403 2212
rect 4436 2007 4443 2443
rect 4476 2287 4483 2493
rect 4496 2446 4503 2573
rect 4556 2476 4563 2573
rect 4576 2507 4583 3256
rect 4596 3227 4603 3293
rect 4616 3287 4623 3313
rect 4647 3303 4660 3307
rect 4647 3296 4663 3303
rect 4696 3296 4703 3333
rect 4736 3307 4743 3373
rect 4647 3293 4660 3296
rect 4676 3260 4683 3263
rect 4673 3247 4687 3260
rect 4756 3263 4763 3433
rect 4736 3256 4763 3263
rect 4636 3008 4643 3213
rect 4607 2963 4620 2967
rect 4607 2956 4623 2963
rect 4607 2953 4620 2956
rect 4656 2887 4663 2963
rect 4716 2947 4723 3033
rect 4596 2727 4603 2793
rect 4636 2776 4643 2813
rect 4676 2776 4683 2913
rect 4713 2787 4727 2793
rect 4656 2727 4663 2743
rect 4596 2627 4603 2653
rect 4596 2476 4603 2613
rect 4496 2256 4503 2293
rect 4476 2187 4483 2223
rect 4356 1787 4363 1973
rect 4396 1956 4403 1973
rect 4476 1967 4483 2173
rect 4556 2127 4563 2193
rect 4456 1867 4463 1923
rect 4496 1787 4503 1993
rect 4516 1787 4523 1973
rect 4556 1956 4563 2053
rect 4576 1987 4583 2443
rect 4596 2147 4603 2293
rect 4636 2287 4643 2533
rect 4656 2447 4663 2713
rect 4716 2587 4723 2733
rect 4736 2727 4743 3256
rect 4796 3047 4803 3483
rect 4856 3387 4863 3514
rect 4896 3487 4903 3673
rect 4973 3528 4987 3533
rect 4956 3480 4963 3483
rect 4953 3467 4967 3480
rect 4813 3308 4827 3313
rect 4856 3296 4863 3373
rect 4956 3347 4963 3453
rect 5036 3387 5043 3513
rect 5056 3487 5063 3713
rect 5076 3486 5083 3633
rect 5107 3523 5120 3527
rect 5107 3516 5123 3523
rect 5107 3513 5120 3516
rect 5196 3527 5203 3553
rect 5180 3483 5193 3487
rect 5176 3476 5193 3483
rect 5180 3473 5193 3476
rect 4836 3247 4843 3263
rect 4827 3236 4843 3247
rect 4827 3233 4840 3236
rect 4956 3047 4963 3252
rect 5016 3227 5023 3263
rect 5076 3187 5083 3313
rect 5133 3300 5147 3313
rect 5136 3296 5143 3300
rect 5176 3296 5183 3453
rect 4833 3000 4847 3013
rect 4836 2996 4843 3000
rect 4776 2783 4783 2963
rect 4816 2960 4823 2963
rect 4813 2947 4827 2960
rect 4816 2807 4823 2933
rect 4756 2776 4783 2783
rect 4756 2627 4763 2776
rect 4836 2776 4843 2873
rect 4876 2863 4883 2973
rect 4896 2887 4903 3013
rect 4996 2996 5003 3033
rect 5036 2987 5043 3173
rect 5116 3047 5123 3263
rect 5216 3227 5223 3693
rect 5236 3547 5243 3913
rect 5316 3847 5323 4053
rect 5353 4040 5367 4053
rect 5356 4036 5363 4040
rect 5376 3947 5383 4003
rect 5416 3967 5423 4003
rect 5476 3927 5483 4252
rect 5496 4006 5503 4193
rect 5516 4036 5523 4273
rect 5556 4267 5563 4453
rect 5576 4307 5583 4512
rect 5636 4348 5643 4554
rect 5656 4467 5663 4793
rect 5676 4767 5683 4823
rect 5716 4763 5723 4854
rect 5736 4807 5743 5313
rect 5756 5207 5763 5373
rect 5773 5327 5787 5333
rect 5816 5247 5823 5343
rect 5856 5327 5863 5343
rect 5756 4867 5763 5153
rect 5796 5088 5803 5113
rect 5836 5107 5843 5253
rect 5856 5127 5863 5313
rect 5876 5107 5883 5333
rect 5896 5267 5903 5413
rect 5836 5076 5843 5093
rect 5776 4856 5783 4913
rect 5856 4867 5863 5043
rect 5796 4820 5803 4823
rect 5793 4807 5807 4820
rect 5796 4767 5803 4793
rect 5716 4756 5743 4763
rect 5676 4387 5683 4673
rect 5736 4568 5743 4756
rect 5773 4560 5787 4573
rect 5776 4556 5783 4560
rect 5716 4347 5723 4512
rect 5756 4487 5763 4523
rect 5816 4507 5823 4773
rect 5836 4527 5843 4812
rect 5853 4787 5867 4793
rect 5896 4687 5903 5193
rect 5916 4587 5923 5593
rect 5976 4868 5983 5173
rect 5996 4887 6003 5513
rect 5956 4820 5963 4823
rect 5936 4587 5943 4813
rect 5953 4807 5967 4820
rect 5616 4300 5623 4303
rect 5613 4287 5627 4300
rect 5656 4247 5663 4303
rect 5576 4036 5583 4113
rect 5287 3843 5300 3847
rect 5287 3833 5303 3843
rect 5256 3786 5263 3833
rect 5296 3816 5303 3833
rect 5336 3816 5343 3893
rect 5396 3783 5403 3913
rect 5516 3828 5523 3873
rect 5356 3727 5363 3783
rect 5376 3776 5403 3783
rect 5376 3743 5383 3776
rect 5416 3767 5423 3814
rect 5376 3736 5403 3743
rect 5296 3516 5303 3613
rect 5236 3487 5243 3512
rect 5376 3467 5383 3514
rect 5396 3443 5403 3736
rect 5456 3528 5463 3783
rect 5496 3528 5503 3751
rect 5556 3727 5563 3853
rect 5576 3786 5583 3893
rect 5576 3747 5583 3772
rect 5596 3723 5603 4193
rect 5696 4087 5703 4293
rect 5716 4207 5723 4312
rect 5616 3827 5623 4053
rect 5636 3907 5643 4073
rect 5736 4067 5743 4373
rect 5756 4267 5763 4413
rect 5776 4347 5783 4493
rect 5836 4487 5843 4513
rect 5816 4247 5823 4303
rect 5740 4043 5753 4047
rect 5736 4036 5753 4043
rect 5740 4033 5753 4036
rect 5636 3816 5643 3853
rect 5656 3847 5663 3993
rect 5676 3967 5683 4003
rect 5716 3947 5723 4003
rect 5716 3867 5723 3933
rect 5676 3816 5683 3853
rect 5776 3827 5783 4133
rect 5856 4087 5863 4573
rect 5933 4560 5947 4573
rect 5936 4556 5943 4560
rect 5956 4363 5963 4523
rect 5956 4356 5983 4363
rect 5976 4336 5983 4356
rect 5996 4347 6003 4813
rect 5876 4063 5883 4333
rect 5956 4267 5963 4303
rect 5876 4056 5903 4063
rect 5896 4048 5903 4056
rect 5796 3887 5803 4033
rect 5836 3887 5843 4003
rect 5856 3828 5863 3973
rect 5876 3947 5883 4003
rect 5576 3716 5603 3723
rect 5376 3436 5403 3443
rect 5316 3308 5323 3353
rect 5236 3266 5243 3293
rect 5093 3000 5107 3013
rect 5096 2996 5103 3000
rect 4876 2856 4903 2863
rect 4896 2747 4903 2856
rect 4936 2783 4943 2963
rect 5156 2963 5163 3033
rect 5116 2956 5163 2963
rect 5176 2927 5183 3213
rect 5216 2996 5223 3033
rect 5256 2996 5263 3293
rect 5336 3247 5343 3263
rect 5327 3233 5333 3247
rect 5376 3147 5383 3436
rect 5436 3387 5443 3483
rect 5476 3480 5483 3483
rect 5473 3467 5487 3480
rect 5536 3407 5543 3514
rect 5556 3467 5563 3613
rect 5576 3527 5583 3716
rect 5596 3627 5603 3693
rect 5616 3567 5623 3773
rect 5696 3687 5703 3772
rect 5653 3520 5667 3533
rect 5656 3516 5663 3520
rect 5576 3383 5583 3473
rect 5636 3463 5643 3483
rect 5660 3463 5673 3467
rect 5636 3456 5673 3463
rect 5556 3376 5583 3383
rect 5656 3453 5673 3456
rect 5396 3247 5403 3294
rect 5236 2943 5243 2963
rect 5216 2936 5243 2943
rect 4916 2776 4943 2783
rect 4956 2776 4963 2813
rect 4716 2476 4723 2533
rect 4736 2327 4743 2443
rect 4656 2256 4663 2313
rect 4756 2187 4763 2413
rect 4776 2367 4783 2433
rect 4796 2427 4803 2713
rect 4816 2407 4823 2693
rect 4856 2583 4863 2732
rect 4836 2576 4863 2583
rect 4836 2487 4843 2576
rect 4916 2547 4923 2776
rect 5176 2776 5183 2873
rect 4976 2727 4983 2743
rect 4973 2707 4987 2713
rect 5016 2607 5023 2732
rect 5076 2627 5083 2774
rect 5116 2740 5123 2743
rect 5113 2727 5127 2740
rect 5116 2667 5123 2713
rect 4876 2476 4883 2533
rect 4816 2256 4823 2353
rect 4896 2327 4903 2443
rect 4936 2367 4943 2433
rect 4936 2256 4943 2313
rect 4956 2287 4963 2533
rect 4976 2447 4983 2593
rect 5036 2476 5043 2533
rect 4596 1956 4603 2133
rect 4716 1956 4723 2033
rect 4656 1927 4663 1954
rect 4576 1920 4583 1923
rect 4573 1907 4587 1920
rect 4736 1867 4743 1923
rect 4776 1847 4783 1923
rect 4796 1823 4803 1853
rect 4776 1816 4803 1823
rect 4376 1667 4383 1703
rect 4367 1656 4383 1667
rect 4367 1653 4380 1656
rect 4316 1516 4343 1523
rect 4316 1367 4323 1493
rect 4116 1296 4163 1303
rect 4116 1256 4123 1296
rect 4156 1216 4183 1223
rect 4036 1183 4043 1213
rect 4036 1176 4063 1183
rect 4176 1127 4183 1216
rect 4216 1186 4223 1313
rect 4276 1216 4283 1253
rect 4336 1223 4343 1516
rect 4436 1467 4443 1773
rect 4596 1706 4603 1773
rect 4373 1440 4387 1453
rect 4413 1440 4427 1453
rect 4456 1447 4463 1533
rect 4516 1527 4523 1703
rect 4376 1436 4383 1440
rect 4416 1436 4423 1440
rect 4336 1216 4363 1223
rect 4056 1087 4063 1113
rect 3816 847 3823 883
rect 3756 696 3783 703
rect 3636 607 3643 693
rect 3707 636 3733 643
rect 3607 543 3620 547
rect 3607 540 3623 543
rect 3607 533 3627 540
rect 3613 527 3627 533
rect 3516 416 3563 423
rect 3456 396 3463 413
rect 3516 396 3523 416
rect 3536 366 3543 393
rect 3556 183 3563 416
rect 3536 176 3563 183
rect 3576 176 3583 473
rect 3616 408 3623 433
rect 3776 427 3783 696
rect 3876 696 3883 853
rect 3896 807 3903 893
rect 3976 847 3983 883
rect 4016 880 4023 883
rect 4013 867 4027 880
rect 4056 863 4063 1073
rect 4076 907 4083 1033
rect 4356 1007 4363 1216
rect 4096 916 4123 923
rect 4316 916 4323 953
rect 4056 856 4073 863
rect 3996 696 4003 793
rect 4076 707 4083 853
rect 4096 847 4103 916
rect 4176 728 4183 843
rect 3856 660 3863 663
rect 3853 647 3867 660
rect 3936 627 3943 694
rect 4016 607 4023 663
rect 4056 627 4063 663
rect 4156 567 4163 663
rect 3653 400 3667 413
rect 3656 396 3663 400
rect 3636 307 3643 363
rect 3616 176 3623 213
rect 3536 146 3543 176
rect 3407 136 3423 143
rect 3476 67 3483 143
rect 3596 140 3603 143
rect 3593 127 3607 140
rect 3696 27 3703 413
rect 3753 400 3767 413
rect 3756 396 3763 400
rect 3776 360 3783 363
rect 3773 347 3787 360
rect 3716 147 3723 273
rect 3856 227 3863 394
rect 3876 367 3883 433
rect 3896 176 3903 493
rect 3976 396 4023 403
rect 4096 396 4103 473
rect 4216 427 4223 713
rect 4236 666 4243 713
rect 4273 700 4287 713
rect 4276 696 4283 700
rect 4316 696 4323 773
rect 4336 727 4343 883
rect 4296 660 4303 663
rect 4336 660 4343 663
rect 4293 647 4307 660
rect 4333 647 4347 660
rect 4376 647 4383 733
rect 4396 507 4403 1353
rect 4476 1267 4483 1473
rect 4556 1448 4563 1671
rect 4596 1436 4603 1473
rect 4496 1387 4503 1433
rect 4527 1403 4540 1407
rect 4527 1396 4543 1403
rect 4527 1393 4540 1396
rect 4496 1327 4503 1373
rect 4493 1220 4507 1233
rect 4496 1216 4503 1220
rect 4556 1216 4563 1253
rect 4576 1247 4583 1403
rect 4616 1267 4623 1393
rect 4636 1247 4643 1613
rect 4676 1487 4683 1703
rect 4716 1700 4723 1703
rect 4713 1687 4727 1700
rect 4656 1267 4663 1433
rect 4696 1400 4703 1403
rect 4693 1387 4707 1400
rect 4736 1267 4743 1353
rect 4587 1236 4603 1243
rect 4436 923 4443 1213
rect 4516 1067 4523 1183
rect 4596 1167 4603 1236
rect 4636 1147 4643 1233
rect 4736 1216 4743 1253
rect 4756 1247 4763 1734
rect 4776 1627 4783 1816
rect 4796 1703 4803 1793
rect 4816 1767 4823 2173
rect 4836 1843 4843 1954
rect 4856 1867 4863 2253
rect 5016 2226 5023 2254
rect 4956 2203 4963 2223
rect 4956 2196 4973 2203
rect 4916 1867 4923 1923
rect 4836 1836 4853 1843
rect 4856 1736 4863 1832
rect 4956 1807 4963 1913
rect 4976 1783 4983 2193
rect 5016 1967 5023 2212
rect 5036 2207 5043 2273
rect 5073 2260 5087 2273
rect 5076 2256 5083 2260
rect 5116 2256 5123 2613
rect 5216 2488 5223 2936
rect 5236 2707 5243 2913
rect 5136 2427 5143 2474
rect 5156 2267 5163 2432
rect 5276 2427 5283 2693
rect 5296 2447 5303 2474
rect 5316 2427 5323 2653
rect 5336 2647 5343 3133
rect 5476 3107 5483 3263
rect 5516 3207 5523 3263
rect 5356 2927 5363 3073
rect 5413 3000 5427 3013
rect 5416 2996 5423 3000
rect 5436 2927 5443 2963
rect 5356 2747 5363 2793
rect 5396 2776 5403 2913
rect 5433 2780 5447 2793
rect 5476 2788 5483 2833
rect 5436 2776 5443 2780
rect 5460 2743 5473 2747
rect 5416 2740 5423 2743
rect 5356 2707 5363 2733
rect 5413 2727 5427 2740
rect 5456 2733 5473 2743
rect 5456 2667 5463 2733
rect 5496 2483 5503 3113
rect 5536 3047 5543 3253
rect 5556 3187 5563 3376
rect 5656 3343 5663 3453
rect 5696 3423 5703 3533
rect 5676 3416 5703 3423
rect 5676 3367 5683 3416
rect 5656 3336 5683 3343
rect 5676 3296 5683 3336
rect 5716 3308 5723 3553
rect 5736 3527 5743 3813
rect 5756 3647 5763 3813
rect 5776 3687 5783 3773
rect 5796 3747 5803 3783
rect 5836 3780 5843 3783
rect 5833 3767 5847 3780
rect 5753 3520 5767 3533
rect 5793 3520 5807 3533
rect 5836 3527 5843 3673
rect 5756 3516 5763 3520
rect 5796 3516 5803 3520
rect 5856 3487 5863 3533
rect 5776 3480 5783 3483
rect 5536 3003 5543 3033
rect 5576 3027 5583 3294
rect 5616 3087 5623 3263
rect 5656 3260 5663 3263
rect 5653 3247 5667 3260
rect 5516 2996 5543 3003
rect 5573 3008 5587 3013
rect 5516 2967 5523 2996
rect 5613 3000 5627 3013
rect 5616 2996 5623 3000
rect 5596 2927 5603 2963
rect 5516 2587 5523 2913
rect 5616 2776 5623 2873
rect 5656 2847 5663 3033
rect 5716 3027 5723 3294
rect 5736 3127 5743 3473
rect 5773 3467 5787 3480
rect 5833 3463 5847 3473
rect 5816 3460 5847 3463
rect 5816 3456 5843 3460
rect 5816 3307 5823 3456
rect 5796 3260 5803 3263
rect 5793 3247 5807 3260
rect 5816 3203 5823 3253
rect 5796 3196 5823 3203
rect 5796 3067 5803 3196
rect 5773 3027 5787 3033
rect 5676 2967 5683 3013
rect 5776 2996 5783 3013
rect 5756 2907 5763 2963
rect 5736 2847 5743 2873
rect 5656 2743 5663 2833
rect 5776 2776 5783 2933
rect 5536 2736 5563 2743
rect 5536 2727 5543 2736
rect 5476 2476 5503 2483
rect 5516 2476 5523 2513
rect 5536 2507 5543 2713
rect 5596 2707 5603 2743
rect 5636 2736 5663 2743
rect 5356 2440 5363 2443
rect 5353 2427 5367 2440
rect 5176 2226 5183 2253
rect 5196 2147 5203 2411
rect 5256 2268 5263 2393
rect 5296 2367 5303 2393
rect 5296 2256 5303 2353
rect 5227 2223 5240 2227
rect 5227 2213 5243 2223
rect 4996 1867 5003 1933
rect 5136 1927 5143 1993
rect 5027 1923 5040 1927
rect 5027 1916 5043 1923
rect 5027 1913 5040 1916
rect 5076 1867 5083 1923
rect 4996 1787 5003 1853
rect 5156 1847 5163 2133
rect 5196 1956 5203 2033
rect 5236 2007 5243 2213
rect 5276 2147 5283 2223
rect 5336 2107 5343 2413
rect 5396 2287 5403 2443
rect 5456 2407 5463 2474
rect 4956 1776 4983 1783
rect 4796 1696 4813 1703
rect 4876 1687 4883 1703
rect 4876 1676 4893 1687
rect 4880 1673 4893 1676
rect 4916 1647 4923 1733
rect 4956 1667 4963 1776
rect 5016 1736 5023 1833
rect 5216 1787 5223 1923
rect 5296 1867 5303 2033
rect 5356 1987 5363 2273
rect 5416 2256 5423 2313
rect 5396 2220 5403 2223
rect 5393 2207 5407 2220
rect 5436 2107 5443 2223
rect 5220 1763 5233 1767
rect 5216 1753 5233 1763
rect 5216 1748 5223 1753
rect 5256 1736 5263 1833
rect 5016 1643 5023 1673
rect 5036 1667 5043 1703
rect 5236 1700 5243 1703
rect 5056 1643 5063 1673
rect 5016 1636 5063 1643
rect 4776 1227 4783 1553
rect 4796 1447 4803 1473
rect 4836 1436 4843 1613
rect 5196 1567 5203 1692
rect 5233 1687 5247 1700
rect 4807 1403 4820 1407
rect 4807 1393 4823 1403
rect 4816 1383 4823 1393
rect 4816 1376 4883 1383
rect 4807 1353 4813 1367
rect 4856 1323 4863 1353
rect 4876 1343 4883 1376
rect 4896 1347 4903 1403
rect 4876 1336 4893 1343
rect 4916 1323 4923 1353
rect 4856 1316 4923 1323
rect 4936 1307 4943 1434
rect 4956 1407 4963 1493
rect 5016 1487 5023 1553
rect 5236 1547 5243 1633
rect 5016 1436 5023 1473
rect 5073 1387 5087 1392
rect 5096 1367 5103 1433
rect 5116 1407 5123 1533
rect 5147 1434 5153 1447
rect 5236 1436 5243 1473
rect 5316 1467 5323 1973
rect 5413 1960 5427 1973
rect 5476 1968 5483 2476
rect 5596 2387 5603 2573
rect 5616 2343 5623 2653
rect 5596 2336 5623 2343
rect 5596 2287 5603 2336
rect 5636 2323 5643 2736
rect 5676 2727 5683 2774
rect 5676 2488 5683 2692
rect 5716 2647 5723 2743
rect 5696 2387 5703 2443
rect 5627 2316 5643 2323
rect 5616 2263 5623 2313
rect 5596 2256 5623 2263
rect 5496 2067 5503 2253
rect 5536 2087 5543 2212
rect 5576 2187 5583 2223
rect 5496 1983 5503 2053
rect 5536 1987 5543 2073
rect 5496 1976 5523 1983
rect 5416 1956 5423 1960
rect 5456 1956 5473 1963
rect 5336 1747 5343 1793
rect 5373 1740 5387 1753
rect 5376 1736 5383 1740
rect 5356 1700 5363 1703
rect 5353 1687 5367 1700
rect 5456 1487 5463 1956
rect 5516 1956 5523 1976
rect 5553 1960 5567 1973
rect 5556 1956 5563 1960
rect 5616 1947 5623 2113
rect 5636 2027 5643 2273
rect 5656 2127 5663 2373
rect 5676 2267 5683 2333
rect 5736 2287 5743 2713
rect 5756 2707 5763 2743
rect 5816 2727 5823 3173
rect 5836 2847 5843 3413
rect 5856 3407 5863 3473
rect 5876 3303 5883 3593
rect 5896 3527 5903 3973
rect 5936 3607 5943 4073
rect 5956 3707 5963 4033
rect 5996 3987 6003 4293
rect 5996 3767 6003 3873
rect 5916 3516 5923 3553
rect 5996 3527 6003 3753
rect 5956 3327 5963 3453
rect 5976 3427 5983 3483
rect 5856 3296 5883 3303
rect 5856 2987 5863 3296
rect 5976 3303 5983 3413
rect 5956 3296 5983 3303
rect 5876 3256 5903 3263
rect 5876 3227 5883 3256
rect 5896 3207 5903 3233
rect 5933 3000 5947 3013
rect 5976 3007 5983 3252
rect 5996 3107 6003 3473
rect 5936 2996 5943 3000
rect 5856 2907 5863 2952
rect 5856 2823 5863 2893
rect 5836 2816 5863 2823
rect 5756 2363 5763 2573
rect 5836 2507 5843 2816
rect 5896 2727 5903 2743
rect 5896 2703 5903 2713
rect 5896 2696 5923 2703
rect 5856 2488 5863 2513
rect 5776 2387 5783 2474
rect 5896 2427 5903 2673
rect 5756 2356 5783 2363
rect 5700 2283 5713 2287
rect 5696 2273 5713 2283
rect 5696 2256 5703 2273
rect 5733 2260 5747 2273
rect 5776 2267 5783 2356
rect 5736 2256 5743 2260
rect 5580 1923 5593 1927
rect 5536 1867 5543 1923
rect 5576 1916 5593 1923
rect 5580 1913 5593 1916
rect 5387 1473 5393 1487
rect 5333 1467 5347 1473
rect 5147 1433 5160 1434
rect 5133 1387 5147 1393
rect 5216 1400 5223 1403
rect 5213 1387 5227 1400
rect 4676 1180 4683 1183
rect 4673 1167 4687 1180
rect 4716 1027 4723 1183
rect 4436 916 4463 923
rect 4416 887 4423 914
rect 4516 827 4523 883
rect 4556 847 4563 953
rect 4636 943 4643 993
rect 4756 987 4763 1173
rect 4796 1067 4803 1253
rect 4816 1047 4823 1293
rect 4876 1267 4883 1293
rect 4913 1243 4927 1253
rect 4896 1240 4927 1243
rect 4896 1236 4923 1240
rect 4847 1223 4860 1227
rect 4847 1216 4863 1223
rect 4896 1216 4903 1236
rect 4847 1213 4860 1216
rect 4836 1147 4843 1172
rect 4876 1107 4883 1133
rect 4916 1107 4923 1172
rect 4636 936 4653 943
rect 4656 916 4663 933
rect 4576 887 4583 914
rect 4736 883 4743 914
rect 4676 767 4683 883
rect 4716 876 4743 883
rect 4716 787 4723 876
rect 4736 807 4743 833
rect 4456 696 4463 753
rect 4676 723 4683 753
rect 4676 716 4703 723
rect 4436 647 4443 663
rect 4427 636 4443 647
rect 4427 633 4440 636
rect 4496 627 4503 693
rect 4576 607 4583 663
rect 3956 360 3963 363
rect 3916 207 3923 353
rect 3953 347 3967 360
rect 4016 307 4023 396
rect 4036 347 4043 373
rect 4176 367 4183 413
rect 4076 307 4083 363
rect 4196 356 4223 363
rect 4116 327 4123 352
rect 3936 176 3943 293
rect 4196 287 4203 356
rect 4216 216 4223 313
rect 4256 247 4263 363
rect 4276 227 4283 353
rect 4296 267 4303 493
rect 4407 433 4413 447
rect 4356 396 4363 433
rect 4393 400 4407 412
rect 4396 396 4403 400
rect 4316 307 4323 393
rect 4376 327 4383 352
rect 4456 327 4463 394
rect 4476 347 4483 433
rect 4556 396 4563 433
rect 4576 427 4583 593
rect 4576 360 4583 363
rect 4533 347 4547 352
rect 4573 347 4587 360
rect 4616 347 4623 663
rect 4676 647 4683 694
rect 4696 607 4703 716
rect 4716 667 4723 773
rect 4756 747 4763 933
rect 4816 916 4823 973
rect 4936 967 4943 1033
rect 4796 880 4803 883
rect 4793 867 4807 880
rect 4756 723 4763 733
rect 4756 716 4783 723
rect 4776 708 4783 716
rect 4816 696 4823 833
rect 4836 787 4843 883
rect 4936 886 4943 953
rect 4956 928 4963 1273
rect 4976 1147 4983 1293
rect 4996 1227 5003 1313
rect 4996 1027 5003 1173
rect 5036 1163 5043 1183
rect 5076 1180 5083 1183
rect 5073 1167 5087 1180
rect 5116 1167 5123 1253
rect 5136 1187 5143 1333
rect 5176 1216 5183 1313
rect 5196 1180 5203 1183
rect 5193 1167 5207 1180
rect 5036 1156 5053 1163
rect 5056 1047 5063 1153
rect 5016 916 5043 923
rect 4876 847 4883 873
rect 4993 867 5007 872
rect 5016 723 5023 773
rect 5036 747 5043 916
rect 5056 847 5063 1033
rect 5156 916 5163 953
rect 5196 847 5203 1093
rect 5236 1047 5243 1183
rect 5256 1007 5263 1173
rect 5276 1167 5283 1453
rect 5296 1387 5303 1453
rect 5393 1440 5407 1452
rect 5396 1436 5403 1440
rect 5436 1407 5443 1473
rect 5316 1347 5323 1393
rect 5336 1307 5343 1403
rect 5296 1067 5303 1293
rect 5376 1228 5383 1273
rect 5456 1243 5463 1452
rect 5476 1447 5483 1773
rect 5616 1748 5623 1933
rect 5636 1926 5643 2013
rect 5636 1887 5643 1912
rect 5656 1743 5663 2073
rect 5676 1967 5683 2213
rect 5796 2223 5803 2393
rect 5713 2187 5727 2191
rect 5756 2167 5763 2223
rect 5776 2216 5803 2223
rect 5696 1956 5703 2093
rect 5726 1993 5727 2000
rect 5713 1987 5727 1993
rect 5736 1956 5743 1993
rect 5776 1967 5783 2216
rect 5816 2207 5823 2373
rect 5836 2267 5843 2313
rect 5856 2256 5863 2413
rect 5916 2347 5923 2696
rect 5936 2327 5943 2933
rect 5893 2260 5907 2273
rect 5896 2256 5903 2260
rect 5696 1847 5703 1893
rect 5636 1736 5663 1743
rect 5676 1736 5683 1793
rect 5713 1740 5727 1753
rect 5716 1736 5723 1740
rect 5636 1707 5643 1736
rect 5580 1703 5593 1707
rect 5536 1667 5543 1703
rect 5576 1696 5593 1703
rect 5580 1693 5593 1696
rect 5596 1607 5603 1693
rect 5496 1467 5503 1593
rect 5567 1453 5573 1467
rect 5513 1440 5527 1453
rect 5616 1447 5623 1553
rect 5636 1447 5643 1672
rect 5696 1667 5703 1692
rect 5736 1607 5743 1703
rect 5667 1463 5680 1467
rect 5667 1453 5683 1463
rect 5560 1446 5580 1447
rect 5560 1443 5573 1446
rect 5516 1436 5523 1440
rect 5556 1436 5573 1443
rect 5560 1433 5573 1436
rect 5676 1436 5683 1453
rect 5436 1236 5463 1243
rect 5356 1180 5363 1183
rect 5353 1167 5367 1180
rect 5396 1107 5403 1183
rect 5436 1167 5443 1236
rect 5476 1227 5483 1253
rect 5536 1247 5543 1403
rect 5596 1263 5603 1413
rect 5616 1367 5623 1433
rect 5656 1400 5663 1403
rect 5696 1400 5703 1403
rect 5653 1387 5667 1400
rect 5693 1387 5707 1400
rect 5736 1387 5743 1473
rect 5776 1467 5783 1733
rect 5796 1706 5803 2193
rect 5816 1747 5823 2053
rect 5836 1987 5843 2213
rect 5873 2207 5887 2212
rect 5916 2167 5923 2223
rect 5956 2167 5963 2633
rect 5976 2407 5983 2774
rect 5996 2587 6003 3053
rect 5876 1956 5883 1993
rect 5916 1988 5923 2153
rect 5936 2007 5943 2093
rect 5976 2047 5983 2273
rect 5967 1993 5973 2007
rect 5996 1983 6003 2474
rect 5976 1976 6003 1983
rect 5856 1787 5863 1912
rect 5896 1887 5903 1923
rect 5907 1876 5923 1883
rect 5876 1700 5883 1703
rect 5873 1687 5887 1700
rect 5887 1676 5903 1683
rect 5776 1387 5783 1453
rect 5813 1440 5827 1453
rect 5816 1436 5823 1440
rect 5856 1436 5863 1473
rect 5836 1367 5843 1403
rect 5576 1256 5603 1263
rect 5553 1227 5567 1233
rect 5456 1186 5463 1213
rect 5496 1180 5503 1183
rect 5273 947 5287 953
rect 5216 887 5223 933
rect 5296 916 5303 1053
rect 5336 916 5383 923
rect 5276 880 5283 883
rect 5316 880 5323 883
rect 5016 716 5043 723
rect 5036 696 5043 716
rect 4756 607 4763 663
rect 4936 660 4943 663
rect 4796 643 4803 652
rect 4933 647 4947 660
rect 4796 636 4823 643
rect 4716 396 4723 513
rect 4636 367 4643 394
rect 4776 367 4783 573
rect 4676 307 4683 333
rect 4696 327 4703 363
rect 4796 347 4803 413
rect 4816 407 4823 636
rect 4996 587 5003 694
rect 5056 607 5063 663
rect 5096 660 5103 663
rect 5093 647 5107 660
rect 4836 396 4843 513
rect 5056 507 5063 593
rect 4873 400 4887 413
rect 4876 396 4883 400
rect 4936 366 4943 473
rect 5013 400 5027 413
rect 5056 408 5063 433
rect 5016 396 5023 400
rect 5096 367 5103 493
rect 5136 443 5143 833
rect 5196 696 5203 793
rect 5216 727 5223 873
rect 5273 867 5287 880
rect 5313 867 5327 880
rect 5376 863 5383 916
rect 5396 887 5403 993
rect 5456 916 5463 953
rect 5476 947 5483 1173
rect 5493 1167 5507 1180
rect 5376 856 5403 863
rect 5356 747 5363 833
rect 5396 807 5403 856
rect 5233 727 5247 733
rect 5233 720 5253 727
rect 5236 716 5253 720
rect 5240 713 5253 716
rect 5216 660 5223 663
rect 5213 647 5227 660
rect 5256 607 5263 663
rect 5116 436 5143 443
rect 4856 360 4863 363
rect 4853 347 4867 360
rect 5116 347 5123 436
rect 5156 396 5163 493
rect 5296 408 5303 713
rect 5396 696 5403 793
rect 5316 527 5323 693
rect 5420 663 5433 667
rect 5376 427 5383 663
rect 5416 656 5433 663
rect 5420 653 5433 656
rect 5456 507 5463 853
rect 5307 396 5323 403
rect 5353 400 5367 413
rect 5356 396 5363 400
rect 5336 360 5343 363
rect 5333 347 5347 360
rect 4367 296 4393 303
rect 5416 287 5423 413
rect 5476 407 5483 851
rect 5516 847 5523 872
rect 5536 767 5543 993
rect 5556 747 5563 953
rect 5576 928 5583 1256
rect 5596 1007 5603 1233
rect 5656 1216 5663 1253
rect 5716 1227 5723 1253
rect 5756 1216 5783 1223
rect 5616 1007 5623 1173
rect 5636 1127 5643 1183
rect 5696 1107 5703 1173
rect 5716 947 5723 1192
rect 5736 1127 5743 1213
rect 5756 1186 5763 1216
rect 5896 1183 5903 1676
rect 5876 1176 5903 1183
rect 5613 928 5627 933
rect 5653 920 5667 933
rect 5656 916 5663 920
rect 5596 847 5603 883
rect 5636 827 5643 883
rect 5516 696 5523 733
rect 5596 707 5603 793
rect 5576 656 5603 663
rect 5596 507 5603 656
rect 5516 396 5523 453
rect 3756 140 3763 143
rect 3753 127 3767 140
rect 3816 47 3823 174
rect 4156 180 4183 183
rect 4153 176 4183 180
rect 3876 47 3883 143
rect 3956 67 3963 113
rect 3976 107 3983 153
rect 3996 47 4003 173
rect 4153 167 4167 176
rect 4476 146 4483 173
rect 4036 140 4043 143
rect 4076 140 4083 143
rect 4276 140 4303 143
rect 4033 127 4047 140
rect 4073 127 4087 140
rect 4276 136 4307 140
rect 4293 127 4307 136
rect 4416 127 4423 143
rect 4036 67 4043 113
rect 4416 87 4423 113
rect 4496 107 4503 253
rect 4516 187 4523 213
rect 4556 176 4563 233
rect 5336 176 5343 213
rect 5436 183 5443 393
rect 5596 347 5603 493
rect 5616 408 5623 733
rect 5636 666 5643 753
rect 5676 743 5683 873
rect 5696 767 5703 933
rect 5756 916 5763 993
rect 5836 886 5843 1093
rect 5776 827 5783 883
rect 5856 847 5863 1113
rect 5916 947 5923 1876
rect 5936 1687 5943 1773
rect 5936 1127 5943 1533
rect 5956 1107 5963 1972
rect 5756 816 5773 823
rect 5676 736 5703 743
rect 5696 696 5703 736
rect 5756 687 5763 816
rect 5676 467 5683 652
rect 5716 547 5723 663
rect 5776 666 5783 753
rect 5876 707 5883 933
rect 5756 656 5773 663
rect 5676 396 5683 453
rect 5716 427 5723 453
rect 5713 400 5727 413
rect 5736 408 5743 653
rect 5716 396 5723 400
rect 5616 227 5623 394
rect 5656 360 5663 363
rect 5653 347 5667 360
rect 5416 176 5443 183
rect 4716 146 4723 173
rect 4407 56 4433 63
rect 4576 47 4583 143
rect 4616 107 4623 143
rect 4856 107 4863 143
rect 3116 -24 3123 13
rect 3776 -24 3783 13
rect 5196 -17 5203 143
rect 5216 47 5223 173
rect 5316 67 5323 143
rect 5396 87 5403 173
rect 5416 146 5423 176
rect 5456 140 5463 143
rect 5416 107 5423 132
rect 5453 127 5467 140
rect 5496 123 5503 143
rect 5536 127 5543 213
rect 5636 203 5643 293
rect 5616 196 5643 203
rect 5616 176 5623 196
rect 5676 147 5683 273
rect 5756 203 5763 656
rect 5856 547 5863 663
rect 5776 247 5783 533
rect 5876 396 5883 453
rect 5856 247 5863 363
rect 5736 196 5763 203
rect 5736 176 5743 196
rect 5776 176 5783 233
rect 5916 188 5923 833
rect 5476 116 5503 123
rect 5476 107 5483 116
rect 5460 106 5483 107
rect 5467 96 5483 106
rect 5467 93 5480 96
rect 5596 67 5603 143
rect 5636 140 5643 143
rect 5633 127 5647 140
rect 5876 140 5883 143
rect 5873 127 5887 140
rect 5936 67 5943 693
rect 5976 307 5983 1976
rect 5996 1227 6003 1833
rect 5996 127 6003 1093
rect 5176 -24 5203 -17
<< m3contact >>
rect 373 5993 387 6007
rect 413 5993 427 6007
rect 873 5993 887 6007
rect 153 5933 167 5947
rect 273 5894 287 5908
rect 353 5893 367 5907
rect 113 5852 127 5866
rect 173 5853 187 5867
rect 113 5594 127 5608
rect 13 5573 27 5587
rect 13 5533 27 5547
rect 93 5533 107 5547
rect 253 5852 267 5866
rect 293 5653 307 5667
rect 433 5894 447 5908
rect 473 5894 487 5908
rect 1193 5993 1207 6007
rect 1013 5973 1027 5987
rect 1053 5973 1067 5987
rect 653 5852 667 5866
rect 793 5852 807 5866
rect 873 5852 887 5866
rect 913 5852 927 5866
rect 1073 5894 1087 5908
rect 1113 5894 1127 5908
rect 593 5833 607 5847
rect 953 5813 967 5827
rect 793 5673 807 5687
rect 513 5653 527 5667
rect 673 5653 687 5667
rect 193 5593 207 5607
rect 233 5594 247 5608
rect 273 5594 287 5608
rect 353 5594 367 5608
rect 413 5594 427 5608
rect 453 5593 467 5607
rect 553 5594 567 5608
rect 713 5594 727 5608
rect 793 5594 807 5608
rect 853 5594 867 5608
rect 893 5594 907 5608
rect 173 5513 187 5527
rect 133 5413 147 5427
rect 173 5413 187 5427
rect 93 5374 107 5388
rect 253 5453 267 5467
rect 353 5413 367 5427
rect 213 5373 227 5387
rect 253 5374 267 5388
rect 293 5374 307 5388
rect 113 5332 127 5346
rect 93 5074 107 5088
rect 113 4933 127 4947
rect 133 4873 147 4887
rect 193 5332 207 5346
rect 233 5333 247 5347
rect 213 5293 227 5307
rect 273 5313 287 5327
rect 253 5293 267 5307
rect 233 5113 247 5127
rect 273 5113 287 5127
rect 233 5074 247 5088
rect 533 5552 547 5566
rect 453 5533 467 5547
rect 533 5513 547 5527
rect 513 5413 527 5427
rect 393 5374 407 5388
rect 453 5374 467 5388
rect 493 5374 507 5388
rect 693 5552 707 5566
rect 733 5513 747 5527
rect 693 5493 707 5507
rect 613 5453 627 5467
rect 633 5433 647 5447
rect 853 5513 867 5527
rect 793 5473 807 5487
rect 573 5393 587 5407
rect 633 5393 647 5407
rect 553 5373 567 5387
rect 433 5313 447 5327
rect 533 5313 547 5327
rect 513 5253 527 5267
rect 453 5074 467 5088
rect 293 5032 307 5046
rect 353 5032 367 5046
rect 253 4973 267 4987
rect 393 4933 407 4947
rect 173 4873 187 4887
rect 153 4853 167 4867
rect 93 4812 107 4826
rect 153 4813 167 4827
rect 293 4793 307 4807
rect 93 4653 107 4667
rect 153 4653 167 4667
rect 193 4593 207 4607
rect 13 4553 27 4567
rect 93 4554 107 4568
rect 113 4512 127 4526
rect 113 4493 127 4507
rect 173 4513 187 4527
rect 153 4413 167 4427
rect 153 4334 167 4348
rect 13 4293 27 4307
rect 13 4253 27 4267
rect 133 4292 147 4306
rect 253 4554 267 4568
rect 293 4554 307 4568
rect 233 4513 247 4527
rect 193 4253 207 4267
rect 93 4213 107 4227
rect 313 4512 327 4526
rect 393 4812 407 4826
rect 373 4533 387 4547
rect 273 4473 287 4487
rect 253 4373 267 4387
rect 253 4334 267 4348
rect 273 4292 287 4306
rect 473 5032 487 5046
rect 533 5013 547 5027
rect 493 4893 507 4907
rect 833 5433 847 5447
rect 713 5373 727 5387
rect 753 5374 767 5388
rect 793 5374 807 5388
rect 913 5552 927 5566
rect 1473 5933 1487 5947
rect 1293 5852 1307 5866
rect 1353 5852 1367 5866
rect 1413 5833 1427 5847
rect 1353 5813 1367 5827
rect 1213 5793 1227 5807
rect 1293 5793 1307 5807
rect 1193 5693 1207 5707
rect 1253 5673 1267 5687
rect 973 5633 987 5647
rect 1013 5594 1027 5608
rect 1193 5594 1207 5608
rect 973 5553 987 5567
rect 953 5513 967 5527
rect 873 5493 887 5507
rect 973 5473 987 5487
rect 853 5413 867 5427
rect 613 5332 627 5346
rect 653 5332 667 5346
rect 693 5332 707 5346
rect 573 5293 587 5307
rect 593 5074 607 5088
rect 653 5074 667 5088
rect 693 5074 707 5088
rect 873 5374 887 5388
rect 913 5374 927 5388
rect 773 5332 787 5346
rect 813 5332 827 5346
rect 853 5332 867 5346
rect 1193 5533 1207 5547
rect 1073 5513 1087 5527
rect 1153 5473 1167 5487
rect 1033 5433 1047 5447
rect 1133 5433 1147 5447
rect 993 5413 1007 5427
rect 933 5332 947 5346
rect 972 5333 986 5347
rect 1033 5374 1047 5388
rect 1073 5374 1087 5388
rect 993 5332 1007 5346
rect 1053 5332 1067 5346
rect 873 5313 887 5327
rect 1173 5433 1187 5447
rect 1213 5473 1227 5487
rect 1193 5393 1207 5407
rect 1173 5373 1187 5387
rect 1273 5413 1287 5427
rect 1193 5332 1207 5346
rect 1153 5293 1167 5307
rect 1253 5293 1267 5307
rect 1173 5273 1187 5287
rect 893 5233 907 5247
rect 1173 5233 1187 5247
rect 873 5153 887 5167
rect 573 5033 587 5047
rect 733 5074 747 5088
rect 673 5032 687 5046
rect 593 4913 607 4927
rect 633 4913 647 4927
rect 653 4893 667 4907
rect 553 4873 567 4887
rect 593 4873 607 4887
rect 473 4812 487 4826
rect 513 4812 527 4826
rect 413 4773 427 4787
rect 693 4854 707 4868
rect 593 4812 607 4826
rect 633 4812 647 4826
rect 813 5074 827 5088
rect 793 5032 807 5046
rect 833 5013 847 5027
rect 753 4893 767 4907
rect 753 4853 767 4867
rect 873 5032 887 5046
rect 853 4953 867 4967
rect 633 4773 647 4787
rect 733 4773 747 4787
rect 473 4753 487 4767
rect 552 4753 566 4767
rect 573 4753 587 4767
rect 473 4613 487 4627
rect 513 4613 527 4627
rect 433 4593 447 4607
rect 453 4512 467 4526
rect 393 4473 407 4487
rect 373 4413 387 4427
rect 413 4334 427 4348
rect 593 4554 607 4568
rect 573 4512 587 4526
rect 533 4413 547 4427
rect 233 4213 247 4227
rect 13 4093 27 4107
rect 93 4034 107 4048
rect 173 3913 187 3927
rect 133 3853 147 3867
rect 93 3772 107 3786
rect 93 3514 107 3528
rect 133 3472 147 3486
rect 173 3472 187 3486
rect 393 4292 407 4306
rect 433 4292 447 4306
rect 473 4292 487 4306
rect 613 4292 627 4306
rect 493 4093 507 4107
rect 553 4093 567 4107
rect 353 4073 367 4087
rect 393 4073 407 4087
rect 253 4033 267 4047
rect 293 4034 307 4048
rect 253 3913 267 3927
rect 253 3873 267 3887
rect 233 3373 247 3387
rect 13 3333 27 3347
rect 73 3293 87 3307
rect 133 3294 147 3308
rect 173 3294 187 3308
rect 13 3253 27 3267
rect 433 4033 447 4047
rect 493 4034 507 4048
rect 473 3992 487 4006
rect 673 4753 687 4767
rect 653 4553 667 4567
rect 1153 5193 1167 5207
rect 933 5153 947 5167
rect 1113 5113 1127 5127
rect 993 5073 1007 5087
rect 1073 5074 1087 5088
rect 913 4993 927 5007
rect 853 4812 867 4826
rect 893 4812 907 4826
rect 773 4793 787 4807
rect 813 4793 827 4807
rect 753 4653 767 4667
rect 733 4554 747 4568
rect 673 4512 687 4526
rect 713 4512 727 4526
rect 853 4613 867 4627
rect 893 4593 907 4607
rect 853 4554 867 4568
rect 973 4993 987 5007
rect 953 4933 967 4947
rect 993 4973 1007 4987
rect 1013 4854 1027 4868
rect 953 4753 967 4767
rect 973 4693 987 4707
rect 953 4673 967 4687
rect 913 4553 927 4567
rect 773 4493 787 4507
rect 693 4373 707 4387
rect 733 4373 747 4387
rect 673 4292 687 4306
rect 873 4512 887 4526
rect 953 4652 967 4666
rect 1093 5032 1107 5046
rect 1073 4933 1087 4947
rect 1133 4913 1147 4927
rect 1093 4873 1107 4887
rect 1073 4813 1087 4827
rect 1053 4753 1067 4767
rect 993 4593 1007 4607
rect 1053 4554 1067 4568
rect 953 4512 967 4526
rect 993 4512 1007 4526
rect 833 4473 847 4487
rect 933 4473 947 4487
rect 1073 4513 1087 4527
rect 1073 4453 1087 4467
rect 1033 4413 1047 4427
rect 873 4373 887 4387
rect 1013 4373 1027 4387
rect 793 4333 807 4347
rect 833 4334 847 4348
rect 1053 4334 1067 4348
rect 813 4293 827 4307
rect 793 4273 807 4287
rect 893 4292 907 4306
rect 853 4273 867 4287
rect 1033 4292 1047 4306
rect 813 4233 827 4247
rect 773 4173 787 4187
rect 873 4133 887 4147
rect 633 4073 647 4087
rect 853 4073 867 4087
rect 573 4033 587 4047
rect 613 4034 627 4048
rect 653 4034 667 4048
rect 693 4034 707 4048
rect 793 4034 807 4048
rect 573 3992 587 4006
rect 633 3973 647 3987
rect 553 3933 567 3947
rect 633 3933 647 3947
rect 513 3893 527 3907
rect 553 3873 567 3887
rect 433 3833 447 3847
rect 473 3833 487 3847
rect 513 3833 527 3847
rect 353 3772 367 3786
rect 393 3773 407 3787
rect 273 3713 287 3727
rect 493 3713 507 3727
rect 593 3653 607 3667
rect 533 3533 547 3547
rect 293 3514 307 3528
rect 353 3514 367 3528
rect 593 3514 607 3528
rect 413 3472 427 3486
rect 733 4013 747 4027
rect 693 3893 707 3907
rect 773 3973 787 3987
rect 913 4073 927 4087
rect 993 4053 1007 4067
rect 873 4033 887 4047
rect 953 4034 967 4048
rect 793 3953 807 3967
rect 853 3953 867 3967
rect 733 3833 747 3847
rect 673 3772 687 3786
rect 733 3653 747 3667
rect 753 3553 767 3567
rect 933 3992 947 4006
rect 993 3973 1007 3987
rect 933 3933 947 3947
rect 853 3873 867 3887
rect 893 3873 907 3887
rect 813 3833 827 3847
rect 893 3814 907 3828
rect 933 3814 947 3828
rect 1213 5113 1227 5127
rect 1313 5693 1327 5707
rect 1293 5193 1307 5207
rect 1253 5074 1267 5088
rect 1233 4993 1247 5007
rect 1253 4933 1267 4947
rect 1153 4873 1167 4887
rect 1173 4854 1187 4868
rect 1113 4812 1127 4826
rect 1153 4812 1167 4826
rect 1193 4812 1207 4826
rect 1193 4693 1207 4707
rect 1213 4673 1227 4687
rect 1133 4653 1147 4667
rect 1193 4653 1207 4667
rect 1133 4553 1147 4567
rect 1173 4554 1187 4568
rect 1153 4512 1167 4526
rect 1113 4493 1127 4507
rect 1213 4493 1227 4507
rect 1193 4473 1207 4487
rect 1113 4373 1127 4387
rect 1112 4333 1126 4347
rect 1133 4334 1147 4348
rect 1173 4334 1187 4348
rect 1353 5673 1367 5687
rect 1393 5633 1407 5647
rect 1433 5594 1447 5608
rect 1413 5473 1427 5487
rect 1373 5413 1387 5427
rect 1353 5374 1367 5388
rect 1393 5374 1407 5388
rect 1453 5373 1467 5387
rect 1333 5333 1347 5347
rect 1333 5153 1347 5167
rect 1413 5332 1427 5346
rect 1413 5293 1427 5307
rect 2293 5953 2307 5967
rect 1673 5913 1687 5927
rect 1533 5894 1547 5908
rect 1653 5894 1667 5908
rect 1693 5852 1707 5866
rect 1653 5833 1667 5847
rect 1573 5633 1587 5647
rect 1493 5594 1507 5608
rect 1533 5594 1547 5608
rect 1753 5633 1767 5647
rect 1713 5594 1727 5608
rect 1873 5894 1887 5908
rect 1913 5894 1927 5908
rect 2153 5894 2167 5908
rect 2293 5894 2307 5908
rect 2373 5953 2387 5967
rect 1933 5833 1947 5847
rect 1973 5813 1987 5827
rect 1873 5773 1887 5787
rect 1933 5773 1947 5787
rect 1853 5693 1867 5707
rect 1993 5693 2007 5707
rect 1933 5633 1947 5647
rect 1793 5594 1807 5608
rect 1893 5594 1907 5608
rect 1973 5594 1987 5608
rect 1653 5573 1667 5587
rect 1553 5552 1567 5566
rect 1493 5473 1507 5487
rect 1533 5374 1547 5388
rect 1573 5373 1587 5387
rect 1513 5332 1527 5346
rect 1553 5333 1567 5347
rect 1553 5293 1567 5307
rect 1513 5273 1527 5287
rect 1473 5233 1487 5247
rect 1453 5213 1467 5227
rect 1493 5173 1507 5187
rect 1413 5093 1427 5107
rect 1373 5073 1387 5087
rect 1553 5253 1567 5267
rect 1553 5193 1567 5207
rect 1513 5153 1527 5167
rect 1573 5113 1587 5127
rect 1693 5552 1707 5566
rect 1733 5453 1747 5467
rect 1733 5432 1747 5446
rect 1773 5433 1787 5447
rect 1673 5413 1687 5427
rect 1633 5374 1647 5388
rect 1753 5373 1767 5387
rect 1613 5313 1627 5327
rect 1693 5332 1707 5346
rect 1733 5332 1747 5346
rect 1853 5413 1867 5427
rect 1913 5453 1927 5467
rect 1813 5374 1827 5388
rect 2073 5833 2087 5847
rect 2333 5833 2347 5847
rect 2053 5673 2067 5687
rect 2313 5813 2327 5827
rect 2493 5913 2507 5927
rect 2413 5893 2427 5907
rect 2453 5894 2467 5908
rect 2553 5893 2567 5907
rect 2513 5833 2527 5847
rect 2533 5852 2547 5866
rect 2413 5773 2427 5787
rect 2373 5733 2387 5747
rect 2453 5733 2467 5747
rect 2433 5673 2447 5687
rect 2333 5653 2347 5667
rect 2313 5633 2327 5647
rect 2033 5594 2047 5608
rect 2073 5594 2087 5608
rect 2192 5593 2206 5607
rect 2213 5594 2227 5608
rect 2253 5594 2267 5608
rect 1993 5552 2007 5566
rect 1933 5433 1947 5447
rect 1973 5433 1987 5447
rect 2093 5552 2107 5566
rect 2133 5552 2147 5566
rect 2373 5552 2387 5566
rect 2433 5552 2447 5566
rect 2213 5533 2227 5547
rect 2313 5533 2327 5547
rect 2073 5493 2087 5507
rect 2193 5493 2207 5507
rect 2053 5473 2067 5487
rect 1993 5413 2007 5427
rect 2033 5413 2047 5427
rect 1933 5373 1947 5387
rect 1993 5374 2007 5388
rect 1773 5332 1787 5346
rect 1833 5332 1847 5346
rect 1873 5332 1887 5346
rect 1933 5332 1947 5346
rect 2133 5453 2147 5467
rect 2093 5433 2107 5447
rect 3093 5993 3107 6007
rect 2753 5973 2767 5987
rect 2793 5973 2807 5987
rect 2613 5894 2627 5908
rect 2653 5894 2667 5908
rect 2713 5894 2727 5908
rect 2573 5853 2587 5867
rect 2633 5852 2647 5866
rect 2673 5833 2687 5847
rect 2813 5894 2827 5908
rect 2853 5894 2867 5908
rect 2733 5793 2747 5807
rect 2753 5773 2767 5787
rect 2733 5753 2747 5767
rect 2713 5733 2727 5747
rect 2553 5693 2567 5707
rect 2553 5653 2567 5667
rect 2713 5653 2727 5667
rect 2553 5632 2567 5646
rect 2493 5594 2507 5608
rect 3033 5793 3047 5807
rect 2953 5653 2967 5667
rect 2853 5593 2867 5607
rect 2613 5552 2627 5566
rect 2693 5552 2707 5566
rect 2413 5473 2427 5487
rect 2453 5473 2467 5487
rect 2133 5374 2147 5388
rect 2013 5332 2027 5346
rect 2072 5332 2086 5346
rect 2093 5333 2107 5347
rect 2153 5332 2167 5346
rect 1753 5313 1767 5327
rect 1653 5273 1667 5287
rect 1873 5273 1887 5287
rect 1953 5273 1967 5287
rect 1653 5233 1667 5247
rect 1713 5233 1727 5247
rect 1613 5193 1627 5207
rect 1613 5112 1627 5126
rect 1593 5093 1607 5107
rect 1393 5032 1407 5046
rect 1433 5032 1447 5046
rect 1493 5033 1507 5047
rect 1333 4953 1347 4967
rect 1313 4933 1327 4947
rect 1273 4893 1287 4907
rect 1373 4853 1387 4867
rect 1273 4812 1287 4826
rect 1333 4812 1347 4826
rect 1373 4812 1387 4826
rect 1253 4493 1267 4507
rect 1233 4473 1247 4487
rect 1573 5032 1587 5046
rect 1533 4993 1547 5007
rect 1493 4953 1507 4967
rect 1493 4893 1507 4907
rect 1453 4854 1467 4868
rect 1393 4733 1407 4747
rect 1453 4753 1467 4767
rect 1433 4673 1447 4687
rect 1313 4593 1327 4607
rect 1293 4573 1307 4587
rect 1373 4554 1387 4568
rect 1533 4813 1547 4827
rect 1473 4713 1487 4727
rect 1493 4573 1507 4587
rect 1573 4913 1587 4927
rect 1673 5193 1687 5207
rect 1673 5033 1687 5047
rect 1653 4933 1667 4947
rect 1633 4873 1647 4887
rect 2153 5233 2167 5247
rect 1953 5153 1967 5167
rect 2053 5093 2067 5107
rect 1833 5074 1847 5088
rect 1873 5074 1887 5088
rect 1913 5074 1927 5088
rect 1973 5074 1987 5088
rect 2373 5332 2387 5346
rect 2373 5233 2387 5247
rect 2473 5413 2487 5427
rect 2713 5533 2727 5547
rect 2713 5413 2727 5427
rect 2613 5374 2627 5388
rect 2873 5552 2887 5566
rect 2853 5513 2867 5527
rect 2913 5513 2927 5527
rect 2913 5473 2927 5487
rect 2993 5473 3007 5487
rect 2733 5393 2747 5407
rect 2773 5374 2787 5388
rect 2853 5374 2867 5388
rect 2973 5374 2987 5388
rect 3033 5374 3047 5388
rect 2453 5332 2467 5346
rect 2593 5313 2607 5327
rect 2633 5313 2647 5327
rect 2493 5293 2507 5307
rect 2433 5273 2447 5287
rect 2233 5213 2247 5227
rect 2413 5213 2427 5227
rect 2213 5193 2227 5207
rect 2213 5153 2227 5167
rect 2193 5133 2207 5147
rect 2453 5253 2467 5267
rect 2393 5113 2407 5127
rect 2433 5113 2447 5127
rect 2313 5087 2327 5088
rect 1933 5032 1947 5046
rect 1733 5013 1747 5027
rect 1833 5013 1847 5027
rect 1872 5013 1886 5027
rect 1893 5013 1907 5027
rect 1853 4953 1867 4967
rect 1733 4933 1747 4947
rect 1653 4854 1667 4868
rect 1633 4812 1647 4826
rect 1713 4812 1727 4826
rect 1553 4773 1567 4787
rect 1673 4773 1687 4787
rect 1653 4713 1667 4727
rect 1673 4693 1687 4707
rect 1693 4673 1707 4687
rect 1693 4573 1707 4587
rect 1533 4554 1547 4568
rect 1653 4554 1667 4568
rect 1813 4913 1827 4927
rect 1773 4873 1787 4887
rect 1893 4973 1907 4987
rect 1873 4933 1887 4947
rect 1873 4893 1887 4907
rect 1933 4893 1947 4907
rect 1853 4873 1867 4887
rect 1813 4854 1827 4868
rect 1793 4812 1807 4826
rect 1833 4733 1847 4747
rect 1753 4713 1767 4727
rect 1753 4653 1767 4667
rect 1793 4653 1807 4667
rect 1293 4512 1307 4526
rect 1293 4473 1307 4487
rect 1453 4512 1467 4526
rect 1513 4512 1527 4526
rect 1333 4453 1347 4467
rect 1673 4512 1687 4526
rect 1713 4512 1727 4526
rect 2313 5074 2327 5087
rect 2353 5074 2367 5088
rect 2033 5032 2047 5046
rect 2213 5032 2227 5046
rect 2173 5013 2187 5027
rect 2513 5233 2527 5247
rect 2473 5213 2487 5227
rect 2373 5032 2387 5046
rect 2413 5032 2427 5046
rect 2453 5033 2467 5047
rect 2313 4993 2327 5007
rect 2373 4973 2387 4987
rect 2553 5074 2567 5088
rect 2393 4953 2407 4967
rect 2473 4953 2487 4967
rect 2273 4933 2287 4947
rect 2073 4913 2087 4927
rect 2053 4853 2067 4867
rect 1893 4793 1907 4807
rect 1873 4673 1887 4687
rect 1833 4633 1847 4647
rect 1853 4593 1867 4607
rect 2053 4812 2067 4826
rect 1993 4793 2007 4807
rect 1953 4653 1967 4667
rect 2013 4653 2027 4667
rect 1933 4633 1947 4647
rect 1913 4554 1927 4568
rect 1893 4533 1907 4547
rect 1793 4513 1807 4527
rect 1573 4493 1587 4507
rect 1613 4493 1627 4507
rect 1753 4493 1767 4507
rect 1813 4493 1827 4507
rect 1893 4493 1907 4507
rect 1553 4433 1567 4447
rect 1273 4413 1287 4427
rect 1533 4373 1547 4387
rect 1113 4292 1127 4306
rect 1413 4333 1427 4347
rect 1493 4334 1507 4348
rect 1533 4334 1547 4348
rect 1193 4292 1207 4306
rect 1353 4273 1367 4287
rect 1173 4233 1187 4247
rect 1233 4233 1247 4247
rect 1273 4233 1287 4247
rect 1373 4233 1387 4247
rect 1133 4193 1147 4207
rect 1113 4173 1127 4187
rect 1153 4153 1167 4167
rect 1033 4073 1047 4087
rect 1113 4072 1127 4086
rect 1073 4034 1087 4048
rect 1053 3973 1067 3987
rect 1153 3993 1167 4007
rect 1333 4213 1347 4227
rect 1313 4153 1327 4167
rect 1213 4093 1227 4107
rect 1233 4073 1247 4087
rect 1273 4034 1287 4048
rect 1213 3992 1227 4006
rect 1173 3953 1187 3967
rect 1253 3953 1267 3967
rect 1093 3933 1107 3947
rect 1013 3913 1027 3927
rect 1133 3913 1147 3927
rect 1053 3853 1067 3867
rect 873 3772 887 3786
rect 933 3773 947 3787
rect 1013 3772 1027 3786
rect 813 3573 827 3587
rect 893 3573 907 3587
rect 1073 3573 1087 3587
rect 813 3533 827 3547
rect 933 3514 947 3528
rect 973 3514 987 3528
rect 1033 3514 1047 3528
rect 773 3472 787 3486
rect 813 3472 827 3486
rect 913 3472 927 3486
rect 733 3433 747 3447
rect 873 3433 887 3447
rect 593 3373 607 3387
rect 633 3373 647 3387
rect 433 3333 447 3347
rect 533 3333 547 3347
rect 253 3253 267 3267
rect 293 3252 307 3266
rect 13 3213 27 3227
rect 293 3153 307 3167
rect 373 3073 387 3087
rect 293 3053 307 3067
rect 113 2994 127 3008
rect 493 3294 507 3308
rect 1053 3472 1067 3486
rect 1093 3472 1107 3486
rect 1273 3893 1287 3907
rect 1153 3693 1167 3707
rect 1273 3753 1287 3767
rect 1233 3653 1247 3667
rect 1193 3533 1207 3547
rect 1293 3533 1307 3547
rect 933 3353 947 3367
rect 973 3353 987 3367
rect 673 3333 687 3347
rect 613 3293 627 3307
rect 713 3294 727 3308
rect 773 3293 787 3307
rect 813 3294 827 3308
rect 973 3294 987 3308
rect 553 3252 567 3266
rect 593 3252 607 3266
rect 513 3213 527 3227
rect 653 3252 667 3266
rect 613 3113 627 3127
rect 713 3113 727 3127
rect 513 3073 527 3087
rect 613 3073 627 3087
rect 433 3013 447 3027
rect 13 2953 27 2967
rect 153 2952 167 2966
rect 193 2952 207 2966
rect 13 2853 27 2867
rect 273 2833 287 2847
rect 433 2833 447 2847
rect 13 2813 27 2827
rect 73 2773 87 2787
rect 133 2774 147 2788
rect 413 2793 427 2807
rect 453 2774 467 2788
rect 13 2733 27 2747
rect 373 2732 387 2746
rect 233 2713 247 2727
rect 553 3013 567 3027
rect 1033 3273 1047 3287
rect 833 3252 847 3266
rect 953 3252 967 3266
rect 973 3233 987 3247
rect 773 3033 787 3047
rect 833 3033 847 3047
rect 773 2994 787 3008
rect 893 2994 907 3008
rect 933 2994 947 3008
rect 713 2952 727 2966
rect 753 2952 767 2966
rect 833 2952 847 2966
rect 873 2952 887 2966
rect 913 2913 927 2927
rect 693 2793 707 2807
rect 1053 3233 1067 3247
rect 1033 3113 1047 3127
rect 1213 3472 1227 3486
rect 1193 3373 1207 3387
rect 1133 3073 1147 3087
rect 1073 3033 1087 3047
rect 993 2932 1007 2946
rect 973 2913 987 2927
rect 1093 2933 1107 2947
rect 1373 4193 1387 4207
rect 1393 4173 1407 4187
rect 1513 4273 1527 4287
rect 1473 4233 1487 4247
rect 1413 4133 1427 4147
rect 1393 4073 1407 4087
rect 1433 4033 1447 4047
rect 1513 4034 1527 4048
rect 1393 3992 1407 4006
rect 1433 3992 1447 4006
rect 1533 3992 1547 4006
rect 1493 3973 1507 3987
rect 1413 3793 1427 3807
rect 1513 3814 1527 3828
rect 1533 3813 1547 3827
rect 1553 3814 1567 3828
rect 1373 3772 1387 3786
rect 1433 3773 1447 3787
rect 1493 3753 1507 3767
rect 1333 3653 1347 3667
rect 1553 3613 1567 3627
rect 1513 3593 1527 3607
rect 1453 3533 1467 3547
rect 1473 3453 1487 3467
rect 1313 3333 1327 3347
rect 1253 3252 1267 3266
rect 1293 3252 1307 3266
rect 1233 2994 1247 3008
rect 1213 2933 1227 2947
rect 1053 2913 1067 2927
rect 1133 2913 1147 2927
rect 573 2713 587 2727
rect 753 2713 767 2727
rect 813 2713 827 2727
rect 633 2673 647 2687
rect 593 2613 607 2627
rect 713 2533 727 2547
rect 93 2513 107 2527
rect 353 2513 367 2527
rect 513 2513 527 2527
rect 593 2513 607 2527
rect 293 2474 307 2488
rect 533 2474 547 2488
rect 953 2733 967 2747
rect 1313 3233 1327 3247
rect 1353 3353 1367 3367
rect 1333 3133 1347 3147
rect 1433 3294 1447 3308
rect 1493 3294 1507 3308
rect 1493 3253 1507 3267
rect 1393 3233 1407 3247
rect 1453 3153 1467 3167
rect 1393 3073 1407 3087
rect 1353 3033 1367 3047
rect 1413 3033 1427 3047
rect 1393 2952 1407 2966
rect 1333 2893 1347 2907
rect 1333 2853 1347 2867
rect 1393 2774 1407 2788
rect 1493 3073 1507 3087
rect 1793 4473 1807 4487
rect 1653 4334 1667 4348
rect 1713 4333 1727 4347
rect 1873 4453 1887 4467
rect 1833 4334 1847 4348
rect 1673 4173 1687 4187
rect 1613 4073 1627 4087
rect 1593 4034 1607 4048
rect 1653 4034 1667 4048
rect 1773 4292 1787 4306
rect 1873 4293 1887 4307
rect 1873 4272 1887 4286
rect 1813 4233 1827 4247
rect 1753 4193 1767 4207
rect 1733 4073 1747 4087
rect 1593 3973 1607 3987
rect 1673 3933 1687 3947
rect 1633 3913 1647 3927
rect 1693 3913 1707 3927
rect 1633 3873 1647 3887
rect 1693 3814 1707 3828
rect 1613 3772 1627 3786
rect 1633 3753 1647 3767
rect 1613 3693 1627 3707
rect 1573 3533 1587 3547
rect 1653 3733 1667 3747
rect 1573 3472 1587 3486
rect 1633 3472 1647 3486
rect 1653 3433 1667 3447
rect 1573 3294 1587 3308
rect 1633 3293 1647 3307
rect 1553 3252 1567 3266
rect 1533 3233 1547 3247
rect 1593 3233 1607 3247
rect 1633 3213 1647 3227
rect 1853 4113 1867 4127
rect 1873 4033 1887 4047
rect 1753 4013 1767 4027
rect 1793 3992 1807 4006
rect 1873 3973 1887 3987
rect 1833 3953 1847 3967
rect 1773 3814 1787 3828
rect 1813 3814 1827 3828
rect 1793 3772 1807 3786
rect 1833 3772 1847 3786
rect 1733 3753 1747 3767
rect 1973 4554 1987 4568
rect 2133 4873 2147 4887
rect 2173 4854 2187 4868
rect 2233 4853 2247 4867
rect 2313 4913 2327 4927
rect 2373 4854 2387 4868
rect 2113 4812 2127 4826
rect 2233 4812 2247 4826
rect 2293 4812 2307 4826
rect 2173 4793 2187 4807
rect 2333 4793 2347 4807
rect 2373 4793 2387 4807
rect 2153 4713 2167 4727
rect 2113 4593 2127 4607
rect 2073 4553 2087 4567
rect 1913 4413 1927 4427
rect 2033 4493 2047 4507
rect 1993 4433 2007 4447
rect 2573 5013 2587 5027
rect 2613 4973 2627 4987
rect 2533 4933 2547 4947
rect 2533 4912 2547 4926
rect 2453 4854 2467 4868
rect 2493 4854 2507 4868
rect 2213 4773 2227 4787
rect 2473 4773 2487 4787
rect 2233 4693 2247 4707
rect 2213 4673 2227 4687
rect 2213 4554 2227 4568
rect 2153 4493 2167 4507
rect 2173 4473 2187 4487
rect 2213 4473 2227 4487
rect 2113 4373 2127 4387
rect 2093 4353 2107 4367
rect 2153 4353 2167 4367
rect 1973 4273 1987 4287
rect 2073 4253 2087 4267
rect 1933 4073 1947 4087
rect 1913 3993 1927 4007
rect 1893 3873 1907 3887
rect 2033 4053 2047 4067
rect 1993 4034 2007 4048
rect 1973 3992 1987 4006
rect 1953 3953 1967 3967
rect 1933 3933 1947 3947
rect 2013 3933 2027 3947
rect 1973 3873 1987 3887
rect 1953 3833 1967 3847
rect 1913 3813 1927 3827
rect 2033 3813 2047 3827
rect 1873 3753 1887 3767
rect 1833 3733 1847 3747
rect 1993 3772 2007 3786
rect 2033 3753 2047 3767
rect 2113 4273 2127 4287
rect 2373 4713 2387 4727
rect 2353 4633 2367 4647
rect 2313 4573 2327 4587
rect 2273 4554 2287 4568
rect 2293 4334 2307 4348
rect 2393 4593 2407 4607
rect 2493 4573 2507 4587
rect 2453 4554 2467 4568
rect 2393 4513 2407 4527
rect 2433 4512 2447 4526
rect 2473 4512 2487 4526
rect 2413 4453 2427 4467
rect 2373 4433 2387 4447
rect 2373 4353 2387 4367
rect 2173 4253 2187 4267
rect 2213 4253 2227 4267
rect 2153 4193 2167 4207
rect 2173 4173 2187 4187
rect 2133 4073 2147 4087
rect 2213 4053 2227 4067
rect 2173 4034 2187 4048
rect 2113 3993 2127 4007
rect 2093 3873 2107 3887
rect 2153 3992 2167 4006
rect 2133 3973 2147 3987
rect 2193 3973 2207 3987
rect 2233 3973 2247 3987
rect 2293 4292 2307 4306
rect 2333 4213 2347 4227
rect 2293 4113 2307 4127
rect 2353 4073 2367 4087
rect 2293 4034 2307 4048
rect 2313 3992 2327 4006
rect 2273 3973 2287 3987
rect 2253 3953 2267 3967
rect 2293 3953 2307 3967
rect 2133 3893 2147 3907
rect 2253 3853 2267 3867
rect 2313 3833 2327 3847
rect 2333 3793 2347 3807
rect 2093 3772 2107 3786
rect 2233 3772 2247 3786
rect 2433 4292 2447 4306
rect 2413 4273 2427 4287
rect 2513 4553 2527 4567
rect 2513 4512 2527 4526
rect 2553 4853 2567 4867
rect 2653 5293 2667 5307
rect 2713 5233 2727 5247
rect 2653 5113 2667 5127
rect 2673 5074 2687 5088
rect 2733 5153 2747 5167
rect 2773 5293 2787 5307
rect 2853 5293 2867 5307
rect 2853 5272 2867 5286
rect 2793 5253 2807 5267
rect 2953 5333 2967 5347
rect 2893 5253 2907 5267
rect 2853 5173 2867 5187
rect 2773 5153 2787 5167
rect 2753 5133 2767 5147
rect 2733 5113 2747 5127
rect 2793 5074 2807 5088
rect 2893 5074 2907 5088
rect 2693 5032 2707 5046
rect 2653 5013 2667 5027
rect 2633 4913 2647 4927
rect 2693 4933 2707 4947
rect 2713 4913 2727 4927
rect 2773 4993 2787 5007
rect 2833 5032 2847 5046
rect 2873 5032 2887 5046
rect 3093 5373 3107 5387
rect 3293 5993 3307 6007
rect 3333 5993 3347 6007
rect 3973 5993 3987 6007
rect 4013 5993 4027 6007
rect 4053 5993 4067 6007
rect 3193 5973 3207 5987
rect 3233 5973 3247 5987
rect 3153 5833 3167 5847
rect 3213 5793 3227 5807
rect 3153 5773 3167 5787
rect 3173 5653 3187 5667
rect 3153 5613 3167 5627
rect 3133 5333 3147 5347
rect 3093 5233 3107 5247
rect 2993 5193 3007 5207
rect 3113 5193 3127 5207
rect 2973 5133 2987 5147
rect 3033 5113 3047 5127
rect 2993 5074 3007 5088
rect 3013 5032 3027 5046
rect 2953 4993 2967 5007
rect 3013 4993 3027 5007
rect 2793 4973 2807 4987
rect 2773 4953 2787 4967
rect 2733 4854 2747 4868
rect 2793 4913 2807 4927
rect 2873 4873 2887 4887
rect 2953 4873 2967 4887
rect 2813 4854 2827 4868
rect 2553 4812 2567 4826
rect 2593 4812 2607 4826
rect 2893 4853 2907 4867
rect 2933 4854 2947 4868
rect 3033 4913 3047 4927
rect 2973 4853 2987 4867
rect 2633 4773 2647 4787
rect 2733 4593 2747 4607
rect 2673 4554 2687 4568
rect 2553 4512 2567 4526
rect 2733 4512 2747 4526
rect 2673 4453 2687 4467
rect 2593 4433 2607 4447
rect 2533 4373 2547 4387
rect 2833 4812 2847 4826
rect 2873 4812 2887 4826
rect 2893 4773 2907 4787
rect 2793 4713 2807 4727
rect 2993 4812 3007 4826
rect 2893 4693 2907 4707
rect 2953 4693 2967 4707
rect 2773 4554 2787 4568
rect 2873 4512 2887 4526
rect 3213 5613 3227 5627
rect 3173 5552 3187 5566
rect 3853 5913 3867 5927
rect 3353 5894 3367 5908
rect 3393 5894 3407 5908
rect 3813 5894 3827 5908
rect 3573 5852 3587 5866
rect 3633 5852 3647 5866
rect 3453 5613 3467 5627
rect 3393 5594 3407 5608
rect 3273 5552 3287 5566
rect 3693 5833 3707 5847
rect 3573 5613 3587 5627
rect 3793 5613 3807 5627
rect 3593 5594 3607 5608
rect 3653 5594 3667 5608
rect 3753 5594 3767 5608
rect 3833 5594 3847 5608
rect 3493 5513 3507 5527
rect 3273 5493 3287 5507
rect 3573 5493 3587 5507
rect 3153 5153 3167 5167
rect 3253 5153 3267 5167
rect 3193 5113 3207 5127
rect 3153 5074 3167 5088
rect 3113 5032 3127 5046
rect 3173 5032 3187 5046
rect 3193 4993 3207 5007
rect 3093 4913 3107 4927
rect 3133 4913 3147 4927
rect 3053 4873 3067 4887
rect 3133 4854 3147 4868
rect 3113 4812 3127 4826
rect 3073 4773 3087 4787
rect 3053 4753 3067 4767
rect 3033 4633 3047 4647
rect 3013 4593 3027 4607
rect 2913 4554 2927 4568
rect 2973 4554 2987 4568
rect 2833 4473 2847 4487
rect 2893 4473 2907 4487
rect 3113 4753 3127 4767
rect 3153 4693 3167 4707
rect 3433 5473 3447 5487
rect 3333 5374 3347 5388
rect 3373 5374 3387 5388
rect 3413 5374 3427 5388
rect 3493 5453 3507 5467
rect 3713 5513 3727 5527
rect 3653 5433 3667 5447
rect 3613 5413 3627 5427
rect 3493 5393 3507 5407
rect 3593 5393 3607 5407
rect 3473 5374 3487 5388
rect 3513 5374 3527 5388
rect 3573 5374 3587 5388
rect 3433 5332 3447 5346
rect 3493 5332 3507 5346
rect 3413 5313 3427 5327
rect 3333 5293 3347 5307
rect 3313 5113 3327 5127
rect 3533 5273 3547 5287
rect 3373 5133 3387 5147
rect 3513 5133 3527 5147
rect 3333 5093 3347 5107
rect 3473 5093 3487 5107
rect 3273 5033 3287 5047
rect 3313 5032 3327 5046
rect 3593 5332 3607 5346
rect 3633 5332 3647 5346
rect 3253 5013 3267 5027
rect 3353 5013 3367 5027
rect 3493 5013 3507 5027
rect 3253 4973 3267 4987
rect 3213 4933 3227 4947
rect 3233 4853 3247 4867
rect 3333 4933 3347 4947
rect 3373 4933 3387 4947
rect 3293 4873 3307 4887
rect 3353 4913 3367 4927
rect 3333 4853 3347 4867
rect 3213 4812 3227 4826
rect 3273 4812 3287 4826
rect 3313 4812 3327 4826
rect 3353 4812 3367 4826
rect 3433 4913 3447 4927
rect 3473 4873 3487 4887
rect 3413 4812 3427 4826
rect 3253 4753 3267 4767
rect 3373 4753 3387 4767
rect 3193 4633 3207 4647
rect 2993 4512 3007 4526
rect 3073 4512 3087 4526
rect 3153 4493 3167 4507
rect 3193 4493 3207 4507
rect 2913 4453 2927 4467
rect 3473 4653 3487 4667
rect 3373 4633 3387 4647
rect 3413 4633 3427 4647
rect 3273 4553 3287 4567
rect 3313 4554 3327 4568
rect 3513 4993 3527 5007
rect 3533 4893 3547 4907
rect 3633 5293 3647 5307
rect 3673 5293 3687 5307
rect 3773 5493 3787 5507
rect 3733 5473 3747 5487
rect 3833 5433 3847 5447
rect 3733 5413 3747 5427
rect 3713 5132 3727 5146
rect 3693 5074 3707 5088
rect 3613 4993 3627 5007
rect 3673 4993 3687 5007
rect 3673 4953 3687 4967
rect 3593 4933 3607 4947
rect 3653 4933 3667 4947
rect 3613 4893 3627 4907
rect 3653 4893 3667 4907
rect 3553 4854 3567 4868
rect 3593 4854 3607 4868
rect 3493 4613 3507 4627
rect 3413 4593 3427 4607
rect 3273 4493 3287 4507
rect 3433 4493 3447 4507
rect 3573 4812 3587 4826
rect 3613 4813 3627 4827
rect 3533 4693 3547 4707
rect 3613 4653 3627 4667
rect 3613 4593 3627 4607
rect 3553 4554 3567 4568
rect 3953 5894 3967 5908
rect 4093 5913 4107 5927
rect 4133 5913 4147 5927
rect 5233 5993 5247 6007
rect 5113 5973 5127 5987
rect 4733 5933 4747 5947
rect 5073 5933 5087 5947
rect 4133 5894 4147 5908
rect 4253 5894 4267 5908
rect 4373 5894 4387 5908
rect 4433 5894 4447 5908
rect 4473 5894 4487 5908
rect 4093 5833 4107 5847
rect 4053 5753 4067 5767
rect 4553 5893 4567 5907
rect 4613 5894 4627 5908
rect 4793 5894 4807 5908
rect 4873 5894 4887 5908
rect 4193 5733 4207 5747
rect 4293 5733 4307 5747
rect 4173 5673 4187 5687
rect 4113 5633 4127 5647
rect 3913 5613 3927 5627
rect 3953 5594 3967 5608
rect 3793 5393 3807 5407
rect 3853 5393 3867 5407
rect 3833 5374 3847 5388
rect 3813 5313 3827 5327
rect 3873 5333 3887 5347
rect 3773 5293 3787 5307
rect 3853 5293 3867 5307
rect 3833 5273 3847 5287
rect 3813 5074 3827 5088
rect 4033 5594 4047 5608
rect 4073 5594 4087 5608
rect 3993 5513 4007 5527
rect 3933 5493 3947 5507
rect 4133 5552 4147 5566
rect 4173 5552 4187 5566
rect 4093 5513 4107 5527
rect 4173 5513 4187 5527
rect 4033 5453 4047 5467
rect 4173 5453 4187 5467
rect 3953 5433 3967 5447
rect 3913 5393 3927 5407
rect 3893 5193 3907 5207
rect 3793 5032 3807 5046
rect 3833 5032 3847 5046
rect 3773 4993 3787 5007
rect 3753 4953 3767 4967
rect 3753 4913 3767 4927
rect 3733 4893 3747 4907
rect 3793 4953 3807 4967
rect 3773 4853 3787 4867
rect 3693 4812 3707 4826
rect 3653 4753 3667 4767
rect 3753 4753 3767 4767
rect 3633 4573 3647 4587
rect 3673 4554 3687 4568
rect 3993 5393 4007 5407
rect 4053 5393 4067 5407
rect 3973 5332 3987 5346
rect 4013 5293 4027 5307
rect 4093 5374 4107 5388
rect 4133 5374 4147 5388
rect 4093 5293 4107 5307
rect 4053 5213 4067 5227
rect 4033 5113 4047 5127
rect 4093 5113 4107 5127
rect 3973 5093 3987 5107
rect 3953 4993 3967 5007
rect 4253 5633 4267 5647
rect 4333 5633 4347 5647
rect 4293 5594 4307 5608
rect 4233 5552 4247 5566
rect 4333 5553 4347 5567
rect 4293 5433 4307 5447
rect 4213 5413 4227 5427
rect 4273 5413 4287 5427
rect 4193 5313 4207 5327
rect 4253 5374 4267 5388
rect 4273 5332 4287 5346
rect 4313 5332 4327 5346
rect 4213 5273 4227 5287
rect 4133 5093 4147 5107
rect 4373 5833 4387 5847
rect 4453 5813 4467 5827
rect 4413 5773 4427 5787
rect 4453 5673 4467 5687
rect 4593 5833 4607 5847
rect 4753 5852 4767 5866
rect 4713 5833 4727 5847
rect 4932 5893 4946 5907
rect 4953 5893 4967 5907
rect 5013 5894 5027 5908
rect 4853 5852 4867 5866
rect 4793 5813 4807 5827
rect 4893 5813 4907 5827
rect 4773 5693 4787 5707
rect 4553 5653 4567 5667
rect 4733 5653 4747 5667
rect 4453 5633 4467 5647
rect 4433 5613 4447 5627
rect 4533 5613 4547 5627
rect 4413 5594 4427 5608
rect 4573 5594 4587 5608
rect 4612 5594 4626 5608
rect 4633 5594 4647 5608
rect 4693 5594 4707 5608
rect 4393 5513 4407 5527
rect 4373 5473 4387 5487
rect 4513 5493 4527 5507
rect 4553 5473 4567 5487
rect 4593 5453 4607 5467
rect 4433 5433 4447 5447
rect 4393 5373 4407 5387
rect 4473 5374 4487 5388
rect 4673 5552 4687 5566
rect 4753 5553 4767 5567
rect 4953 5852 4967 5866
rect 5033 5852 5047 5866
rect 4993 5753 5007 5767
rect 4933 5693 4947 5707
rect 4853 5653 4867 5667
rect 4893 5653 4907 5667
rect 4893 5594 4907 5608
rect 4973 5633 4987 5647
rect 4953 5613 4967 5627
rect 4833 5552 4847 5566
rect 4873 5552 4887 5566
rect 4933 5552 4947 5566
rect 4753 5473 4767 5487
rect 4633 5453 4647 5467
rect 4893 5453 4907 5467
rect 4613 5433 4627 5447
rect 4713 5433 4727 5447
rect 4833 5433 4847 5447
rect 4813 5413 4827 5427
rect 4753 5374 4767 5388
rect 4373 5332 4387 5346
rect 4413 5332 4427 5346
rect 4493 5333 4507 5347
rect 4833 5374 4847 5388
rect 4533 5313 4547 5327
rect 4573 5313 4587 5327
rect 4493 5293 4507 5307
rect 4233 5074 4247 5088
rect 4033 4913 4047 4927
rect 4193 5032 4207 5046
rect 4253 5032 4267 5046
rect 4293 5032 4307 5046
rect 4113 4993 4127 5007
rect 4373 5074 4387 5088
rect 4433 5074 4447 5088
rect 4513 5074 4527 5088
rect 4233 4973 4247 4987
rect 4333 4973 4347 4987
rect 4093 4913 4107 4927
rect 3913 4873 3927 4887
rect 3953 4873 3967 4887
rect 4073 4873 4087 4887
rect 3813 4853 3827 4867
rect 3853 4854 3867 4868
rect 3873 4812 3887 4826
rect 3873 4773 3887 4787
rect 3913 4713 3927 4727
rect 3913 4613 3927 4627
rect 3813 4573 3827 4587
rect 3873 4573 3887 4587
rect 3433 4472 3447 4486
rect 3513 4473 3527 4487
rect 2753 4433 2767 4447
rect 2933 4433 2947 4447
rect 3253 4433 3267 4447
rect 2733 4373 2747 4387
rect 2833 4373 2847 4387
rect 2573 4353 2587 4367
rect 2673 4353 2687 4367
rect 2533 4334 2547 4348
rect 2773 4334 2787 4348
rect 2753 4292 2767 4306
rect 2593 4253 2607 4267
rect 2713 4253 2727 4267
rect 2553 4233 2567 4247
rect 2493 4193 2507 4207
rect 2413 4133 2427 4147
rect 2453 4073 2467 4087
rect 2273 3753 2287 3767
rect 2353 3753 2367 3767
rect 2133 3733 2147 3747
rect 1933 3713 1947 3727
rect 2053 3713 2067 3727
rect 2153 3713 2167 3727
rect 1733 3613 1747 3627
rect 1913 3553 1927 3567
rect 1733 3514 1747 3528
rect 1793 3513 1807 3527
rect 1853 3514 1867 3528
rect 1693 3473 1707 3487
rect 1673 3293 1687 3307
rect 1793 3472 1807 3486
rect 1833 3472 1847 3486
rect 1713 3433 1727 3447
rect 1913 3433 1927 3447
rect 1793 3353 1807 3367
rect 1873 3353 1887 3367
rect 1653 3153 1667 3167
rect 1573 3133 1587 3147
rect 1533 3093 1547 3107
rect 1453 2994 1467 3008
rect 1473 2952 1487 2966
rect 1453 2893 1467 2907
rect 1513 2893 1527 2907
rect 1013 2732 1027 2746
rect 1253 2732 1267 2746
rect 1293 2732 1307 2746
rect 973 2673 987 2687
rect 1133 2673 1147 2687
rect 873 2613 887 2627
rect 713 2493 727 2507
rect 633 2474 647 2488
rect 133 2432 147 2446
rect 173 2432 187 2446
rect 413 2432 427 2446
rect 733 2432 747 2446
rect 633 2353 647 2367
rect 813 2474 827 2488
rect 873 2474 887 2488
rect 913 2474 927 2488
rect 813 2433 827 2447
rect 793 2333 807 2347
rect 653 2313 667 2327
rect 753 2313 767 2327
rect 153 2273 167 2287
rect 13 2253 27 2267
rect 293 2254 307 2268
rect 333 2254 347 2268
rect 693 2273 707 2287
rect 113 2212 127 2226
rect 13 2173 27 2187
rect 253 2173 267 2187
rect 513 2193 527 2207
rect 573 2193 587 2207
rect 73 2033 87 2047
rect 313 2033 327 2047
rect 193 1954 207 1968
rect 353 1993 367 2007
rect 353 1954 367 1968
rect 473 1954 487 1968
rect 513 1954 527 1968
rect 853 2373 867 2387
rect 813 2273 827 2287
rect 933 2432 947 2446
rect 933 2333 947 2347
rect 753 2133 767 2147
rect 633 1954 647 1968
rect 693 1954 707 1968
rect 733 1954 747 1968
rect 53 1793 67 1807
rect 113 1793 127 1807
rect 153 1813 167 1827
rect 233 1813 247 1827
rect 133 1773 147 1787
rect 193 1773 207 1787
rect 213 1753 227 1767
rect 53 1693 67 1707
rect 173 1692 187 1706
rect 213 1693 227 1707
rect 133 1653 147 1667
rect 193 1434 207 1448
rect 93 1392 107 1406
rect 133 1353 147 1367
rect 113 1313 127 1327
rect 273 1753 287 1767
rect 293 1692 307 1706
rect 232 1434 246 1448
rect 253 1434 267 1448
rect 293 1434 307 1448
rect 393 1912 407 1926
rect 453 1912 467 1926
rect 353 1773 367 1787
rect 393 1773 407 1787
rect 433 1734 447 1748
rect 593 1793 607 1807
rect 653 1933 667 1947
rect 633 1773 647 1787
rect 713 1912 727 1926
rect 713 1793 727 1807
rect 773 1793 787 1807
rect 653 1753 667 1767
rect 593 1734 607 1748
rect 633 1734 647 1748
rect 753 1734 767 1748
rect 873 2193 887 2207
rect 913 2033 927 2047
rect 893 1993 907 2007
rect 813 1913 827 1927
rect 873 1853 887 1867
rect 1373 2653 1387 2667
rect 1073 2553 1087 2567
rect 1313 2513 1327 2527
rect 1373 2513 1387 2527
rect 1073 2493 1087 2507
rect 1133 2493 1147 2507
rect 1033 2474 1047 2488
rect 993 2453 1007 2467
rect 1113 2453 1127 2467
rect 1053 2432 1067 2446
rect 993 2293 1007 2307
rect 1113 2413 1127 2427
rect 1193 2474 1207 2488
rect 1232 2473 1246 2487
rect 1253 2474 1267 2488
rect 1353 2474 1367 2488
rect 1533 2773 1547 2787
rect 1513 2732 1527 2746
rect 1453 2553 1467 2567
rect 1533 2533 1547 2547
rect 1233 2432 1247 2446
rect 1173 2413 1187 2427
rect 1393 2453 1407 2467
rect 1173 2373 1187 2387
rect 1253 2373 1267 2387
rect 1133 2333 1147 2347
rect 1133 2273 1147 2287
rect 933 1833 947 1847
rect 973 2193 987 2207
rect 1013 1993 1027 2007
rect 1013 1954 1027 1968
rect 1213 2293 1227 2307
rect 1293 2432 1307 2446
rect 1293 2333 1307 2347
rect 1233 2212 1247 2226
rect 1193 2013 1207 2027
rect 1193 1992 1207 2006
rect 1153 1954 1167 1968
rect 1093 1933 1107 1947
rect 1273 2212 1287 2226
rect 1273 2133 1287 2147
rect 1013 1873 1027 1887
rect 953 1813 967 1827
rect 653 1713 667 1727
rect 413 1692 427 1706
rect 473 1693 487 1707
rect 453 1673 467 1687
rect 353 1653 367 1667
rect 453 1493 467 1507
rect 573 1692 587 1706
rect 633 1693 647 1707
rect 693 1692 707 1706
rect 733 1692 747 1706
rect 773 1693 787 1707
rect 733 1493 747 1507
rect 593 1434 607 1448
rect 653 1434 667 1448
rect 693 1434 707 1448
rect 313 1373 327 1387
rect 553 1393 567 1407
rect 633 1392 647 1406
rect 593 1373 607 1387
rect 413 1353 427 1367
rect 253 1313 267 1327
rect 313 1273 327 1287
rect 253 1233 267 1247
rect 293 1233 307 1247
rect 133 1172 147 1186
rect 193 1172 207 1186
rect 233 1172 247 1186
rect 513 1353 527 1367
rect 553 1353 567 1367
rect 473 1233 487 1247
rect 373 1214 387 1228
rect 453 1213 467 1227
rect 973 1692 987 1706
rect 913 1673 927 1687
rect 1133 1912 1147 1926
rect 1073 1833 1087 1847
rect 1113 1833 1127 1847
rect 1153 1833 1167 1847
rect 1033 1813 1047 1827
rect 1073 1734 1087 1748
rect 1133 1734 1147 1748
rect 1253 1912 1267 1926
rect 1393 2413 1407 2427
rect 1333 2293 1347 2307
rect 1373 2254 1387 2268
rect 1653 3013 1667 3027
rect 1833 3294 1847 3308
rect 1873 3294 1887 3308
rect 1793 3253 1807 3267
rect 1853 3252 1867 3266
rect 1893 3213 1907 3227
rect 1853 3173 1867 3187
rect 2093 3673 2107 3687
rect 2073 3613 2087 3627
rect 2013 3593 2027 3607
rect 1973 3514 1987 3528
rect 2033 3472 2047 3486
rect 2073 3472 2087 3486
rect 1993 3453 2007 3467
rect 2013 3413 2027 3427
rect 2073 3273 2087 3287
rect 2033 3252 2047 3266
rect 1993 3213 2007 3227
rect 2013 3133 2027 3147
rect 1933 3093 1947 3107
rect 1913 3073 1927 3087
rect 1733 3053 1747 3067
rect 1793 3053 1807 3067
rect 1753 2994 1767 3008
rect 1633 2952 1647 2966
rect 1693 2952 1707 2966
rect 1793 2833 1807 2847
rect 1773 2813 1787 2827
rect 1753 2793 1767 2807
rect 1693 2774 1707 2788
rect 1753 2774 1767 2788
rect 1853 2813 1867 2827
rect 1733 2693 1747 2707
rect 1633 2593 1647 2607
rect 1653 2553 1667 2567
rect 1693 2553 1707 2567
rect 1473 2373 1487 2387
rect 1533 2373 1547 2387
rect 1593 2474 1607 2488
rect 1452 2293 1466 2307
rect 1473 2293 1487 2307
rect 1553 2293 1567 2307
rect 1353 2212 1367 2226
rect 1413 2113 1427 2127
rect 1293 2073 1307 2087
rect 1313 2013 1327 2027
rect 1393 1993 1407 2007
rect 1353 1954 1367 1968
rect 1393 1954 1407 1968
rect 1333 1853 1347 1867
rect 1273 1813 1287 1827
rect 1333 1813 1347 1827
rect 1253 1773 1267 1787
rect 1033 1692 1047 1706
rect 1053 1653 1067 1667
rect 1013 1573 1027 1587
rect 833 1493 847 1507
rect 773 1434 787 1448
rect 873 1434 887 1448
rect 933 1434 947 1448
rect 813 1392 827 1406
rect 1033 1392 1047 1406
rect 873 1353 887 1367
rect 673 1333 687 1347
rect 733 1333 747 1347
rect 1093 1693 1107 1707
rect 1073 1613 1087 1627
rect 1013 1313 1027 1327
rect 1053 1313 1067 1327
rect 693 1273 707 1287
rect 753 1273 767 1287
rect 993 1273 1007 1287
rect 573 1233 587 1247
rect 313 1173 327 1187
rect 593 1213 607 1227
rect 653 1214 667 1228
rect 573 1193 587 1207
rect 393 1172 407 1186
rect 453 1172 467 1186
rect 493 1172 507 1186
rect 713 1172 727 1186
rect 73 913 87 927
rect 393 914 407 928
rect 473 914 487 928
rect 593 914 607 928
rect 133 833 147 847
rect 233 833 247 847
rect 313 833 327 847
rect 153 713 167 727
rect 73 693 87 707
rect 113 694 127 708
rect 173 652 187 666
rect 73 613 87 627
rect 113 394 127 408
rect 333 753 347 767
rect 293 713 307 727
rect 493 872 507 886
rect 573 872 587 886
rect 453 773 467 787
rect 833 1233 847 1247
rect 873 1214 887 1228
rect 953 1214 967 1228
rect 793 1172 807 1186
rect 753 953 767 967
rect 713 914 727 928
rect 853 1133 867 1147
rect 933 1073 947 1087
rect 813 913 827 927
rect 873 914 887 928
rect 653 833 667 847
rect 533 773 547 787
rect 493 733 507 747
rect 373 713 387 727
rect 273 652 287 666
rect 393 692 407 706
rect 453 694 467 708
rect 393 613 407 627
rect 333 573 347 587
rect 373 573 387 587
rect 313 493 327 507
rect 273 453 287 467
rect 233 394 247 408
rect 173 353 187 367
rect 213 353 227 367
rect 133 293 147 307
rect 113 174 127 188
rect 173 174 187 188
rect 133 132 147 146
rect 173 133 187 147
rect 253 352 267 366
rect 273 174 287 188
rect 233 132 247 146
rect 393 493 407 507
rect 333 394 347 408
rect 733 872 747 886
rect 793 873 807 887
rect 833 873 847 887
rect 813 793 827 807
rect 693 753 707 767
rect 713 753 727 767
rect 593 694 607 708
rect 753 694 767 708
rect 613 652 627 666
rect 733 652 747 666
rect 773 652 787 666
rect 813 652 827 666
rect 473 633 487 647
rect 533 633 547 647
rect 412 453 426 467
rect 433 453 447 467
rect 453 413 467 427
rect 433 394 447 408
rect 493 453 507 467
rect 713 453 727 467
rect 333 353 347 367
rect 413 352 427 366
rect 473 353 487 367
rect 553 413 567 427
rect 633 394 647 408
rect 673 394 687 408
rect 713 394 727 408
rect 613 353 627 367
rect 413 293 427 307
rect 633 293 647 307
rect 373 173 387 187
rect 733 352 747 366
rect 1073 1172 1087 1186
rect 953 1033 967 1047
rect 1013 1033 1027 1047
rect 953 953 967 967
rect 933 793 947 807
rect 893 753 907 767
rect 973 913 987 927
rect 1073 914 1087 928
rect 873 733 887 747
rect 953 733 967 747
rect 913 713 927 727
rect 953 712 967 726
rect 893 694 907 708
rect 873 652 887 666
rect 993 733 1007 747
rect 1113 1573 1127 1587
rect 1293 1734 1307 1748
rect 1493 2253 1507 2267
rect 1553 2254 1567 2268
rect 1493 2212 1507 2226
rect 1533 2212 1547 2226
rect 1473 2173 1487 2187
rect 1573 2173 1587 2187
rect 1513 2133 1527 2147
rect 1473 2093 1487 2107
rect 1513 2073 1527 2087
rect 1553 2033 1567 2047
rect 1413 1873 1427 1887
rect 1513 1954 1527 1968
rect 1433 1853 1447 1867
rect 1473 1853 1487 1867
rect 1433 1813 1447 1827
rect 1373 1793 1387 1807
rect 1353 1773 1367 1787
rect 1393 1773 1407 1787
rect 1273 1692 1287 1706
rect 1333 1692 1347 1706
rect 1233 1673 1247 1687
rect 1393 1734 1407 1748
rect 1413 1692 1427 1706
rect 1473 1673 1487 1687
rect 1353 1653 1367 1667
rect 1553 1773 1567 1787
rect 1893 2994 1907 3008
rect 1973 3013 1987 3027
rect 1973 2994 1987 3008
rect 1893 2953 1907 2967
rect 1933 2952 1947 2966
rect 1933 2893 1947 2907
rect 1953 2853 1967 2867
rect 1933 2813 1947 2827
rect 1913 2793 1927 2807
rect 1873 2733 1887 2747
rect 1773 2653 1787 2667
rect 1773 2513 1787 2527
rect 1733 2493 1747 2507
rect 1813 2474 1827 2488
rect 1693 2393 1707 2407
rect 1793 2393 1807 2407
rect 1753 2373 1767 2387
rect 1713 2254 1727 2268
rect 1793 2253 1807 2267
rect 1833 2254 1847 2268
rect 1933 2653 1947 2667
rect 1973 2653 1987 2667
rect 1893 2513 1907 2527
rect 2073 3213 2087 3227
rect 2033 3073 2047 3087
rect 2433 3992 2447 4006
rect 2433 3833 2447 3847
rect 2453 3772 2467 3786
rect 2352 3673 2366 3687
rect 2373 3673 2387 3687
rect 2893 4334 2907 4348
rect 3293 4353 3307 4367
rect 3373 4353 3387 4367
rect 2973 4333 2987 4347
rect 3033 4334 3047 4348
rect 3073 4334 3087 4348
rect 3133 4334 3147 4348
rect 3213 4334 3227 4348
rect 2913 4292 2927 4306
rect 2973 4292 2987 4306
rect 3053 4292 3067 4306
rect 2833 4273 2847 4287
rect 2753 4233 2767 4247
rect 2713 4193 2727 4207
rect 2633 4173 2647 4187
rect 2513 4073 2527 4087
rect 2553 4073 2567 4087
rect 2613 4073 2627 4087
rect 2573 4034 2587 4048
rect 2793 4153 2807 4167
rect 2653 4073 2667 4087
rect 2753 4073 2767 4087
rect 2513 3993 2527 4007
rect 2593 3933 2607 3947
rect 2553 3893 2567 3907
rect 2573 3853 2587 3867
rect 2613 3814 2627 3828
rect 2673 4034 2687 4048
rect 2713 4034 2727 4048
rect 2573 3733 2587 3747
rect 2493 3713 2507 3727
rect 2553 3713 2567 3727
rect 2653 3772 2667 3786
rect 2733 3992 2747 4006
rect 2713 3973 2727 3987
rect 2773 3814 2787 3828
rect 2593 3673 2607 3687
rect 2733 3772 2747 3786
rect 2773 3773 2787 3787
rect 2913 4253 2927 4267
rect 2873 4034 2887 4048
rect 2813 3993 2827 4007
rect 2853 3992 2867 4006
rect 3073 4213 3087 4227
rect 2973 4034 2987 4048
rect 3013 4034 3027 4048
rect 3053 4034 3067 4048
rect 3273 4333 3287 4347
rect 3193 4273 3207 4287
rect 3273 4292 3287 4306
rect 3333 4334 3347 4348
rect 3573 4373 3587 4387
rect 3913 4554 3927 4568
rect 3773 4512 3787 4526
rect 3813 4512 3827 4526
rect 3753 4453 3767 4467
rect 3513 4334 3527 4348
rect 3353 4292 3367 4306
rect 3393 4292 3407 4306
rect 3433 4293 3447 4307
rect 3233 4233 3247 4247
rect 3293 4233 3307 4247
rect 3493 4273 3507 4287
rect 3393 4213 3407 4227
rect 3133 4173 3147 4187
rect 3333 4173 3347 4187
rect 3533 4173 3547 4187
rect 3133 4133 3147 4147
rect 3173 4073 3187 4087
rect 3093 4034 3107 4048
rect 3133 4034 3147 4048
rect 3173 4034 3187 4048
rect 3233 4034 3247 4048
rect 3293 4034 3307 4048
rect 3033 3992 3047 4006
rect 3073 3993 3087 4007
rect 2993 3933 3007 3947
rect 2973 3893 2987 3907
rect 2873 3814 2887 3828
rect 2913 3814 2927 3828
rect 2973 3814 2987 3828
rect 2813 3753 2827 3767
rect 2893 3772 2907 3786
rect 2793 3733 2807 3747
rect 2833 3733 2847 3747
rect 2913 3753 2927 3767
rect 2893 3713 2907 3727
rect 2813 3673 2827 3687
rect 2693 3653 2707 3667
rect 2593 3633 2607 3647
rect 2573 3613 2587 3627
rect 2393 3553 2407 3567
rect 2153 3514 2167 3528
rect 2233 3514 2247 3528
rect 2293 3514 2307 3528
rect 2333 3514 2347 3528
rect 2373 3514 2387 3528
rect 2233 3453 2247 3467
rect 2333 3453 2347 3467
rect 2313 3433 2327 3447
rect 2173 3393 2187 3407
rect 2233 3373 2247 3387
rect 2153 3313 2167 3327
rect 2213 3313 2227 3327
rect 2133 3213 2147 3227
rect 2193 3213 2207 3227
rect 2053 2993 2067 3007
rect 2093 2994 2107 3008
rect 2133 2994 2147 3008
rect 2173 2994 2187 3008
rect 2113 2913 2127 2927
rect 2133 2813 2147 2827
rect 2173 2813 2187 2827
rect 2073 2733 2087 2747
rect 2053 2673 2067 2687
rect 1913 2474 1927 2488
rect 1973 2474 1987 2488
rect 1953 2393 1967 2407
rect 1913 2313 1927 2327
rect 1733 2212 1747 2226
rect 1773 2212 1787 2226
rect 1693 2193 1707 2207
rect 1693 2093 1707 2107
rect 1613 2033 1627 2047
rect 1673 2033 1687 2047
rect 2093 2732 2107 2746
rect 2153 2653 2167 2667
rect 2113 2593 2127 2607
rect 2173 2593 2187 2607
rect 2113 2533 2127 2547
rect 1993 2333 2007 2347
rect 1953 2293 1967 2307
rect 1993 2254 2007 2268
rect 2093 2413 2107 2427
rect 2133 2373 2147 2387
rect 2273 3313 2287 3327
rect 2233 3293 2247 3307
rect 2353 3353 2367 3367
rect 2253 3252 2267 3266
rect 2293 3252 2307 3266
rect 2333 3252 2347 3266
rect 2433 3533 2447 3547
rect 2633 3533 2647 3547
rect 2433 3514 2447 3528
rect 2473 3514 2487 3528
rect 2532 3514 2546 3528
rect 2553 3514 2567 3528
rect 2593 3514 2607 3528
rect 2413 3473 2427 3487
rect 2453 3433 2467 3447
rect 2392 3353 2406 3367
rect 2413 3353 2427 3367
rect 2373 3333 2387 3347
rect 2533 3472 2547 3486
rect 2613 3472 2627 3486
rect 2653 3472 2667 3486
rect 2553 3433 2567 3447
rect 2533 3413 2547 3427
rect 2613 3373 2627 3387
rect 2713 3514 2727 3528
rect 2773 3514 2787 3528
rect 3013 3772 3027 3786
rect 3053 3772 3067 3786
rect 3213 3973 3227 3987
rect 3153 3933 3167 3947
rect 3153 3814 3167 3828
rect 3133 3772 3147 3786
rect 3173 3753 3187 3767
rect 3093 3733 3107 3747
rect 3133 3733 3147 3747
rect 3113 3713 3127 3727
rect 3213 3673 3227 3687
rect 3113 3633 3127 3647
rect 3173 3633 3187 3647
rect 2873 3613 2887 3627
rect 2973 3613 2987 3627
rect 3033 3613 3047 3627
rect 2713 3473 2727 3487
rect 2753 3472 2767 3486
rect 2453 3333 2467 3347
rect 2493 3333 2507 3347
rect 2473 3313 2487 3327
rect 2433 3252 2447 3266
rect 2353 3213 2367 3227
rect 2393 3213 2407 3227
rect 2413 3173 2427 3187
rect 2213 3133 2227 3147
rect 2233 3093 2247 3107
rect 2273 3093 2287 3107
rect 2313 3033 2327 3047
rect 2333 2994 2347 3008
rect 2373 2994 2387 3008
rect 2493 3294 2507 3308
rect 2573 3294 2587 3308
rect 2613 3294 2627 3308
rect 2493 3253 2507 3267
rect 2473 3233 2487 3247
rect 2433 3093 2447 3107
rect 2313 2953 2327 2967
rect 2253 2813 2267 2827
rect 2213 2774 2227 2788
rect 2293 2774 2307 2788
rect 2313 2713 2327 2727
rect 2393 2952 2407 2966
rect 2433 2873 2447 2887
rect 2473 2813 2487 2827
rect 2433 2774 2447 2788
rect 2413 2713 2427 2727
rect 2253 2673 2267 2687
rect 2453 2653 2467 2667
rect 2553 3213 2567 3227
rect 2633 3252 2647 3266
rect 2633 3213 2647 3227
rect 2593 3173 2607 3187
rect 2533 3113 2547 3127
rect 2733 3353 2747 3367
rect 2693 3313 2707 3327
rect 2853 3453 2867 3467
rect 2793 3433 2807 3447
rect 2973 3592 2987 3606
rect 2933 3514 2947 3528
rect 2993 3513 3007 3527
rect 3013 3493 3027 3507
rect 2913 3472 2927 3486
rect 2953 3472 2967 3486
rect 2873 3413 2887 3427
rect 2993 3413 3007 3427
rect 2853 3393 2867 3407
rect 2893 3353 2907 3367
rect 2953 3353 2967 3367
rect 2813 3333 2827 3347
rect 2873 3333 2887 3347
rect 2753 3313 2767 3327
rect 2813 3293 2827 3307
rect 2913 3333 2927 3347
rect 2893 3313 2907 3327
rect 2753 3252 2767 3266
rect 2792 3253 2806 3267
rect 2973 3293 2987 3307
rect 2953 3273 2967 3287
rect 2813 3252 2827 3266
rect 2853 3252 2867 3266
rect 2893 3213 2907 3227
rect 2753 3193 2767 3207
rect 2833 3193 2847 3207
rect 2693 3173 2707 3187
rect 2793 3153 2807 3167
rect 2753 3113 2767 3127
rect 2633 3053 2647 3067
rect 2533 3033 2547 3047
rect 2573 3013 2587 3027
rect 2593 2952 2607 2966
rect 2633 2952 2647 2966
rect 2613 2913 2627 2927
rect 2553 2853 2567 2867
rect 2553 2813 2567 2827
rect 2513 2773 2527 2787
rect 2513 2713 2527 2727
rect 2353 2613 2367 2627
rect 2493 2613 2507 2627
rect 2533 2613 2547 2627
rect 2253 2553 2267 2567
rect 2193 2493 2207 2507
rect 2473 2573 2487 2587
rect 2533 2573 2547 2587
rect 2393 2553 2407 2567
rect 2213 2473 2227 2487
rect 2253 2474 2267 2488
rect 2173 2413 2187 2427
rect 1853 2212 1867 2226
rect 1913 2213 1927 2227
rect 1613 1993 1627 2007
rect 1693 1973 1707 1987
rect 1753 1973 1767 1987
rect 1633 1912 1647 1926
rect 1673 1912 1687 1926
rect 2073 2253 2087 2267
rect 2273 2333 2287 2347
rect 2173 2293 2187 2307
rect 2233 2293 2247 2307
rect 2013 2212 2027 2226
rect 2053 2212 2067 2226
rect 1973 2133 1987 2147
rect 1993 2033 2007 2047
rect 1933 2013 1947 2027
rect 1933 1992 1947 2006
rect 1853 1954 1867 1968
rect 1893 1954 1907 1968
rect 1733 1912 1747 1926
rect 1773 1912 1787 1926
rect 1813 1912 1827 1926
rect 1693 1833 1707 1847
rect 1613 1793 1627 1807
rect 1573 1753 1587 1767
rect 1553 1734 1567 1748
rect 1693 1753 1707 1767
rect 1553 1673 1567 1687
rect 1413 1513 1427 1527
rect 1493 1513 1507 1527
rect 1193 1473 1207 1487
rect 1233 1473 1247 1487
rect 1353 1473 1367 1487
rect 1393 1473 1407 1487
rect 1153 1434 1167 1448
rect 1293 1434 1307 1448
rect 1333 1434 1347 1448
rect 1173 1392 1187 1406
rect 1233 1392 1247 1406
rect 1313 1392 1327 1406
rect 1333 1353 1347 1367
rect 1273 1273 1287 1287
rect 1193 1233 1207 1247
rect 1233 1214 1247 1228
rect 1293 1253 1307 1267
rect 1213 1172 1227 1186
rect 1273 1173 1287 1187
rect 1133 1073 1147 1087
rect 1353 1253 1367 1267
rect 1473 1473 1487 1487
rect 1493 1392 1507 1406
rect 1613 1693 1627 1707
rect 1673 1692 1687 1706
rect 1853 1833 1867 1847
rect 1833 1813 1847 1827
rect 1833 1753 1847 1767
rect 2033 2013 2047 2027
rect 2113 2212 2127 2226
rect 2193 2193 2207 2207
rect 2153 2153 2167 2167
rect 2253 2253 2267 2267
rect 2253 2153 2267 2167
rect 2233 2133 2247 2147
rect 2553 2553 2567 2567
rect 2473 2533 2487 2547
rect 2493 2513 2507 2527
rect 2433 2493 2447 2507
rect 2393 2293 2407 2307
rect 2313 2253 2327 2267
rect 2373 2254 2387 2268
rect 2333 2173 2347 2187
rect 2293 2113 2307 2127
rect 2373 2113 2387 2127
rect 2293 2073 2307 2087
rect 2273 2033 2287 2047
rect 2553 2493 2567 2507
rect 2493 2474 2507 2488
rect 2573 2473 2587 2487
rect 2453 2453 2467 2467
rect 2453 2413 2467 2427
rect 2733 3033 2747 3047
rect 2693 3013 2707 3027
rect 2673 2993 2687 3007
rect 2653 2873 2667 2887
rect 2713 2952 2727 2966
rect 2813 3113 2827 3127
rect 2753 2873 2767 2887
rect 2673 2853 2687 2867
rect 2693 2833 2707 2847
rect 2733 2793 2747 2807
rect 2673 2713 2687 2727
rect 2713 2732 2727 2746
rect 2673 2673 2687 2687
rect 2693 2653 2707 2667
rect 2653 2533 2667 2547
rect 2733 2553 2747 2567
rect 2613 2432 2627 2446
rect 2573 2413 2587 2427
rect 2513 2373 2527 2387
rect 2953 3053 2967 3067
rect 2873 3033 2887 3047
rect 2913 3033 2927 3047
rect 2833 2993 2847 3007
rect 2873 2994 2887 3008
rect 2832 2953 2846 2967
rect 2853 2952 2867 2966
rect 2833 2913 2847 2927
rect 2813 2853 2827 2867
rect 2793 2833 2807 2847
rect 2793 2732 2807 2746
rect 2913 2853 2927 2867
rect 2853 2793 2867 2807
rect 2893 2793 2907 2807
rect 2873 2774 2887 2788
rect 2853 2732 2867 2746
rect 2953 2693 2967 2707
rect 2893 2673 2907 2687
rect 3053 3553 3067 3567
rect 3093 3514 3107 3528
rect 3273 3933 3287 3947
rect 3273 3893 3287 3907
rect 3593 4334 3607 4348
rect 3633 4334 3647 4348
rect 3893 4453 3907 4467
rect 3773 4292 3787 4306
rect 3513 4133 3527 4147
rect 3572 4133 3586 4147
rect 3593 4133 3607 4147
rect 3693 4133 3707 4147
rect 3833 4413 3847 4427
rect 3873 4373 3887 4387
rect 3833 4334 3847 4348
rect 3913 4334 3927 4348
rect 3853 4292 3867 4306
rect 3893 4273 3907 4287
rect 3493 4113 3507 4127
rect 3473 4073 3487 4087
rect 3453 4034 3467 4048
rect 3433 3992 3447 4006
rect 3493 3993 3507 4007
rect 3393 3973 3407 3987
rect 3353 3953 3367 3967
rect 3373 3913 3387 3927
rect 3353 3813 3367 3827
rect 3493 3893 3507 3907
rect 3393 3814 3407 3828
rect 3433 3814 3447 3828
rect 3333 3733 3347 3747
rect 3373 3733 3387 3747
rect 3453 3772 3467 3786
rect 3273 3693 3287 3707
rect 3393 3693 3407 3707
rect 3493 3733 3507 3747
rect 3453 3653 3467 3667
rect 3373 3633 3387 3647
rect 3253 3553 3267 3567
rect 3353 3553 3367 3567
rect 3133 3513 3147 3527
rect 3193 3513 3207 3527
rect 3053 3453 3067 3467
rect 3033 3433 3047 3447
rect 3033 3353 3047 3367
rect 3013 3333 3027 3347
rect 3153 3472 3167 3486
rect 3193 3373 3207 3387
rect 3233 3533 3247 3547
rect 3273 3472 3287 3486
rect 3333 3473 3347 3487
rect 3313 3393 3327 3407
rect 3353 3453 3367 3467
rect 3433 3613 3447 3627
rect 3453 3593 3467 3607
rect 3473 3573 3487 3587
rect 3453 3553 3467 3567
rect 3413 3514 3427 3528
rect 3473 3472 3487 3486
rect 3333 3373 3347 3387
rect 3133 3333 3147 3347
rect 3192 3333 3206 3347
rect 3213 3333 3227 3347
rect 3313 3333 3327 3347
rect 3113 3313 3127 3327
rect 3073 3294 3087 3308
rect 3173 3294 3187 3308
rect 3093 3252 3107 3266
rect 3133 3252 3147 3266
rect 3253 3294 3267 3308
rect 3173 3213 3187 3227
rect 3053 3193 3067 3207
rect 3153 3193 3167 3207
rect 2993 3153 3007 3167
rect 3153 3133 3167 3147
rect 3173 3113 3187 3127
rect 3133 3073 3147 3087
rect 3073 3053 3087 3067
rect 3033 2994 3047 3008
rect 3013 2952 3027 2966
rect 3053 2952 3067 2966
rect 3113 2953 3127 2967
rect 3113 2913 3127 2927
rect 3113 2873 3127 2887
rect 3053 2813 3067 2827
rect 3013 2793 3027 2807
rect 3113 2753 3127 2767
rect 3033 2732 3047 2746
rect 3053 2673 3067 2687
rect 2973 2653 2987 2667
rect 2933 2613 2947 2627
rect 2993 2613 3007 2627
rect 2953 2593 2967 2607
rect 2813 2493 2827 2507
rect 2793 2474 2807 2488
rect 3033 2553 3047 2567
rect 2993 2493 3007 2507
rect 2793 2393 2807 2407
rect 2933 2432 2947 2446
rect 2953 2393 2967 2407
rect 2833 2373 2847 2387
rect 2733 2353 2747 2367
rect 2893 2333 2907 2347
rect 2513 2313 2527 2327
rect 2613 2313 2627 2327
rect 2673 2313 2687 2327
rect 2793 2313 2807 2327
rect 2453 2254 2467 2268
rect 2413 2193 2427 2207
rect 2493 2153 2507 2167
rect 2653 2293 2667 2307
rect 2633 2254 2647 2268
rect 2673 2254 2687 2268
rect 2713 2254 2727 2268
rect 2613 2212 2627 2226
rect 2593 2173 2607 2187
rect 2853 2293 2867 2307
rect 2933 2253 2947 2267
rect 2693 2212 2707 2226
rect 2633 2153 2647 2167
rect 2693 2153 2707 2167
rect 2553 2133 2567 2147
rect 2633 2113 2647 2127
rect 2293 2013 2307 2027
rect 2333 2013 2347 2027
rect 2393 2013 2407 2027
rect 2533 2013 2547 2027
rect 2073 1993 2087 2007
rect 2153 1993 2167 2007
rect 2093 1954 2107 1968
rect 2033 1912 2047 1926
rect 2053 1913 2067 1927
rect 2213 1973 2227 1987
rect 2273 1953 2287 1967
rect 1953 1893 1967 1907
rect 1993 1893 2007 1907
rect 2013 1833 2027 1847
rect 1913 1752 1927 1766
rect 1953 1733 1967 1747
rect 1793 1653 1807 1667
rect 1873 1692 1887 1706
rect 1953 1692 1967 1706
rect 1813 1533 1827 1547
rect 2073 1912 2087 1926
rect 2153 1912 2167 1926
rect 2193 1912 2207 1926
rect 2273 1893 2287 1907
rect 2153 1753 2167 1767
rect 2053 1734 2067 1748
rect 2093 1734 2107 1748
rect 2253 1734 2267 1748
rect 2373 1973 2387 1987
rect 2493 1973 2507 1987
rect 2793 2212 2807 2226
rect 2833 2212 2847 2226
rect 2733 2113 2747 2127
rect 2733 1954 2747 1968
rect 2793 1954 2807 1968
rect 2873 2193 2887 2207
rect 2933 2153 2947 2167
rect 2933 2073 2947 2087
rect 2913 2013 2927 2027
rect 2773 1933 2787 1947
rect 2353 1893 2367 1907
rect 2513 1912 2527 1926
rect 2433 1893 2447 1907
rect 2393 1853 2407 1867
rect 2493 1853 2507 1867
rect 2433 1833 2447 1847
rect 2333 1813 2347 1827
rect 2393 1813 2407 1827
rect 2313 1733 2327 1747
rect 2173 1713 2187 1727
rect 2013 1692 2027 1706
rect 2073 1692 2087 1706
rect 2113 1692 2127 1706
rect 2153 1692 2167 1706
rect 2233 1673 2247 1687
rect 2173 1533 2187 1547
rect 1973 1513 1987 1527
rect 2073 1513 2087 1527
rect 1813 1473 1827 1487
rect 1573 1453 1587 1467
rect 1673 1453 1687 1467
rect 1733 1434 1747 1448
rect 1773 1434 1787 1448
rect 1993 1453 2007 1467
rect 1893 1434 1907 1448
rect 1413 1353 1427 1367
rect 1453 1353 1467 1367
rect 1553 1353 1567 1367
rect 1413 1313 1427 1327
rect 1393 1233 1407 1247
rect 1333 1214 1347 1228
rect 1453 1273 1467 1287
rect 1593 1273 1607 1287
rect 1573 1233 1587 1247
rect 1493 1214 1507 1228
rect 1553 1213 1567 1227
rect 1353 1172 1367 1186
rect 1393 1173 1407 1187
rect 1473 1153 1487 1167
rect 1333 1133 1347 1147
rect 1133 914 1147 928
rect 1173 914 1187 928
rect 1233 914 1247 928
rect 1153 833 1167 847
rect 1093 753 1107 767
rect 1173 753 1187 767
rect 973 652 987 666
rect 1113 652 1127 666
rect 1293 913 1307 927
rect 1513 1113 1527 1127
rect 1653 1353 1667 1367
rect 1993 1434 2007 1448
rect 1833 1392 1847 1406
rect 1893 1393 1907 1407
rect 2373 1653 2387 1667
rect 2333 1593 2347 1607
rect 2213 1473 2227 1487
rect 2133 1453 2147 1467
rect 2173 1434 2187 1448
rect 1793 1353 1807 1367
rect 1733 1313 1747 1327
rect 1613 1233 1627 1247
rect 1733 1233 1747 1247
rect 1793 1233 1807 1247
rect 1653 1214 1667 1228
rect 1713 1213 1727 1227
rect 1573 1172 1587 1186
rect 1633 1172 1647 1186
rect 1553 1093 1567 1107
rect 1693 1033 1707 1047
rect 1653 953 1667 967
rect 1413 913 1427 927
rect 1473 914 1487 928
rect 1553 914 1567 928
rect 1613 914 1627 928
rect 1253 873 1267 887
rect 1253 833 1267 847
rect 1393 873 1407 887
rect 1313 793 1327 807
rect 1233 694 1247 708
rect 1273 652 1287 666
rect 1173 633 1187 647
rect 793 453 807 467
rect 833 453 847 467
rect 1333 753 1347 767
rect 1393 694 1407 708
rect 1333 652 1347 666
rect 1433 653 1447 667
rect 1373 613 1387 627
rect 833 394 847 408
rect 893 394 907 408
rect 973 394 987 408
rect 793 352 807 366
rect 773 333 787 347
rect 853 333 867 347
rect 853 293 867 307
rect 813 253 827 267
rect 693 233 707 247
rect 753 233 767 247
rect 493 173 507 187
rect 693 174 707 188
rect 813 174 827 188
rect 993 352 1007 366
rect 893 253 907 267
rect 913 174 927 188
rect 1113 394 1127 408
rect 1253 393 1267 407
rect 1293 394 1307 408
rect 1053 293 1067 307
rect 1133 293 1147 307
rect 1113 233 1127 247
rect 1073 174 1087 188
rect 1313 352 1327 366
rect 1393 353 1407 367
rect 1833 1213 1847 1227
rect 1773 1172 1787 1186
rect 1733 1113 1747 1127
rect 1773 1053 1787 1067
rect 1713 933 1727 947
rect 1973 1333 1987 1347
rect 1993 1253 2007 1267
rect 1893 1214 1907 1228
rect 1933 1214 1947 1228
rect 1853 1173 1867 1187
rect 1953 1172 1967 1186
rect 1913 1093 1927 1107
rect 2073 1392 2087 1406
rect 2073 1333 2087 1347
rect 2153 1392 2167 1406
rect 2113 1253 2127 1267
rect 2153 1233 2167 1247
rect 2013 1214 2027 1228
rect 2073 1214 2087 1228
rect 2113 1214 2127 1228
rect 2173 1213 2187 1227
rect 2153 1193 2167 1207
rect 2093 1172 2107 1186
rect 2053 1093 2067 1107
rect 1873 1053 1887 1067
rect 1993 1053 2007 1067
rect 1833 993 1847 1007
rect 1853 973 1867 987
rect 1813 953 1827 967
rect 1813 914 1827 928
rect 1853 914 1867 928
rect 1633 872 1647 886
rect 1693 872 1707 886
rect 1593 833 1607 847
rect 1493 813 1507 827
rect 1553 813 1567 827
rect 1693 813 1707 827
rect 1573 753 1587 767
rect 1493 694 1507 708
rect 1533 694 1547 708
rect 1653 694 1667 708
rect 2053 993 2067 1007
rect 2133 993 2147 1007
rect 1913 953 1927 967
rect 1933 933 1947 947
rect 1973 914 1987 928
rect 1873 872 1887 886
rect 1953 872 1967 886
rect 2093 933 2107 947
rect 2133 914 2147 928
rect 2233 1434 2247 1448
rect 2273 1434 2287 1448
rect 2253 1393 2267 1407
rect 2293 1392 2307 1406
rect 2253 1233 2267 1247
rect 2453 1692 2467 1706
rect 2413 1553 2427 1567
rect 2433 1513 2447 1527
rect 2473 1553 2487 1567
rect 2453 1473 2467 1487
rect 2473 1433 2487 1447
rect 2633 1912 2647 1926
rect 2673 1912 2687 1926
rect 2553 1773 2567 1787
rect 2653 1773 2667 1787
rect 2513 1734 2527 1748
rect 2573 1734 2587 1748
rect 2613 1734 2627 1748
rect 2553 1653 2567 1667
rect 2673 1733 2687 1747
rect 2713 1734 2727 1748
rect 2653 1653 2667 1667
rect 2593 1633 2607 1647
rect 2693 1653 2707 1667
rect 2673 1593 2687 1607
rect 2553 1553 2567 1567
rect 2593 1553 2607 1567
rect 2513 1533 2527 1547
rect 2533 1493 2547 1507
rect 2353 1392 2367 1406
rect 2273 1214 2287 1228
rect 2333 1214 2347 1228
rect 2193 1113 2207 1127
rect 2193 953 2207 967
rect 2293 1172 2307 1186
rect 2413 1373 2427 1387
rect 2453 1333 2467 1347
rect 2393 1214 2407 1228
rect 2433 1214 2447 1228
rect 2393 1173 2407 1187
rect 2353 993 2367 1007
rect 2253 973 2267 987
rect 2233 933 2247 947
rect 2293 953 2307 967
rect 2373 933 2387 947
rect 2113 872 2127 886
rect 2053 833 2067 847
rect 1793 793 1807 807
rect 2153 773 2167 787
rect 1933 753 1947 767
rect 1733 694 1747 708
rect 1493 653 1507 667
rect 1613 652 1627 666
rect 1553 613 1567 627
rect 1593 613 1607 627
rect 1453 533 1467 547
rect 1353 313 1367 327
rect 1253 174 1267 188
rect 1313 173 1327 187
rect 1793 693 1807 707
rect 1873 694 1887 708
rect 1713 652 1727 666
rect 1753 652 1767 666
rect 1653 613 1667 627
rect 1753 533 1767 547
rect 1693 394 1707 408
rect 2293 914 2307 928
rect 2273 833 2287 847
rect 2233 793 2247 807
rect 1973 733 1987 747
rect 2033 733 2047 747
rect 2193 733 2207 747
rect 1893 652 1907 666
rect 1933 652 1947 666
rect 1853 613 1867 627
rect 1493 273 1507 287
rect 1613 273 1627 287
rect 1593 213 1607 227
rect 1753 352 1767 366
rect 1833 394 1847 408
rect 1993 694 2007 708
rect 2353 853 2367 867
rect 2253 773 2267 787
rect 2313 773 2327 787
rect 2233 673 2247 687
rect 2093 652 2107 666
rect 1973 613 1987 627
rect 2133 633 2147 647
rect 2193 633 2207 647
rect 2113 533 2127 547
rect 1913 433 1927 447
rect 1973 433 1987 447
rect 2113 433 2127 447
rect 1813 352 1827 366
rect 1873 353 1887 367
rect 1713 333 1727 347
rect 1773 333 1787 347
rect 2313 713 2327 727
rect 2353 713 2367 727
rect 2253 613 2267 627
rect 2273 553 2287 567
rect 2353 553 2367 567
rect 2133 413 2147 427
rect 2193 413 2207 427
rect 2293 493 2307 507
rect 2153 394 2167 408
rect 2053 373 2067 387
rect 1953 352 1967 366
rect 2133 352 2147 366
rect 2513 1392 2527 1406
rect 2593 1513 2607 1527
rect 2553 1433 2567 1447
rect 2673 1434 2687 1448
rect 2573 1392 2587 1406
rect 2533 1333 2547 1347
rect 2833 1912 2847 1926
rect 2913 1813 2927 1827
rect 2793 1733 2807 1747
rect 2853 1734 2867 1748
rect 2913 1734 2927 1748
rect 2773 1673 2787 1687
rect 3073 2653 3087 2667
rect 3153 3033 3167 3047
rect 3153 2993 3167 3007
rect 3293 3113 3307 3127
rect 3213 2993 3227 3007
rect 3273 2993 3287 3007
rect 3193 2952 3207 2966
rect 3233 2952 3247 2966
rect 3193 2873 3207 2887
rect 3333 3294 3347 3308
rect 3373 3413 3387 3427
rect 3353 3173 3367 3187
rect 3333 3113 3347 3127
rect 3333 3073 3347 3087
rect 3413 3313 3427 3327
rect 3433 3294 3447 3308
rect 3473 3293 3487 3307
rect 3453 3252 3467 3266
rect 3393 3173 3407 3187
rect 3373 3053 3387 3067
rect 3333 2994 3347 3008
rect 3433 2993 3447 3007
rect 3613 4093 3627 4107
rect 3593 4072 3607 4086
rect 3673 4073 3687 4087
rect 3793 4113 3807 4127
rect 3733 4093 3747 4107
rect 3613 4052 3627 4066
rect 3573 4033 3587 4047
rect 3652 3993 3666 4007
rect 3693 4053 3707 4067
rect 3593 3973 3607 3987
rect 3553 3953 3567 3967
rect 3553 3833 3567 3847
rect 3533 3813 3547 3827
rect 3593 3814 3607 3828
rect 3533 3772 3547 3786
rect 3613 3772 3627 3786
rect 3673 3992 3687 4006
rect 3713 3992 3727 4006
rect 3793 3973 3807 3987
rect 3753 3933 3767 3947
rect 3893 4113 3907 4127
rect 3933 4113 3947 4127
rect 3833 4073 3847 4087
rect 3853 4053 3867 4067
rect 3893 4053 3907 4067
rect 3913 4034 3927 4048
rect 3833 3992 3847 4006
rect 3893 3933 3907 3947
rect 3813 3913 3827 3927
rect 3673 3873 3687 3887
rect 3793 3873 3807 3887
rect 3653 3733 3667 3747
rect 3553 3713 3567 3727
rect 3613 3693 3627 3707
rect 3653 3613 3667 3627
rect 3633 3593 3647 3607
rect 3592 3573 3606 3587
rect 3613 3573 3627 3587
rect 3633 3553 3647 3567
rect 3593 3514 3607 3528
rect 3553 3453 3567 3467
rect 3613 3453 3627 3467
rect 3573 3433 3587 3447
rect 3533 3333 3547 3347
rect 3633 3333 3647 3347
rect 3613 3313 3627 3327
rect 3513 3293 3527 3307
rect 3573 3294 3587 3308
rect 3713 3833 3727 3847
rect 3693 3813 3707 3827
rect 3753 3833 3767 3847
rect 3693 3773 3707 3787
rect 3853 3853 3867 3867
rect 3833 3833 3847 3847
rect 3853 3813 3867 3827
rect 3973 4854 3987 4868
rect 4033 4854 4047 4868
rect 4113 4873 4127 4887
rect 4013 4812 4027 4826
rect 3973 4773 3987 4787
rect 4053 4713 4067 4727
rect 4133 4854 4147 4868
rect 4173 4854 4187 4868
rect 4133 4813 4147 4827
rect 4133 4613 4147 4627
rect 3973 4553 3987 4567
rect 3973 4512 3987 4526
rect 4033 4512 4047 4526
rect 4053 4373 4067 4387
rect 4113 4554 4127 4568
rect 4193 4812 4207 4826
rect 4253 4953 4267 4967
rect 4313 4953 4327 4967
rect 4413 4993 4427 5007
rect 4393 4953 4407 4967
rect 4233 4613 4247 4627
rect 4293 4933 4307 4947
rect 4273 4913 4287 4927
rect 4273 4853 4287 4867
rect 4333 4893 4347 4907
rect 4413 4933 4427 4947
rect 4393 4853 4407 4867
rect 4313 4812 4327 4826
rect 4353 4812 4367 4826
rect 4393 4812 4407 4826
rect 4773 5332 4787 5346
rect 4812 5332 4826 5346
rect 4833 5333 4847 5347
rect 4873 5332 4887 5346
rect 4733 5313 4747 5327
rect 4613 5273 4627 5287
rect 5293 5894 5307 5908
rect 5353 5893 5367 5907
rect 5393 5893 5407 5907
rect 5453 5894 5467 5908
rect 5533 5894 5547 5908
rect 5573 5894 5587 5908
rect 5613 5894 5627 5908
rect 5653 5894 5667 5908
rect 5753 5894 5767 5908
rect 5793 5894 5807 5908
rect 5173 5852 5187 5866
rect 5233 5853 5247 5867
rect 5273 5852 5287 5866
rect 5173 5813 5187 5827
rect 5233 5813 5247 5827
rect 5133 5753 5147 5767
rect 5113 5613 5127 5627
rect 5033 5594 5047 5608
rect 5073 5594 5087 5608
rect 5113 5592 5127 5606
rect 4973 5553 4987 5567
rect 5013 5552 5027 5566
rect 5033 5533 5047 5547
rect 5013 5493 5027 5507
rect 4993 5453 5007 5467
rect 5053 5453 5067 5467
rect 5093 5453 5107 5467
rect 5033 5433 5047 5447
rect 5053 5413 5067 5427
rect 5013 5393 5027 5407
rect 5033 5374 5047 5388
rect 5013 5332 5027 5346
rect 5053 5332 5067 5346
rect 5093 5332 5107 5346
rect 5193 5653 5207 5667
rect 5353 5852 5367 5866
rect 5313 5813 5327 5827
rect 5273 5673 5287 5687
rect 5233 5594 5247 5608
rect 5133 5552 5147 5566
rect 5213 5552 5227 5566
rect 5213 5513 5227 5527
rect 5173 5493 5187 5507
rect 5173 5413 5187 5427
rect 5173 5374 5187 5388
rect 5353 5653 5367 5667
rect 5433 5852 5447 5866
rect 5433 5713 5447 5727
rect 5533 5813 5547 5827
rect 5653 5833 5667 5847
rect 5593 5813 5607 5827
rect 5573 5673 5587 5687
rect 5473 5653 5487 5667
rect 5393 5593 5407 5607
rect 5293 5533 5307 5547
rect 5373 5513 5387 5527
rect 5393 5493 5407 5507
rect 5333 5453 5347 5467
rect 5373 5453 5387 5467
rect 5113 5313 5127 5327
rect 5153 5273 5167 5287
rect 4693 5253 4707 5267
rect 4953 5253 4967 5267
rect 4613 5193 4627 5207
rect 4573 5074 4587 5088
rect 4613 5074 4627 5088
rect 4553 5033 4567 5047
rect 5133 5213 5147 5227
rect 5133 5113 5147 5127
rect 4753 5074 4767 5088
rect 4833 5073 4847 5087
rect 4893 5074 4907 5088
rect 4933 5074 4947 5088
rect 4993 5073 5007 5087
rect 5073 5074 5087 5088
rect 4573 4993 4587 5007
rect 4553 4973 4567 4987
rect 4533 4933 4547 4947
rect 4493 4913 4507 4927
rect 4453 4893 4467 4907
rect 4513 4893 4527 4907
rect 4553 4893 4567 4907
rect 4493 4873 4507 4887
rect 4473 4854 4487 4868
rect 4413 4753 4427 4767
rect 4293 4713 4307 4727
rect 4253 4573 4267 4587
rect 4213 4554 4227 4568
rect 4533 4813 4547 4827
rect 4593 4953 4607 4967
rect 4673 4993 4687 5007
rect 4593 4893 4607 4907
rect 4633 4893 4647 4907
rect 4633 4854 4647 4868
rect 4693 4953 4707 4967
rect 4693 4873 4707 4887
rect 4553 4793 4567 4807
rect 4533 4773 4547 4787
rect 4473 4753 4487 4767
rect 4373 4653 4387 4667
rect 4453 4653 4467 4667
rect 4413 4613 4427 4627
rect 4453 4573 4467 4587
rect 4453 4533 4467 4547
rect 4173 4413 4187 4427
rect 4033 4292 4047 4306
rect 4093 4293 4107 4307
rect 3993 4273 4007 4287
rect 3993 4173 4007 4187
rect 3973 4033 3987 4047
rect 3953 3813 3967 3827
rect 3773 3772 3787 3786
rect 3813 3772 3827 3786
rect 3873 3772 3887 3786
rect 3953 3773 3967 3787
rect 3733 3733 3747 3747
rect 3773 3733 3787 3747
rect 3813 3733 3827 3747
rect 3693 3693 3707 3707
rect 3693 3514 3707 3528
rect 3913 3613 3927 3627
rect 3853 3573 3867 3587
rect 3773 3513 3787 3527
rect 3813 3514 3827 3528
rect 3913 3553 3927 3567
rect 3893 3533 3907 3547
rect 3793 3493 3807 3507
rect 3673 3473 3687 3487
rect 3693 3453 3707 3467
rect 3673 3433 3687 3447
rect 3673 3373 3687 3387
rect 3513 3272 3527 3286
rect 3493 3253 3507 3267
rect 3553 3252 3567 3266
rect 3573 3233 3587 3247
rect 3353 2952 3367 2966
rect 3293 2873 3307 2887
rect 3393 2873 3407 2887
rect 3533 2993 3547 3007
rect 3633 3233 3647 3247
rect 3633 3193 3647 3207
rect 3593 3033 3607 3047
rect 3873 3472 3887 3486
rect 3713 3433 3727 3447
rect 3813 3433 3827 3447
rect 3733 3373 3747 3387
rect 3733 3294 3747 3308
rect 3773 3294 3787 3308
rect 3793 3252 3807 3266
rect 3833 3252 3847 3266
rect 3913 3252 3927 3266
rect 3693 3233 3707 3247
rect 3753 3233 3767 3247
rect 3773 3213 3787 3227
rect 3833 3193 3847 3207
rect 3673 3173 3687 3187
rect 3713 3173 3727 3187
rect 3813 3173 3827 3187
rect 3673 2994 3687 3008
rect 3233 2813 3247 2827
rect 3273 2813 3287 2827
rect 3213 2732 3227 2746
rect 3273 2732 3287 2746
rect 3153 2693 3167 2707
rect 3353 2774 3367 2788
rect 3333 2732 3347 2746
rect 3373 2732 3387 2746
rect 3413 2713 3427 2727
rect 3373 2693 3387 2707
rect 3413 2613 3427 2627
rect 3413 2573 3427 2587
rect 3293 2553 3307 2567
rect 3133 2533 3147 2547
rect 3393 2533 3407 2547
rect 3153 2474 3167 2488
rect 3373 2453 3387 2467
rect 3053 2432 3067 2446
rect 3133 2432 3147 2446
rect 3033 2393 3047 2407
rect 2973 2353 2987 2367
rect 3093 2353 3107 2367
rect 3013 2293 3027 2307
rect 3053 2254 3067 2268
rect 3033 2212 3047 2226
rect 2993 2193 3007 2207
rect 3053 2093 3067 2107
rect 3033 1993 3047 2007
rect 2973 1954 2987 1968
rect 3073 2033 3087 2047
rect 3013 1893 3027 1907
rect 3053 1893 3067 1907
rect 3153 2333 3167 2347
rect 3313 2413 3327 2427
rect 3293 2393 3307 2407
rect 3253 2333 3267 2347
rect 3233 2313 3247 2327
rect 3153 2273 3167 2287
rect 3113 2253 3127 2267
rect 3193 2254 3207 2268
rect 3133 2213 3147 2227
rect 3113 2173 3127 2187
rect 3213 2212 3227 2226
rect 3173 2133 3187 2147
rect 3273 2254 3287 2268
rect 3333 2273 3347 2287
rect 3573 2952 3587 2966
rect 3613 2952 3627 2966
rect 3653 2952 3667 2966
rect 3693 2933 3707 2947
rect 3673 2873 3687 2887
rect 3493 2633 3507 2647
rect 3593 2713 3607 2727
rect 3593 2653 3607 2667
rect 3573 2633 3587 2647
rect 3513 2593 3527 2607
rect 3553 2593 3567 2607
rect 3513 2493 3527 2507
rect 3453 2474 3467 2488
rect 3493 2473 3507 2487
rect 3413 2413 3427 2427
rect 3453 2353 3467 2367
rect 3393 2333 3407 2347
rect 3433 2273 3447 2287
rect 3273 2212 3287 2226
rect 3313 2212 3327 2226
rect 3293 2192 3307 2206
rect 3353 2193 3367 2207
rect 3313 2153 3327 2167
rect 3293 2133 3307 2147
rect 3353 2133 3367 2147
rect 3273 2053 3287 2067
rect 3253 2033 3267 2047
rect 3093 1973 3107 1987
rect 3133 1972 3147 1986
rect 3093 1952 3107 1966
rect 3233 1993 3247 2007
rect 3213 1953 3227 1967
rect 2973 1813 2987 1827
rect 3073 1813 3087 1827
rect 2953 1753 2967 1767
rect 3033 1773 3047 1787
rect 2993 1753 3007 1767
rect 2813 1692 2827 1706
rect 2933 1692 2947 1706
rect 3073 1734 3087 1748
rect 3153 1893 3167 1907
rect 3173 1833 3187 1847
rect 3153 1793 3167 1807
rect 3113 1773 3127 1787
rect 3013 1692 3027 1706
rect 2833 1653 2847 1667
rect 2993 1653 3007 1667
rect 2753 1553 2767 1567
rect 2733 1533 2747 1547
rect 2813 1613 2827 1627
rect 2933 1513 2947 1527
rect 2773 1473 2787 1487
rect 2893 1473 2907 1487
rect 2773 1434 2787 1448
rect 2853 1433 2867 1447
rect 2793 1392 2807 1406
rect 2833 1393 2847 1407
rect 2693 1353 2707 1367
rect 2753 1353 2767 1367
rect 2753 1332 2767 1346
rect 2673 1293 2687 1307
rect 2613 1253 2627 1267
rect 2753 1253 2767 1267
rect 2773 1233 2787 1247
rect 2593 1214 2607 1228
rect 2633 1214 2647 1228
rect 2672 1213 2686 1227
rect 2693 1214 2707 1228
rect 2733 1214 2747 1228
rect 2473 1133 2487 1147
rect 2413 1113 2427 1127
rect 2473 914 2487 928
rect 2393 873 2407 887
rect 2413 833 2427 847
rect 2493 853 2507 867
rect 2453 713 2467 727
rect 2473 693 2487 707
rect 2393 653 2407 667
rect 2433 652 2447 666
rect 2453 553 2467 567
rect 2373 413 2387 427
rect 2413 413 2427 427
rect 2293 333 2307 347
rect 1993 313 2007 327
rect 2052 313 2066 327
rect 2073 313 2087 327
rect 1913 233 1927 247
rect 2213 233 2227 247
rect 1773 213 1787 227
rect 1673 173 1687 187
rect 1773 173 1787 187
rect 1813 174 1827 188
rect 1873 174 1887 188
rect 2113 174 2127 188
rect 1293 153 1307 167
rect 393 132 407 146
rect 433 132 447 146
rect 472 132 486 146
rect 493 132 507 146
rect 533 132 547 146
rect 333 113 347 127
rect 713 132 727 146
rect 753 132 767 146
rect 833 132 847 146
rect 913 133 927 147
rect 953 132 967 146
rect 1093 132 1107 146
rect 1133 132 1147 146
rect 1233 132 1247 146
rect 1313 132 1327 146
rect 1373 132 1387 146
rect 1653 132 1667 146
rect 673 113 687 127
rect 1753 132 1767 146
rect 1693 113 1707 127
rect 313 93 327 107
rect 573 93 587 107
rect 1933 132 1947 146
rect 1933 113 1947 127
rect 1813 73 1827 87
rect 2013 73 2027 87
rect 2573 1133 2587 1147
rect 2573 914 2587 928
rect 2753 1172 2767 1186
rect 2693 1133 2707 1147
rect 2713 1033 2727 1047
rect 2713 973 2727 987
rect 2593 853 2607 867
rect 2513 833 2527 847
rect 2553 733 2567 747
rect 2513 693 2527 707
rect 2613 713 2627 727
rect 2573 613 2587 627
rect 2513 513 2527 527
rect 2573 513 2587 527
rect 2613 513 2627 527
rect 2493 413 2507 427
rect 2533 394 2547 408
rect 2453 353 2467 367
rect 2513 333 2527 347
rect 2493 313 2507 327
rect 2533 313 2547 327
rect 2493 292 2507 306
rect 2413 233 2427 247
rect 2453 233 2467 247
rect 2373 193 2387 207
rect 2413 193 2427 207
rect 2233 174 2247 188
rect 2453 133 2467 147
rect 2753 914 2767 928
rect 2793 914 2807 928
rect 2913 1392 2927 1406
rect 2873 1353 2887 1367
rect 2853 1333 2867 1347
rect 2913 1273 2927 1287
rect 3033 1573 3047 1587
rect 3073 1553 3087 1567
rect 3053 1433 3067 1447
rect 3133 1753 3147 1767
rect 3193 1813 3207 1827
rect 3253 1973 3267 1987
rect 3313 1954 3327 1968
rect 3393 2093 3407 2107
rect 3553 2393 3567 2407
rect 3593 2593 3607 2607
rect 3653 2773 3667 2787
rect 3753 3153 3767 3167
rect 3733 2994 3747 3008
rect 3773 2994 3787 3008
rect 4153 4292 4167 4306
rect 4193 4292 4207 4306
rect 4113 4093 4127 4107
rect 4173 4193 4187 4207
rect 4033 4053 4047 4067
rect 4073 4053 4087 4067
rect 4133 4053 4147 4067
rect 4053 3992 4067 4006
rect 4093 3992 4107 4006
rect 4033 3853 4047 3867
rect 4073 3814 4087 3828
rect 4213 4133 4227 4147
rect 4293 4513 4307 4527
rect 4353 4512 4367 4526
rect 4533 4633 4547 4647
rect 4573 4593 4587 4607
rect 4813 5013 4827 5027
rect 4773 4993 4787 5007
rect 4733 4953 4747 4967
rect 4773 4854 4787 4868
rect 4993 5032 5007 5046
rect 5053 5032 5067 5046
rect 4833 4993 4847 5007
rect 4873 4993 4887 5007
rect 4833 4913 4847 4927
rect 4833 4873 4847 4887
rect 4753 4813 4767 4827
rect 4653 4793 4667 4807
rect 4653 4633 4667 4647
rect 4613 4573 4627 4587
rect 4793 4812 4807 4826
rect 4833 4812 4847 4826
rect 4873 4812 4887 4826
rect 4793 4673 4807 4687
rect 4753 4593 4767 4607
rect 4713 4573 4727 4587
rect 4393 4453 4407 4467
rect 4373 4393 4387 4407
rect 4253 4373 4267 4387
rect 4313 4334 4327 4348
rect 4393 4333 4407 4347
rect 4433 4334 4447 4348
rect 4253 4292 4267 4306
rect 4333 4292 4347 4306
rect 4373 4293 4387 4307
rect 4333 4233 4347 4247
rect 4313 4213 4327 4227
rect 4293 4173 4307 4187
rect 4293 4093 4307 4107
rect 4153 3993 4167 4007
rect 4233 3992 4247 4006
rect 4293 3853 4307 3867
rect 4153 3814 4167 3828
rect 4213 3814 4227 3828
rect 4013 3773 4027 3787
rect 3993 3753 4007 3767
rect 4093 3772 4107 3786
rect 4153 3773 4167 3787
rect 4233 3733 4247 3747
rect 4193 3693 4207 3707
rect 4273 3633 4287 3647
rect 4013 3593 4027 3607
rect 4193 3593 4207 3607
rect 4113 3573 4127 3587
rect 3993 3514 4007 3528
rect 4033 3514 4047 3528
rect 4093 3514 4107 3528
rect 3973 3453 3987 3467
rect 4093 3453 4107 3467
rect 4013 3433 4027 3447
rect 4093 3333 4107 3347
rect 3993 3293 4007 3307
rect 4053 3294 4067 3308
rect 4153 3514 4167 3528
rect 4213 3472 4227 3486
rect 4173 3413 4187 3427
rect 4153 3353 4167 3367
rect 4213 3353 4227 3367
rect 3973 3233 3987 3247
rect 4073 3233 4087 3247
rect 3993 3213 4007 3227
rect 3993 3053 4007 3067
rect 3793 2952 3807 2966
rect 3733 2913 3747 2927
rect 3813 2913 3827 2927
rect 3713 2793 3727 2807
rect 3793 2793 3807 2807
rect 3673 2732 3687 2746
rect 3713 2732 3727 2746
rect 3773 2732 3787 2746
rect 3653 2713 3667 2727
rect 3733 2713 3747 2727
rect 3773 2693 3787 2707
rect 3773 2653 3787 2667
rect 3633 2573 3647 2587
rect 3733 2553 3747 2567
rect 3593 2533 3607 2547
rect 3713 2474 3727 2488
rect 3573 2353 3587 2367
rect 3513 2273 3527 2287
rect 3533 2254 3547 2268
rect 3513 2212 3527 2226
rect 3553 2173 3567 2187
rect 3453 2133 3467 2147
rect 3493 2113 3507 2127
rect 3493 2073 3507 2087
rect 3513 2053 3527 2067
rect 3393 1954 3407 1968
rect 3273 1913 3287 1927
rect 3253 1893 3267 1907
rect 3253 1813 3267 1827
rect 3233 1753 3247 1767
rect 3173 1734 3187 1748
rect 3213 1734 3227 1748
rect 3333 1912 3347 1926
rect 3393 1913 3407 1927
rect 3313 1893 3327 1907
rect 3293 1833 3307 1847
rect 3293 1793 3307 1807
rect 3273 1752 3287 1766
rect 3153 1693 3167 1707
rect 3233 1692 3247 1706
rect 3193 1673 3207 1687
rect 3153 1593 3167 1607
rect 3273 1692 3287 1706
rect 3253 1573 3267 1587
rect 3133 1533 3147 1547
rect 3113 1473 3127 1487
rect 3193 1473 3207 1487
rect 3253 1473 3267 1487
rect 3173 1413 3187 1427
rect 3033 1392 3047 1406
rect 3093 1392 3107 1406
rect 3173 1353 3187 1367
rect 3133 1253 3147 1267
rect 2993 1233 3007 1247
rect 3113 1233 3127 1247
rect 2973 1213 2987 1227
rect 2893 1172 2907 1186
rect 2933 1172 2947 1186
rect 2973 1172 2987 1186
rect 3053 1214 3067 1228
rect 3333 1772 3347 1786
rect 3373 1753 3387 1767
rect 3333 1734 3347 1748
rect 3433 1993 3447 2007
rect 3473 1993 3487 2007
rect 3473 1954 3487 1968
rect 3553 2033 3567 2047
rect 3653 2393 3667 2407
rect 3613 2273 3627 2287
rect 3713 2273 3727 2287
rect 3673 2254 3687 2268
rect 3753 2493 3767 2507
rect 3753 2432 3767 2446
rect 3732 2253 3746 2267
rect 3753 2253 3767 2267
rect 3693 2212 3707 2226
rect 3753 2212 3767 2226
rect 3653 2173 3667 2187
rect 3593 1973 3607 1987
rect 3433 1912 3447 1926
rect 3533 1912 3547 1926
rect 3593 1893 3607 1907
rect 3493 1873 3507 1887
rect 3573 1873 3587 1887
rect 3673 2153 3687 2167
rect 3673 2113 3687 2127
rect 3713 2173 3727 2187
rect 3693 2093 3707 2107
rect 3713 2033 3727 2047
rect 3673 1993 3687 2007
rect 3633 1973 3647 1987
rect 3653 1954 3667 1968
rect 3733 1993 3747 2007
rect 3853 2833 3867 2847
rect 3813 2673 3827 2687
rect 3793 2573 3807 2587
rect 3953 2993 3967 3007
rect 4033 2993 4047 3007
rect 3933 2913 3947 2927
rect 3913 2873 3927 2887
rect 3893 2793 3907 2807
rect 3953 2793 3967 2807
rect 3873 2732 3887 2746
rect 3893 2673 3907 2687
rect 3833 2553 3847 2567
rect 3873 2474 3887 2488
rect 3933 2533 3947 2547
rect 4393 4073 4407 4087
rect 4513 4512 4527 4526
rect 4553 4453 4567 4467
rect 4513 4413 4527 4427
rect 4613 4413 4627 4427
rect 4573 4373 4587 4387
rect 4613 4334 4627 4348
rect 4653 4334 4667 4348
rect 4513 4273 4527 4287
rect 4553 4273 4567 4287
rect 4493 4213 4507 4227
rect 4593 4153 4607 4167
rect 4373 4034 4387 4048
rect 4413 4034 4427 4048
rect 4453 4033 4467 4047
rect 4453 4012 4467 4026
rect 4353 3992 4367 4006
rect 4453 3953 4467 3967
rect 4393 3893 4407 3907
rect 4393 3853 4407 3867
rect 4313 3813 4327 3827
rect 4353 3814 4367 3828
rect 4333 3753 4347 3767
rect 4333 3653 4347 3667
rect 4513 4034 4527 4048
rect 4553 3933 4567 3947
rect 4533 3893 4547 3907
rect 4533 3853 4547 3867
rect 4493 3814 4507 3828
rect 4493 3773 4507 3787
rect 4573 3772 4587 3786
rect 4473 3753 4487 3767
rect 4373 3593 4387 3607
rect 4533 3693 4547 3707
rect 4573 3693 4587 3707
rect 4313 3553 4327 3567
rect 4413 3553 4427 3567
rect 4293 3514 4307 3528
rect 4413 3532 4427 3546
rect 4453 3533 4467 3547
rect 4353 3514 4367 3528
rect 4313 3433 4327 3447
rect 4273 3313 4287 3327
rect 4253 3294 4267 3308
rect 4153 3252 4167 3266
rect 4193 3252 4207 3266
rect 4233 3153 4247 3167
rect 4253 3113 4267 3127
rect 4133 3053 4147 3067
rect 4233 3053 4247 3067
rect 4173 3013 4187 3027
rect 4133 2994 4147 3008
rect 4073 2953 4087 2967
rect 4033 2933 4047 2947
rect 4033 2912 4047 2926
rect 4073 2774 4087 2788
rect 4153 2952 4167 2966
rect 4193 2952 4207 2966
rect 4093 2732 4107 2746
rect 4053 2713 4067 2727
rect 4053 2573 4067 2587
rect 3973 2513 3987 2527
rect 3913 2493 3927 2507
rect 3953 2493 3967 2507
rect 3813 2432 3827 2446
rect 3873 2433 3887 2447
rect 4013 2474 4027 2488
rect 3913 2373 3927 2387
rect 3993 2432 4007 2446
rect 3953 2393 3967 2407
rect 4153 2774 4167 2788
rect 4233 2853 4247 2867
rect 4493 3514 4507 3528
rect 4473 3472 4487 3486
rect 4413 3393 4427 3407
rect 4473 3333 4487 3347
rect 4373 3313 4387 3327
rect 4453 3293 4467 3307
rect 4433 3273 4447 3287
rect 4333 3193 4347 3207
rect 4433 3213 4447 3227
rect 4393 3173 4407 3187
rect 4693 4512 4707 4526
rect 4773 4513 4787 4527
rect 4753 4473 4767 4487
rect 4733 4453 4747 4467
rect 4693 4393 4707 4407
rect 4813 4633 4827 4647
rect 4913 5013 4927 5027
rect 4913 4973 4927 4987
rect 5093 4993 5107 5007
rect 5073 4973 5087 4987
rect 5053 4913 5067 4927
rect 4993 4854 5007 4868
rect 5053 4854 5067 4868
rect 4913 4812 4927 4826
rect 4893 4593 4907 4607
rect 4833 4553 4847 4567
rect 4913 4554 4927 4568
rect 4973 4812 4987 4826
rect 5053 4813 5067 4827
rect 5013 4713 5027 4727
rect 5133 4993 5147 5007
rect 5193 5074 5207 5088
rect 5213 5013 5227 5027
rect 5153 4973 5167 4987
rect 5333 5374 5347 5388
rect 5373 5374 5387 5388
rect 5273 5333 5287 5347
rect 5553 5594 5567 5608
rect 5533 5552 5547 5566
rect 5533 5533 5547 5547
rect 5493 5493 5507 5507
rect 5453 5453 5467 5467
rect 5433 5413 5447 5427
rect 5313 5332 5327 5346
rect 5353 5332 5367 5346
rect 5393 5332 5407 5346
rect 5273 5293 5287 5307
rect 5433 5373 5447 5387
rect 5573 5393 5587 5407
rect 5513 5374 5527 5388
rect 5553 5374 5567 5388
rect 5453 5332 5467 5346
rect 5473 5293 5487 5307
rect 5573 5233 5587 5247
rect 5473 5173 5487 5187
rect 5373 5113 5387 5127
rect 5413 5113 5427 5127
rect 5333 5074 5347 5088
rect 5413 5074 5427 5088
rect 5313 5013 5327 5027
rect 5153 4913 5167 4927
rect 5113 4893 5127 4907
rect 5193 4854 5207 4868
rect 5093 4733 5107 4747
rect 5073 4673 5087 4687
rect 5193 4733 5207 4747
rect 5193 4653 5207 4667
rect 5173 4633 5187 4647
rect 4953 4593 4967 4607
rect 4893 4512 4907 4526
rect 4793 4493 4807 4507
rect 4853 4493 4867 4507
rect 4713 4292 4727 4306
rect 4813 4233 4827 4247
rect 4653 4153 4667 4167
rect 4793 4133 4807 4147
rect 4713 4073 4727 4087
rect 4753 4034 4767 4048
rect 4653 3993 4667 4007
rect 4693 3992 4707 4006
rect 4713 3953 4727 3967
rect 4653 3813 4667 3827
rect 4793 3993 4807 4007
rect 4733 3933 4747 3947
rect 4753 3814 4767 3828
rect 4793 3813 4807 3827
rect 4573 3653 4587 3667
rect 4633 3653 4647 3667
rect 4733 3772 4747 3786
rect 4693 3753 4707 3767
rect 4673 3653 4687 3667
rect 4653 3573 4667 3587
rect 4653 3533 4667 3547
rect 4593 3514 4607 3528
rect 4573 3413 4587 3427
rect 4513 3294 4527 3308
rect 4473 3273 4487 3287
rect 4953 4393 4967 4407
rect 5053 4554 5067 4568
rect 5093 4554 5107 4568
rect 5133 4553 5147 4567
rect 5173 4553 5187 4567
rect 5253 4893 5267 4907
rect 5233 4613 5247 4627
rect 5353 4873 5367 4887
rect 5293 4854 5307 4868
rect 5273 4813 5287 4827
rect 5253 4573 5267 4587
rect 5353 4812 5367 4826
rect 5313 4753 5327 4767
rect 5413 4913 5427 4927
rect 5513 5113 5527 5127
rect 5692 5653 5706 5667
rect 5713 5653 5727 5667
rect 5653 5594 5667 5608
rect 5693 5594 5707 5608
rect 5753 5833 5767 5847
rect 5673 5552 5687 5566
rect 5693 5393 5707 5407
rect 5733 5553 5747 5567
rect 5813 5833 5827 5847
rect 5753 5513 5767 5527
rect 5813 5713 5827 5727
rect 5853 5653 5867 5667
rect 5853 5594 5867 5608
rect 5953 5594 5967 5608
rect 5793 5453 5807 5467
rect 5873 5453 5887 5467
rect 5793 5413 5807 5427
rect 5833 5413 5847 5427
rect 5753 5373 5767 5387
rect 5833 5374 5847 5388
rect 5893 5413 5907 5427
rect 5873 5373 5887 5387
rect 5673 5332 5687 5346
rect 5713 5333 5727 5347
rect 5633 5313 5647 5327
rect 5733 5313 5747 5327
rect 5613 5153 5627 5167
rect 5653 5093 5667 5107
rect 5553 5033 5567 5047
rect 5593 5033 5607 5047
rect 5533 4993 5547 5007
rect 5493 4913 5507 4927
rect 5453 4873 5467 4887
rect 5433 4853 5447 4867
rect 5412 4812 5426 4826
rect 5433 4793 5447 4807
rect 5473 4812 5487 4826
rect 5673 5032 5687 5046
rect 5633 4993 5647 5007
rect 5593 4913 5607 4927
rect 5573 4854 5587 4868
rect 5653 4854 5667 4868
rect 5713 4854 5727 4868
rect 5553 4773 5567 4787
rect 5473 4753 5487 4767
rect 5413 4713 5427 4727
rect 5373 4653 5387 4667
rect 5313 4613 5327 4627
rect 5293 4573 5307 4587
rect 5273 4553 5287 4567
rect 5073 4512 5087 4526
rect 5113 4513 5127 4527
rect 5033 4473 5047 4487
rect 5093 4393 5107 4407
rect 4993 4373 5007 4387
rect 4933 4292 4947 4306
rect 4853 4233 4867 4247
rect 5153 4512 5167 4526
rect 5213 4512 5227 4526
rect 5253 4512 5267 4526
rect 5233 4453 5247 4467
rect 5133 4353 5147 4367
rect 5173 4334 5187 4348
rect 5253 4333 5267 4347
rect 5453 4573 5467 4587
rect 5413 4554 5427 4568
rect 5393 4512 5407 4526
rect 5353 4453 5367 4467
rect 5333 4413 5347 4427
rect 5313 4353 5327 4367
rect 5393 4353 5407 4367
rect 5233 4313 5247 4327
rect 5153 4292 5167 4306
rect 5093 4273 5107 4287
rect 5193 4273 5207 4287
rect 4833 4173 4847 4187
rect 5053 4173 5067 4187
rect 4913 4073 4927 4087
rect 4973 4073 4987 4087
rect 5053 4073 5067 4087
rect 5193 4073 5207 4087
rect 4873 4034 4887 4048
rect 4953 4034 4967 4048
rect 4853 3992 4867 4006
rect 4953 3993 4967 4007
rect 4893 3933 4907 3947
rect 4873 3853 4887 3867
rect 4933 3853 4947 3867
rect 5093 4034 5107 4048
rect 5133 4034 5147 4048
rect 5313 4292 5327 4306
rect 5313 4193 5327 4207
rect 5393 4133 5407 4147
rect 5453 4493 5467 4507
rect 5433 4333 5447 4347
rect 5553 4633 5567 4647
rect 5513 4573 5527 4587
rect 5633 4812 5647 4826
rect 5653 4793 5667 4807
rect 5593 4554 5607 4568
rect 5633 4554 5647 4568
rect 5573 4512 5587 4526
rect 5553 4453 5567 4467
rect 5473 4413 5487 4427
rect 5493 4334 5507 4348
rect 5473 4252 5487 4266
rect 5353 4113 5367 4127
rect 5413 4113 5427 4127
rect 5273 4073 5287 4087
rect 5233 4034 5247 4048
rect 5293 4034 5307 4048
rect 5033 3992 5047 4006
rect 5073 3992 5087 4006
rect 5173 3992 5187 4006
rect 5073 3893 5087 3907
rect 5133 3893 5147 3907
rect 5013 3814 5027 3828
rect 4853 3772 4867 3786
rect 4933 3772 4947 3786
rect 5033 3772 5047 3786
rect 4993 3733 5007 3747
rect 5053 3713 5067 3727
rect 5153 3853 5167 3867
rect 5213 3953 5227 3967
rect 5253 3953 5267 3967
rect 5233 3913 5247 3927
rect 5293 3913 5307 3927
rect 5093 3813 5107 3827
rect 5133 3814 5147 3828
rect 5173 3814 5187 3828
rect 5153 3753 5167 3767
rect 5093 3733 5107 3747
rect 5213 3773 5227 3787
rect 5213 3733 5227 3747
rect 5193 3713 5207 3727
rect 4813 3693 4827 3707
rect 4893 3673 4907 3687
rect 4793 3633 4807 3647
rect 4773 3553 4787 3567
rect 4693 3533 4707 3547
rect 4673 3433 4687 3447
rect 4633 3393 4647 3407
rect 4813 3514 4827 3528
rect 4853 3514 4867 3528
rect 4753 3472 4767 3486
rect 4753 3433 4767 3447
rect 4693 3373 4707 3387
rect 4733 3373 4747 3387
rect 4693 3333 4707 3347
rect 4613 3313 4627 3327
rect 4653 3313 4667 3327
rect 4493 3173 4507 3187
rect 4453 3113 4467 3127
rect 4313 3053 4327 3067
rect 4292 3013 4306 3027
rect 4313 3013 4327 3027
rect 4413 3013 4427 3027
rect 4453 3013 4467 3027
rect 4473 3013 4487 3027
rect 4393 2994 4407 3008
rect 4293 2933 4307 2947
rect 4513 2994 4527 3008
rect 4553 2993 4567 3007
rect 4413 2973 4427 2987
rect 4393 2933 4407 2947
rect 4333 2913 4347 2927
rect 4353 2853 4367 2867
rect 4313 2833 4327 2847
rect 4253 2793 4267 2807
rect 4293 2793 4307 2807
rect 4233 2774 4247 2788
rect 4213 2732 4227 2746
rect 4253 2732 4267 2746
rect 4153 2653 4167 2667
rect 4253 2713 4267 2727
rect 4253 2673 4267 2687
rect 4233 2653 4247 2667
rect 4213 2613 4227 2627
rect 4213 2553 4227 2567
rect 4153 2513 4167 2527
rect 4073 2473 4087 2487
rect 4113 2474 4127 2488
rect 4193 2493 4207 2507
rect 4053 2333 4067 2347
rect 3953 2313 3967 2327
rect 3913 2273 3927 2287
rect 3853 2254 3867 2268
rect 3893 2254 3907 2268
rect 3933 2253 3947 2267
rect 3813 2033 3827 2047
rect 3673 1912 3687 1926
rect 3713 1913 3727 1927
rect 3653 1873 3667 1887
rect 3613 1833 3627 1847
rect 3553 1773 3567 1787
rect 3533 1753 3547 1767
rect 3393 1653 3407 1667
rect 3353 1633 3367 1647
rect 3273 1453 3287 1467
rect 3293 1434 3307 1448
rect 3333 1434 3347 1448
rect 3233 1392 3247 1406
rect 3253 1373 3267 1387
rect 3193 1333 3207 1347
rect 3213 1293 3227 1307
rect 3213 1233 3227 1247
rect 3233 1213 3247 1227
rect 3193 1172 3207 1186
rect 3453 1734 3467 1748
rect 3593 1733 3607 1747
rect 3653 1734 3667 1748
rect 3553 1713 3567 1727
rect 3513 1673 3527 1687
rect 3553 1673 3567 1687
rect 3473 1653 3487 1667
rect 3453 1593 3467 1607
rect 3393 1473 3407 1487
rect 3433 1473 3447 1487
rect 3373 1453 3387 1467
rect 3353 1393 3367 1407
rect 3333 1373 3347 1387
rect 3273 1333 3287 1347
rect 3313 1333 3327 1347
rect 3453 1434 3467 1448
rect 3513 1533 3527 1547
rect 3533 1473 3547 1487
rect 3573 1473 3587 1487
rect 3413 1392 3427 1406
rect 3473 1392 3487 1406
rect 3513 1392 3527 1406
rect 3673 1692 3687 1706
rect 3693 1653 3707 1667
rect 3633 1633 3647 1647
rect 3693 1573 3707 1587
rect 3673 1533 3687 1547
rect 3613 1473 3627 1487
rect 3573 1434 3587 1448
rect 3593 1392 3607 1406
rect 3633 1392 3647 1406
rect 3373 1293 3387 1307
rect 3533 1293 3547 1307
rect 3413 1253 3427 1267
rect 3553 1253 3567 1267
rect 3353 1233 3367 1247
rect 3393 1233 3407 1247
rect 3253 1173 3267 1187
rect 3293 1172 3307 1186
rect 3373 1173 3387 1187
rect 3073 1133 3087 1147
rect 3233 993 3247 1007
rect 3193 953 3207 967
rect 2893 914 2907 928
rect 2953 914 2967 928
rect 2993 914 3007 928
rect 3033 914 3047 928
rect 3073 914 3087 928
rect 2733 872 2747 886
rect 2813 872 2827 886
rect 2813 833 2827 847
rect 2793 813 2807 827
rect 2693 793 2707 807
rect 2673 773 2687 787
rect 2873 773 2887 787
rect 2993 853 3007 867
rect 2713 753 2727 767
rect 2953 753 2967 767
rect 2833 733 2847 747
rect 2933 733 2947 747
rect 2753 694 2767 708
rect 2813 694 2827 708
rect 2693 653 2707 667
rect 2673 633 2687 647
rect 2773 652 2787 666
rect 2753 633 2767 647
rect 2733 553 2747 567
rect 2593 453 2607 467
rect 2653 453 2667 467
rect 2693 453 2707 467
rect 2573 273 2587 287
rect 2533 174 2547 188
rect 2573 113 2587 127
rect 2613 413 2627 427
rect 2613 353 2627 367
rect 2593 73 2607 87
rect 2733 352 2747 366
rect 2673 273 2687 287
rect 2633 174 2647 188
rect 2713 193 2727 207
rect 2633 133 2647 147
rect 2673 132 2687 146
rect 2893 694 2907 708
rect 2973 693 2987 707
rect 2833 652 2847 666
rect 2873 633 2887 647
rect 2913 593 2927 607
rect 2833 553 2847 567
rect 2933 473 2947 487
rect 2873 394 2887 408
rect 3113 913 3127 927
rect 3153 914 3167 928
rect 3393 1093 3407 1107
rect 3373 973 3387 987
rect 3273 953 3287 967
rect 3093 893 3107 907
rect 3293 914 3307 928
rect 3373 914 3387 928
rect 3213 872 3227 886
rect 3273 872 3287 886
rect 3293 853 3307 867
rect 3013 833 3027 847
rect 3173 833 3187 847
rect 3093 793 3107 807
rect 3253 793 3267 807
rect 3053 694 3067 708
rect 3313 773 3327 787
rect 3353 773 3367 787
rect 3153 753 3167 767
rect 3253 753 3267 767
rect 3133 693 3147 707
rect 3033 633 3047 647
rect 2993 533 3007 547
rect 3073 533 3087 547
rect 2893 352 2907 366
rect 2933 352 2947 366
rect 3013 352 3027 366
rect 2853 313 2867 327
rect 2773 233 2787 247
rect 3013 213 3027 227
rect 2873 193 2887 207
rect 2953 193 2967 207
rect 2833 132 2847 146
rect 2953 132 2967 146
rect 2993 132 3007 146
rect 3033 132 3047 146
rect 2753 113 2767 127
rect 2893 113 2907 127
rect 3033 113 3047 127
rect 3133 613 3147 627
rect 3113 593 3127 607
rect 3093 473 3107 487
rect 3133 553 3147 567
rect 3233 733 3247 747
rect 3193 694 3207 708
rect 3233 694 3247 708
rect 3493 1233 3507 1247
rect 3453 1214 3467 1228
rect 3873 2113 3887 2127
rect 4013 2254 4027 2268
rect 3993 2212 4007 2226
rect 4033 2212 4047 2226
rect 3953 2173 3967 2187
rect 3893 2033 3907 2047
rect 3933 2033 3947 2047
rect 3813 1912 3827 1926
rect 3813 1873 3827 1887
rect 3813 1852 3827 1866
rect 3773 1833 3787 1847
rect 3873 1893 3887 1907
rect 3853 1793 3867 1807
rect 3853 1733 3867 1747
rect 3733 1692 3747 1706
rect 3733 1593 3747 1607
rect 3713 1473 3727 1487
rect 3693 1433 3707 1447
rect 3673 1233 3687 1247
rect 3593 1214 3607 1228
rect 3633 1214 3647 1228
rect 3513 1172 3527 1186
rect 3553 1172 3567 1186
rect 3473 1133 3487 1147
rect 3473 993 3487 1007
rect 3513 993 3527 1007
rect 3513 953 3527 967
rect 3453 913 3467 927
rect 3653 1033 3667 1047
rect 3953 1954 3967 1968
rect 4093 2353 4107 2367
rect 4093 2212 4107 2226
rect 4013 2053 4027 2067
rect 3993 1953 4007 1967
rect 3913 1912 3927 1926
rect 3973 1912 3987 1926
rect 4033 1953 4047 1967
rect 4013 1853 4027 1867
rect 3993 1773 4007 1787
rect 3933 1753 3947 1767
rect 3893 1733 3907 1747
rect 4073 2133 4087 2147
rect 4133 2393 4147 2407
rect 4273 2553 4287 2567
rect 4233 2473 4247 2487
rect 4293 2493 4307 2507
rect 4253 2432 4267 2446
rect 4213 2393 4227 2407
rect 4193 2353 4207 2367
rect 4233 2333 4247 2347
rect 4173 2254 4187 2268
rect 4353 2774 4367 2788
rect 4453 2933 4467 2947
rect 4493 2913 4507 2927
rect 4533 2813 4547 2827
rect 4493 2774 4507 2788
rect 4373 2732 4387 2746
rect 4413 2733 4427 2747
rect 4373 2673 4387 2687
rect 4333 2613 4347 2627
rect 4473 2713 4487 2727
rect 4553 2733 4567 2747
rect 4553 2613 4567 2627
rect 4413 2573 4427 2587
rect 4493 2573 4507 2587
rect 4553 2573 4567 2587
rect 4413 2552 4427 2566
rect 4473 2493 4487 2507
rect 4333 2432 4347 2446
rect 4393 2432 4407 2446
rect 4253 2254 4267 2268
rect 4153 2173 4167 2187
rect 4133 2113 4147 2127
rect 4113 2053 4127 2067
rect 4253 2213 4267 2227
rect 4233 2053 4247 2067
rect 4213 1953 4227 1967
rect 4313 2273 4327 2287
rect 4393 2273 4407 2287
rect 4353 2212 4367 2226
rect 4393 2212 4407 2226
rect 4293 2193 4307 2207
rect 4333 2193 4347 2207
rect 4293 2153 4307 2167
rect 4293 2113 4307 2127
rect 4253 1993 4267 2007
rect 4293 1954 4307 1968
rect 4113 1912 4127 1926
rect 4153 1912 4167 1926
rect 4233 1913 4247 1927
rect 4273 1912 4287 1926
rect 4213 1893 4227 1907
rect 4233 1833 4247 1847
rect 3993 1713 4007 1727
rect 3873 1692 3887 1706
rect 3913 1692 3927 1706
rect 3913 1653 3927 1667
rect 3953 1653 3967 1667
rect 3853 1533 3867 1547
rect 3793 1453 3807 1467
rect 3893 1453 3907 1467
rect 3753 1434 3767 1448
rect 3733 1393 3747 1407
rect 3793 1392 3807 1406
rect 3833 1392 3847 1406
rect 4093 1734 4107 1748
rect 4313 1753 4327 1767
rect 4293 1734 4307 1748
rect 4133 1693 4147 1707
rect 4073 1653 4087 1667
rect 4013 1633 4027 1647
rect 4013 1473 4027 1487
rect 3953 1434 3967 1448
rect 4073 1392 4087 1406
rect 4213 1692 4227 1706
rect 4253 1692 4267 1706
rect 4293 1692 4307 1706
rect 4253 1653 4267 1667
rect 4253 1493 4267 1507
rect 4253 1453 4267 1467
rect 4153 1434 4167 1448
rect 4193 1434 4207 1448
rect 4013 1313 4027 1327
rect 4133 1313 4147 1327
rect 3913 1273 3927 1287
rect 3893 1253 3907 1267
rect 3713 1233 3727 1247
rect 3753 1214 3767 1228
rect 3953 1214 3967 1228
rect 3993 1213 4007 1227
rect 3713 1153 3727 1167
rect 3773 1133 3787 1147
rect 3893 1153 3907 1167
rect 3933 1153 3947 1167
rect 3853 1073 3867 1087
rect 3933 993 3947 1007
rect 3953 973 3967 987
rect 3693 933 3707 947
rect 3753 933 3767 947
rect 3653 913 3667 927
rect 3593 873 3607 887
rect 3673 872 3687 886
rect 3733 853 3747 867
rect 3493 813 3507 827
rect 3533 813 3547 827
rect 3613 813 3627 827
rect 3533 753 3547 767
rect 3413 713 3427 727
rect 3473 713 3487 727
rect 3373 694 3387 708
rect 3233 633 3247 647
rect 3153 513 3167 527
rect 3193 473 3207 487
rect 3113 453 3127 467
rect 3113 394 3127 408
rect 3153 394 3167 408
rect 3313 652 3327 666
rect 3393 652 3407 666
rect 3353 633 3367 647
rect 3373 553 3387 567
rect 3333 493 3347 507
rect 3333 453 3347 467
rect 3293 394 3307 408
rect 3113 353 3127 367
rect 3173 352 3187 366
rect 3233 353 3247 367
rect 3313 352 3327 366
rect 3453 513 3467 527
rect 3433 453 3447 467
rect 3393 433 3407 447
rect 3373 253 3387 267
rect 3293 193 3307 207
rect 3373 193 3387 207
rect 3153 174 3167 188
rect 3233 173 3247 187
rect 3133 73 3147 87
rect 3233 132 3247 146
rect 3273 132 3287 146
rect 3313 132 3327 146
rect 3493 693 3507 707
rect 3573 694 3587 708
rect 3513 652 3527 666
rect 3553 652 3567 666
rect 3533 633 3547 647
rect 3693 753 3707 767
rect 3633 693 3647 707
rect 3733 694 3747 708
rect 3793 914 3807 928
rect 3833 914 3847 928
rect 3953 914 3967 928
rect 4353 2173 4367 2187
rect 4733 3293 4747 3307
rect 4613 3273 4627 3287
rect 4713 3252 4727 3266
rect 4713 3033 4727 3047
rect 4633 2994 4647 3008
rect 4673 2994 4687 3008
rect 4713 2933 4727 2947
rect 4673 2913 4687 2927
rect 4653 2873 4667 2887
rect 4633 2813 4647 2827
rect 4713 2773 4727 2787
rect 4693 2732 4707 2746
rect 4593 2713 4607 2727
rect 4593 2653 4607 2667
rect 4593 2613 4607 2627
rect 4573 2493 4587 2507
rect 4633 2533 4647 2547
rect 4493 2432 4507 2446
rect 4533 2432 4547 2446
rect 4493 2293 4507 2307
rect 4473 2273 4487 2287
rect 4513 2212 4527 2226
rect 4553 2193 4567 2207
rect 4473 2173 4487 2187
rect 4433 1993 4447 2007
rect 4353 1973 4367 1987
rect 4393 1973 4407 1987
rect 4433 1954 4447 1968
rect 4553 2113 4567 2127
rect 4553 2053 4567 2067
rect 4493 1993 4507 2007
rect 4473 1953 4487 1967
rect 4413 1912 4427 1926
rect 4453 1853 4467 1867
rect 4513 1973 4527 1987
rect 4593 2293 4607 2307
rect 4973 3533 4987 3547
rect 4933 3514 4947 3528
rect 4973 3514 4987 3528
rect 4893 3473 4907 3487
rect 4993 3472 5007 3486
rect 4953 3453 4967 3467
rect 4853 3373 4867 3387
rect 4813 3294 4827 3308
rect 5213 3693 5227 3707
rect 5073 3633 5087 3647
rect 5052 3473 5066 3487
rect 5193 3553 5207 3567
rect 5153 3514 5167 3528
rect 5073 3472 5087 3486
rect 5133 3472 5147 3486
rect 5193 3473 5207 3487
rect 5173 3453 5187 3467
rect 5033 3373 5047 3387
rect 4953 3333 4967 3347
rect 5073 3313 5087 3327
rect 5133 3313 5147 3327
rect 4973 3294 4987 3308
rect 4953 3252 4967 3266
rect 5013 3213 5027 3227
rect 5033 3173 5047 3187
rect 5073 3173 5087 3187
rect 4793 3033 4807 3047
rect 4953 3033 4967 3047
rect 4993 3033 5007 3047
rect 4793 2994 4807 3008
rect 4873 2973 4887 2987
rect 4813 2933 4827 2947
rect 4833 2873 4847 2887
rect 4813 2793 4827 2807
rect 4733 2713 4747 2727
rect 4793 2774 4807 2788
rect 4953 2994 4967 3008
rect 5153 3252 5167 3266
rect 5393 4034 5407 4048
rect 5413 3953 5427 3967
rect 5373 3933 5387 3947
rect 5493 4193 5507 4207
rect 5673 4753 5687 4767
rect 5773 5313 5787 5327
rect 5873 5333 5887 5347
rect 5853 5313 5867 5327
rect 5833 5253 5847 5267
rect 5813 5233 5827 5247
rect 5753 5193 5767 5207
rect 5753 5153 5767 5167
rect 5793 5113 5807 5127
rect 5853 5113 5867 5127
rect 5893 5253 5907 5267
rect 5893 5193 5907 5207
rect 5873 5093 5887 5107
rect 5793 5074 5807 5088
rect 5813 5032 5827 5046
rect 5773 4913 5787 4927
rect 5753 4853 5767 4867
rect 5813 4854 5827 4868
rect 5853 4853 5867 4867
rect 5833 4812 5847 4826
rect 5733 4793 5747 4807
rect 5813 4773 5827 4787
rect 5673 4673 5687 4687
rect 5653 4453 5667 4467
rect 5793 4753 5807 4767
rect 5773 4573 5787 4587
rect 5733 4554 5747 4568
rect 5713 4512 5727 4526
rect 5673 4373 5687 4387
rect 5633 4334 5647 4348
rect 5673 4334 5687 4348
rect 5853 4773 5867 4787
rect 5893 4673 5907 4687
rect 5973 5552 5987 5566
rect 5993 5513 6007 5527
rect 5973 5173 5987 5187
rect 5993 4873 6007 4887
rect 5973 4854 5987 4868
rect 5933 4813 5947 4827
rect 5993 4813 6007 4827
rect 5953 4793 5967 4807
rect 5933 4573 5947 4587
rect 5833 4513 5847 4527
rect 5773 4493 5787 4507
rect 5813 4493 5827 4507
rect 5753 4473 5767 4487
rect 5753 4413 5767 4427
rect 5733 4373 5747 4387
rect 5713 4333 5727 4347
rect 5553 4253 5567 4267
rect 5693 4293 5707 4307
rect 5653 4233 5667 4247
rect 5593 4193 5607 4207
rect 5573 4113 5587 4127
rect 5493 3992 5507 4006
rect 5533 3992 5547 4006
rect 5393 3913 5407 3927
rect 5473 3913 5487 3927
rect 5333 3893 5347 3907
rect 5253 3833 5267 3847
rect 5313 3833 5327 3847
rect 5253 3772 5267 3786
rect 5313 3772 5327 3786
rect 5573 3893 5587 3907
rect 5513 3873 5527 3887
rect 5553 3853 5567 3867
rect 5413 3814 5427 3828
rect 5473 3814 5487 3828
rect 5513 3814 5527 3828
rect 5353 3713 5367 3727
rect 5293 3613 5307 3627
rect 5233 3533 5247 3547
rect 5333 3514 5347 3528
rect 5373 3514 5387 3528
rect 5233 3473 5247 3487
rect 5273 3472 5287 3486
rect 5313 3472 5327 3486
rect 5373 3453 5387 3467
rect 5493 3772 5507 3786
rect 5573 3772 5587 3786
rect 5573 3733 5587 3747
rect 5553 3713 5567 3727
rect 5713 4193 5727 4207
rect 5633 4073 5647 4087
rect 5693 4073 5707 4087
rect 5613 4053 5627 4067
rect 5833 4473 5847 4487
rect 5793 4334 5807 4348
rect 5753 4253 5767 4267
rect 5813 4233 5827 4247
rect 5773 4133 5787 4147
rect 5733 4053 5747 4067
rect 5693 4034 5707 4048
rect 5753 4033 5767 4047
rect 5653 3993 5667 4007
rect 5633 3893 5647 3907
rect 5633 3853 5647 3867
rect 5673 3953 5687 3967
rect 5713 3933 5727 3947
rect 5673 3853 5687 3867
rect 5713 3853 5727 3867
rect 5653 3833 5667 3847
rect 5893 4554 5907 4568
rect 5913 4512 5927 4526
rect 5873 4333 5887 4347
rect 5933 4334 5947 4348
rect 5993 4333 6007 4347
rect 5853 4073 5867 4087
rect 5913 4292 5927 4306
rect 5993 4293 6007 4307
rect 5953 4253 5967 4267
rect 5933 4073 5947 4087
rect 5793 4033 5807 4047
rect 5853 4034 5867 4048
rect 5893 4034 5907 4048
rect 5853 3973 5867 3987
rect 5793 3873 5807 3887
rect 5833 3873 5847 3887
rect 5893 3973 5907 3987
rect 5873 3933 5887 3947
rect 5753 3813 5767 3827
rect 5813 3814 5827 3828
rect 5853 3814 5867 3828
rect 5553 3613 5567 3627
rect 5453 3514 5467 3528
rect 5493 3514 5507 3528
rect 5533 3514 5547 3528
rect 5313 3353 5327 3367
rect 5232 3293 5246 3307
rect 5253 3293 5267 3307
rect 5313 3294 5327 3308
rect 5233 3252 5247 3266
rect 5173 3213 5187 3227
rect 5213 3213 5227 3227
rect 5113 3033 5127 3047
rect 5153 3033 5167 3047
rect 5093 3013 5107 3027
rect 5033 2973 5047 2987
rect 4893 2873 4907 2887
rect 4973 2952 4987 2966
rect 5213 3033 5227 3047
rect 5293 3252 5307 3266
rect 5313 3233 5327 3247
rect 5473 3453 5487 3467
rect 5593 3693 5607 3707
rect 5593 3613 5607 3627
rect 5653 3772 5667 3786
rect 5693 3772 5707 3786
rect 5693 3673 5707 3687
rect 5613 3553 5627 3567
rect 5713 3553 5727 3567
rect 5613 3514 5627 3528
rect 5553 3453 5567 3467
rect 5533 3393 5547 3407
rect 5433 3373 5447 3387
rect 5593 3472 5607 3486
rect 5393 3294 5407 3308
rect 5453 3294 5467 3308
rect 5493 3294 5507 3308
rect 5433 3252 5447 3266
rect 5333 3133 5347 3147
rect 5373 3133 5387 3147
rect 5273 2952 5287 2966
rect 5173 2913 5187 2927
rect 5173 2873 5187 2887
rect 4953 2813 4967 2827
rect 4813 2732 4827 2746
rect 4853 2732 4867 2746
rect 4893 2733 4907 2747
rect 4793 2713 4807 2727
rect 4753 2613 4767 2627
rect 4713 2573 4727 2587
rect 4713 2533 4727 2547
rect 4753 2474 4767 2488
rect 4653 2433 4667 2447
rect 4693 2432 4707 2446
rect 4773 2433 4787 2447
rect 4653 2313 4667 2327
rect 4733 2313 4747 2327
rect 4633 2273 4647 2287
rect 4693 2254 4707 2268
rect 4633 2212 4647 2226
rect 4673 2212 4687 2226
rect 4813 2693 4827 2707
rect 4993 2774 5007 2788
rect 5073 2774 5087 2788
rect 5133 2774 5147 2788
rect 5013 2732 5027 2746
rect 4973 2693 4987 2707
rect 5153 2732 5167 2746
rect 5113 2653 5127 2667
rect 5073 2613 5087 2627
rect 5113 2613 5127 2627
rect 4973 2593 4987 2607
rect 5013 2593 5027 2607
rect 4873 2533 4887 2547
rect 4913 2533 4927 2547
rect 4953 2533 4967 2547
rect 4833 2473 4847 2487
rect 4913 2474 4927 2488
rect 4853 2432 4867 2446
rect 4813 2393 4827 2407
rect 4773 2353 4787 2367
rect 4813 2353 4827 2367
rect 4933 2433 4947 2447
rect 4933 2353 4947 2367
rect 4893 2313 4907 2327
rect 4933 2313 4947 2327
rect 4853 2253 4867 2267
rect 5033 2533 5047 2547
rect 5073 2474 5087 2488
rect 4973 2433 4987 2447
rect 5013 2432 5027 2446
rect 5053 2432 5067 2446
rect 4953 2273 4967 2287
rect 5033 2273 5047 2287
rect 5073 2273 5087 2287
rect 4973 2254 4987 2268
rect 5013 2254 5027 2268
rect 4793 2212 4807 2226
rect 4753 2173 4767 2187
rect 4813 2173 4827 2187
rect 4593 2133 4607 2147
rect 4573 1973 4587 1987
rect 4713 2033 4727 2047
rect 4653 1954 4667 1968
rect 4753 1954 4767 1968
rect 4613 1912 4627 1926
rect 4653 1913 4667 1927
rect 4573 1893 4587 1907
rect 4733 1853 4747 1867
rect 4773 1833 4787 1847
rect 4353 1773 4367 1787
rect 4433 1773 4447 1787
rect 4492 1773 4506 1787
rect 4513 1773 4527 1787
rect 4593 1773 4607 1787
rect 4393 1734 4407 1748
rect 4333 1673 4347 1687
rect 4313 1493 4327 1507
rect 4293 1393 4307 1407
rect 4313 1353 4327 1367
rect 4213 1313 4227 1327
rect 4033 1213 4047 1227
rect 4013 1153 4027 1167
rect 4273 1253 4287 1267
rect 4313 1214 4327 1228
rect 4493 1734 4507 1748
rect 4533 1734 4547 1748
rect 4653 1734 4667 1748
rect 4693 1734 4707 1748
rect 4753 1734 4767 1748
rect 4453 1533 4467 1547
rect 4373 1453 4387 1467
rect 4433 1453 4447 1467
rect 4553 1692 4567 1706
rect 4593 1692 4607 1706
rect 4553 1671 4567 1685
rect 4513 1513 4527 1527
rect 4473 1473 4487 1487
rect 4453 1433 4467 1447
rect 4393 1392 4407 1406
rect 4433 1392 4447 1406
rect 4393 1353 4407 1367
rect 4213 1172 4227 1186
rect 4253 1172 4267 1186
rect 4293 1172 4307 1186
rect 4053 1113 4067 1127
rect 4173 1113 4187 1127
rect 4053 1073 4067 1087
rect 3893 893 3907 907
rect 3873 853 3887 867
rect 3813 833 3827 847
rect 3673 652 3687 666
rect 3713 652 3727 666
rect 3693 633 3707 647
rect 3733 633 3747 647
rect 3633 593 3647 607
rect 3613 553 3627 567
rect 3593 533 3607 547
rect 3613 513 3627 527
rect 3573 473 3587 487
rect 3553 453 3567 467
rect 3473 433 3487 447
rect 3453 413 3467 427
rect 3533 393 3547 407
rect 3433 353 3447 367
rect 3493 352 3507 366
rect 3533 352 3547 366
rect 3453 174 3467 188
rect 3613 433 3627 447
rect 3833 694 3847 708
rect 4013 853 4027 867
rect 4073 1033 4087 1047
rect 4353 993 4367 1007
rect 4313 953 4327 967
rect 4073 893 4087 907
rect 4073 853 4087 867
rect 3973 833 3987 847
rect 3893 793 3907 807
rect 3993 793 4007 807
rect 3933 694 3947 708
rect 4033 694 4047 708
rect 4353 914 4367 928
rect 4213 872 4227 886
rect 4093 833 4107 847
rect 4313 773 4327 787
rect 4233 713 4247 727
rect 4273 713 4287 727
rect 3893 652 3907 666
rect 3853 633 3867 647
rect 4073 693 4087 707
rect 4173 693 4187 707
rect 3933 613 3947 627
rect 4053 613 4067 627
rect 4013 593 4027 607
rect 4153 553 4167 567
rect 3893 493 3907 507
rect 3873 433 3887 447
rect 3653 413 3667 427
rect 3753 413 3767 427
rect 3613 394 3627 408
rect 3633 293 3647 307
rect 3613 213 3627 227
rect 3393 132 3407 146
rect 3373 93 3387 107
rect 3533 132 3547 146
rect 3633 132 3647 146
rect 3593 113 3607 127
rect 3473 53 3487 67
rect 3793 394 3807 408
rect 3853 394 3867 408
rect 3813 352 3827 366
rect 3773 333 3787 347
rect 3713 273 3727 287
rect 3873 353 3887 367
rect 3853 213 3867 227
rect 3773 174 3787 188
rect 3813 174 3827 188
rect 4093 473 4107 487
rect 3933 394 3947 408
rect 4373 733 4387 747
rect 4333 713 4347 727
rect 4233 652 4247 666
rect 4333 633 4347 647
rect 4373 633 4387 647
rect 4633 1613 4647 1627
rect 4593 1473 4607 1487
rect 4493 1433 4507 1447
rect 4553 1434 4567 1448
rect 4493 1373 4507 1387
rect 4493 1313 4507 1327
rect 4473 1253 4487 1267
rect 4433 1213 4447 1227
rect 4613 1393 4627 1407
rect 4713 1673 4727 1687
rect 4673 1473 4687 1487
rect 4653 1433 4667 1447
rect 4713 1434 4727 1448
rect 4693 1373 4707 1387
rect 4653 1253 4667 1267
rect 4733 1253 4747 1267
rect 4573 1233 4587 1247
rect 4413 914 4427 928
rect 4453 1172 4467 1186
rect 4693 1214 4707 1228
rect 4793 1793 4807 1807
rect 4833 1954 4847 1968
rect 4913 2212 4927 2226
rect 5013 2212 5027 2226
rect 4893 1954 4907 1968
rect 4933 1954 4947 1968
rect 4953 1913 4967 1927
rect 4913 1853 4927 1867
rect 4853 1832 4867 1846
rect 4813 1753 4827 1767
rect 4953 1793 4967 1807
rect 5233 2913 5247 2927
rect 5293 2774 5307 2788
rect 5273 2732 5287 2746
rect 5233 2693 5247 2707
rect 5273 2693 5287 2707
rect 5133 2474 5147 2488
rect 5173 2474 5187 2488
rect 5213 2474 5227 2488
rect 5153 2432 5167 2446
rect 5193 2432 5207 2446
rect 5233 2432 5247 2446
rect 5313 2653 5327 2667
rect 5293 2474 5307 2488
rect 5293 2433 5307 2447
rect 5533 3253 5547 3267
rect 5513 3193 5527 3207
rect 5493 3113 5507 3127
rect 5473 3093 5487 3107
rect 5353 3073 5367 3087
rect 5413 3013 5427 3027
rect 5453 2994 5467 3008
rect 5393 2952 5407 2966
rect 5353 2913 5367 2927
rect 5393 2913 5407 2927
rect 5433 2913 5447 2927
rect 5353 2793 5367 2807
rect 5473 2833 5487 2847
rect 5433 2793 5447 2807
rect 5473 2774 5487 2788
rect 5353 2733 5367 2747
rect 5413 2713 5427 2727
rect 5473 2733 5487 2747
rect 5353 2693 5367 2707
rect 5453 2653 5467 2667
rect 5333 2633 5347 2647
rect 5373 2474 5387 2488
rect 5413 2474 5427 2488
rect 5453 2474 5467 2488
rect 5673 3353 5687 3367
rect 5573 3294 5587 3308
rect 5633 3294 5647 3308
rect 5773 3773 5787 3787
rect 5833 3753 5847 3767
rect 5793 3733 5807 3747
rect 5773 3673 5787 3687
rect 5833 3673 5847 3687
rect 5753 3633 5767 3647
rect 5753 3533 5767 3547
rect 5733 3513 5747 3527
rect 5873 3593 5887 3607
rect 5853 3533 5867 3547
rect 5833 3513 5847 3527
rect 5733 3473 5747 3487
rect 5713 3294 5727 3308
rect 5553 3173 5567 3187
rect 5533 3033 5547 3047
rect 5653 3233 5667 3247
rect 5613 3073 5627 3087
rect 5653 3033 5667 3047
rect 5573 2994 5587 3008
rect 5613 3013 5627 3027
rect 5513 2953 5527 2967
rect 5553 2952 5567 2966
rect 5513 2913 5527 2927
rect 5593 2913 5607 2927
rect 5613 2873 5627 2887
rect 5573 2774 5587 2788
rect 5813 3472 5827 3486
rect 5853 3473 5867 3487
rect 5773 3294 5787 3308
rect 5833 3413 5847 3427
rect 5813 3293 5827 3307
rect 5813 3253 5827 3267
rect 5793 3233 5807 3247
rect 5733 3113 5747 3127
rect 5813 3173 5827 3187
rect 5793 3053 5807 3067
rect 5773 3033 5787 3047
rect 5713 3013 5727 3027
rect 5733 2994 5747 3008
rect 5673 2953 5687 2967
rect 5713 2952 5727 2966
rect 5773 2933 5787 2947
rect 5753 2893 5767 2907
rect 5733 2873 5747 2887
rect 5653 2833 5667 2847
rect 5733 2833 5747 2847
rect 5673 2774 5687 2788
rect 5733 2774 5747 2788
rect 5533 2713 5547 2727
rect 5513 2573 5527 2587
rect 5513 2513 5527 2527
rect 5593 2693 5607 2707
rect 5613 2653 5627 2667
rect 5593 2573 5607 2587
rect 5533 2493 5547 2507
rect 5313 2413 5327 2427
rect 5353 2413 5367 2427
rect 5173 2253 5187 2267
rect 5093 2212 5107 2226
rect 5133 2212 5147 2226
rect 5173 2212 5187 2226
rect 5253 2393 5267 2407
rect 5293 2393 5307 2407
rect 5293 2353 5307 2367
rect 5253 2254 5267 2268
rect 5153 2133 5167 2147
rect 5193 2133 5207 2147
rect 5133 1993 5147 2007
rect 5053 1954 5067 1968
rect 5093 1954 5107 1968
rect 4993 1933 5007 1947
rect 5133 1913 5147 1927
rect 4993 1853 5007 1867
rect 5073 1853 5087 1867
rect 5193 2033 5207 2047
rect 5273 2133 5287 2147
rect 5453 2393 5467 2407
rect 5413 2313 5427 2327
rect 5353 2273 5367 2287
rect 5393 2273 5407 2287
rect 5333 2093 5347 2107
rect 5293 2033 5307 2047
rect 5233 1993 5247 2007
rect 5233 1954 5247 1968
rect 5013 1833 5027 1847
rect 5153 1833 5167 1847
rect 4913 1733 4927 1747
rect 4813 1692 4827 1706
rect 4993 1773 5007 1787
rect 5253 1912 5267 1926
rect 5393 2193 5407 2207
rect 5433 2093 5447 2107
rect 5313 1973 5327 1987
rect 5353 1973 5367 1987
rect 5413 1973 5427 1987
rect 5293 1853 5307 1867
rect 5253 1833 5267 1847
rect 5213 1773 5227 1787
rect 5233 1753 5247 1767
rect 5053 1734 5067 1748
rect 5213 1734 5227 1748
rect 4993 1692 5007 1706
rect 4953 1653 4967 1667
rect 4913 1633 4927 1647
rect 5073 1692 5087 1706
rect 5193 1692 5207 1706
rect 5053 1673 5067 1687
rect 5033 1653 5047 1667
rect 4773 1613 4787 1627
rect 4833 1613 4847 1627
rect 4773 1553 4787 1567
rect 4753 1233 4767 1247
rect 4793 1473 4807 1487
rect 4793 1433 4807 1447
rect 5233 1673 5247 1687
rect 5233 1633 5247 1647
rect 5013 1553 5027 1567
rect 5193 1553 5207 1567
rect 4953 1493 4967 1507
rect 4873 1434 4887 1448
rect 4933 1434 4947 1448
rect 4793 1393 4807 1407
rect 4853 1392 4867 1406
rect 4813 1353 4827 1367
rect 4853 1353 4867 1367
rect 4913 1353 4927 1367
rect 4893 1333 4907 1347
rect 5113 1533 5127 1547
rect 5233 1533 5247 1547
rect 5013 1473 5027 1487
rect 5053 1434 5067 1448
rect 5093 1447 5107 1448
rect 5093 1434 5107 1447
rect 4953 1393 4967 1407
rect 4993 1392 5007 1406
rect 5033 1392 5047 1406
rect 5073 1392 5087 1406
rect 5233 1473 5247 1487
rect 5153 1434 5167 1448
rect 5193 1434 5207 1448
rect 5373 1954 5387 1968
rect 5553 2474 5567 2488
rect 5533 2432 5547 2446
rect 5613 2313 5627 2327
rect 5673 2713 5687 2727
rect 5733 2713 5747 2727
rect 5713 2633 5727 2647
rect 5673 2474 5687 2488
rect 5693 2373 5707 2387
rect 5593 2273 5607 2287
rect 5493 2253 5507 2267
rect 5553 2254 5567 2268
rect 5633 2273 5647 2287
rect 5533 2212 5547 2226
rect 5573 2173 5587 2187
rect 5613 2113 5627 2127
rect 5533 2073 5547 2087
rect 5493 2053 5507 2067
rect 5353 1912 5367 1926
rect 5393 1912 5407 1926
rect 5333 1793 5347 1807
rect 5373 1753 5387 1767
rect 5333 1733 5347 1747
rect 5413 1734 5427 1748
rect 5393 1692 5407 1706
rect 5353 1673 5367 1687
rect 5473 1954 5487 1968
rect 5533 1973 5547 1987
rect 5673 2333 5687 2347
rect 5853 3393 5867 3407
rect 5953 4033 5967 4047
rect 5993 3973 6007 3987
rect 5993 3873 6007 3887
rect 5993 3753 6007 3767
rect 5953 3693 5967 3707
rect 5933 3593 5947 3607
rect 5913 3553 5927 3567
rect 5953 3514 5967 3528
rect 5993 3513 6007 3527
rect 5933 3472 5947 3486
rect 5953 3453 5967 3467
rect 5993 3473 6007 3487
rect 5973 3413 5987 3427
rect 5953 3313 5967 3327
rect 5913 3294 5927 3308
rect 5933 3252 5947 3266
rect 5973 3252 5987 3266
rect 5893 3233 5907 3247
rect 5873 3213 5887 3227
rect 5893 3193 5907 3207
rect 5893 2994 5907 3008
rect 5993 3093 6007 3107
rect 5993 3053 6007 3067
rect 5973 2993 5987 3007
rect 5853 2952 5867 2966
rect 5913 2952 5927 2966
rect 5953 2952 5967 2966
rect 5853 2893 5867 2907
rect 5833 2833 5847 2847
rect 5813 2713 5827 2727
rect 5753 2573 5767 2587
rect 5873 2774 5887 2788
rect 5893 2713 5907 2727
rect 5893 2673 5907 2687
rect 5853 2513 5867 2527
rect 5833 2493 5847 2507
rect 5773 2474 5787 2488
rect 5813 2474 5827 2488
rect 5853 2474 5867 2488
rect 5833 2432 5847 2446
rect 5853 2413 5867 2427
rect 5893 2413 5907 2427
rect 5793 2393 5807 2407
rect 5773 2373 5787 2387
rect 5733 2273 5747 2287
rect 5673 2253 5687 2267
rect 5773 2253 5787 2267
rect 5673 2213 5687 2227
rect 5653 2113 5667 2127
rect 5653 2073 5667 2087
rect 5633 2013 5647 2027
rect 5613 1933 5627 1947
rect 5533 1853 5547 1867
rect 5473 1773 5487 1787
rect 5333 1473 5347 1487
rect 5373 1473 5387 1487
rect 5453 1473 5467 1487
rect 5273 1453 5287 1467
rect 5313 1453 5327 1467
rect 5113 1393 5127 1407
rect 5173 1392 5187 1406
rect 5133 1373 5147 1387
rect 5213 1373 5227 1387
rect 5093 1353 5107 1367
rect 5133 1333 5147 1347
rect 4993 1313 5007 1327
rect 4813 1293 4827 1307
rect 4873 1293 4887 1307
rect 4933 1293 4947 1307
rect 4973 1293 4987 1307
rect 4793 1253 4807 1267
rect 4633 1133 4647 1147
rect 4513 1053 4527 1067
rect 4753 1173 4767 1187
rect 4713 1013 4727 1027
rect 4633 993 4647 1007
rect 4553 953 4567 967
rect 4493 914 4507 928
rect 4413 873 4427 887
rect 4473 872 4487 886
rect 4793 1053 4807 1067
rect 4953 1273 4967 1287
rect 4873 1253 4887 1267
rect 4913 1253 4927 1267
rect 4833 1172 4847 1186
rect 4873 1172 4887 1186
rect 4913 1172 4927 1186
rect 4833 1133 4847 1147
rect 4873 1133 4887 1147
rect 4873 1093 4887 1107
rect 4913 1093 4927 1107
rect 4813 1033 4827 1047
rect 4933 1033 4947 1047
rect 4753 973 4767 987
rect 4813 973 4827 987
rect 4573 914 4587 928
rect 4693 914 4707 928
rect 4733 914 4747 928
rect 4573 873 4587 887
rect 4633 872 4647 886
rect 4553 833 4567 847
rect 4513 813 4527 827
rect 4733 833 4747 847
rect 4733 793 4747 807
rect 4713 773 4727 787
rect 4453 753 4467 767
rect 4673 753 4687 767
rect 4493 693 4507 707
rect 4593 694 4607 708
rect 4633 694 4647 708
rect 4673 694 4687 708
rect 4493 613 4507 627
rect 4573 593 4587 607
rect 4293 493 4307 507
rect 4393 493 4407 507
rect 4173 413 4187 427
rect 4213 413 4227 427
rect 3913 353 3927 367
rect 3953 333 3967 347
rect 4033 373 4047 387
rect 4233 394 4247 408
rect 4033 333 4047 347
rect 4113 352 4127 366
rect 4173 353 4187 367
rect 4113 313 4127 327
rect 3933 293 3947 307
rect 4013 293 4027 307
rect 4073 293 4087 307
rect 3913 193 3927 207
rect 4213 313 4227 327
rect 4193 273 4207 287
rect 4273 353 4287 367
rect 4253 233 4267 247
rect 4353 433 4367 447
rect 4413 433 4427 447
rect 4473 433 4487 447
rect 4553 433 4567 447
rect 4313 393 4327 407
rect 4393 412 4407 426
rect 4453 394 4467 408
rect 4373 352 4387 366
rect 4413 352 4427 366
rect 4513 394 4527 408
rect 4573 413 4587 427
rect 4533 352 4547 366
rect 4673 633 4687 647
rect 4933 953 4947 967
rect 4853 914 4867 928
rect 4793 853 4807 867
rect 4813 833 4827 847
rect 4753 733 4767 747
rect 4773 694 4787 708
rect 4873 873 4887 887
rect 5113 1253 5127 1267
rect 5013 1214 5027 1228
rect 5053 1214 5067 1228
rect 4973 1133 4987 1147
rect 5173 1313 5187 1327
rect 5213 1214 5227 1228
rect 5133 1173 5147 1187
rect 5073 1153 5087 1167
rect 5193 1153 5207 1167
rect 5193 1093 5207 1107
rect 5053 1033 5067 1047
rect 4993 1013 5007 1027
rect 4953 914 4967 928
rect 4933 872 4947 886
rect 4993 872 5007 886
rect 4993 853 5007 867
rect 4873 833 4887 847
rect 4833 773 4847 787
rect 5013 773 5027 787
rect 5153 953 5167 967
rect 5113 914 5127 928
rect 5133 872 5147 886
rect 5253 1173 5267 1187
rect 5233 1033 5247 1047
rect 5393 1452 5407 1466
rect 5353 1434 5367 1448
rect 5313 1393 5327 1407
rect 5293 1373 5307 1387
rect 5313 1333 5327 1347
rect 5373 1392 5387 1406
rect 5433 1393 5447 1407
rect 5293 1293 5307 1307
rect 5333 1293 5347 1307
rect 5273 1153 5287 1167
rect 5373 1273 5387 1287
rect 5633 1912 5647 1926
rect 5633 1873 5647 1887
rect 5513 1734 5527 1748
rect 5553 1734 5567 1748
rect 5613 1734 5627 1748
rect 5713 2212 5727 2226
rect 5813 2373 5827 2387
rect 5713 2173 5727 2187
rect 5753 2153 5767 2167
rect 5693 2093 5707 2107
rect 5712 1993 5726 2007
rect 5733 1993 5747 2007
rect 5833 2313 5847 2327
rect 5913 2333 5927 2347
rect 5973 2774 5987 2788
rect 5953 2633 5967 2647
rect 5933 2313 5947 2327
rect 5893 2273 5907 2287
rect 5833 2213 5847 2227
rect 5813 2193 5827 2207
rect 5773 1953 5787 1967
rect 5713 1912 5727 1926
rect 5753 1912 5767 1926
rect 5693 1833 5707 1847
rect 5673 1793 5687 1807
rect 5713 1753 5727 1767
rect 5533 1653 5547 1667
rect 5693 1692 5707 1706
rect 5633 1672 5647 1686
rect 5493 1593 5507 1607
rect 5593 1593 5607 1607
rect 5613 1553 5627 1567
rect 5513 1453 5527 1467
rect 5553 1453 5567 1467
rect 5473 1433 5487 1447
rect 5693 1653 5707 1667
rect 5733 1593 5747 1607
rect 5733 1473 5747 1487
rect 5633 1433 5647 1447
rect 5593 1413 5607 1427
rect 5493 1392 5507 1406
rect 5473 1253 5487 1267
rect 5333 1214 5347 1228
rect 5373 1214 5387 1228
rect 5653 1373 5667 1387
rect 5813 2053 5827 2067
rect 5873 2212 5887 2226
rect 5873 2193 5887 2207
rect 5993 2573 6007 2587
rect 5993 2474 6007 2488
rect 5973 2393 5987 2407
rect 5973 2273 5987 2287
rect 5913 2153 5927 2167
rect 5953 2153 5967 2167
rect 5873 1993 5887 2007
rect 5833 1973 5847 1987
rect 5933 2093 5947 2107
rect 5973 2033 5987 2047
rect 5933 1993 5947 2007
rect 5973 1993 5987 2007
rect 5913 1953 5927 1967
rect 5853 1912 5867 1926
rect 5893 1873 5907 1887
rect 5853 1773 5867 1787
rect 5853 1734 5867 1748
rect 5793 1692 5807 1706
rect 5833 1692 5847 1706
rect 5853 1473 5867 1487
rect 5733 1373 5747 1387
rect 5613 1353 5627 1367
rect 5833 1353 5847 1367
rect 5553 1233 5567 1247
rect 5453 1213 5467 1227
rect 5513 1214 5527 1228
rect 5453 1172 5467 1186
rect 5393 1093 5407 1107
rect 5293 1053 5307 1067
rect 5253 993 5267 1007
rect 5273 953 5287 967
rect 5253 914 5267 928
rect 5393 993 5407 1007
rect 5213 873 5227 887
rect 5053 833 5067 847
rect 5133 833 5147 847
rect 5193 833 5207 847
rect 5033 733 5047 747
rect 4913 694 4927 708
rect 4993 694 5007 708
rect 5073 694 5087 708
rect 4713 653 4727 667
rect 4793 652 4807 666
rect 4693 593 4707 607
rect 4753 593 4767 607
rect 4773 573 4787 587
rect 4713 513 4727 527
rect 4633 394 4647 408
rect 4673 394 4687 408
rect 4793 413 4807 427
rect 4633 353 4647 367
rect 4573 333 4587 347
rect 4613 333 4627 347
rect 4673 333 4687 347
rect 4373 313 4387 327
rect 4453 313 4467 327
rect 4733 352 4747 366
rect 4773 353 4787 367
rect 4933 633 4947 647
rect 5093 633 5107 647
rect 5053 593 5067 607
rect 4993 573 5007 587
rect 4833 513 4847 527
rect 4813 393 4827 407
rect 5053 493 5067 507
rect 5093 493 5107 507
rect 4933 473 4947 487
rect 4873 413 4887 427
rect 5053 433 5067 447
rect 5013 413 5027 427
rect 5053 394 5067 408
rect 5193 793 5207 807
rect 5273 853 5287 867
rect 5313 853 5327 867
rect 5453 953 5467 967
rect 5533 1172 5547 1186
rect 5533 993 5547 1007
rect 5493 914 5507 928
rect 5393 873 5407 887
rect 5433 872 5447 886
rect 5473 872 5487 886
rect 5513 872 5527 886
rect 5353 833 5367 847
rect 5453 853 5467 867
rect 5393 793 5407 807
rect 5233 733 5247 747
rect 5353 733 5367 747
rect 5253 713 5267 727
rect 5233 694 5247 708
rect 5213 633 5227 647
rect 5253 593 5267 607
rect 5153 493 5167 507
rect 4893 352 4907 366
rect 4933 352 4947 366
rect 4993 352 5007 366
rect 5033 352 5047 366
rect 5093 353 5107 367
rect 5313 693 5327 707
rect 5353 694 5367 708
rect 5313 513 5327 527
rect 5433 653 5447 667
rect 5453 493 5467 507
rect 5353 413 5367 427
rect 5373 413 5387 427
rect 5413 413 5427 427
rect 5193 394 5207 408
rect 5293 394 5307 408
rect 5173 352 5187 366
rect 5213 352 5227 366
rect 5373 352 5387 366
rect 4793 333 4807 347
rect 4853 333 4867 347
rect 5113 333 5127 347
rect 5333 333 5347 347
rect 4693 313 4707 327
rect 4313 293 4327 307
rect 4353 293 4367 307
rect 4393 293 4407 307
rect 4673 293 4687 307
rect 5513 833 5527 847
rect 5553 953 5567 967
rect 5533 753 5547 767
rect 5653 1253 5667 1267
rect 5713 1253 5727 1267
rect 5813 1253 5827 1267
rect 5733 1213 5747 1227
rect 5713 1192 5727 1206
rect 5673 1172 5687 1186
rect 5633 1113 5647 1127
rect 5693 1093 5707 1107
rect 5592 993 5606 1007
rect 5613 993 5627 1007
rect 5753 1172 5767 1186
rect 5733 1113 5747 1127
rect 5853 1113 5867 1127
rect 5833 1093 5847 1107
rect 5753 993 5767 1007
rect 5573 914 5587 928
rect 5613 914 5627 928
rect 5653 933 5667 947
rect 5713 933 5727 947
rect 5593 833 5607 847
rect 5673 873 5687 887
rect 5633 813 5647 827
rect 5593 793 5607 807
rect 5513 733 5527 747
rect 5553 733 5567 747
rect 5553 694 5567 708
rect 5633 753 5647 767
rect 5613 733 5627 747
rect 5593 693 5607 707
rect 5533 652 5547 666
rect 5593 493 5607 507
rect 5513 453 5527 467
rect 5433 393 5447 407
rect 5473 393 5487 407
rect 5553 394 5567 408
rect 5413 273 5427 287
rect 4293 253 4307 267
rect 4493 253 4507 267
rect 4273 213 4287 227
rect 3713 133 3727 147
rect 3753 113 3767 127
rect 3993 173 4007 187
rect 4053 174 4067 188
rect 3973 153 3987 167
rect 3913 132 3927 146
rect 3973 93 3987 107
rect 3953 53 3967 67
rect 4393 174 4407 188
rect 4473 173 4487 187
rect 4153 153 4167 167
rect 4073 113 4087 127
rect 4373 132 4387 146
rect 4473 132 4487 146
rect 4293 113 4307 127
rect 4413 113 4427 127
rect 4553 233 4567 247
rect 4513 213 4527 227
rect 4513 173 4527 187
rect 5333 213 5347 227
rect 4713 173 4727 187
rect 4793 174 4807 188
rect 5033 174 5047 188
rect 5153 174 5167 188
rect 5213 173 5227 187
rect 5293 174 5307 188
rect 5393 173 5407 187
rect 5493 352 5507 366
rect 5533 352 5547 366
rect 5793 914 5807 928
rect 5833 872 5847 886
rect 5933 1773 5947 1787
rect 5933 1533 5947 1547
rect 5933 1113 5947 1127
rect 5953 1093 5967 1107
rect 5853 833 5867 847
rect 5693 753 5707 767
rect 5773 813 5787 827
rect 5773 753 5787 767
rect 5633 652 5647 666
rect 5673 652 5687 666
rect 5833 694 5847 708
rect 5933 914 5947 928
rect 5913 872 5927 886
rect 5913 833 5927 847
rect 5873 693 5887 707
rect 5713 533 5727 547
rect 5673 453 5687 467
rect 5713 453 5727 467
rect 5613 394 5627 408
rect 5713 413 5727 427
rect 5733 394 5747 408
rect 5593 333 5607 347
rect 5693 352 5707 366
rect 5653 333 5667 347
rect 5633 293 5647 307
rect 5533 213 5547 227
rect 5613 213 5627 227
rect 4533 132 4547 146
rect 4493 93 4507 107
rect 4413 73 4427 87
rect 4033 53 4047 67
rect 4393 53 4407 67
rect 4433 53 4447 67
rect 4673 132 4687 146
rect 4713 132 4727 146
rect 4913 132 4927 146
rect 4613 93 4627 107
rect 4853 93 4867 107
rect 3813 33 3827 47
rect 3873 33 3887 47
rect 3993 33 4007 47
rect 4573 33 4587 47
rect 3073 13 3087 27
rect 3113 13 3127 27
rect 3173 13 3187 27
rect 3693 13 3707 27
rect 3773 13 3787 27
rect 5353 132 5367 146
rect 5473 174 5487 188
rect 5413 132 5427 146
rect 5453 113 5467 127
rect 5673 273 5687 287
rect 5773 652 5787 666
rect 5813 652 5827 666
rect 5773 533 5787 547
rect 5853 533 5867 547
rect 5873 453 5887 467
rect 5833 394 5847 408
rect 5773 233 5787 247
rect 5853 233 5867 247
rect 5933 693 5947 707
rect 5913 174 5927 188
rect 5533 113 5547 127
rect 5393 73 5407 87
rect 5673 133 5687 147
rect 5753 132 5767 146
rect 5633 113 5647 127
rect 5873 113 5887 127
rect 5993 1833 6007 1847
rect 5993 1213 6007 1227
rect 5993 1093 6007 1107
rect 5973 293 5987 307
rect 5993 113 6007 127
rect 5313 53 5327 67
rect 5593 53 5607 67
rect 5933 53 5947 67
rect 5213 33 5227 47
<< metal3 >>
rect 387 5996 413 6004
rect 887 5996 1193 6004
rect 1207 5996 3093 6004
rect 3307 5996 3333 6004
rect 3987 5996 4013 6004
rect 4067 5996 5233 6004
rect 1027 5976 1053 5984
rect 2767 5976 2793 5984
rect 3207 5976 3233 5984
rect 3247 5976 5113 5984
rect 2307 5956 2373 5964
rect 167 5936 1473 5944
rect 4747 5936 5073 5944
rect 2507 5916 2664 5924
rect 287 5896 353 5904
rect 447 5896 473 5904
rect 1087 5896 1113 5904
rect 1547 5896 1653 5904
rect 127 5856 173 5864
rect 187 5856 253 5864
rect 667 5856 793 5864
rect 887 5855 913 5863
rect 1307 5856 1353 5864
rect 1676 5864 1684 5913
rect 2656 5908 2664 5916
rect 3867 5916 4093 5924
rect 4107 5916 4133 5924
rect 1887 5897 1913 5905
rect 2167 5896 2293 5904
rect 2427 5896 2453 5904
rect 2567 5896 2613 5904
rect 2667 5897 2713 5905
rect 2827 5896 2853 5904
rect 3367 5896 3393 5904
rect 3827 5896 3953 5904
rect 4147 5896 4253 5904
rect 4387 5897 4433 5905
rect 4487 5896 4553 5904
rect 4627 5897 4793 5905
rect 4887 5896 4932 5904
rect 4967 5896 5013 5904
rect 5307 5896 5353 5904
rect 5407 5896 5453 5904
rect 5547 5897 5573 5905
rect 5627 5897 5653 5905
rect 5767 5897 5793 5905
rect 1676 5856 1693 5864
rect 2547 5855 2573 5863
rect 2587 5855 2633 5863
rect 3587 5856 3633 5864
rect 4767 5856 4853 5864
rect 4867 5855 4953 5863
rect 5047 5856 5173 5864
rect 5247 5856 5273 5864
rect 5367 5855 5433 5863
rect 607 5836 644 5844
rect 636 5824 644 5836
rect 1427 5836 1653 5844
rect 1947 5836 2073 5844
rect 2347 5836 2513 5844
rect 2527 5836 2673 5844
rect 2687 5836 3153 5844
rect 3707 5836 4093 5844
rect 4107 5836 4373 5844
rect 4607 5836 4713 5844
rect 5667 5836 5753 5844
rect 5767 5836 5813 5844
rect 636 5816 953 5824
rect 1367 5816 1973 5824
rect 1987 5816 2313 5824
rect 4596 5824 4604 5833
rect 4467 5816 4604 5824
rect 4807 5816 4893 5824
rect 5187 5816 5233 5824
rect 5247 5816 5313 5824
rect 5547 5816 5593 5824
rect 1227 5796 1293 5804
rect 1307 5796 2733 5804
rect 3047 5796 3213 5804
rect 1887 5776 1933 5784
rect 1947 5776 2413 5784
rect 2427 5776 2753 5784
rect 3167 5776 4413 5784
rect 2747 5756 4053 5764
rect 4596 5756 4993 5764
rect 2387 5736 2453 5744
rect 2727 5736 4193 5744
rect 4596 5744 4604 5756
rect 5007 5756 5133 5764
rect 4307 5736 4604 5744
rect 5447 5716 5813 5724
rect 1207 5696 1313 5704
rect 1867 5696 1993 5704
rect 2007 5696 2553 5704
rect 4787 5696 4933 5704
rect 807 5676 1253 5684
rect 1267 5676 1353 5684
rect 2067 5676 2433 5684
rect 4187 5676 4453 5684
rect 5287 5676 5573 5684
rect 307 5656 513 5664
rect 527 5656 673 5664
rect 687 5656 2333 5664
rect 2567 5656 2713 5664
rect 2967 5656 3173 5664
rect 4567 5656 4733 5664
rect 4747 5656 4853 5664
rect 4907 5656 5193 5664
rect 5207 5656 5353 5664
rect 5487 5656 5692 5664
rect 5727 5656 5853 5664
rect 987 5636 1393 5644
rect 1407 5636 1573 5644
rect 1767 5636 1933 5644
rect 2327 5636 2553 5644
rect 4127 5636 4253 5644
rect 4267 5636 4333 5644
rect 4467 5636 4973 5644
rect 3167 5616 3213 5624
rect 3227 5616 3453 5624
rect 3467 5616 3573 5624
rect 3807 5616 3913 5624
rect 4447 5616 4533 5624
rect 4967 5616 5113 5624
rect -24 5584 -16 5604
rect 127 5596 193 5604
rect 207 5596 233 5604
rect 287 5597 353 5605
rect 427 5596 453 5604
rect 467 5596 553 5604
rect 567 5596 713 5604
rect 807 5597 853 5605
rect 907 5596 1013 5604
rect 1507 5597 1533 5605
rect 1727 5597 1793 5605
rect 1807 5596 1893 5604
rect 1987 5597 2033 5605
rect 2087 5596 2192 5604
rect -24 5576 13 5584
rect 547 5556 693 5564
rect 927 5556 973 5564
rect 1196 5547 1204 5594
rect 1436 5564 1444 5594
rect 2227 5597 2253 5605
rect 2507 5596 2853 5604
rect 3407 5596 3593 5604
rect 3667 5597 3753 5605
rect 3847 5597 3953 5605
rect 4047 5597 4073 5605
rect 4307 5596 4413 5604
rect 4587 5597 4612 5605
rect 4647 5597 4693 5605
rect 4707 5596 4893 5604
rect 5087 5596 5113 5604
rect 1667 5576 2144 5584
rect 2136 5566 2144 5576
rect 1436 5556 1553 5564
rect 1567 5556 1693 5564
rect 2007 5555 2093 5563
rect 2387 5555 2433 5563
rect 2627 5555 2693 5563
rect 2856 5556 2873 5564
rect 27 5536 93 5544
rect 107 5536 453 5544
rect 2227 5536 2313 5544
rect 2856 5544 2864 5556
rect 3187 5555 3273 5563
rect 4147 5555 4173 5563
rect 4187 5556 4233 5564
rect 4347 5556 4673 5564
rect 4767 5556 4833 5564
rect 4887 5555 4933 5563
rect 4987 5556 5013 5564
rect 5036 5547 5044 5594
rect 5247 5596 5393 5604
rect 5407 5596 5553 5604
rect 5567 5596 5653 5604
rect 5867 5596 5953 5604
rect 5696 5584 5704 5594
rect 5696 5576 5724 5584
rect 5147 5555 5213 5563
rect 5547 5556 5673 5564
rect 5716 5564 5724 5576
rect 5716 5556 5733 5564
rect 5747 5556 5973 5564
rect 5987 5556 6044 5564
rect 2727 5536 2864 5544
rect 5307 5536 5533 5544
rect 187 5516 533 5524
rect 747 5516 853 5524
rect 967 5516 1073 5524
rect 2867 5516 2913 5524
rect 3507 5516 3713 5524
rect 4007 5516 4093 5524
rect 4187 5516 4393 5524
rect 5227 5516 5373 5524
rect 5767 5516 5993 5524
rect 707 5496 873 5504
rect 2087 5496 2193 5504
rect 3287 5496 3573 5504
rect 3787 5496 3933 5504
rect 3947 5496 4513 5504
rect 5027 5496 5173 5504
rect 5407 5496 5493 5504
rect 807 5476 973 5484
rect 1167 5476 1213 5484
rect 1427 5476 1493 5484
rect 1507 5476 2053 5484
rect 2427 5476 2453 5484
rect 2927 5476 2993 5484
rect 3447 5476 3733 5484
rect 4387 5476 4553 5484
rect 4567 5476 4753 5484
rect 267 5456 613 5464
rect 1747 5456 1913 5464
rect 1927 5456 2133 5464
rect 3507 5456 4033 5464
rect 4047 5456 4173 5464
rect 4607 5456 4633 5464
rect 4647 5456 4893 5464
rect 4907 5456 4993 5464
rect 5067 5456 5093 5464
rect 5107 5456 5333 5464
rect 5387 5456 5453 5464
rect 5807 5456 5873 5464
rect 647 5436 833 5444
rect 847 5436 1033 5444
rect 1047 5436 1133 5444
rect 1187 5436 1733 5444
rect 1747 5436 1773 5444
rect 1947 5436 1973 5444
rect 1987 5436 2093 5444
rect 3667 5436 3833 5444
rect 3847 5436 3953 5444
rect 4307 5436 4433 5444
rect 4447 5436 4613 5444
rect 4627 5436 4713 5444
rect 4847 5436 5033 5444
rect 147 5416 173 5424
rect 367 5416 513 5424
rect 867 5416 993 5424
rect 1287 5416 1373 5424
rect 1687 5416 1853 5424
rect 2007 5416 2033 5424
rect 2487 5416 2713 5424
rect 3627 5416 3733 5424
rect 4227 5416 4273 5424
rect 4827 5416 5053 5424
rect 5187 5416 5433 5424
rect 5447 5416 5793 5424
rect 5847 5416 5893 5424
rect 587 5396 633 5404
rect 2747 5396 3493 5404
rect 3607 5396 3793 5404
rect 3867 5396 3913 5404
rect 4007 5396 4053 5404
rect 5587 5396 5693 5404
rect 107 5376 213 5384
rect 236 5376 253 5384
rect 236 5347 244 5376
rect 307 5376 393 5384
rect 407 5377 453 5385
rect 507 5376 553 5384
rect 727 5376 753 5384
rect 776 5376 793 5384
rect 776 5364 784 5376
rect 887 5377 913 5385
rect 927 5376 1033 5384
rect 1087 5376 1173 5384
rect 616 5356 784 5364
rect 127 5335 193 5343
rect 616 5346 624 5356
rect 667 5335 693 5343
rect 707 5336 773 5344
rect 827 5335 853 5343
rect 947 5336 972 5344
rect 1196 5346 1204 5393
rect 1336 5376 1353 5384
rect 1336 5347 1344 5376
rect 1407 5376 1453 5384
rect 1536 5347 1544 5374
rect 1587 5376 1633 5384
rect 1767 5376 1813 5384
rect 1947 5376 1993 5384
rect 2147 5376 2613 5384
rect 2787 5377 2853 5385
rect 2987 5377 3033 5385
rect 3107 5376 3333 5384
rect 3387 5377 3413 5385
rect 3427 5376 3473 5384
rect 3527 5377 3573 5385
rect 4107 5377 4133 5385
rect 4156 5376 4253 5384
rect 1007 5335 1053 5343
rect 1427 5336 1513 5344
rect 1536 5336 1553 5347
rect 1540 5333 1553 5336
rect 1707 5335 1733 5343
rect 1787 5335 1833 5343
rect 1887 5335 1933 5343
rect 2027 5335 2072 5343
rect 2107 5336 2153 5344
rect 2387 5335 2453 5343
rect 2967 5336 3133 5344
rect 3447 5335 3493 5343
rect 3607 5335 3633 5343
rect 3836 5344 3844 5374
rect 4156 5364 4164 5376
rect 4407 5384 4420 5387
rect 4407 5373 4424 5384
rect 4767 5377 4833 5385
rect 4416 5364 4424 5373
rect 4116 5356 4164 5364
rect 4276 5356 4424 5364
rect 3836 5336 3873 5344
rect 4116 5344 4124 5356
rect 4276 5346 4284 5356
rect 4416 5346 4424 5356
rect 4476 5347 4484 5374
rect 3987 5336 4124 5344
rect 4327 5335 4373 5343
rect 4476 5336 4493 5347
rect 4480 5333 4493 5336
rect 4787 5335 4812 5343
rect 5016 5346 5024 5393
rect 5187 5376 5324 5384
rect 5036 5364 5044 5374
rect 5036 5356 5184 5364
rect 4847 5336 4873 5344
rect 5067 5335 5093 5343
rect 5176 5344 5184 5356
rect 5176 5336 5273 5344
rect 5316 5346 5324 5376
rect 5347 5377 5373 5385
rect 5447 5384 5460 5387
rect 5447 5373 5464 5384
rect 5527 5377 5553 5385
rect 5767 5376 5833 5384
rect 5456 5346 5464 5373
rect 5876 5347 5884 5373
rect 5367 5335 5393 5343
rect 5687 5336 5713 5344
rect 287 5316 433 5324
rect 447 5316 533 5324
rect 547 5316 873 5324
rect 1627 5316 1753 5324
rect 2607 5316 2633 5324
rect 3427 5316 3813 5324
rect 4207 5316 4533 5324
rect 4547 5316 4573 5324
rect 4747 5316 5113 5324
rect 5647 5316 5733 5324
rect 5787 5316 5853 5324
rect 227 5296 253 5304
rect 587 5296 1153 5304
rect 1267 5296 1413 5304
rect 1567 5296 2493 5304
rect 2667 5296 2773 5304
rect 2867 5296 3333 5304
rect 3647 5296 3673 5304
rect 3687 5296 3773 5304
rect 3867 5296 4013 5304
rect 4027 5296 4093 5304
rect 4107 5296 4493 5304
rect 5287 5296 5473 5304
rect 1187 5276 1513 5284
rect 1667 5276 1873 5284
rect 1967 5276 2433 5284
rect 2867 5276 3533 5284
rect 3847 5276 4213 5284
rect 4627 5276 5153 5284
rect 527 5256 1553 5264
rect 2467 5256 2793 5264
rect 2807 5256 2893 5264
rect 4707 5256 4953 5264
rect 5847 5256 5893 5264
rect 907 5236 1173 5244
rect 1487 5236 1653 5244
rect 1727 5236 2153 5244
rect 2167 5236 2373 5244
rect 2527 5236 2713 5244
rect 2727 5236 3093 5244
rect 5587 5236 5813 5244
rect 1467 5216 2233 5224
rect 2427 5216 2473 5224
rect 4067 5216 5133 5224
rect 1167 5196 1293 5204
rect 1567 5196 1613 5204
rect 1687 5196 2213 5204
rect 3007 5196 3113 5204
rect 3127 5196 3893 5204
rect 4076 5196 4613 5204
rect 1507 5176 2853 5184
rect 4076 5184 4084 5196
rect 5767 5196 5893 5204
rect 2896 5176 4084 5184
rect 887 5156 933 5164
rect 947 5156 1333 5164
rect 1527 5156 1953 5164
rect 2227 5156 2733 5164
rect 2896 5164 2904 5176
rect 5487 5176 5973 5184
rect 2787 5156 2904 5164
rect 3167 5156 3253 5164
rect 5627 5156 5753 5164
rect 2207 5136 2753 5144
rect 2767 5136 2973 5144
rect 3387 5136 3513 5144
rect 3527 5136 3713 5144
rect 247 5116 273 5124
rect 1127 5116 1213 5124
rect 1227 5116 1573 5124
rect 1587 5116 1613 5124
rect 2336 5116 2393 5124
rect 1427 5096 1593 5104
rect 2336 5104 2344 5116
rect 2447 5116 2653 5124
rect 2747 5116 3033 5124
rect 3047 5116 3193 5124
rect 3207 5116 3313 5124
rect 4047 5116 4093 5124
rect 5147 5116 5373 5124
rect 5427 5116 5513 5124
rect 5807 5116 5853 5124
rect 2067 5096 2344 5104
rect 3347 5096 3473 5104
rect 3987 5096 4133 5104
rect 5667 5096 5873 5104
rect 107 5076 233 5084
rect 467 5077 593 5085
rect 707 5077 733 5085
rect 756 5076 813 5084
rect 656 5064 664 5074
rect 756 5064 764 5076
rect 827 5076 993 5084
rect 1087 5076 1253 5084
rect 1267 5076 1373 5084
rect 1847 5077 1873 5085
rect 1927 5077 1973 5085
rect 2327 5077 2353 5085
rect 2567 5076 2673 5084
rect 2687 5077 2793 5085
rect 2907 5076 2993 5084
rect 3016 5076 3153 5084
rect 476 5056 764 5064
rect 476 5046 484 5056
rect 307 5035 353 5043
rect 587 5036 673 5044
rect 807 5035 873 5043
rect 1107 5036 1393 5044
rect 1447 5036 1493 5044
rect 1587 5036 1673 5044
rect 1947 5036 2033 5044
rect 2227 5036 2373 5044
rect 2427 5036 2453 5044
rect 3016 5046 3024 5076
rect 3167 5076 3344 5084
rect 3336 5064 3344 5076
rect 3707 5076 3813 5084
rect 3827 5076 4233 5084
rect 4387 5077 4433 5085
rect 4527 5077 4573 5085
rect 4627 5076 4753 5084
rect 4847 5076 4893 5084
rect 4947 5076 4993 5084
rect 5087 5076 5193 5084
rect 5347 5077 5413 5085
rect 5676 5076 5793 5084
rect 3336 5056 3524 5064
rect 2707 5036 2833 5044
rect 2887 5036 3013 5044
rect 3127 5035 3173 5043
rect 3287 5036 3313 5044
rect 3516 5044 3524 5056
rect 3516 5036 3793 5044
rect 3847 5036 4193 5044
rect 4207 5035 4253 5043
rect 4307 5036 4553 5044
rect 5007 5035 5053 5043
rect 5567 5036 5593 5044
rect 5676 5046 5684 5076
rect 5816 5046 5824 5096
rect 547 5016 833 5024
rect 1747 5016 1833 5024
rect 1847 5016 1872 5024
rect 1907 5016 2173 5024
rect 2587 5016 2653 5024
rect 3240 5024 3253 5027
rect 3236 5013 3253 5024
rect 3367 5016 3493 5024
rect 4827 5016 4913 5024
rect 4927 5016 5213 5024
rect 5227 5016 5313 5024
rect 796 4996 913 5004
rect 796 4984 804 4996
rect 927 4996 973 5004
rect 1247 4996 1533 5004
rect 2327 4996 2773 5004
rect 2967 4996 3013 5004
rect 3236 5004 3244 5013
rect 3207 4996 3244 5004
rect 3527 4996 3613 5004
rect 3687 4996 3773 5004
rect 3787 4996 3953 5004
rect 4127 4996 4413 5004
rect 4587 4996 4673 5004
rect 4687 4996 4773 5004
rect 4847 4996 4873 5004
rect 5107 4996 5133 5004
rect 5547 4996 5633 5004
rect 267 4976 804 4984
rect 1007 4976 1893 4984
rect 2387 4976 2613 4984
rect 2807 4976 3253 4984
rect 4247 4976 4333 4984
rect 4567 4976 4913 4984
rect 5087 4976 5153 4984
rect 867 4956 1333 4964
rect 1507 4956 1853 4964
rect 2407 4956 2473 4964
rect 2787 4956 3673 4964
rect 3767 4956 3793 4964
rect 4267 4956 4313 4964
rect 4407 4956 4593 4964
rect 4707 4956 4733 4964
rect 127 4936 393 4944
rect 967 4936 1073 4944
rect 1267 4936 1313 4944
rect 1667 4936 1733 4944
rect 1887 4936 2273 4944
rect 2547 4936 2693 4944
rect 3227 4936 3333 4944
rect 3387 4936 3593 4944
rect 3607 4936 3653 4944
rect 3776 4936 4293 4944
rect 3776 4927 3784 4936
rect 4427 4936 4533 4944
rect 607 4916 633 4924
rect 647 4916 1133 4924
rect 1587 4916 1813 4924
rect 2087 4916 2313 4924
rect 2547 4916 2633 4924
rect 2727 4916 2793 4924
rect 3047 4916 3093 4924
rect 3147 4916 3353 4924
rect 3367 4916 3433 4924
rect 3767 4916 3784 4927
rect 3767 4913 3780 4916
rect 4047 4916 4093 4924
rect 4287 4916 4493 4924
rect 4847 4916 5053 4924
rect 5067 4916 5153 4924
rect 5427 4916 5493 4924
rect 5607 4916 5773 4924
rect 507 4896 653 4904
rect 667 4896 753 4904
rect 1287 4896 1493 4904
rect 1887 4896 1933 4904
rect 3547 4896 3613 4904
rect 3667 4896 3733 4904
rect 4347 4896 4453 4904
rect 4527 4896 4553 4904
rect 4607 4896 4633 4904
rect 5127 4896 5253 4904
rect 147 4876 173 4884
rect 567 4876 593 4884
rect 1107 4876 1153 4884
rect 1647 4876 1773 4884
rect 1867 4876 2133 4884
rect 2887 4876 2953 4884
rect 3067 4876 3144 4884
rect 3136 4868 3144 4876
rect 3307 4876 3473 4884
rect 3927 4876 3953 4884
rect 4087 4876 4113 4884
rect 4507 4876 4693 4884
rect 4820 4884 4833 4887
rect 4816 4873 4833 4884
rect 5056 4876 5353 4884
rect 707 4856 753 4864
rect 1027 4856 1173 4864
rect 1187 4856 1373 4864
rect 1387 4856 1453 4864
rect 1536 4856 1653 4864
rect 156 4827 164 4853
rect 1536 4827 1544 4856
rect 1827 4856 2053 4864
rect 2187 4856 2233 4864
rect 2387 4857 2453 4865
rect 2507 4856 2553 4864
rect 2747 4857 2813 4865
rect 2907 4856 2933 4864
rect 2987 4856 3133 4864
rect 3247 4856 3284 4864
rect -24 4816 93 4824
rect 407 4815 473 4823
rect 527 4816 593 4824
rect 607 4815 633 4823
rect 867 4815 893 4823
rect 1087 4816 1113 4824
rect 1127 4815 1153 4823
rect 1207 4815 1273 4823
rect 1347 4815 1373 4823
rect 3276 4826 3284 4856
rect 3347 4856 3553 4864
rect 3607 4856 3624 4864
rect 3616 4827 3624 4856
rect 3827 4856 3853 4864
rect 3987 4857 4033 4865
rect 4147 4857 4173 4865
rect 4407 4856 4473 4864
rect 4536 4856 4633 4864
rect 1647 4816 1713 4824
rect 1727 4815 1793 4823
rect 2067 4815 2113 4823
rect 2247 4815 2293 4823
rect 2567 4815 2593 4823
rect 2847 4815 2873 4823
rect 3007 4816 3113 4824
rect 3127 4815 3213 4823
rect 3327 4815 3353 4823
rect 3427 4816 3573 4824
rect 3776 4824 3784 4853
rect 3707 4816 3784 4824
rect 3887 4816 4013 4824
rect 4027 4816 4133 4824
rect 4276 4824 4284 4853
rect 4536 4827 4544 4856
rect 4756 4856 4773 4864
rect 4756 4827 4764 4856
rect 4816 4864 4824 4873
rect 5056 4868 5064 4876
rect 5367 4876 5453 4884
rect 6007 4884 6020 4887
rect 6007 4873 6024 4884
rect 4796 4856 4824 4864
rect 4207 4816 4313 4824
rect 4367 4815 4393 4823
rect 4796 4826 4804 4856
rect 5007 4857 5053 4865
rect 5207 4856 5293 4864
rect 5447 4856 5544 4864
rect 5536 4844 5544 4856
rect 5587 4857 5653 4865
rect 5727 4857 5753 4865
rect 5767 4857 5813 4865
rect 5536 4836 5644 4844
rect 4847 4815 4873 4823
rect 4927 4815 4973 4823
rect 5067 4816 5273 4824
rect 5636 4826 5644 4836
rect 5367 4815 5412 4823
rect 5436 4820 5473 4824
rect 5433 4816 5473 4820
rect 5433 4807 5447 4816
rect 5856 4824 5864 4853
rect 5847 4816 5864 4824
rect 5976 4824 5984 4854
rect 6016 4827 6024 4873
rect 5947 4816 5984 4824
rect 6007 4816 6024 4827
rect 6007 4813 6020 4816
rect 307 4796 773 4804
rect 787 4796 813 4804
rect 1907 4796 1993 4804
rect 2187 4796 2333 4804
rect 2347 4796 2373 4804
rect 4567 4796 4653 4804
rect 5667 4796 5733 4804
rect 5856 4800 5953 4804
rect 5853 4796 5953 4800
rect 5853 4787 5867 4796
rect 427 4776 633 4784
rect 647 4776 733 4784
rect 1567 4776 1673 4784
rect 2227 4776 2473 4784
rect 2647 4776 2893 4784
rect 3087 4776 3873 4784
rect 3987 4776 4533 4784
rect 5567 4776 5813 4784
rect 487 4756 552 4764
rect 587 4756 673 4764
rect 687 4756 953 4764
rect 1067 4756 1453 4764
rect 3067 4756 3113 4764
rect 3267 4756 3373 4764
rect 3667 4756 3753 4764
rect 4427 4756 4473 4764
rect 5327 4756 5473 4764
rect 5687 4756 5793 4764
rect 1407 4736 1833 4744
rect 5107 4736 5193 4744
rect 1487 4716 1653 4724
rect 1767 4716 2153 4724
rect 2387 4716 2793 4724
rect 3927 4716 4053 4724
rect 4067 4716 4293 4724
rect 5027 4716 5413 4724
rect 987 4696 1193 4704
rect 1687 4696 2233 4704
rect 2907 4696 2953 4704
rect 2967 4696 3153 4704
rect 3167 4696 3533 4704
rect 967 4676 1213 4684
rect 1227 4676 1433 4684
rect 1707 4676 1873 4684
rect 1887 4676 2213 4684
rect 4807 4676 5073 4684
rect 5687 4676 5893 4684
rect 107 4656 153 4664
rect 767 4656 953 4664
rect 967 4656 1133 4664
rect 1207 4656 1753 4664
rect 1807 4656 1953 4664
rect 1967 4656 2013 4664
rect 3487 4656 3524 4664
rect 1847 4636 1933 4644
rect 2367 4636 3033 4644
rect 3207 4636 3373 4644
rect 3387 4636 3413 4644
rect 3516 4644 3524 4656
rect 3627 4656 4373 4664
rect 4387 4656 4453 4664
rect 5207 4656 5373 4664
rect 3516 4636 4533 4644
rect 4667 4636 4813 4644
rect 5187 4636 5553 4644
rect 487 4616 513 4624
rect 527 4616 853 4624
rect 3507 4616 3913 4624
rect 4147 4616 4233 4624
rect 4427 4616 4484 4624
rect 207 4596 433 4604
rect 907 4596 993 4604
rect 1007 4596 1313 4604
rect 1867 4596 2113 4604
rect 2407 4596 2733 4604
rect 2747 4596 3013 4604
rect 3427 4596 3613 4604
rect 4476 4604 4484 4616
rect 5247 4616 5313 4624
rect 4476 4596 4573 4604
rect 4587 4596 4753 4604
rect 4907 4596 4953 4604
rect 1307 4576 1493 4584
rect 1507 4576 1693 4584
rect 2327 4576 2493 4584
rect 3647 4576 3813 4584
rect 3827 4576 3873 4584
rect 4267 4576 4453 4584
rect 4627 4576 4713 4584
rect 5267 4576 5293 4584
rect 5467 4576 5513 4584
rect 5787 4576 5933 4584
rect -24 4556 13 4564
rect 607 4556 653 4564
rect 96 4544 104 4554
rect 96 4536 144 4544
rect -24 4516 113 4524
rect 136 4524 144 4536
rect 256 4527 264 4554
rect 296 4544 304 4554
rect 747 4556 853 4564
rect 876 4556 913 4564
rect 296 4536 373 4544
rect 136 4516 173 4524
rect 247 4516 264 4527
rect 876 4526 884 4556
rect 1056 4527 1064 4554
rect 1547 4556 1653 4564
rect 1927 4557 1973 4565
rect 1987 4556 2073 4564
rect 1133 4544 1147 4553
rect 1133 4540 1164 4544
rect 1136 4536 1164 4540
rect 247 4513 260 4516
rect 327 4516 453 4524
rect 467 4516 573 4524
rect 687 4515 713 4523
rect 967 4515 993 4523
rect 1056 4516 1073 4527
rect 1060 4513 1073 4516
rect 1156 4526 1164 4536
rect 1176 4524 1184 4554
rect 1376 4544 1384 4554
rect 2227 4557 2273 4565
rect 2467 4556 2513 4564
rect 2687 4557 2773 4565
rect 2927 4557 2973 4565
rect 3287 4556 3313 4564
rect 3567 4557 3673 4565
rect 3927 4557 3973 4565
rect 3987 4557 4113 4565
rect 4776 4556 4833 4564
rect 1376 4536 1893 4544
rect 4216 4544 4224 4554
rect 4216 4536 4384 4544
rect 1176 4516 1293 4524
rect 1467 4515 1513 4523
rect 1527 4516 1673 4524
rect 1727 4516 1793 4524
rect 2407 4516 2433 4524
rect 2447 4515 2473 4523
rect 2527 4515 2553 4523
rect 2747 4515 2873 4523
rect 3007 4515 3073 4523
rect 3787 4515 3813 4523
rect 3987 4515 4033 4523
rect 4307 4516 4353 4524
rect 4376 4524 4384 4536
rect 4467 4536 4564 4544
rect 4376 4516 4513 4524
rect 4556 4524 4564 4536
rect 4776 4527 4784 4556
rect 4927 4556 5053 4564
rect 5107 4556 5133 4564
rect 5187 4556 5264 4564
rect 4556 4516 4693 4524
rect 4907 4516 5073 4524
rect 5087 4516 5113 4524
rect 5256 4526 5264 4556
rect 5427 4556 5464 4564
rect 5167 4515 5213 4523
rect 5276 4524 5284 4553
rect 5276 4516 5393 4524
rect 5456 4507 5464 4556
rect 5607 4557 5633 4565
rect 5747 4556 5893 4564
rect 5587 4516 5713 4524
rect 5847 4516 5913 4524
rect 127 4496 773 4504
rect 1127 4496 1213 4504
rect 1267 4496 1573 4504
rect 1627 4496 1753 4504
rect 1767 4496 1813 4504
rect 1907 4496 2033 4504
rect 2047 4496 2153 4504
rect 3167 4496 3193 4504
rect 3287 4496 3433 4504
rect 4807 4496 4853 4504
rect 5787 4496 5813 4504
rect 287 4476 393 4484
rect 847 4476 933 4484
rect 1207 4476 1233 4484
rect 1307 4476 1793 4484
rect 2187 4476 2213 4484
rect 2847 4476 2893 4484
rect 1296 4464 1304 4473
rect 3447 4476 3513 4484
rect 4767 4476 5033 4484
rect 5767 4476 5833 4484
rect 1087 4456 1304 4464
rect 1347 4456 1873 4464
rect 1887 4456 2413 4464
rect 2687 4456 2913 4464
rect 3767 4456 3893 4464
rect 4407 4456 4553 4464
rect 4567 4456 4733 4464
rect 5247 4456 5353 4464
rect 5567 4456 5653 4464
rect 1567 4436 1864 4444
rect 167 4416 373 4424
rect 387 4416 533 4424
rect 1047 4416 1273 4424
rect 1856 4424 1864 4436
rect 2007 4436 2373 4444
rect 2607 4436 2753 4444
rect 2947 4436 3253 4444
rect 1856 4416 1913 4424
rect 3847 4416 4173 4424
rect 4527 4416 4613 4424
rect 5347 4416 5473 4424
rect 5487 4416 5753 4424
rect 4387 4396 4693 4404
rect 4967 4396 5093 4404
rect 267 4376 693 4384
rect 747 4376 873 4384
rect 887 4376 1013 4384
rect 1127 4376 1533 4384
rect 2127 4376 2533 4384
rect 2547 4376 2733 4384
rect 2747 4376 2833 4384
rect 3587 4376 3873 4384
rect 4067 4376 4253 4384
rect 4267 4376 4573 4384
rect 5007 4384 5020 4387
rect 5007 4373 5024 4384
rect 5687 4376 5733 4384
rect 2016 4356 2093 4364
rect 167 4336 253 4344
rect 427 4336 793 4344
rect 816 4336 833 4344
rect 816 4307 824 4336
rect 1067 4336 1112 4344
rect 1147 4337 1173 4345
rect 1427 4336 1493 4344
rect 1547 4336 1653 4344
rect 1727 4336 1833 4344
rect 2016 4344 2024 4356
rect 2167 4356 2373 4364
rect 2587 4356 2673 4364
rect 3307 4356 3373 4364
rect 5016 4364 5024 4373
rect 5016 4356 5133 4364
rect 5327 4356 5393 4364
rect 1847 4336 2024 4344
rect 2307 4337 2533 4345
rect 2787 4336 2893 4344
rect 2987 4336 3033 4344
rect 3087 4337 3133 4345
rect 3227 4336 3273 4344
rect 3527 4337 3593 4345
rect 3647 4336 3833 4344
rect 4327 4336 4393 4344
rect 3336 4324 3344 4334
rect 2876 4316 3344 4324
rect 27 4296 133 4304
rect 287 4296 393 4304
rect 447 4295 473 4303
rect 627 4295 673 4303
rect 907 4296 1033 4304
rect 1127 4295 1193 4303
rect 1787 4295 1873 4303
rect 2307 4295 2433 4303
rect 2876 4304 2884 4316
rect 2767 4296 2884 4304
rect 2927 4295 2973 4303
rect 3067 4296 3273 4304
rect 3287 4295 3353 4303
rect 3407 4296 3433 4304
rect 3787 4295 3853 4303
rect 3916 4304 3924 4334
rect 4407 4336 4433 4344
rect 4627 4337 4653 4345
rect 5187 4336 5253 4344
rect 5507 4336 5633 4344
rect 5156 4316 5233 4324
rect 3916 4296 4033 4304
rect 4107 4296 4153 4304
rect 4207 4295 4253 4303
rect 4347 4296 4373 4304
rect 5156 4306 5164 4316
rect 4727 4296 4933 4304
rect 5436 4304 5444 4333
rect 5676 4324 5684 4334
rect 5727 4336 5793 4344
rect 5676 4320 5704 4324
rect 5676 4316 5707 4320
rect 5327 4296 5444 4304
rect 5693 4307 5707 4316
rect 5796 4304 5804 4334
rect 5887 4336 5933 4344
rect 5996 4307 6004 4333
rect 5796 4296 5913 4304
rect 807 4276 853 4284
rect 1367 4276 1513 4284
rect 1887 4276 1973 4284
rect 2127 4276 2413 4284
rect 2847 4276 3193 4284
rect 3207 4276 3493 4284
rect 3907 4276 3993 4284
rect 4527 4276 4553 4284
rect 5107 4276 5193 4284
rect 27 4256 193 4264
rect 2087 4256 2173 4264
rect 2227 4256 2593 4264
rect 2727 4256 2913 4264
rect 827 4236 1173 4244
rect 1187 4236 1233 4244
rect 1247 4236 1273 4244
rect 1387 4236 1473 4244
rect 1487 4236 1813 4244
rect 2567 4236 2753 4244
rect 2916 4244 2924 4253
rect 5487 4256 5553 4264
rect 5767 4256 5953 4264
rect 2916 4236 3233 4244
rect 3307 4236 4333 4244
rect 4827 4236 4853 4244
rect 5667 4236 5813 4244
rect 107 4216 233 4224
rect 247 4216 1333 4224
rect 1347 4216 2333 4224
rect 3087 4216 3393 4224
rect 4327 4216 4493 4224
rect 1147 4196 1373 4204
rect 1767 4196 2153 4204
rect 2507 4196 2713 4204
rect 4187 4196 5313 4204
rect 5327 4196 5493 4204
rect 5607 4196 5713 4204
rect 787 4176 1113 4184
rect 1407 4176 1673 4184
rect 2187 4176 2633 4184
rect 3147 4176 3333 4184
rect 3347 4176 3533 4184
rect 3547 4176 3993 4184
rect 4307 4176 4833 4184
rect 4847 4176 5053 4184
rect 1167 4156 1313 4164
rect 4296 4164 4304 4173
rect 2807 4156 4304 4164
rect 4607 4156 4653 4164
rect 887 4136 1413 4144
rect 2427 4136 3133 4144
rect 3527 4136 3572 4144
rect 3607 4136 3693 4144
rect 4227 4136 4793 4144
rect 5407 4136 5773 4144
rect 1867 4116 2293 4124
rect 3507 4116 3793 4124
rect 3807 4116 3893 4124
rect 3947 4116 5353 4124
rect 5367 4116 5413 4124
rect 5427 4116 5573 4124
rect -24 4096 13 4104
rect 507 4096 553 4104
rect 1227 4096 2364 4104
rect 2356 4087 2364 4096
rect 3627 4096 3733 4104
rect 4127 4096 4293 4104
rect 367 4076 393 4084
rect 647 4076 824 4084
rect 816 4064 824 4076
rect 867 4076 913 4084
rect 1047 4076 1113 4084
rect 1247 4076 1393 4084
rect 1627 4076 1733 4084
rect 1947 4076 2133 4084
rect 2367 4076 2453 4084
rect 2527 4076 2553 4084
rect 2567 4076 2613 4084
rect 2667 4076 2753 4084
rect 2767 4076 3173 4084
rect 3487 4076 3593 4084
rect 3687 4076 3833 4084
rect 4407 4076 4713 4084
rect 4727 4076 4913 4084
rect 4927 4076 4973 4084
rect 5067 4076 5193 4084
rect 5207 4076 5273 4084
rect 5647 4076 5693 4084
rect 5867 4076 5933 4084
rect 816 4056 993 4064
rect 2047 4056 2213 4064
rect 3627 4056 3693 4064
rect 3707 4056 3853 4064
rect 3907 4056 4033 4064
rect 4087 4056 4133 4064
rect 5627 4056 5733 4064
rect -24 4036 93 4044
rect 267 4036 293 4044
rect 447 4036 493 4044
rect 587 4036 613 4044
rect 667 4037 693 4045
rect 796 4024 804 4034
rect 887 4036 944 4044
rect 747 4016 804 4024
rect 936 4006 944 4036
rect 967 4036 1073 4044
rect 1287 4036 1433 4044
rect 1447 4036 1513 4044
rect 1607 4037 1653 4045
rect 2007 4036 2173 4044
rect 2196 4036 2293 4044
rect 1696 4016 1753 4024
rect -24 3996 473 4004
rect 487 3995 573 4003
rect 1167 3996 1213 4004
rect 1407 3995 1433 4003
rect 1696 4004 1704 4016
rect 1547 3996 1704 4004
rect 1876 4004 1884 4033
rect 2176 4024 2184 4034
rect 2136 4016 2184 4024
rect 2136 4007 2144 4016
rect 1807 3996 1884 4004
rect 1927 3996 1973 4004
rect 2127 3996 2144 4007
rect 2127 3993 2140 3996
rect 2196 4004 2204 4036
rect 2587 4037 2673 4045
rect 2887 4036 2973 4044
rect 3027 4037 3053 4045
rect 3107 4037 3133 4045
rect 3187 4037 3233 4045
rect 3307 4036 3453 4044
rect 2167 3996 2204 4004
rect 2276 4000 2313 4004
rect 2273 3996 2313 4000
rect 2273 3987 2287 3996
rect 2447 3996 2513 4004
rect 2716 3987 2724 4034
rect 3927 4036 3973 4044
rect 4427 4037 4453 4045
rect 2747 3996 2813 4004
rect 2827 3996 2853 4004
rect 3047 3996 3073 4004
rect 3447 3996 3493 4004
rect 3576 4004 3584 4033
rect 4376 4024 4384 4034
rect 4767 4036 4873 4044
rect 4887 4037 4953 4045
rect 5107 4037 5133 4045
rect 5247 4037 5293 4045
rect 5307 4036 5393 4044
rect 4376 4016 4453 4024
rect 4516 4024 4524 4034
rect 4467 4016 4524 4024
rect 3576 3996 3652 4004
rect 3687 3995 3713 4003
rect 3847 3995 4053 4003
rect 4107 3996 4153 4004
rect 4247 3996 4353 4004
rect 4667 3996 4693 4004
rect 4807 3996 4853 4004
rect 4967 3996 5033 4004
rect 5087 3995 5173 4003
rect 5507 3995 5533 4003
rect 5696 4004 5704 4034
rect 5767 4036 5793 4044
rect 5907 4036 5953 4044
rect 5667 3996 5704 4004
rect 5856 3987 5864 4034
rect 647 3976 773 3984
rect 1007 3976 1053 3984
rect 1507 3976 1593 3984
rect 1607 3976 1873 3984
rect 1887 3976 2133 3984
rect 2207 3976 2233 3984
rect 3227 3976 3393 3984
rect 3607 3976 3793 3984
rect 5907 3976 5993 3984
rect 807 3956 853 3964
rect 1187 3956 1253 3964
rect 1847 3956 1953 3964
rect 2267 3956 2293 3964
rect 3367 3956 3553 3964
rect 4467 3956 4713 3964
rect 4727 3956 5213 3964
rect 5267 3956 5413 3964
rect 5427 3956 5673 3964
rect 567 3936 633 3944
rect 947 3936 1093 3944
rect 1687 3936 1933 3944
rect 1947 3936 2013 3944
rect 2607 3936 2993 3944
rect 3167 3936 3273 3944
rect 3767 3936 3893 3944
rect 3907 3936 4553 3944
rect 4747 3936 4893 3944
rect 4907 3936 5373 3944
rect 5727 3936 5873 3944
rect 187 3916 253 3924
rect 1027 3916 1133 3924
rect 1647 3916 1693 3924
rect 3387 3916 3813 3924
rect 5247 3916 5293 3924
rect 5407 3916 5473 3924
rect 527 3896 693 3904
rect 707 3896 1273 3904
rect 2147 3896 2553 3904
rect 2567 3896 2973 3904
rect 3287 3896 3493 3904
rect 4407 3896 4533 3904
rect 5087 3896 5133 3904
rect 5147 3896 5333 3904
rect 5587 3896 5633 3904
rect 267 3876 553 3884
rect 867 3876 893 3884
rect 1647 3876 1893 3884
rect 1987 3876 2093 3884
rect 3687 3876 3793 3884
rect 5527 3876 5793 3884
rect 5847 3876 5993 3884
rect 147 3856 1053 3864
rect 2267 3856 2573 3864
rect 3867 3856 4033 3864
rect 4307 3856 4393 3864
rect 4547 3856 4873 3864
rect 4887 3856 4933 3864
rect 4947 3856 5153 3864
rect 5567 3856 5633 3864
rect 5687 3856 5713 3864
rect 447 3836 473 3844
rect 527 3836 733 3844
rect 747 3836 813 3844
rect 2256 3844 2264 3853
rect 1967 3836 2264 3844
rect 2327 3836 2433 3844
rect 3567 3836 3713 3844
rect 3767 3836 3833 3844
rect 5267 3836 5313 3844
rect 907 3817 933 3825
rect 1527 3817 1533 3825
rect 1547 3817 1553 3825
rect 1707 3817 1773 3825
rect 1827 3816 1913 3824
rect 1927 3816 2033 3824
rect 2627 3817 2773 3825
rect 2887 3817 2913 3825
rect 2987 3817 3153 3825
rect 3167 3816 3353 3824
rect 3407 3817 3433 3825
rect 3607 3816 3693 3824
rect 3867 3824 3880 3827
rect 3867 3813 3884 3824
rect 4016 3816 4073 3824
rect 1427 3796 1504 3804
rect -24 3776 93 3784
rect 367 3776 393 3784
rect 687 3776 873 3784
rect 947 3776 1013 3784
rect 1387 3776 1433 3784
rect 1496 3784 1504 3796
rect 2236 3796 2333 3804
rect 2236 3786 2244 3796
rect 3533 3804 3547 3813
rect 3516 3800 3547 3804
rect 3516 3796 3544 3800
rect 1496 3776 1613 3784
rect 1847 3776 1993 3784
rect 2007 3776 2093 3784
rect 2467 3775 2653 3783
rect 2747 3776 2773 3784
rect 2907 3776 3013 3784
rect 3067 3775 3133 3783
rect 3516 3784 3524 3796
rect 3467 3776 3524 3784
rect 3547 3775 3613 3783
rect 3627 3776 3693 3784
rect 3876 3786 3884 3813
rect 3956 3787 3964 3813
rect 4016 3787 4024 3816
rect 4167 3817 4213 3825
rect 4327 3816 4353 3824
rect 4367 3817 4493 3825
rect 4667 3816 4753 3824
rect 4807 3816 5013 3824
rect 5107 3816 5133 3824
rect 5427 3817 5473 3825
rect 5653 3824 5667 3833
rect 5527 3816 5644 3824
rect 5653 3820 5684 3824
rect 5656 3816 5684 3820
rect 3787 3775 3813 3783
rect 3836 3776 3873 3784
rect 1287 3756 1493 3764
rect 1647 3756 1733 3764
rect 1796 3764 1804 3772
rect 1796 3756 1873 3764
rect 2047 3756 2273 3764
rect 2367 3756 2813 3764
rect 2927 3756 3173 3764
rect 3836 3764 3844 3776
rect 4107 3776 4153 3784
rect 4507 3776 4573 3784
rect 4747 3776 4853 3784
rect 4947 3775 5033 3783
rect 5176 3784 5184 3814
rect 5176 3776 5213 3784
rect 5267 3775 5313 3783
rect 5507 3775 5573 3783
rect 5636 3784 5644 3816
rect 5676 3804 5684 3816
rect 5767 3816 5813 3824
rect 5676 3796 5704 3804
rect 5696 3786 5704 3796
rect 5636 3776 5653 3784
rect 5856 3784 5864 3814
rect 5787 3776 5864 3784
rect 3636 3756 3844 3764
rect 1667 3736 1833 3744
rect 2147 3736 2564 3744
rect 2556 3727 2564 3736
rect 2587 3736 2793 3744
rect 2847 3736 3093 3744
rect 3147 3736 3333 3744
rect 3347 3736 3373 3744
rect 3636 3744 3644 3756
rect 4007 3756 4333 3764
rect 4487 3756 4693 3764
rect 5256 3764 5264 3772
rect 5167 3756 5264 3764
rect 5847 3756 5993 3764
rect 3507 3736 3644 3744
rect 3667 3736 3733 3744
rect 3747 3736 3773 3744
rect 3827 3736 4233 3744
rect 5007 3736 5093 3744
rect 5227 3736 5364 3744
rect 5356 3727 5364 3736
rect 5587 3736 5793 3744
rect 287 3716 493 3724
rect 1947 3716 2053 3724
rect 2167 3716 2493 3724
rect 2567 3716 2893 3724
rect 3127 3716 3553 3724
rect 5067 3716 5193 3724
rect 5367 3716 5553 3724
rect 1167 3696 1613 3704
rect 1627 3696 3273 3704
rect 3287 3696 3393 3704
rect 3407 3696 3613 3704
rect 3707 3696 4193 3704
rect 4547 3696 4573 3704
rect 4827 3696 5213 3704
rect 5607 3696 5953 3704
rect 2107 3676 2352 3684
rect 2387 3676 2593 3684
rect 2827 3676 3213 3684
rect 4907 3676 5693 3684
rect 5787 3676 5833 3684
rect 607 3656 733 3664
rect 747 3656 1233 3664
rect 1247 3656 1333 3664
rect 2707 3656 3453 3664
rect 4347 3656 4573 3664
rect 4647 3656 4673 3664
rect 2607 3636 3113 3644
rect 3187 3636 3373 3644
rect 4287 3636 4793 3644
rect 5087 3636 5753 3644
rect 1567 3616 1733 3624
rect 2087 3616 2573 3624
rect 2887 3616 2973 3624
rect 3047 3616 3433 3624
rect 3667 3616 3913 3624
rect 5307 3616 5553 3624
rect 5567 3616 5593 3624
rect 1527 3596 2013 3604
rect 2987 3596 3453 3604
rect 3647 3596 4013 3604
rect 4207 3596 4373 3604
rect 5887 3596 5933 3604
rect 827 3576 893 3584
rect 907 3576 1073 3584
rect 3487 3576 3592 3584
rect 3627 3576 3853 3584
rect 4127 3576 4653 3584
rect 576 3556 753 3564
rect 576 3544 584 3556
rect 1927 3556 2393 3564
rect 3067 3556 3253 3564
rect 3267 3556 3353 3564
rect 3467 3556 3633 3564
rect 3927 3556 4313 3564
rect 4327 3556 4413 3564
rect 4787 3556 5193 3564
rect 5627 3556 5713 3564
rect 5727 3556 5913 3564
rect 547 3536 584 3544
rect 827 3536 1193 3544
rect 1307 3536 1453 3544
rect 1467 3536 1573 3544
rect 2447 3536 2633 3544
rect 3247 3536 3893 3544
rect 4427 3536 4453 3544
rect 4667 3536 4693 3544
rect 4707 3536 4973 3544
rect 5767 3536 5853 3544
rect -24 3516 93 3524
rect 307 3516 344 3524
rect 336 3504 344 3516
rect 367 3516 593 3524
rect 947 3517 973 3525
rect 987 3516 1033 3524
rect 1747 3516 1793 3524
rect 1867 3516 1973 3524
rect 1987 3516 2153 3524
rect 2247 3517 2293 3525
rect 2347 3517 2373 3525
rect 2487 3517 2532 3525
rect 2567 3517 2593 3525
rect 2727 3517 2773 3525
rect 2787 3516 2933 3524
rect 336 3496 424 3504
rect 416 3486 424 3496
rect 2436 3487 2444 3514
rect 3036 3516 3093 3524
rect 147 3476 173 3484
rect 787 3475 813 3483
rect 927 3476 1053 3484
rect 1107 3476 1213 3484
rect 1587 3475 1633 3483
rect 1647 3476 1693 3484
rect 1807 3475 1833 3483
rect 2047 3475 2073 3483
rect 2427 3476 2444 3487
rect 2427 3473 2440 3476
rect 2547 3475 2613 3483
rect 2667 3476 2713 3484
rect 2767 3476 2913 3484
rect 2996 3484 3004 3513
rect 3036 3507 3044 3516
rect 3147 3516 3193 3524
rect 3336 3516 3413 3524
rect 3027 3496 3044 3507
rect 3027 3493 3040 3496
rect 3336 3487 3344 3516
rect 3607 3516 3693 3524
rect 3827 3517 3993 3525
rect 4107 3517 4153 3525
rect 4307 3517 4353 3525
rect 4456 3516 4493 3524
rect 2967 3476 3004 3484
rect 3167 3476 3273 3484
rect 3487 3476 3673 3484
rect 1487 3456 1993 3464
rect 2007 3456 2233 3464
rect 2247 3456 2333 3464
rect 2867 3456 3053 3464
rect 3367 3456 3544 3464
rect 747 3436 873 3444
rect 1667 3436 1713 3444
rect 1727 3436 1913 3444
rect 2327 3436 2453 3444
rect 2467 3436 2553 3444
rect 2807 3436 3033 3444
rect 3536 3444 3544 3456
rect 3567 3456 3613 3464
rect 3776 3464 3784 3513
rect 4036 3504 4044 3514
rect 4456 3504 4464 3516
rect 4507 3516 4593 3524
rect 4827 3517 4853 3525
rect 4867 3516 4933 3524
rect 4987 3516 5153 3524
rect 5236 3504 5244 3533
rect 5347 3517 5373 3525
rect 5387 3516 5453 3524
rect 5547 3517 5613 3525
rect 3807 3496 4464 3504
rect 5216 3496 5244 3504
rect 5216 3487 5224 3496
rect 3887 3476 4213 3484
rect 4487 3476 4753 3484
rect 4767 3476 4893 3484
rect 5007 3476 5052 3484
rect 5087 3475 5133 3483
rect 5207 3476 5224 3487
rect 5207 3473 5220 3476
rect 5247 3476 5273 3484
rect 5496 3484 5504 3514
rect 5736 3487 5744 3513
rect 5833 3504 5847 3513
rect 5816 3500 5847 3504
rect 5816 3496 5844 3500
rect 5327 3476 5593 3484
rect 5816 3486 5824 3496
rect 5867 3476 5933 3484
rect 3707 3456 3784 3464
rect 3987 3456 4093 3464
rect 5076 3464 5084 3472
rect 5956 3467 5964 3514
rect 5996 3487 6004 3513
rect 4967 3456 5084 3464
rect 5187 3456 5373 3464
rect 5487 3456 5553 3464
rect 3536 3436 3573 3444
rect 3687 3436 3713 3444
rect 3727 3436 3813 3444
rect 4027 3436 4313 3444
rect 4687 3436 4753 3444
rect 6036 3444 6044 3524
rect 5656 3436 6044 3444
rect 2027 3416 2533 3424
rect 2887 3416 2993 3424
rect 3387 3416 4173 3424
rect 5656 3424 5664 3436
rect 4587 3416 5664 3424
rect 5847 3416 5973 3424
rect 2187 3396 2853 3404
rect 3327 3396 4413 3404
rect 4427 3396 4633 3404
rect 5547 3396 5853 3404
rect 247 3376 593 3384
rect 647 3376 1193 3384
rect 2247 3376 2613 3384
rect 3207 3376 3333 3384
rect 3687 3376 3733 3384
rect 4707 3376 4733 3384
rect 4867 3376 5033 3384
rect 5047 3376 5433 3384
rect 947 3356 973 3364
rect 1367 3356 1793 3364
rect 1807 3356 1873 3364
rect 2367 3356 2392 3364
rect 2427 3356 2733 3364
rect 2796 3356 2893 3364
rect 27 3336 433 3344
rect 447 3336 533 3344
rect 547 3336 673 3344
rect 687 3336 1313 3344
rect 2387 3336 2453 3344
rect 2796 3344 2804 3356
rect 2967 3356 3033 3364
rect 4167 3356 4213 3364
rect 5327 3356 5673 3364
rect 2507 3336 2804 3344
rect 2827 3336 2873 3344
rect 2927 3336 3013 3344
rect 3027 3336 3133 3344
rect 3147 3336 3192 3344
rect 3227 3336 3313 3344
rect 3547 3336 3633 3344
rect 4107 3336 4473 3344
rect 4707 3336 4953 3344
rect 2167 3316 2213 3324
rect 2287 3316 2473 3324
rect 2707 3316 2753 3324
rect 2907 3316 3113 3324
rect 3127 3316 3413 3324
rect 3627 3316 4044 3324
rect -24 3296 73 3304
rect 147 3296 173 3304
rect 507 3296 613 3304
rect 727 3296 773 3304
rect 787 3296 813 3304
rect 1447 3297 1493 3305
rect 1587 3296 1633 3304
rect 976 3284 984 3294
rect 1687 3296 1833 3304
rect 1887 3296 2233 3304
rect 2507 3297 2573 3305
rect 2627 3296 2813 3304
rect 2987 3296 3073 3304
rect 3187 3297 3253 3305
rect 3347 3297 3433 3305
rect 3487 3296 3513 3304
rect 3596 3296 3733 3304
rect 976 3276 1033 3284
rect 2087 3276 2953 3284
rect 3576 3284 3584 3294
rect 3527 3276 3584 3284
rect -24 3256 13 3264
rect 267 3256 293 3264
rect 567 3255 593 3263
rect 607 3256 653 3264
rect 847 3256 953 3264
rect 1267 3255 1293 3263
rect 1507 3256 1553 3264
rect 1807 3256 1853 3264
rect 2047 3256 2253 3264
rect 2307 3255 2333 3263
rect 2447 3256 2493 3264
rect 2536 3256 2633 3264
rect 987 3236 1053 3244
rect 1327 3236 1393 3244
rect 1407 3236 1533 3244
rect 1547 3236 1593 3244
rect 2536 3244 2544 3256
rect 2767 3256 2792 3264
rect 2827 3255 2853 3263
rect 3107 3255 3133 3263
rect 3467 3256 3493 3264
rect 3507 3256 3553 3264
rect 3596 3264 3604 3296
rect 3787 3296 3993 3304
rect 4036 3304 4044 3316
rect 4287 3316 4373 3324
rect 4627 3316 4653 3324
rect 5087 3316 5133 3324
rect 4036 3296 4053 3304
rect 3576 3260 3604 3264
rect 3573 3256 3604 3260
rect 2487 3236 2544 3244
rect 3573 3247 3587 3256
rect 3807 3255 3833 3263
rect 4036 3264 4044 3296
rect 4267 3296 4424 3304
rect 4416 3287 4424 3296
rect 4467 3296 4513 3304
rect 4720 3304 4733 3307
rect 4716 3293 4733 3304
rect 4827 3297 4973 3305
rect 4987 3296 5232 3304
rect 5267 3296 5313 3304
rect 5407 3297 5453 3305
rect 5587 3297 5633 3305
rect 5727 3297 5773 3305
rect 4416 3276 4433 3287
rect 4420 3273 4433 3276
rect 4487 3276 4613 3284
rect 4716 3266 4724 3293
rect 3927 3256 4044 3264
rect 4167 3255 4193 3263
rect 4967 3256 5153 3264
rect 5247 3255 5293 3263
rect 5307 3256 5433 3264
rect 5496 3264 5504 3294
rect 5896 3296 5913 3304
rect 5816 3267 5824 3293
rect 5496 3256 5533 3264
rect 5896 3247 5904 3296
rect 5956 3263 5964 3313
rect 5947 3255 5973 3263
rect 3647 3236 3693 3244
rect 3707 3236 3753 3244
rect 3987 3236 4073 3244
rect 5016 3236 5313 3244
rect 5016 3227 5024 3236
rect 5667 3236 5793 3244
rect 27 3216 513 3224
rect 1647 3216 1893 3224
rect 1907 3216 1993 3224
rect 2007 3216 2073 3224
rect 2147 3216 2193 3224
rect 2367 3216 2393 3224
rect 2407 3216 2553 3224
rect 2647 3216 2893 3224
rect 2907 3216 3173 3224
rect 3787 3216 3993 3224
rect 4447 3216 5013 3224
rect 5187 3216 5213 3224
rect 5796 3224 5804 3233
rect 5796 3216 5873 3224
rect 2767 3196 2833 3204
rect 2847 3196 3053 3204
rect 3167 3196 3633 3204
rect 3847 3196 4333 3204
rect 5527 3196 5893 3204
rect 1867 3176 2413 3184
rect 2607 3176 2693 3184
rect 3367 3176 3393 3184
rect 3407 3176 3673 3184
rect 3687 3176 3713 3184
rect 3827 3176 4393 3184
rect 4407 3176 4493 3184
rect 5047 3176 5073 3184
rect 5516 3184 5524 3193
rect 5087 3176 5524 3184
rect 5567 3176 5813 3184
rect 307 3156 1453 3164
rect 1467 3156 1653 3164
rect 2807 3156 2993 3164
rect 3767 3156 4233 3164
rect 1347 3136 1573 3144
rect 2027 3136 2213 3144
rect 2227 3136 3153 3144
rect 5347 3136 5373 3144
rect 627 3116 713 3124
rect 727 3116 1033 3124
rect 2547 3116 2753 3124
rect 2827 3116 3173 3124
rect 3187 3116 3293 3124
rect 3347 3116 4253 3124
rect 4267 3116 4453 3124
rect 5507 3116 5733 3124
rect 1547 3096 1933 3104
rect 1947 3096 2233 3104
rect 2287 3096 2433 3104
rect 5487 3096 5993 3104
rect 387 3076 513 3084
rect 527 3076 613 3084
rect 627 3076 1133 3084
rect 1407 3076 1493 3084
rect 1927 3076 2033 3084
rect 3147 3076 3333 3084
rect 5367 3076 5613 3084
rect -24 3056 293 3064
rect 1747 3056 1793 3064
rect 2536 3056 2633 3064
rect 2536 3047 2544 3056
rect 2967 3056 3073 3064
rect 3087 3056 3373 3064
rect 4007 3056 4133 3064
rect 4247 3056 4313 3064
rect 5807 3056 5993 3064
rect 787 3036 833 3044
rect 847 3036 1073 3044
rect 1367 3036 1413 3044
rect 2327 3036 2533 3044
rect 2747 3036 2873 3044
rect 2927 3036 3153 3044
rect 3167 3036 3593 3044
rect 4727 3036 4793 3044
rect 4967 3036 4993 3044
rect 5127 3036 5153 3044
rect 5167 3036 5213 3044
rect 5227 3036 5533 3044
rect 5667 3036 5773 3044
rect 447 3016 553 3024
rect 1667 3016 1973 3024
rect 2587 3016 2693 3024
rect 4187 3016 4292 3024
rect 4327 3016 4413 3024
rect 4467 3013 4473 3027
rect 5016 3016 5093 3024
rect -24 2996 113 3004
rect 787 2996 893 3004
rect 1247 2996 1453 3004
rect 1767 2997 1893 3005
rect 1987 2996 2053 3004
rect -24 2956 13 2964
rect 167 2956 193 2964
rect 727 2955 753 2963
rect 847 2955 873 2963
rect 936 2944 944 2994
rect 2067 2996 2093 3004
rect 2147 2997 2173 3005
rect 2347 2997 2373 3005
rect 2616 2996 2673 3004
rect 1407 2955 1473 2963
rect 1647 2955 1693 2963
rect 1907 2956 1933 2964
rect 2327 2956 2393 2964
rect 2616 2964 2624 2996
rect 2887 2996 3033 3004
rect 3167 2996 3204 3004
rect 2836 2967 2844 2993
rect 2607 2956 2624 2964
rect 2647 2955 2713 2963
rect 2867 2956 3013 2964
rect 3067 2956 3113 2964
rect 3196 2966 3204 2996
rect 3287 2997 3333 3005
rect 3447 2996 3533 3004
rect 3687 2996 3733 3004
rect 3747 2997 3773 3005
rect 3967 2996 4033 3004
rect 4147 2997 4393 3005
rect 936 2936 993 2944
rect 1007 2936 1093 2944
rect 1107 2936 1213 2944
rect 927 2916 973 2924
rect 1067 2916 1133 2924
rect 2127 2916 2613 2924
rect 2627 2916 2833 2924
rect 3216 2924 3224 2993
rect 4516 2984 4524 2994
rect 4567 2996 4633 3004
rect 4687 2996 4793 3004
rect 5016 3004 5024 3016
rect 5427 3016 5613 3024
rect 5627 3016 5713 3024
rect 4967 2996 5024 3004
rect 5467 2996 5573 3004
rect 5747 2996 5893 3004
rect 4427 2976 4524 2984
rect 4796 2984 4804 2994
rect 4796 2976 4873 2984
rect 4976 2976 5033 2984
rect 3247 2956 3353 2964
rect 3587 2955 3613 2963
rect 3667 2960 3704 2964
rect 3667 2956 3707 2960
rect 3693 2947 3707 2956
rect 3807 2956 4073 2964
rect 4976 2966 4984 2976
rect 4167 2955 4193 2963
rect 5287 2956 5393 2964
rect 5527 2956 5553 2964
rect 5687 2956 5713 2964
rect 4047 2936 4293 2944
rect 4407 2936 4453 2944
rect 4727 2936 4813 2944
rect 5736 2944 5744 2994
rect 5867 2955 5913 2963
rect 5976 2964 5984 2993
rect 5967 2956 5984 2964
rect 5736 2936 5773 2944
rect 3127 2916 3224 2924
rect 3747 2916 3813 2924
rect 3947 2916 4033 2924
rect 4347 2916 4493 2924
rect 4507 2916 4673 2924
rect 5187 2916 5233 2924
rect 5367 2916 5393 2924
rect 5407 2916 5433 2924
rect 5447 2916 5513 2924
rect 5527 2916 5593 2924
rect 1347 2896 1453 2904
rect 1467 2896 1513 2904
rect 1527 2896 1933 2904
rect 5767 2896 5853 2904
rect 2447 2876 2653 2884
rect 2767 2876 3113 2884
rect 3207 2876 3293 2884
rect 3407 2876 3673 2884
rect 3687 2876 3913 2884
rect 4667 2876 4833 2884
rect 4847 2876 4893 2884
rect 4907 2876 5173 2884
rect 5627 2876 5733 2884
rect 27 2856 1333 2864
rect 1967 2856 2553 2864
rect 2567 2856 2673 2864
rect 2827 2856 2913 2864
rect 4247 2856 4353 2864
rect 287 2836 433 2844
rect 1807 2836 2693 2844
rect 2707 2836 2793 2844
rect 3867 2836 4313 2844
rect 5487 2836 5653 2844
rect 5747 2836 5833 2844
rect -24 2816 13 2824
rect 1787 2816 1853 2824
rect 1947 2816 2133 2824
rect 2147 2816 2173 2824
rect 2267 2816 2473 2824
rect 2487 2816 2553 2824
rect 3067 2816 3233 2824
rect 3247 2816 3273 2824
rect 4547 2816 4633 2824
rect 4647 2816 4953 2824
rect 427 2796 693 2804
rect 1767 2796 1913 2804
rect 2747 2796 2853 2804
rect 2907 2796 3004 2804
rect -24 2776 73 2784
rect 147 2776 453 2784
rect 1407 2776 1533 2784
rect 1707 2777 1753 2785
rect 2227 2777 2293 2785
rect 2447 2776 2513 2784
rect 2996 2784 3004 2796
rect 3027 2796 3264 2804
rect 2996 2776 3044 2784
rect 2876 2764 2884 2774
rect 2776 2756 2884 2764
rect -24 2724 -16 2744
rect 27 2736 373 2744
rect 967 2736 1013 2744
rect 1267 2735 1293 2743
rect 1307 2736 1513 2744
rect 1887 2735 2073 2743
rect 2087 2735 2093 2743
rect 2776 2744 2784 2756
rect 3036 2746 3044 2776
rect 3256 2764 3264 2796
rect 3727 2796 3793 2804
rect 3907 2796 3953 2804
rect 4267 2796 4293 2804
rect 5367 2796 5433 2804
rect 3367 2776 3653 2784
rect 4087 2776 4153 2784
rect 4167 2777 4233 2785
rect 4256 2776 4353 2784
rect 3127 2756 3224 2764
rect 3256 2756 3384 2764
rect 3216 2746 3224 2756
rect 3376 2746 3384 2756
rect 4256 2746 4264 2776
rect 4507 2776 4564 2784
rect 4556 2747 4564 2776
rect 4727 2776 4793 2784
rect 4816 2764 4824 2793
rect 5007 2776 5073 2784
rect 5087 2777 5133 2785
rect 5307 2777 5473 2785
rect 5687 2777 5733 2785
rect 5887 2777 5973 2785
rect 4696 2756 4824 2764
rect 2727 2736 2784 2744
rect 2807 2735 2853 2743
rect 3287 2735 3333 2743
rect 3687 2735 3713 2743
rect 3787 2735 3873 2743
rect 4107 2736 4213 2744
rect 4387 2736 4413 2744
rect 4696 2746 4704 2756
rect 4816 2746 4824 2756
rect 4867 2736 4893 2744
rect 5027 2736 5153 2744
rect 5287 2736 5353 2744
rect 5576 2744 5584 2774
rect 5487 2736 5584 2744
rect -24 2716 233 2724
rect 587 2716 753 2724
rect 2327 2716 2413 2724
rect 2527 2716 2673 2724
rect 3427 2716 3593 2724
rect 3667 2716 3733 2724
rect 4067 2716 4253 2724
rect 4487 2716 4593 2724
rect 4747 2716 4793 2724
rect 5427 2716 5533 2724
rect 5687 2716 5733 2724
rect 5827 2716 5893 2724
rect 813 2704 827 2713
rect 813 2700 1733 2704
rect 816 2696 1733 2700
rect 2967 2696 3153 2704
rect 3387 2696 3773 2704
rect 4827 2696 4973 2704
rect 5247 2696 5273 2704
rect 5367 2696 5593 2704
rect 647 2676 973 2684
rect 987 2676 1133 2684
rect 2067 2676 2253 2684
rect 2687 2676 2893 2684
rect 2907 2676 3053 2684
rect 3827 2676 3893 2684
rect 4267 2676 4373 2684
rect 5616 2676 5893 2684
rect 5616 2667 5624 2676
rect 1387 2656 1773 2664
rect 1787 2656 1933 2664
rect 1987 2656 2153 2664
rect 2167 2656 2453 2664
rect 2467 2656 2693 2664
rect 2987 2656 3073 2664
rect 3607 2656 3773 2664
rect 4167 2656 4233 2664
rect 4247 2656 4593 2664
rect 5127 2656 5313 2664
rect 5467 2656 5613 2664
rect 3507 2636 3573 2644
rect 5347 2636 5713 2644
rect 5727 2636 5953 2644
rect 607 2616 873 2624
rect 2367 2616 2493 2624
rect 2547 2616 2933 2624
rect 3007 2616 3413 2624
rect 4227 2616 4333 2624
rect 4347 2616 4553 2624
rect 4607 2616 4753 2624
rect 5087 2616 5113 2624
rect 1647 2596 2113 2604
rect 2187 2596 2953 2604
rect 3527 2596 3553 2604
rect 3607 2596 3804 2604
rect 3796 2587 3804 2596
rect 4987 2596 5013 2604
rect 2487 2576 2533 2584
rect 3427 2576 3633 2584
rect 3807 2576 4053 2584
rect 4427 2576 4493 2584
rect 4567 2576 4713 2584
rect 5527 2576 5593 2584
rect 5767 2576 5993 2584
rect -24 2556 1073 2564
rect 1467 2556 1653 2564
rect 1667 2556 1693 2564
rect 2267 2556 2393 2564
rect 2567 2556 2704 2564
rect 727 2536 1533 2544
rect 2127 2536 2473 2544
rect 2536 2536 2653 2544
rect -24 2516 93 2524
rect 367 2516 513 2524
rect 527 2516 593 2524
rect 1327 2516 1373 2524
rect 1787 2516 1893 2524
rect 2536 2524 2544 2536
rect 2696 2544 2704 2556
rect 2747 2556 3033 2564
rect 3307 2556 3733 2564
rect 3847 2556 4213 2564
rect 4287 2556 4413 2564
rect 2696 2536 3133 2544
rect 3407 2536 3593 2544
rect 3947 2536 4633 2544
rect 4647 2536 4713 2544
rect 4727 2536 4873 2544
rect 4927 2536 4953 2544
rect 4967 2536 5033 2544
rect 2507 2516 2544 2524
rect 3987 2516 4153 2524
rect 5527 2516 5853 2524
rect -24 2496 713 2504
rect -24 2476 -16 2496
rect 1087 2496 1133 2504
rect 1747 2496 2193 2504
rect 2207 2496 2433 2504
rect 2447 2496 2553 2504
rect 2827 2496 2993 2504
rect 3527 2496 3753 2504
rect 3927 2496 3953 2504
rect 4207 2496 4293 2504
rect 4487 2496 4573 2504
rect 307 2476 424 2484
rect 416 2446 424 2476
rect 547 2477 633 2485
rect 827 2477 873 2485
rect 1207 2476 1232 2484
rect 916 2464 924 2474
rect 916 2456 993 2464
rect 1036 2464 1044 2474
rect 1267 2477 1353 2485
rect 1827 2476 1913 2484
rect 1987 2476 2213 2484
rect 1036 2456 1113 2464
rect 1596 2464 1604 2474
rect 1916 2464 1924 2474
rect 2267 2476 2493 2484
rect 2587 2476 2793 2484
rect 3167 2476 3453 2484
rect 3727 2477 3873 2485
rect 4027 2476 4073 2484
rect 4087 2476 4113 2484
rect 4247 2484 4260 2487
rect 4247 2473 4264 2484
rect 1407 2456 2453 2464
rect 3496 2464 3504 2473
rect 3387 2456 3504 2464
rect 147 2436 173 2444
rect 747 2436 813 2444
rect 947 2436 1053 2444
rect 1247 2435 1293 2443
rect 2627 2435 2933 2443
rect 3067 2435 3133 2443
rect 3767 2435 3813 2443
rect 4256 2446 4264 2473
rect 4756 2447 4764 2474
rect 5087 2476 5133 2484
rect 5147 2477 5173 2485
rect 5307 2477 5373 2485
rect 5427 2477 5453 2485
rect 5533 2484 5547 2493
rect 5516 2480 5547 2484
rect 5516 2476 5544 2480
rect 3887 2436 3993 2444
rect 4347 2435 4393 2443
rect 4507 2435 4533 2443
rect 4667 2436 4693 2444
rect 4756 2436 4773 2447
rect 4760 2433 4773 2436
rect 4836 2444 4844 2473
rect 4916 2447 4924 2474
rect 4836 2436 4853 2444
rect 4916 2436 4933 2447
rect 4920 2433 4933 2436
rect 4987 2436 5013 2444
rect 5067 2436 5153 2444
rect 5167 2435 5193 2443
rect 1127 2416 1173 2424
rect 1187 2416 1393 2424
rect 2107 2416 2173 2424
rect 2467 2416 2573 2424
rect 3327 2416 3413 2424
rect 1707 2396 1793 2404
rect 1807 2396 1953 2404
rect 2807 2396 2953 2404
rect 3047 2396 3293 2404
rect 3567 2396 3653 2404
rect 3967 2396 4133 2404
rect 4227 2396 4813 2404
rect 5216 2404 5224 2474
rect 5247 2436 5293 2444
rect 5516 2444 5524 2476
rect 5567 2476 5673 2484
rect 5787 2477 5813 2485
rect 5836 2446 5844 2493
rect 5867 2477 5993 2485
rect 5516 2436 5533 2444
rect 5327 2416 5353 2424
rect 5867 2416 5893 2424
rect 5216 2396 5253 2404
rect 5307 2396 5453 2404
rect 5807 2396 5973 2404
rect 867 2376 1173 2384
rect 1187 2376 1253 2384
rect 1267 2376 1473 2384
rect 1547 2376 1753 2384
rect 1767 2376 2133 2384
rect 2147 2376 2513 2384
rect 2847 2376 3913 2384
rect 5707 2376 5773 2384
rect 5787 2376 5813 2384
rect 647 2356 2733 2364
rect 2987 2356 3093 2364
rect 3467 2356 3573 2364
rect 4107 2356 4193 2364
rect 4787 2356 4813 2364
rect 4827 2356 4933 2364
rect 4947 2356 5293 2364
rect 807 2336 933 2344
rect 1147 2336 1293 2344
rect 2007 2336 2273 2344
rect 2907 2336 3153 2344
rect 3267 2336 3393 2344
rect 4067 2336 4233 2344
rect 5687 2336 5913 2344
rect 667 2316 753 2324
rect 1927 2316 2513 2324
rect 2527 2316 2613 2324
rect 2687 2316 2793 2324
rect 3247 2316 3953 2324
rect 4667 2316 4733 2324
rect 4747 2316 4893 2324
rect 4907 2316 4933 2324
rect 5427 2316 5613 2324
rect 5847 2316 5933 2324
rect 1007 2296 1213 2304
rect 1347 2296 1452 2304
rect 1487 2296 1553 2304
rect 1967 2296 2173 2304
rect 2247 2296 2393 2304
rect 2667 2296 2853 2304
rect 2867 2296 3013 2304
rect 4507 2296 4593 2304
rect 167 2276 693 2284
rect 827 2276 1133 2284
rect 3167 2276 3333 2284
rect 3447 2276 3513 2284
rect 3627 2276 3713 2284
rect 3927 2276 4313 2284
rect 4407 2276 4473 2284
rect 4940 2284 4953 2287
rect 4936 2273 4953 2284
rect 5047 2276 5073 2284
rect 5367 2276 5393 2284
rect 5580 2284 5593 2287
rect 5576 2273 5593 2284
rect 5647 2276 5733 2284
rect 5747 2276 5893 2284
rect 5907 2276 5973 2284
rect -24 2256 13 2264
rect 307 2256 333 2264
rect 1236 2256 1373 2264
rect 1236 2226 1244 2256
rect 1507 2256 1553 2264
rect 1727 2256 1793 2264
rect 1807 2256 1833 2264
rect 2007 2256 2073 2264
rect 2267 2256 2313 2264
rect 2387 2257 2453 2265
rect 2647 2257 2673 2265
rect 2727 2256 2933 2264
rect 3067 2256 3113 2264
rect 3176 2256 3193 2264
rect 3176 2244 3184 2256
rect 3287 2257 3533 2265
rect 1536 2236 1784 2244
rect 3136 2240 3184 2244
rect 1536 2226 1544 2236
rect 1776 2226 1784 2236
rect 3133 2236 3184 2240
rect 3133 2227 3147 2236
rect -24 2216 113 2224
rect 1287 2216 1353 2224
rect 1367 2215 1493 2223
rect 1747 2215 1773 2223
rect 1867 2216 1913 2224
rect 2027 2215 2053 2223
rect 2067 2216 2113 2224
rect 2627 2215 2693 2223
rect 2807 2215 2833 2223
rect 2847 2216 3033 2224
rect 3227 2215 3273 2223
rect 3327 2215 3513 2223
rect 3676 2224 3684 2254
rect 3746 2253 3747 2260
rect 3767 2256 3853 2264
rect 3907 2256 3933 2264
rect 3947 2256 4013 2264
rect 4187 2257 4253 2265
rect 3733 2244 3747 2253
rect 3733 2240 4004 2244
rect 3736 2236 4004 2240
rect 3996 2226 4004 2236
rect 3527 2216 3684 2224
rect 3707 2215 3753 2223
rect 4047 2215 4093 2223
rect 4636 2226 4644 2273
rect 4707 2256 4853 2264
rect 4936 2264 4944 2273
rect 4916 2256 4944 2264
rect 4916 2226 4924 2256
rect 4987 2257 5013 2265
rect 5187 2256 5253 2264
rect 5507 2256 5553 2264
rect 5576 2244 5584 2273
rect 5536 2236 5584 2244
rect 5536 2226 5544 2236
rect 5676 2227 5684 2253
rect 5773 2244 5787 2253
rect 5773 2240 5804 2244
rect 5776 2236 5804 2240
rect 4267 2216 4353 2224
rect 4407 2215 4513 2223
rect 4687 2216 4793 2224
rect 5027 2215 5093 2223
rect 5147 2215 5173 2223
rect 5796 2224 5804 2236
rect 5727 2216 5744 2224
rect 5796 2216 5833 2224
rect 527 2196 573 2204
rect 587 2196 873 2204
rect 887 2196 973 2204
rect 1707 2196 2193 2204
rect 2207 2196 2413 2204
rect 2887 2196 2993 2204
rect 3307 2196 3353 2204
rect 4307 2196 4333 2204
rect 4567 2196 5393 2204
rect 5736 2204 5744 2216
rect 5887 2216 6044 2224
rect 5736 2196 5813 2204
rect 5827 2196 5873 2204
rect 27 2176 253 2184
rect 1487 2176 1573 2184
rect 2347 2176 2593 2184
rect 3127 2176 3553 2184
rect 3567 2176 3653 2184
rect 3727 2176 3953 2184
rect 3967 2176 4153 2184
rect 4367 2176 4473 2184
rect 4767 2176 4813 2184
rect 5587 2176 5713 2184
rect 2167 2156 2253 2164
rect 2267 2156 2493 2164
rect 2507 2156 2633 2164
rect 2647 2156 2693 2164
rect 2947 2156 3313 2164
rect 3687 2156 4293 2164
rect 5767 2156 5913 2164
rect 5927 2156 5953 2164
rect 767 2136 1273 2144
rect 1527 2136 1973 2144
rect 1987 2136 2233 2144
rect 2567 2136 3173 2144
rect 3187 2136 3293 2144
rect 3367 2136 3453 2144
rect 3467 2136 4073 2144
rect 4087 2136 4593 2144
rect 5167 2136 5193 2144
rect 5207 2136 5273 2144
rect 1427 2116 2293 2124
rect 2387 2116 2633 2124
rect 2647 2116 2733 2124
rect 3507 2116 3673 2124
rect 3887 2116 4133 2124
rect 4307 2116 4553 2124
rect 5627 2116 5653 2124
rect 1487 2096 1693 2104
rect 3067 2096 3364 2104
rect 1307 2076 1513 2084
rect 2307 2076 2933 2084
rect 3356 2084 3364 2096
rect 3407 2096 3693 2104
rect 5347 2096 5433 2104
rect 5447 2096 5693 2104
rect 5707 2096 5933 2104
rect 3356 2076 3493 2084
rect 5547 2076 5653 2084
rect 3287 2056 3513 2064
rect 4027 2056 4113 2064
rect 4247 2056 4553 2064
rect 5507 2056 5813 2064
rect 87 2036 313 2044
rect 327 2036 913 2044
rect 1567 2036 1613 2044
rect 1627 2036 1673 2044
rect 2007 2036 2273 2044
rect 3087 2036 3253 2044
rect 3567 2036 3713 2044
rect 3827 2036 3893 2044
rect 3947 2036 4713 2044
rect 5207 2036 5293 2044
rect 5987 2036 6044 2044
rect 1207 2016 1313 2024
rect 1947 2016 2033 2024
rect 2307 2016 2333 2024
rect 2347 2016 2393 2024
rect 2407 2016 2533 2024
rect 2927 2016 5633 2024
rect 367 1996 893 2004
rect 1027 1996 1193 2004
rect 1407 1996 1613 2004
rect 1627 1996 1933 2004
rect 2087 1996 2153 2004
rect 3047 1996 3233 2004
rect 3247 1996 3433 2004
rect 3487 1996 3673 2004
rect 3747 1996 4253 2004
rect 4447 1996 4493 2004
rect 5147 1996 5233 2004
rect 5747 1996 5873 2004
rect 5947 2004 5960 2007
rect 5947 1993 5964 2004
rect 5987 1996 6044 2004
rect 1707 1976 1753 1984
rect 2227 1976 2373 1984
rect 2387 1976 2493 1984
rect 3107 1976 3133 1984
rect 3267 1976 3593 1984
rect 3607 1976 3633 1984
rect 4367 1976 4393 1984
rect 4527 1976 4573 1984
rect 5327 1976 5353 1984
rect 5427 1976 5533 1984
rect 5715 1984 5723 1993
rect 5715 1976 5833 1984
rect 207 1956 353 1964
rect 487 1957 513 1965
rect 647 1957 693 1965
rect 716 1956 733 1964
rect 716 1944 724 1956
rect 747 1956 1013 1964
rect 1196 1956 1353 1964
rect 667 1936 724 1944
rect 1156 1944 1164 1954
rect 1196 1944 1204 1956
rect 1367 1957 1393 1965
rect 1527 1956 1644 1964
rect 1107 1936 1204 1944
rect 407 1915 453 1923
rect 727 1916 813 1924
rect 1636 1926 1644 1956
rect 1867 1957 1893 1965
rect 2107 1956 2273 1964
rect 2287 1956 2364 1964
rect 2356 1944 2364 1956
rect 2747 1957 2793 1965
rect 2356 1936 2484 1944
rect 1147 1915 1253 1923
rect 1687 1915 1733 1923
rect 1787 1915 1813 1923
rect 2047 1915 2053 1923
rect 2067 1915 2073 1923
rect 2167 1915 2193 1923
rect 2476 1924 2484 1936
rect 2976 1944 2984 1954
rect 3107 1956 3213 1964
rect 3407 1957 3473 1965
rect 3916 1956 3953 1964
rect 2787 1936 2984 1944
rect 2476 1916 2513 1924
rect 2647 1915 2673 1923
rect 2687 1916 2833 1924
rect 2976 1924 2984 1936
rect 2976 1916 3273 1924
rect 3316 1907 3324 1954
rect 3347 1916 3393 1924
rect 3447 1915 3533 1923
rect 3656 1924 3664 1954
rect 3916 1944 3924 1956
rect 4007 1956 4033 1964
rect 4227 1956 4293 1964
rect 4396 1956 4433 1964
rect 3816 1936 3924 1944
rect 3547 1916 3664 1924
rect 3687 1916 3713 1924
rect 3816 1926 3824 1936
rect 3927 1915 3973 1923
rect 4127 1915 4153 1923
rect 4247 1916 4273 1924
rect 4396 1924 4404 1956
rect 4460 1964 4473 1967
rect 4456 1953 4473 1964
rect 4667 1957 4753 1965
rect 4847 1957 4893 1965
rect 5107 1956 5233 1964
rect 5387 1957 5473 1965
rect 5715 1964 5723 1976
rect 5956 1984 5964 1993
rect 5956 1976 6044 1984
rect 5715 1956 5744 1964
rect 4456 1944 4464 1953
rect 4416 1936 4464 1944
rect 4416 1926 4424 1936
rect 4936 1927 4944 1954
rect 5056 1944 5064 1954
rect 5007 1936 5064 1944
rect 5236 1944 5244 1954
rect 5236 1936 5284 1944
rect 4287 1916 4404 1924
rect 4627 1916 4653 1924
rect 4936 1916 4953 1927
rect 4940 1913 4953 1916
rect 5147 1916 5253 1924
rect 5276 1924 5284 1936
rect 5416 1936 5613 1944
rect 5276 1916 5353 1924
rect 5416 1924 5424 1936
rect 5736 1944 5744 1956
rect 6036 1964 6044 1976
rect 5927 1956 6044 1964
rect 5773 1944 5787 1953
rect 5736 1936 5764 1944
rect 5773 1940 5804 1944
rect 5776 1936 5804 1940
rect 5756 1926 5764 1936
rect 5407 1916 5424 1924
rect 5647 1915 5713 1923
rect 5796 1924 5804 1936
rect 5796 1916 5853 1924
rect 1967 1896 1993 1904
rect 2287 1896 2353 1904
rect 2447 1896 3013 1904
rect 3027 1896 3053 1904
rect 3167 1896 3253 1904
rect 3607 1896 3873 1904
rect 4227 1896 4573 1904
rect 1027 1876 1413 1884
rect 3507 1876 3573 1884
rect 3667 1876 3813 1884
rect 5647 1876 5893 1884
rect 887 1856 1333 1864
rect 1447 1856 1473 1864
rect 2407 1856 2493 1864
rect 3827 1856 4013 1864
rect 4467 1856 4733 1864
rect 4927 1856 4993 1864
rect 5087 1856 5293 1864
rect 5307 1856 5533 1864
rect 947 1836 1073 1844
rect 1127 1836 1153 1844
rect 1707 1836 1853 1844
rect 1867 1836 2013 1844
rect 2196 1836 2433 1844
rect 167 1816 233 1824
rect 967 1816 1033 1824
rect 1287 1816 1333 1824
rect 1347 1816 1433 1824
rect 2196 1824 2204 1836
rect 3187 1836 3293 1844
rect 3627 1836 3773 1844
rect 3787 1836 4233 1844
rect 4787 1836 4853 1844
rect 4867 1836 5013 1844
rect 5167 1836 5253 1844
rect 5707 1836 5993 1844
rect 1847 1816 2204 1824
rect 2347 1816 2393 1824
rect 2407 1816 2913 1824
rect 2987 1816 3073 1824
rect 3207 1816 3253 1824
rect 67 1796 113 1804
rect 127 1796 593 1804
rect 727 1796 773 1804
rect 1387 1796 1613 1804
rect 1627 1796 3153 1804
rect 3167 1796 3293 1804
rect 3867 1796 4793 1804
rect 4807 1796 4953 1804
rect 5347 1796 5673 1804
rect 147 1776 193 1784
rect 367 1776 393 1784
rect 407 1776 633 1784
rect 1267 1776 1353 1784
rect 1407 1776 1553 1784
rect 2567 1776 2653 1784
rect 3047 1776 3113 1784
rect 3347 1776 3553 1784
rect 4007 1776 4353 1784
rect 4447 1776 4492 1784
rect 4527 1776 4593 1784
rect 5007 1776 5213 1784
rect 5227 1776 5473 1784
rect 5867 1776 5933 1784
rect 227 1756 273 1764
rect 287 1756 653 1764
rect 1587 1756 1693 1764
rect 1707 1756 1833 1764
rect 1927 1756 2153 1764
rect 2967 1756 2993 1764
rect 3007 1756 3104 1764
rect 607 1737 633 1745
rect 767 1736 784 1744
rect -24 1696 53 1704
rect 187 1695 213 1703
rect 307 1696 413 1704
rect 436 1687 444 1734
rect 667 1716 744 1724
rect 487 1696 573 1704
rect 736 1706 744 1716
rect 776 1707 784 1736
rect 1087 1737 1133 1745
rect 1307 1736 1393 1744
rect 1556 1724 1564 1734
rect 1967 1736 2053 1744
rect 2107 1736 2164 1744
rect 1456 1716 1564 1724
rect 2156 1727 2164 1736
rect 2267 1736 2313 1744
rect 2527 1737 2573 1745
rect 2627 1736 2673 1744
rect 2727 1736 2793 1744
rect 2867 1737 2913 1745
rect 3096 1744 3104 1756
rect 3147 1756 3204 1764
rect 3096 1736 3173 1744
rect 3196 1744 3204 1756
rect 3247 1756 3273 1764
rect 3387 1756 3533 1764
rect 3947 1756 4313 1764
rect 5247 1756 5373 1764
rect 5387 1756 5444 1764
rect 3196 1736 3213 1744
rect 3347 1737 3453 1745
rect 2156 1716 2173 1727
rect 647 1696 693 1704
rect 987 1695 1033 1703
rect 1047 1696 1093 1704
rect 1287 1695 1333 1703
rect 1456 1704 1464 1716
rect 2160 1713 2173 1716
rect 3076 1724 3084 1734
rect 3607 1736 3653 1744
rect 3867 1736 3893 1744
rect 4107 1736 4144 1744
rect 3076 1720 3164 1724
rect 3076 1716 3167 1720
rect 3153 1707 3167 1716
rect 3567 1716 3993 1724
rect 4136 1707 4144 1736
rect 4307 1737 4393 1745
rect 4416 1736 4493 1744
rect 4416 1724 4424 1736
rect 4547 1736 4653 1744
rect 4707 1737 4753 1745
rect 4813 1744 4827 1753
rect 4813 1740 4913 1744
rect 4816 1736 4913 1740
rect 5067 1736 5213 1744
rect 5347 1736 5404 1744
rect 4216 1716 4424 1724
rect 1427 1696 1464 1704
rect 1627 1696 1673 1704
rect 1887 1695 1953 1703
rect 2027 1695 2073 1703
rect 2127 1695 2153 1703
rect 2467 1695 2813 1703
rect 2947 1695 3013 1703
rect 3027 1696 3144 1704
rect 436 1676 453 1687
rect 440 1673 453 1676
rect 1247 1676 1473 1684
rect 1487 1676 1553 1684
rect 1956 1684 1964 1692
rect 1956 1676 2233 1684
rect 2476 1676 2773 1684
rect 147 1656 353 1664
rect 913 1664 927 1673
rect 913 1660 1053 1664
rect 916 1656 1053 1660
rect 1367 1656 1793 1664
rect 2476 1664 2484 1676
rect 3136 1684 3144 1696
rect 3247 1695 3273 1703
rect 3687 1695 3733 1703
rect 3887 1695 3913 1703
rect 4216 1706 4224 1716
rect 5396 1706 5404 1736
rect 5436 1744 5444 1756
rect 5616 1756 5713 1764
rect 5616 1748 5624 1756
rect 5436 1736 5513 1744
rect 5567 1737 5613 1745
rect 5696 1736 5853 1744
rect 5416 1724 5424 1734
rect 5416 1716 5644 1724
rect 4267 1695 4293 1703
rect 4567 1695 4593 1703
rect 4827 1696 4993 1704
rect 5087 1696 5193 1704
rect 3136 1676 3193 1684
rect 3527 1676 3553 1684
rect 4347 1676 4553 1684
rect 4567 1676 4713 1684
rect 5067 1676 5233 1684
rect 5247 1676 5353 1684
rect 5636 1686 5644 1716
rect 5696 1706 5704 1736
rect 5807 1695 5833 1703
rect 2387 1656 2484 1664
rect 2567 1656 2653 1664
rect 2667 1656 2693 1664
rect 2847 1656 2993 1664
rect 3007 1656 3393 1664
rect 3407 1656 3473 1664
rect 3707 1656 3913 1664
rect 3927 1656 3953 1664
rect 4087 1656 4253 1664
rect 4967 1656 5033 1664
rect 5547 1656 5693 1664
rect 2607 1636 3353 1644
rect 3376 1636 3633 1644
rect 3376 1624 3384 1636
rect 3647 1636 4013 1644
rect 4927 1636 5233 1644
rect 2827 1616 3384 1624
rect 4647 1616 4773 1624
rect 4787 1616 4833 1624
rect 1073 1604 1087 1613
rect 1073 1600 2333 1604
rect 1076 1596 2333 1600
rect 2687 1596 2804 1604
rect 1027 1576 1113 1584
rect 2796 1584 2804 1596
rect 3167 1596 3453 1604
rect 3747 1596 5493 1604
rect 5607 1596 5733 1604
rect 2796 1576 3033 1584
rect 3267 1576 3693 1584
rect 2427 1556 2473 1564
rect 2567 1556 2593 1564
rect 2767 1556 3073 1564
rect 4787 1556 5013 1564
rect 5207 1556 5613 1564
rect 1827 1536 2164 1544
rect 1427 1516 1493 1524
rect 1987 1516 2073 1524
rect 2156 1524 2164 1536
rect 2187 1536 2513 1544
rect 2527 1536 2733 1544
rect 3147 1536 3513 1544
rect 3687 1536 3853 1544
rect 4467 1536 5113 1544
rect 5247 1536 5933 1544
rect 2156 1516 2433 1524
rect 2447 1516 2593 1524
rect 2656 1516 2933 1524
rect 467 1496 733 1504
rect 747 1496 833 1504
rect 2656 1504 2664 1516
rect 4527 1516 4624 1524
rect 2547 1496 2664 1504
rect 4267 1496 4313 1504
rect 4616 1504 4624 1516
rect 4616 1496 4953 1504
rect 1207 1476 1233 1484
rect 1367 1476 1393 1484
rect 1407 1476 1473 1484
rect 1676 1476 1813 1484
rect 1676 1467 1684 1476
rect 2227 1476 2453 1484
rect 2787 1476 2893 1484
rect 3127 1476 3193 1484
rect 3267 1476 3393 1484
rect 3447 1476 3533 1484
rect 3587 1476 3613 1484
rect 3727 1476 4013 1484
rect 4487 1476 4593 1484
rect 4607 1476 4673 1484
rect 4687 1476 4793 1484
rect 5027 1476 5233 1484
rect 5347 1476 5373 1484
rect 5467 1476 5733 1484
rect 5747 1476 5853 1484
rect 1587 1456 1673 1464
rect 2007 1456 2133 1464
rect 3287 1456 3373 1464
rect 3387 1456 3444 1464
rect -24 1404 -16 1444
rect 207 1437 232 1445
rect 267 1437 293 1445
rect 607 1437 653 1445
rect 707 1437 773 1445
rect 887 1437 933 1445
rect 1167 1436 1293 1444
rect 1747 1437 1773 1445
rect 1907 1437 1993 1445
rect 2187 1437 2233 1445
rect 2256 1436 2273 1444
rect 1336 1424 1344 1434
rect 1336 1416 1504 1424
rect -24 1396 93 1404
rect 1496 1406 1504 1416
rect 2256 1407 2264 1436
rect 2487 1436 2553 1444
rect 2687 1437 2773 1445
rect 2867 1436 3053 1444
rect 3307 1437 3333 1445
rect 3436 1444 3444 1456
rect 3807 1456 3893 1464
rect 4016 1464 4024 1473
rect 4016 1456 4253 1464
rect 4387 1456 4433 1464
rect 5287 1456 5313 1464
rect 5327 1456 5393 1464
rect 5527 1456 5553 1464
rect 3436 1436 3453 1444
rect 3476 1436 3573 1444
rect 3476 1424 3484 1436
rect 3707 1436 3753 1444
rect 3967 1436 4084 1444
rect 3187 1416 3484 1424
rect 567 1396 633 1404
rect 827 1396 1033 1404
rect 1187 1395 1233 1403
rect 1247 1396 1313 1404
rect 1847 1396 1893 1404
rect 2087 1395 2153 1403
rect 2307 1395 2353 1403
rect 2527 1395 2573 1403
rect 2807 1396 2833 1404
rect 2847 1396 2913 1404
rect 3047 1395 3093 1403
rect 3247 1396 3353 1404
rect 3427 1395 3473 1403
rect 3527 1395 3593 1403
rect 3647 1396 3733 1404
rect 4076 1406 4084 1436
rect 4167 1437 4193 1445
rect 4440 1444 4453 1447
rect 4436 1433 4453 1444
rect 4507 1436 4553 1444
rect 4667 1436 4713 1444
rect 4807 1444 4820 1447
rect 4807 1433 4824 1444
rect 4887 1437 4933 1445
rect 5067 1437 5093 1445
rect 5167 1437 5193 1445
rect 3807 1396 3833 1404
rect 4436 1406 4444 1433
rect 4307 1396 4393 1404
rect 4627 1396 4793 1404
rect 4816 1404 4824 1433
rect 4816 1396 4853 1404
rect 4967 1396 4993 1404
rect 5047 1395 5073 1403
rect 5127 1396 5173 1404
rect 5356 1404 5364 1434
rect 5487 1444 5500 1447
rect 5487 1433 5504 1444
rect 5596 1440 5633 1444
rect 5327 1396 5364 1404
rect 5387 1396 5433 1404
rect 5496 1406 5504 1433
rect 5593 1436 5633 1440
rect 5593 1427 5607 1436
rect 327 1376 593 1384
rect 2516 1384 2524 1392
rect 2427 1376 2524 1384
rect 3267 1376 3333 1384
rect 4507 1376 4693 1384
rect 5147 1376 5213 1384
rect 5227 1376 5293 1384
rect 5667 1376 5733 1384
rect 147 1356 413 1364
rect 527 1356 553 1364
rect 596 1364 604 1373
rect 596 1356 873 1364
rect 1347 1356 1413 1364
rect 1427 1356 1453 1364
rect 1567 1356 1653 1364
rect 1667 1356 1793 1364
rect 2707 1356 2753 1364
rect 2887 1356 3173 1364
rect 4327 1356 4393 1364
rect 4827 1356 4853 1364
rect 4927 1356 5093 1364
rect 5627 1356 5833 1364
rect 687 1336 733 1344
rect 1987 1336 2073 1344
rect 2467 1336 2533 1344
rect 2767 1336 2853 1344
rect 3207 1336 3273 1344
rect 3287 1336 3313 1344
rect 4907 1336 5133 1344
rect 5147 1336 5313 1344
rect 127 1316 253 1324
rect 1027 1316 1053 1324
rect 1427 1316 1733 1324
rect 4027 1316 4133 1324
rect 4227 1316 4493 1324
rect 5007 1316 5173 1324
rect 2687 1296 2784 1304
rect 327 1276 693 1284
rect 767 1276 993 1284
rect 1287 1276 1453 1284
rect 1467 1276 1593 1284
rect 2776 1284 2784 1296
rect 3227 1296 3373 1304
rect 3547 1296 4813 1304
rect 4887 1296 4933 1304
rect 4987 1296 5284 1304
rect 2776 1276 2913 1284
rect 3927 1276 4953 1284
rect 5276 1284 5284 1296
rect 5307 1296 5333 1304
rect 5276 1276 5373 1284
rect 1307 1256 1353 1264
rect 2007 1256 2113 1264
rect 2627 1256 2753 1264
rect 3147 1256 3413 1264
rect 3567 1256 3893 1264
rect 4287 1256 4473 1264
rect 4667 1256 4733 1264
rect 4807 1256 4873 1264
rect 4927 1256 5113 1264
rect 5487 1256 5653 1264
rect 5727 1256 5813 1264
rect 267 1236 293 1244
rect 307 1236 473 1244
rect 587 1236 833 1244
rect 1207 1236 1393 1244
rect 1587 1236 1613 1244
rect 1747 1236 1793 1244
rect 2167 1236 2253 1244
rect 2787 1236 2993 1244
rect 3127 1236 3213 1244
rect 3367 1236 3393 1244
rect 3507 1236 3673 1244
rect 3687 1236 3713 1244
rect 4587 1236 4753 1244
rect 4767 1236 4804 1244
rect 387 1216 453 1224
rect 607 1216 653 1224
rect 887 1217 953 1225
rect 1247 1216 1333 1224
rect 1507 1216 1553 1224
rect 1667 1216 1713 1224
rect 1847 1216 1893 1224
rect 1947 1216 2013 1224
rect 2027 1217 2073 1225
rect 2127 1216 2173 1224
rect 2287 1217 2333 1225
rect 2407 1217 2433 1225
rect 2447 1216 2593 1224
rect 2647 1216 2672 1224
rect 2707 1217 2733 1225
rect 2987 1216 3053 1224
rect 3067 1216 3233 1224
rect 3416 1216 3453 1224
rect 396 1196 573 1204
rect 147 1175 193 1183
rect 247 1176 313 1184
rect 396 1186 404 1196
rect 1956 1196 2153 1204
rect 467 1175 493 1183
rect 727 1175 793 1183
rect 1227 1176 1273 1184
rect 1367 1176 1393 1184
rect 1587 1175 1633 1183
rect 1787 1176 1853 1184
rect 1956 1186 1964 1196
rect 2096 1186 2104 1196
rect 3416 1204 3424 1216
rect 3607 1217 3633 1225
rect 3647 1216 3753 1224
rect 3967 1216 3993 1224
rect 4007 1216 4033 1224
rect 4327 1216 4433 1224
rect 4796 1224 4804 1236
rect 4707 1216 4744 1224
rect 4796 1216 5013 1224
rect 3376 1200 3424 1204
rect 3373 1196 3424 1200
rect 3373 1187 3387 1196
rect 2307 1176 2393 1184
rect 2767 1176 2893 1184
rect 2947 1175 2973 1183
rect 3207 1176 3253 1184
rect 3267 1176 3293 1184
rect 4736 1187 4744 1216
rect 5116 1216 5213 1224
rect 5056 1204 5064 1214
rect 5116 1204 5124 1216
rect 5347 1216 5364 1224
rect 5056 1196 5124 1204
rect 5356 1204 5364 1216
rect 5387 1216 5453 1224
rect 5553 1224 5567 1233
rect 5527 1220 5567 1224
rect 5527 1216 5564 1220
rect 5747 1216 5993 1224
rect 5356 1196 5713 1204
rect 3527 1175 3553 1183
rect 4227 1175 4253 1183
rect 4307 1176 4453 1184
rect 4736 1176 4753 1187
rect 4740 1173 4753 1176
rect 4847 1175 4873 1183
rect 5056 1184 5064 1196
rect 4927 1176 5064 1184
rect 5147 1176 5253 1184
rect 5467 1175 5533 1183
rect 5687 1175 5753 1183
rect 5767 1176 5884 1184
rect 1076 1144 1084 1172
rect 1576 1164 1584 1172
rect 1487 1156 1584 1164
rect 3727 1156 3893 1164
rect 3947 1156 4013 1164
rect 5087 1156 5193 1164
rect 5207 1156 5273 1164
rect 5876 1164 5884 1176
rect 5976 1176 6044 1184
rect 5976 1164 5984 1176
rect 5876 1156 5984 1164
rect 867 1136 1333 1144
rect 2487 1136 2573 1144
rect 2587 1136 2693 1144
rect 2707 1136 3073 1144
rect 3487 1136 3773 1144
rect 4647 1136 4833 1144
rect 4887 1136 4973 1144
rect 1527 1116 1733 1124
rect 1747 1116 2193 1124
rect 2207 1116 2413 1124
rect 4067 1116 4173 1124
rect 5647 1116 5733 1124
rect 5867 1116 5933 1124
rect 1567 1096 1913 1104
rect 1927 1096 2053 1104
rect 3407 1096 4873 1104
rect 4927 1096 5193 1104
rect 5407 1096 5693 1104
rect 5707 1096 5833 1104
rect 5967 1096 5993 1104
rect 947 1076 1133 1084
rect 3867 1076 4053 1084
rect 1787 1056 1873 1064
rect 1887 1056 1993 1064
rect 4527 1056 4793 1064
rect 4807 1056 5293 1064
rect 967 1036 1013 1044
rect 1707 1036 2713 1044
rect 3667 1036 4073 1044
rect 4827 1036 4933 1044
rect 5067 1036 5233 1044
rect 4727 1016 4993 1024
rect 1847 996 2053 1004
rect 2147 996 2353 1004
rect 3247 996 3473 1004
rect 3527 996 3933 1004
rect 4367 996 4633 1004
rect 5267 996 5393 1004
rect 5547 996 5592 1004
rect 5627 996 5753 1004
rect 1867 976 2253 984
rect 2727 976 3373 984
rect 3967 976 4324 984
rect 4316 967 4324 976
rect 4767 976 4813 984
rect 767 956 953 964
rect 1667 956 1813 964
rect 1927 956 2193 964
rect 2307 956 3193 964
rect 3287 956 3513 964
rect 4327 956 4553 964
rect 4947 956 5153 964
rect 5287 956 5453 964
rect 5567 956 5664 964
rect 5656 947 5664 956
rect 1727 936 1933 944
rect 1947 936 2093 944
rect 2247 936 2373 944
rect 3707 936 3753 944
rect 5667 936 5713 944
rect -24 916 73 924
rect 407 917 473 925
rect 607 916 713 924
rect 727 916 813 924
rect 887 916 973 924
rect 1087 917 1133 925
rect 1187 917 1233 925
rect 1427 916 1473 924
rect 1567 917 1613 925
rect 1827 917 1853 925
rect 1987 916 2133 924
rect 2487 916 2573 924
rect 2767 917 2793 925
rect 2907 917 2953 925
rect 3047 917 3073 925
rect 1296 904 1304 913
rect 2296 904 2304 914
rect 2996 904 3004 914
rect 3127 916 3153 924
rect 3167 917 3293 925
rect 3387 916 3453 924
rect 3847 916 3953 924
rect 4367 917 4413 925
rect 4507 917 4573 925
rect 4707 917 4733 925
rect 4967 916 5113 924
rect 5127 916 5253 924
rect 5587 917 5613 925
rect 5807 916 5933 924
rect 1296 896 1364 904
rect 2296 896 2384 904
rect 2996 896 3093 904
rect 507 875 573 883
rect 747 876 793 884
rect 847 876 1253 884
rect 1356 884 1364 896
rect 2376 887 2384 896
rect 3656 904 3664 913
rect 3796 904 3804 914
rect 3656 896 3893 904
rect 4087 896 4224 904
rect 1356 876 1393 884
rect 1647 875 1693 883
rect 1887 875 1953 883
rect 1967 876 2113 884
rect 2376 876 2393 887
rect 2380 873 2393 876
rect 2747 875 2813 883
rect 3227 875 3273 883
rect 4216 886 4224 896
rect 4856 887 4864 914
rect 5496 904 5504 914
rect 5496 896 5544 904
rect 3607 876 3673 884
rect 4427 876 4473 884
rect 4587 876 4633 884
rect 4856 876 4873 887
rect 4860 873 4873 876
rect 4947 875 4993 883
rect 5147 876 5213 884
rect 5407 876 5433 884
rect 5487 875 5513 883
rect 5536 884 5544 896
rect 5536 876 5673 884
rect 5847 875 5913 883
rect 2367 856 2493 864
rect 2607 856 2993 864
rect 3307 856 3733 864
rect 3747 856 3873 864
rect 4027 856 4073 864
rect 4696 856 4793 864
rect 147 836 233 844
rect 247 836 313 844
rect 667 836 1153 844
rect 1267 836 1593 844
rect 2067 836 2273 844
rect 2427 836 2513 844
rect 2827 836 3013 844
rect 3187 836 3813 844
rect 3987 836 4093 844
rect 4696 844 4704 856
rect 5007 856 5273 864
rect 5327 856 5453 864
rect 4720 844 4733 847
rect 4567 836 4704 844
rect 4716 833 4733 844
rect 4827 836 4873 844
rect 5067 836 5133 844
rect 5207 836 5353 844
rect 5527 836 5593 844
rect 5867 836 5913 844
rect 1507 816 1553 824
rect 1567 816 1693 824
rect 2807 816 3493 824
rect 3547 816 3613 824
rect 4716 824 4724 833
rect 4527 816 4724 824
rect 5647 816 5773 824
rect 827 796 933 804
rect 1327 796 1793 804
rect 2247 796 2693 804
rect 3107 796 3253 804
rect 3907 796 3993 804
rect 4747 796 5193 804
rect 5407 796 5593 804
rect 467 776 533 784
rect 2167 776 2253 784
rect 2327 776 2673 784
rect 2887 776 3313 784
rect 3327 776 3353 784
rect 4327 776 4713 784
rect 4847 776 5013 784
rect 347 756 693 764
rect 707 756 713 764
rect 727 756 893 764
rect 1107 756 1173 764
rect 1347 756 1573 764
rect 1947 756 2713 764
rect 2967 756 3153 764
rect 3267 756 3533 764
rect 3547 756 3693 764
rect 4467 756 4673 764
rect 5547 756 5633 764
rect 5707 756 5773 764
rect 507 736 873 744
rect 967 736 993 744
rect 1987 736 2033 744
rect 2207 736 2553 744
rect 2847 736 2933 744
rect 2947 736 3233 744
rect 4387 736 4753 744
rect 5047 736 5233 744
rect 5367 736 5513 744
rect 5567 736 5613 744
rect 167 716 293 724
rect 307 716 373 724
rect 927 716 953 724
rect 2327 716 2353 724
rect 2467 716 2604 724
rect 87 696 113 704
rect 407 697 453 705
rect 467 696 593 704
rect 767 696 884 704
rect 876 666 884 696
rect 1247 696 1393 704
rect 1507 697 1533 705
rect 1667 697 1733 705
rect 896 684 904 694
rect 1807 696 1873 704
rect 1887 696 1993 704
rect 2487 696 2513 704
rect 2596 704 2604 716
rect 2627 716 2884 724
rect 2596 696 2704 704
rect 896 676 944 684
rect 187 656 273 664
rect 627 656 733 664
rect 787 655 813 663
rect 487 636 533 644
rect 936 644 944 676
rect 2096 676 2233 684
rect 987 655 1113 663
rect 1287 655 1333 663
rect 1447 656 1493 664
rect 2096 666 2104 676
rect 2696 667 2704 696
rect 2767 697 2813 705
rect 2876 704 2884 716
rect 3427 716 3473 724
rect 4247 716 4273 724
rect 4296 716 4333 724
rect 2876 696 2893 704
rect 2907 696 2973 704
rect 2987 696 3053 704
rect 3147 696 3193 704
rect 3247 696 3373 704
rect 3507 704 3520 707
rect 3507 693 3524 704
rect 3587 696 3633 704
rect 3747 696 3833 704
rect 3947 697 4033 705
rect 4087 696 4173 704
rect 4296 704 4304 716
rect 5267 716 5544 724
rect 4187 696 4304 704
rect 4507 696 4593 704
rect 4647 697 4673 705
rect 4787 696 4913 704
rect 5007 697 5073 705
rect 5087 696 5233 704
rect 5327 696 5353 704
rect 5536 704 5544 716
rect 5436 696 5544 704
rect 3516 684 3524 693
rect 3516 676 3724 684
rect 1627 655 1713 663
rect 1767 656 1893 664
rect 1907 655 1933 663
rect 2407 656 2433 664
rect 3516 666 3524 676
rect 3716 666 3724 676
rect 5436 667 5444 696
rect 2787 655 2833 663
rect 3327 655 3393 663
rect 3567 656 3673 664
rect 3907 655 4233 663
rect 4727 656 4793 664
rect 5536 666 5544 696
rect 5567 696 5593 704
rect 5607 696 5833 704
rect 5887 696 5933 704
rect 5647 655 5673 663
rect 5787 655 5813 663
rect 936 636 964 644
rect 87 616 393 624
rect 956 624 964 636
rect 1187 636 2133 644
rect 2687 636 2753 644
rect 2767 636 2873 644
rect 2887 636 3033 644
rect 3247 636 3353 644
rect 3547 636 3693 644
rect 3747 636 3853 644
rect 4347 636 4373 644
rect 4687 636 4933 644
rect 4947 636 5093 644
rect 5107 636 5213 644
rect 956 616 1373 624
rect 1387 616 1553 624
rect 1607 616 1653 624
rect 1667 616 1853 624
rect 2193 624 2207 633
rect 1987 620 2207 624
rect 1987 616 2204 620
rect 2267 616 2573 624
rect 3147 616 3933 624
rect 4067 616 4493 624
rect 2927 596 3113 604
rect 3647 596 4013 604
rect 4587 596 4693 604
rect 4707 596 4753 604
rect 5067 596 5253 604
rect 347 576 373 584
rect 4787 576 4993 584
rect 2287 556 2353 564
rect 2467 556 2733 564
rect 2847 556 3133 564
rect 3387 556 3484 564
rect 1467 536 1753 544
rect 1767 536 2113 544
rect 3007 536 3073 544
rect 3476 544 3484 556
rect 3627 556 4153 564
rect 3476 536 3593 544
rect 5727 536 5773 544
rect 5787 536 5853 544
rect 2527 516 2573 524
rect 2587 516 2613 524
rect 3167 516 3453 524
rect 3476 516 3604 524
rect 327 496 393 504
rect 407 496 2293 504
rect 3476 504 3484 516
rect 3347 496 3484 504
rect 3596 504 3604 516
rect 3627 516 4304 524
rect 4296 507 4304 516
rect 4727 516 4833 524
rect 4847 516 5313 524
rect 3596 496 3893 504
rect 4307 496 4393 504
rect 5067 496 5093 504
rect 5167 496 5453 504
rect 5467 496 5593 504
rect 2947 476 3093 484
rect 3107 476 3193 484
rect 3207 476 3573 484
rect 4107 476 4933 484
rect 287 456 412 464
rect 447 456 493 464
rect 507 456 713 464
rect 807 456 833 464
rect 2607 456 2653 464
rect 2707 456 3064 464
rect 1927 436 1973 444
rect 1987 436 2113 444
rect 3056 444 3064 456
rect 3127 456 3333 464
rect 3447 456 3553 464
rect 5527 456 5673 464
rect 5727 456 5873 464
rect 3056 436 3393 444
rect 3487 436 3613 444
rect 3887 436 4353 444
rect 4427 436 4473 444
rect 4496 436 4553 444
rect 467 416 553 424
rect 2147 416 2193 424
rect 2387 416 2413 424
rect 2507 416 2613 424
rect 3467 416 3653 424
rect 3667 416 3753 424
rect 4187 416 4213 424
rect 4496 424 4504 436
rect 4567 436 5053 444
rect 4407 416 4504 424
rect 4807 416 4873 424
rect 4887 416 5013 424
rect 5367 416 5373 424
rect 5387 416 5413 424
rect 5616 416 5713 424
rect 127 396 233 404
rect 347 397 433 405
rect 647 397 673 405
rect 727 396 833 404
rect 907 397 973 405
rect 976 384 984 394
rect 1116 384 1124 394
rect 1267 396 1293 404
rect 1707 396 1833 404
rect 2887 396 3113 404
rect 3127 397 3153 405
rect 3167 396 3293 404
rect 976 376 1124 384
rect 2156 384 2164 394
rect 2067 376 2164 384
rect 187 356 213 364
rect 267 356 333 364
rect 427 356 473 364
rect 627 356 733 364
rect 747 355 793 363
rect 1007 356 1313 364
rect 1327 356 1393 364
rect 1767 355 1813 363
rect 1887 356 1953 364
rect 2147 356 2453 364
rect 2536 364 2544 394
rect 3547 396 3613 404
rect 3807 397 3853 405
rect 4247 396 4313 404
rect 3936 367 3944 394
rect 4467 397 4513 405
rect 4576 384 4584 413
rect 5616 408 5624 416
rect 4647 397 4673 405
rect 5207 397 5293 405
rect 4047 376 4384 384
rect 2536 356 2613 364
rect 2627 356 2733 364
rect 2907 355 2933 363
rect 3027 356 3113 364
rect 3187 356 3233 364
rect 3327 356 3433 364
rect 3507 355 3533 363
rect 3827 356 3873 364
rect 3927 364 3944 367
rect 3927 356 4113 364
rect 3927 353 3940 356
rect 4187 356 4273 364
rect 4376 366 4384 376
rect 4516 376 4584 384
rect 4516 364 4524 376
rect 4427 356 4524 364
rect 4547 356 4633 364
rect 4747 356 4773 364
rect 787 336 853 344
rect 1727 336 1773 344
rect 2307 336 2513 344
rect 3536 344 3544 352
rect 3536 336 3773 344
rect 3967 336 4033 344
rect 4587 336 4613 344
rect 4687 336 4793 344
rect 4816 344 4824 393
rect 5056 384 5064 394
rect 5447 396 5473 404
rect 5567 397 5613 405
rect 5696 396 5733 404
rect 5056 376 5144 384
rect 4907 355 4933 363
rect 4947 356 4993 364
rect 5047 356 5093 364
rect 5136 364 5144 376
rect 5696 366 5704 396
rect 5747 397 5833 405
rect 5136 356 5173 364
rect 5227 356 5373 364
rect 5387 356 5493 364
rect 5547 356 5693 364
rect 4816 336 4853 344
rect 5127 336 5333 344
rect 5607 336 5653 344
rect 1367 316 1993 324
rect 2007 316 2052 324
rect 2087 316 2493 324
rect 2547 316 2853 324
rect 4127 316 4213 324
rect 4387 316 4453 324
rect 4467 316 4693 324
rect 147 296 413 304
rect 427 296 633 304
rect 867 296 1053 304
rect 1067 296 1133 304
rect 1147 296 2493 304
rect 3647 296 3933 304
rect 3947 296 4013 304
rect 4027 296 4073 304
rect 4327 296 4353 304
rect 4407 296 4673 304
rect 5647 296 5973 304
rect 1507 276 1613 284
rect 2587 276 2673 284
rect 3727 276 4193 284
rect 5427 276 5673 284
rect 827 256 893 264
rect 2696 256 3373 264
rect 707 236 753 244
rect 1127 236 1913 244
rect 2227 236 2413 244
rect 2696 244 2704 256
rect 4307 256 4493 264
rect 2467 236 2704 244
rect 2787 236 2904 244
rect 1607 216 1773 224
rect 2896 224 2904 236
rect 4267 236 4553 244
rect 5787 236 5853 244
rect 2896 216 3013 224
rect 3627 216 3853 224
rect 4256 224 4264 233
rect 3867 216 4264 224
rect 4287 216 4513 224
rect 5347 216 5533 224
rect 5547 216 5613 224
rect 2387 196 2413 204
rect 2727 196 2873 204
rect 2887 196 2953 204
rect 3307 196 3373 204
rect -24 176 113 184
rect -24 136 -16 176
rect 187 177 273 185
rect 287 176 373 184
rect 387 176 493 184
rect 707 176 813 184
rect 927 177 1073 185
rect 1087 176 1244 184
rect 1236 164 1244 176
rect 1267 176 1313 184
rect 1660 184 1673 187
rect 1656 173 1673 184
rect 1760 184 1773 187
rect 1756 173 1773 184
rect 1827 177 1873 185
rect 2127 176 2233 184
rect 2547 177 2633 185
rect 3167 176 3233 184
rect 3247 176 3453 184
rect 3787 177 3813 185
rect 1236 156 1293 164
rect 147 136 173 144
rect 247 136 393 144
rect 447 135 472 143
rect 507 135 533 143
rect 727 135 753 143
rect 847 136 913 144
rect 1656 146 1664 173
rect 1756 146 1764 173
rect 1936 156 1984 164
rect 1936 146 1944 156
rect 967 136 1093 144
rect 1147 136 1233 144
rect 1327 135 1373 143
rect 1976 144 1984 156
rect 1976 136 2453 144
rect 2647 136 2673 144
rect 2687 136 2833 144
rect 2967 135 2993 143
rect 3047 136 3233 144
rect 3247 135 3273 143
rect 3327 135 3393 143
rect 3547 135 3633 143
rect 3647 136 3713 144
rect 3916 146 3924 193
rect 4007 176 4053 184
rect 4407 176 4473 184
rect 4527 176 4713 184
rect 5047 176 5153 184
rect 3987 156 4153 164
rect 4167 156 4384 164
rect 4376 146 4384 156
rect 4487 135 4533 143
rect 4687 135 4713 143
rect 4796 144 4804 174
rect 5227 176 5293 184
rect 5407 176 5473 184
rect 5927 176 6044 184
rect 4796 136 4913 144
rect 5367 135 5413 143
rect 5687 136 5753 144
rect 347 116 673 124
rect 1707 116 1933 124
rect 2587 116 2753 124
rect 2907 116 3033 124
rect 3607 116 3753 124
rect 4087 116 4293 124
rect 4307 116 4413 124
rect 5467 116 5533 124
rect 5647 116 5873 124
rect 5887 116 5993 124
rect 327 96 573 104
rect 3387 96 3973 104
rect 4507 96 4613 104
rect 4627 96 4853 104
rect 1827 76 2013 84
rect 2607 76 3133 84
rect 4427 76 5393 84
rect 3487 56 3953 64
rect 4047 56 4393 64
rect 4447 56 5313 64
rect 5607 56 5933 64
rect 3827 36 3873 44
rect 3887 36 3993 44
rect 4587 36 5213 44
rect 3087 16 3113 24
rect 3127 16 3173 24
rect 3707 16 3773 24
use INVX1  _756_
timestamp 0
transform 1 0 1350 0 -1 3910
box -6 -8 46 268
use INVX1  _757_
timestamp 0
transform 1 0 1710 0 1 3390
box -6 -8 46 268
use NOR2X1  _758_
timestamp 0
transform 1 0 1470 0 -1 3910
box -6 -8 66 268
use NAND2X1  _759_
timestamp 0
transform 1 0 610 0 1 3910
box -6 -8 66 268
use INVX1  _760_
timestamp 0
transform 1 0 770 0 1 3910
box -6 -8 46 268
use NOR2X1  _761_
timestamp 0
transform 1 0 470 0 1 3910
box -6 -8 66 268
use NOR2X1  _762_
timestamp 0
transform 1 0 470 0 -1 3910
box -6 -8 66 268
use NAND2X1  _763_
timestamp 0
transform -1 0 1250 0 1 2870
box -6 -8 66 268
use INVX1  _764_
timestamp 0
transform 1 0 990 0 -1 2870
box -6 -8 46 268
use NAND3X1  _765_
timestamp 0
transform -1 0 570 0 -1 3390
box -6 -8 86 268
use AOI21X1  _766_
timestamp 0
transform 1 0 650 0 -1 3390
box -6 -8 86 268
use INVX1  _767_
timestamp 0
transform 1 0 810 0 -1 3390
box -6 -8 46 268
use NAND3X1  _768_
timestamp 0
transform -1 0 1010 0 -1 3390
box -6 -8 86 268
use INVX1  _769_
timestamp 0
transform 1 0 750 0 1 2870
box -6 -8 46 268
use OAI21X1  _770_
timestamp 0
transform 1 0 870 0 1 2870
box -6 -8 86 268
use NAND3X1  _771_
timestamp 0
transform 1 0 1030 0 1 3390
box -6 -8 86 268
use INVX1  _772_
timestamp 0
transform -1 0 1230 0 1 3390
box -6 -8 46 268
use AOI21X1  _773_
timestamp 0
transform -1 0 950 0 1 3390
box -6 -8 86 268
use NOR2X1  _774_
timestamp 0
transform 1 0 730 0 1 3390
box -6 -8 66 268
use INVX2  _775_
timestamp 0
transform -1 0 3190 0 -1 3910
box -6 -8 46 268
use NOR2X1  _776_
timestamp 0
transform -1 0 1550 0 1 3910
box -6 -8 66 268
use OAI21X1  _777_
timestamp 0
transform -1 0 1110 0 1 2870
box -6 -8 86 268
use NAND2X1  _778_
timestamp 0
transform 1 0 430 0 1 4430
box -6 -8 66 268
use INVX1  _779_
timestamp 0
transform 1 0 570 0 1 4430
box -6 -8 46 268
use NAND3X1  _780_
timestamp 0
transform 1 0 90 0 -1 4430
box -6 -8 86 268
use AOI21X1  _781_
timestamp 0
transform 1 0 90 0 1 4430
box -6 -8 86 268
use INVX1  _782_
timestamp 0
transform 1 0 530 0 -1 4430
box -6 -8 46 268
use NAND3X1  _783_
timestamp 0
transform 1 0 670 0 -1 4430
box -6 -8 86 268
use INVX1  _784_
timestamp 0
transform 1 0 250 0 -1 4430
box -6 -8 46 268
use OAI21X1  _785_
timestamp 0
transform 1 0 370 0 -1 4430
box -6 -8 86 268
use NAND3X1  _786_
timestamp 0
transform -1 0 910 0 -1 4430
box -6 -8 86 268
use AOI21X1  _787_
timestamp 0
transform 1 0 990 0 -1 4430
box -6 -8 86 268
use INVX1  _788_
timestamp 0
transform 1 0 1650 0 -1 4430
box -6 -8 46 268
use NAND3X1  _789_
timestamp 0
transform -1 0 1290 0 1 3910
box -6 -8 86 268
use INVX1  _790_
timestamp 0
transform -1 0 1410 0 1 3910
box -6 -8 46 268
use INVX1  _791_
timestamp 0
transform 1 0 1330 0 -1 4430
box -6 -8 46 268
use OAI21X1  _792_
timestamp 0
transform -1 0 1550 0 -1 4430
box -6 -8 86 268
use NAND3X1  _793_
timestamp 0
transform -1 0 1130 0 1 3910
box -6 -8 86 268
use INVX1  _794_
timestamp 0
transform 1 0 990 0 -1 3910
box -6 -8 46 268
use AOI21X1  _795_
timestamp 0
transform -1 0 970 0 1 3910
box -6 -8 86 268
use NOR2X1  _796_
timestamp 0
transform 1 0 850 0 -1 3910
box -6 -8 66 268
use OAI21X1  _797_
timestamp 0
transform 1 0 1170 0 -1 4430
box -6 -8 86 268
use INVX1  _798_
timestamp 0
transform -1 0 970 0 1 4950
box -6 -8 46 268
use INVX2  _799_
timestamp 0
transform -1 0 3530 0 -1 1830
box -6 -8 46 268
use NAND2X1  _800_
timestamp 0
transform 1 0 2270 0 1 4430
box -6 -8 66 268
use OAI21X1  _801_
timestamp 0
transform 1 0 2370 0 -1 4430
box -6 -8 86 268
use AND2X2  _802_
timestamp 0
transform 1 0 1930 0 -1 3910
box -6 -8 86 268
use NAND2X1  _803_
timestamp 0
transform -1 0 1670 0 -1 3910
box -6 -8 66 268
use AND2X2  _804_
timestamp 0
transform -1 0 1390 0 1 4430
box -6 -8 86 268
use OAI21X1  _805_
timestamp 0
transform -1 0 330 0 1 4430
box -6 -8 86 268
use NAND2X1  _806_
timestamp 0
transform -1 0 870 0 -1 4950
box -6 -8 66 268
use INVX1  _807_
timestamp 0
transform 1 0 910 0 -1 5470
box -6 -8 46 268
use NAND3X1  _808_
timestamp 0
transform 1 0 510 0 1 5470
box -6 -8 86 268
use INVX1  _809_
timestamp 0
transform 1 0 90 0 1 5470
box -6 -8 46 268
use NAND2X1  _810_
timestamp 0
transform -1 0 310 0 -1 5990
box -6 -8 66 268
use NAND2X1  _811_
timestamp 0
transform 1 0 230 0 1 5470
box -6 -8 66 268
use NAND3X1  _812_
timestamp 0
transform -1 0 830 0 -1 5470
box -6 -8 86 268
use NAND2X1  _813_
timestamp 0
transform -1 0 430 0 1 5470
box -6 -8 66 268
use NAND3X1  _814_
timestamp 0
transform -1 0 170 0 -1 5470
box -6 -8 86 268
use NAND3X1  _815_
timestamp 0
transform 1 0 430 0 -1 5470
box -6 -8 86 268
use NAND3X1  _816_
timestamp 0
transform 1 0 470 0 -1 4950
box -6 -8 86 268
use INVX1  _817_
timestamp 0
transform -1 0 130 0 1 4950
box -6 -8 46 268
use AOI21X1  _818_
timestamp 0
transform -1 0 330 0 -1 5470
box -6 -8 86 268
use AOI21X1  _819_
timestamp 0
transform -1 0 670 0 -1 5470
box -6 -8 86 268
use OAI21X1  _820_
timestamp 0
transform -1 0 310 0 1 4950
box -6 -8 86 268
use NAND3X1  _821_
timestamp 0
transform 1 0 950 0 -1 4950
box -6 -8 86 268
use NAND2X1  _822_
timestamp 0
transform 1 0 2070 0 -1 4430
box -6 -8 66 268
use OAI21X1  _823_
timestamp 0
transform -1 0 1850 0 -1 4430
box -6 -8 86 268
use INVX1  _824_
timestamp 0
transform 1 0 710 0 1 4430
box -6 -8 46 268
use AOI21X1  _825_
timestamp 0
transform 1 0 630 0 -1 4950
box -6 -8 86 268
use OAI21X1  _826_
timestamp 0
transform 1 0 990 0 1 4430
box -6 -8 86 268
use NAND2X1  _827_
timestamp 0
transform -1 0 1350 0 -1 4950
box -6 -8 66 268
use NOR2X1  _828_
timestamp 0
transform 1 0 790 0 1 4950
box -6 -8 66 268
use AOI21X1  _829_
timestamp 0
transform -1 0 1210 0 -1 4950
box -6 -8 86 268
use NOR3X1  _830_
timestamp 0
transform 1 0 390 0 1 4950
box -6 -8 166 268
use INVX1  _831_
timestamp 0
transform -1 0 1550 0 -1 5470
box -6 -8 46 268
use OAI21X1  _832_
timestamp 0
transform 1 0 630 0 1 4950
box -6 -8 86 268
use AND2X2  _833_
timestamp 0
transform -1 0 1270 0 -1 5470
box -6 -8 86 268
use INVX1  _834_
timestamp 0
transform 1 0 2150 0 1 4430
box -6 -8 46 268
use OAI21X1  _835_
timestamp 0
transform 1 0 1150 0 1 4430
box -6 -8 86 268
use AOI21X1  _836_
timestamp 0
transform 1 0 670 0 1 5470
box -6 -8 86 268
use OAI21X1  _837_
timestamp 0
transform 1 0 1030 0 -1 5470
box -6 -8 86 268
use NAND3X1  _838_
timestamp 0
transform -1 0 2530 0 -1 5990
box -6 -8 86 268
use AOI21X1  _839_
timestamp 0
transform -1 0 2690 0 -1 5990
box -6 -8 86 268
use INVX1  _840_
timestamp 0
transform -1 0 1830 0 -1 5990
box -6 -8 46 268
use NAND2X1  _841_
timestamp 0
transform -1 0 2650 0 -1 5470
box -6 -8 66 268
use INVX1  _842_
timestamp 0
transform 1 0 2130 0 -1 5470
box -6 -8 46 268
use NAND3X1  _843_
timestamp 0
transform -1 0 1950 0 1 5470
box -6 -8 86 268
use INVX1  _844_
timestamp 0
transform 1 0 1910 0 -1 5990
box -6 -8 46 268
use OAI21X1  _845_
timestamp 0
transform -1 0 2050 0 -1 5470
box -6 -8 86 268
use NAND3X1  _846_
timestamp 0
transform -1 0 1710 0 -1 5470
box -6 -8 86 268
use INVX1  _847_
timestamp 0
transform -1 0 1050 0 1 5470
box -6 -8 46 268
use AOI21X1  _848_
timestamp 0
transform 1 0 850 0 1 5470
box -6 -8 86 268
use OAI21X1  _849_
timestamp 0
transform -1 0 2110 0 1 5470
box -6 -8 86 268
use NAND3X1  _850_
timestamp 0
transform -1 0 1770 0 1 5470
box -6 -8 86 268
use NAND3X1  _851_
timestamp 0
transform -1 0 1450 0 1 5470
box -6 -8 86 268
use NAND2X1  _852_
timestamp 0
transform 1 0 2410 0 -1 3910
box -6 -8 66 268
use AND2X2  _853_
timestamp 0
transform 1 0 2830 0 -1 3910
box -6 -8 86 268
use NAND2X1  _854_
timestamp 0
transform 1 0 2090 0 -1 3910
box -6 -8 66 268
use INVX2  _855_
timestamp 0
transform -1 0 1670 0 1 2870
box -6 -8 46 268
use OAI21X1  _856_
timestamp 0
transform 1 0 1630 0 1 3910
box -6 -8 86 268
use NAND3X1  _857_
timestamp 0
transform -1 0 2050 0 1 3910
box -6 -8 86 268
use INVX1  _858_
timestamp 0
transform -1 0 2330 0 1 3910
box -6 -8 46 268
use INVX1  _859_
timestamp 0
transform 1 0 2710 0 -1 3910
box -6 -8 46 268
use OAI21X1  _860_
timestamp 0
transform -1 0 2630 0 -1 3910
box -6 -8 86 268
use OAI21X1  _861_
timestamp 0
transform 1 0 1770 0 -1 3910
box -6 -8 86 268
use NAND3X1  _862_
timestamp 0
transform -1 0 1870 0 1 3910
box -6 -8 86 268
use NAND2X1  _863_
timestamp 0
transform 1 0 1930 0 -1 4430
box -6 -8 66 268
use NAND3X1  _864_
timestamp 0
transform -1 0 1130 0 1 4950
box -6 -8 86 268
use AOI21X1  _865_
timestamp 0
transform 1 0 1530 0 1 5470
box -6 -8 86 268
use AOI21X1  _866_
timestamp 0
transform -1 0 1890 0 -1 5470
box -6 -8 86 268
use NAND3X1  _867_
timestamp 0
transform 1 0 2130 0 1 3910
box -6 -8 86 268
use NAND3X1  _868_
timestamp 0
transform 1 0 2230 0 -1 3910
box -6 -8 86 268
use NAND2X1  _869_
timestamp 0
transform 1 0 2210 0 -1 4430
box -6 -8 66 268
use OAI21X1  _870_
timestamp 0
transform 1 0 1610 0 -1 4950
box -6 -8 86 268
use NAND3X1  _871_
timestamp 0
transform 1 0 1490 0 1 4430
box -6 -8 86 268
use AOI21X1  _872_
timestamp 0
transform -1 0 910 0 1 4430
box -6 -8 86 268
use OAI21X1  _873_
timestamp 0
transform 1 0 1770 0 -1 4950
box -6 -8 86 268
use NAND3X1  _874_
timestamp 0
transform 1 0 1210 0 1 4950
box -6 -8 86 268
use NAND3X1  _875_
timestamp 0
transform 1 0 2110 0 -1 4950
box -6 -8 86 268
use NAND3X1  _876_
timestamp 0
transform -1 0 2350 0 -1 4950
box -6 -8 86 268
use AOI22X1  _877_
timestamp 0
transform 1 0 1430 0 -1 4950
box -6 -8 106 268
use AOI21X1  _878_
timestamp 0
transform 1 0 1650 0 1 4430
box -6 -8 86 268
use OAI21X1  _879_
timestamp 0
transform 1 0 1930 0 -1 4950
box -6 -8 86 268
use AND2X2  _880_
timestamp 0
transform -1 0 1790 0 1 4950
box -6 -8 86 268
use NAND2X1  _881_
timestamp 0
transform 1 0 2450 0 -1 5470
box -6 -8 66 268
use NAND3X1  _882_
timestamp 0
transform 1 0 1870 0 1 4950
box -6 -8 86 268
use INVX1  _883_
timestamp 0
transform 1 0 2030 0 1 4950
box -6 -8 46 268
use OAI21X1  _884_
timestamp 0
transform -1 0 2050 0 1 4430
box -6 -8 86 268
use INVX1  _885_
timestamp 0
transform 1 0 1330 0 1 2870
box -6 -8 46 268
use NOR2X1  _886_
timestamp 0
transform 1 0 1830 0 1 3390
box -6 -8 66 268
use NAND2X1  _887_
timestamp 0
transform -1 0 2470 0 1 3910
box -6 -8 66 268
use OAI21X1  _888_
timestamp 0
transform 1 0 2530 0 -1 4430
box -6 -8 86 268
use XOR2X1  _889_
timestamp 0
transform 1 0 2770 0 1 4430
box -6 -8 126 268
use OAI21X1  _890_
timestamp 0
transform 1 0 1530 0 1 4950
box -6 -8 86 268
use NAND2X1  _891_
timestamp 0
transform 1 0 2710 0 1 3910
box -6 -8 66 268
use INVX1  _892_
timestamp 0
transform 1 0 2850 0 1 3910
box -6 -8 46 268
use AND2X2  _893_
timestamp 0
transform 1 0 3270 0 -1 3910
box -6 -8 86 268
use NAND2X1  _894_
timestamp 0
transform 1 0 3010 0 -1 3910
box -6 -8 66 268
use INVX1  _895_
timestamp 0
transform 1 0 3430 0 -1 3910
box -6 -8 46 268
use OAI21X1  _896_
timestamp 0
transform 1 0 2550 0 1 3910
box -6 -8 86 268
use NAND3X1  _897_
timestamp 0
transform 1 0 2970 0 1 3910
box -6 -8 86 268
use NAND3X1  _898_
timestamp 0
transform 1 0 2710 0 -1 4430
box -6 -8 86 268
use NAND2X1  _899_
timestamp 0
transform -1 0 3250 0 -1 4430
box -6 -8 66 268
use NAND3X1  _900_
timestamp 0
transform -1 0 3110 0 -1 4430
box -6 -8 86 268
use NAND3X1  _901_
timestamp 0
transform 1 0 2870 0 -1 4430
box -6 -8 86 268
use AND2X2  _902_
timestamp 0
transform 1 0 3630 0 1 4950
box -6 -8 86 268
use OAI21X1  _903_
timestamp 0
transform 1 0 2690 0 1 5470
box -6 -8 86 268
use NAND2X1  _904_
timestamp 0
transform -1 0 4630 0 -1 5470
box -6 -8 66 268
use INVX1  _905_
timestamp 0
transform -1 0 4910 0 -1 5470
box -6 -8 46 268
use NAND3X1  _906_
timestamp 0
transform -1 0 5410 0 1 5470
box -6 -8 86 268
use INVX1  _907_
timestamp 0
transform -1 0 4630 0 -1 5990
box -6 -8 46 268
use NAND2X1  _908_
timestamp 0
transform -1 0 5050 0 -1 5990
box -6 -8 66 268
use NAND2X1  _909_
timestamp 0
transform 1 0 4710 0 -1 5990
box -6 -8 66 268
use NAND3X1  _910_
timestamp 0
transform -1 0 4790 0 -1 5470
box -6 -8 86 268
use NAND2X1  _911_
timestamp 0
transform -1 0 4910 0 -1 5990
box -6 -8 66 268
use NAND3X1  _912_
timestamp 0
transform 1 0 4410 0 -1 5990
box -6 -8 86 268
use NAND3X1  _913_
timestamp 0
transform -1 0 4910 0 1 5470
box -6 -8 86 268
use NAND3X1  _914_
timestamp 0
transform 1 0 4410 0 -1 5470
box -6 -8 86 268
use INVX1  _915_
timestamp 0
transform 1 0 4390 0 1 5470
box -6 -8 46 268
use AOI21X1  _916_
timestamp 0
transform -1 0 4750 0 1 5470
box -6 -8 86 268
use AOI21X1  _917_
timestamp 0
transform -1 0 5090 0 1 5470
box -6 -8 86 268
use OAI21X1  _918_
timestamp 0
transform 1 0 4230 0 1 5470
box -6 -8 86 268
use NAND3X1  _919_
timestamp 0
transform -1 0 3870 0 1 4950
box -6 -8 86 268
use NAND2X1  _920_
timestamp 0
transform 1 0 3630 0 -1 5470
box -6 -8 66 268
use OAI21X1  _921_
timestamp 0
transform -1 0 4150 0 1 5470
box -6 -8 86 268
use NAND3X1  _922_
timestamp 0
transform -1 0 4590 0 1 5470
box -6 -8 86 268
use NAND3X1  _923_
timestamp 0
transform -1 0 3970 0 1 5470
box -6 -8 86 268
use NAND3X1  _924_
timestamp 0
transform 1 0 2990 0 1 4950
box -6 -8 86 268
use AOI21X1  _925_
timestamp 0
transform 1 0 1370 0 1 4950
box -6 -8 86 268
use AOI21X1  _926_
timestamp 0
transform -1 0 3810 0 1 5470
box -6 -8 86 268
use AOI22X1  _927_
timestamp 0
transform 1 0 3770 0 -1 5470
box -6 -8 106 268
use OAI21X1  _928_
timestamp 0
transform 1 0 3470 0 -1 5470
box -6 -8 86 268
use NAND3X1  _929_
timestamp 0
transform -1 0 3170 0 -1 4950
box -6 -8 86 268
use INVX1  _930_
timestamp 0
transform 1 0 2430 0 1 4430
box -6 -8 46 268
use XOR2X1  _931_
timestamp 0
transform -1 0 2670 0 1 4430
box -6 -8 126 268
use OAI21X1  _932_
timestamp 0
transform -1 0 3390 0 -1 5470
box -6 -8 86 268
use NAND3X1  _933_
timestamp 0
transform -1 0 2910 0 1 4950
box -6 -8 86 268
use NAND3X1  _934_
timestamp 0
transform 1 0 2670 0 1 4950
box -6 -8 86 268
use NAND3X1  _935_
timestamp 0
transform -1 0 2850 0 -1 4950
box -6 -8 86 268
use AOI21X1  _936_
timestamp 0
transform 1 0 2430 0 -1 4950
box -6 -8 86 268
use AOI21X1  _937_
timestamp 0
transform 1 0 2510 0 1 4950
box -6 -8 86 268
use AOI21X1  _938_
timestamp 0
transform -1 0 3010 0 -1 4950
box -6 -8 86 268
use OAI21X1  _939_
timestamp 0
transform -1 0 2670 0 -1 4950
box -6 -8 86 268
use NAND3X1  _940_
timestamp 0
transform 1 0 2350 0 1 4950
box -6 -8 86 268
use AOI22X1  _941_
timestamp 0
transform -1 0 2250 0 1 4950
box -6 -8 106 268
use INVX1  _942_
timestamp 0
transform 1 0 3030 0 -1 5470
box -6 -8 46 268
use NAND2X1  _943_
timestamp 0
transform 1 0 2890 0 -1 5470
box -6 -8 66 268
use XOR2X1  _944_
timestamp 0
transform -1 0 2990 0 1 5470
box -6 -8 126 268
use OAI21X1  _945_
timestamp 0
transform 1 0 2730 0 -1 5470
box -6 -8 86 268
use NAND2X1  _946_
timestamp 0
transform -1 0 3030 0 1 4430
box -6 -8 66 268
use AOI21X1  _947_
timestamp 0
transform 1 0 3150 0 1 4950
box -6 -8 86 268
use OAI21X1  _948_
timestamp 0
transform 1 0 3250 0 -1 4950
box -6 -8 86 268
use AND2X2  _949_
timestamp 0
transform 1 0 1390 0 -1 3390
box -6 -8 86 268
use AOI22X1  _950_
timestamp 0
transform 1 0 1450 0 1 2870
box -6 -8 106 268
use AOI21X1  _951_
timestamp 0
transform 1 0 1970 0 1 3390
box -6 -8 86 268
use OAI21X1  _952_
timestamp 0
transform 1 0 3330 0 -1 4430
box -6 -8 86 268
use XNOR2X1  _953_
timestamp 0
transform 1 0 4930 0 -1 4430
box -6 -8 126 268
use AOI21X1  _954_
timestamp 0
transform -1 0 4330 0 -1 5470
box -6 -8 86 268
use OAI21X1  _955_
timestamp 0
transform 1 0 3950 0 -1 5470
box -6 -8 86 268
use NAND2X1  _956_
timestamp 0
transform 1 0 3130 0 1 3910
box -6 -8 66 268
use INVX1  _957_
timestamp 0
transform 1 0 3270 0 1 3910
box -6 -8 46 268
use AND2X2  _958_
timestamp 0
transform 1 0 3390 0 -1 3390
box -6 -8 86 268
use NAND2X1  _959_
timestamp 0
transform -1 0 4250 0 -1 3910
box -6 -8 66 268
use INVX2  _960_
timestamp 0
transform 1 0 2130 0 -1 3390
box -6 -8 46 268
use NAND2X1  _961_
timestamp 0
transform 1 0 3490 0 -1 4430
box -6 -8 66 268
use OAI21X1  _962_
timestamp 0
transform 1 0 3550 0 1 3910
box -6 -8 86 268
use NAND3X1  _963_
timestamp 0
transform 1 0 4030 0 1 3910
box -6 -8 86 268
use OAI21X1  _964_
timestamp 0
transform 1 0 3710 0 -1 3910
box -6 -8 86 268
use OAI21X1  _965_
timestamp 0
transform 1 0 3550 0 -1 3910
box -6 -8 86 268
use NAND3X1  _966_
timestamp 0
transform 1 0 3870 0 -1 3910
box -6 -8 86 268
use NAND2X1  _967_
timestamp 0
transform 1 0 5310 0 -1 4430
box -6 -8 66 268
use AOI21X1  _968_
timestamp 0
transform -1 0 5250 0 1 5470
box -6 -8 86 268
use OAI21X1  _969_
timestamp 0
transform 1 0 4990 0 -1 5470
box -6 -8 86 268
use NAND2X1  _970_
timestamp 0
transform 1 0 5150 0 -1 5470
box -6 -8 66 268
use NAND2X1  _971_
timestamp 0
transform -1 0 5330 0 -1 5990
box -6 -8 66 268
use NAND2X1  _972_
timestamp 0
transform -1 0 5490 0 -1 5990
box -6 -8 66 268
use INVX1  _973_
timestamp 0
transform -1 0 5990 0 1 5470
box -6 -8 46 268
use NAND3X1  _974_
timestamp 0
transform -1 0 5570 0 1 5470
box -6 -8 86 268
use AOI21X1  _975_
timestamp 0
transform -1 0 5370 0 -1 5470
box -6 -8 86 268
use INVX1  _976_
timestamp 0
transform -1 0 5770 0 -1 5990
box -6 -8 46 268
use NAND3X1  _977_
timestamp 0
transform 1 0 5650 0 1 5470
box -6 -8 86 268
use NAND2X1  _978_
timestamp 0
transform -1 0 5870 0 1 5470
box -6 -8 66 268
use AOI21X1  _979_
timestamp 0
transform -1 0 5710 0 1 4950
box -6 -8 86 268
use OAI21X1  _980_
timestamp 0
transform -1 0 5550 0 1 4950
box -6 -8 86 268
use INVX1  _981_
timestamp 0
transform -1 0 5990 0 -1 4950
box -6 -8 46 268
use NAND3X1  _982_
timestamp 0
transform 1 0 5790 0 1 4950
box -6 -8 86 268
use NAND3X1  _983_
timestamp 0
transform 1 0 5450 0 -1 5470
box -6 -8 86 268
use NAND3X1  _984_
timestamp 0
transform -1 0 5850 0 -1 4950
box -6 -8 86 268
use AOI21X1  _985_
timestamp 0
transform -1 0 5370 0 -1 4950
box -6 -8 86 268
use NAND3X1  _986_
timestamp 0
transform -1 0 5790 0 1 4430
box -6 -8 86 268
use OAI21X1  _987_
timestamp 0
transform 1 0 5610 0 -1 4950
box -6 -8 86 268
use AOI22X1  _988_
timestamp 0
transform 1 0 5510 0 1 4430
box -6 -8 106 268
use OAI21X1  _989_
timestamp 0
transform -1 0 5270 0 1 4430
box -6 -8 86 268
use INVX1  _990_
timestamp 0
transform 1 0 4130 0 -1 5470
box -6 -8 46 268
use AOI21X1  _991_
timestamp 0
transform 1 0 4230 0 1 4950
box -6 -8 86 268
use AND2X2  _992_
timestamp 0
transform -1 0 5590 0 1 3910
box -6 -8 86 268
use NAND3X1  _993_
timestamp 0
transform -1 0 5530 0 -1 4430
box -6 -8 86 268
use NAND3X1  _994_
timestamp 0
transform -1 0 5530 0 -1 4950
box -6 -8 86 268
use NAND3X1  _995_
timestamp 0
transform -1 0 5030 0 -1 4950
box -6 -8 86 268
use AOI21X1  _996_
timestamp 0
transform -1 0 4930 0 1 4430
box -6 -8 86 268
use XOR2X1  _997_
timestamp 0
transform 1 0 4710 0 -1 4430
box -6 -8 126 268
use NAND3X1  _998_
timestamp 0
transform -1 0 5390 0 1 4950
box -6 -8 86 268
use OAI21X1  _999_
timestamp 0
transform -1 0 5210 0 -1 4950
box -6 -8 86 268
use AOI21X1  _1000_
timestamp 0
transform -1 0 4950 0 1 4950
box -6 -8 86 268
use OAI21X1  _1001_
timestamp 0
transform -1 0 4690 0 -1 4950
box -6 -8 86 268
use INVX1  _1002_
timestamp 0
transform -1 0 3450 0 -1 4950
box -6 -8 46 268
use AOI21X1  _1003_
timestamp 0
transform 1 0 3530 0 -1 4950
box -6 -8 86 268
use NAND3X1  _1004_
timestamp 0
transform -1 0 4850 0 -1 4950
box -6 -8 86 268
use NAND3X1  _1005_
timestamp 0
transform -1 0 5110 0 1 4430
box -6 -8 86 268
use NAND3X1  _1006_
timestamp 0
transform -1 0 4430 0 1 4430
box -6 -8 86 268
use AOI21X1  _1007_
timestamp 0
transform -1 0 3930 0 -1 4950
box -6 -8 86 268
use INVX1  _1008_
timestamp 0
transform 1 0 4170 0 -1 4950
box -6 -8 46 268
use NAND3X1  _1009_
timestamp 0
transform -1 0 4770 0 1 4430
box -6 -8 86 268
use OAI21X1  _1010_
timestamp 0
transform -1 0 4530 0 -1 4950
box -6 -8 86 268
use AOI21X1  _1011_
timestamp 0
transform -1 0 4370 0 -1 4950
box -6 -8 86 268
use OAI21X1  _1012_
timestamp 0
transform -1 0 3770 0 -1 4950
box -6 -8 86 268
use INVX1  _1013_
timestamp 0
transform 1 0 3950 0 1 4950
box -6 -8 46 268
use NAND3X1  _1014_
timestamp 0
transform -1 0 4490 0 1 4950
box -6 -8 86 268
use NAND3X1  _1015_
timestamp 0
transform 1 0 4010 0 -1 4950
box -6 -8 86 268
use NAND3X1  _1016_
timestamp 0
transform -1 0 4150 0 1 4950
box -6 -8 86 268
use NAND3X1  _1017_
timestamp 0
transform 1 0 3470 0 1 4950
box -6 -8 86 268
use INVX1  _1018_
timestamp 0
transform -1 0 3790 0 1 4430
box -6 -8 46 268
use AOI21X1  _1019_
timestamp 0
transform -1 0 3390 0 1 4950
box -6 -8 86 268
use NOR2X1  _1020_
timestamp 0
transform 1 0 3570 0 1 5470
box -6 -8 66 268
use NAND2X1  _1021_
timestamp 0
transform -1 0 3930 0 1 4430
box -6 -8 66 268
use AOI21X1  _1022_
timestamp 0
transform -1 0 4590 0 1 4430
box -6 -8 86 268
use OAI21X1  _1023_
timestamp 0
transform 1 0 4190 0 1 4430
box -6 -8 86 268
use NAND2X1  _1024_
timestamp 0
transform 1 0 4290 0 -1 4430
box -6 -8 66 268
use INVX1  _1025_
timestamp 0
transform 1 0 4430 0 -1 4430
box -6 -8 46 268
use AOI21X1  _1026_
timestamp 0
transform -1 0 5430 0 1 4430
box -6 -8 86 268
use OAI21X1  _1027_
timestamp 0
transform 1 0 5130 0 -1 4430
box -6 -8 86 268
use NAND2X1  _1028_
timestamp 0
transform -1 0 2210 0 1 3390
box -6 -8 66 268
use INVX1  _1029_
timestamp 0
transform 1 0 3570 0 1 3390
box -6 -8 46 268
use NAND2X1  _1030_
timestamp 0
transform 1 0 2390 0 -1 3390
box -6 -8 66 268
use INVX1  _1031_
timestamp 0
transform 1 0 2730 0 -1 3390
box -6 -8 46 268
use AND2X2  _1032_
timestamp 0
transform -1 0 1990 0 1 2870
box -6 -8 86 268
use NAND2X1  _1033_
timestamp 0
transform -1 0 2310 0 -1 3390
box -6 -8 66 268
use NAND2X1  _1034_
timestamp 0
transform -1 0 1610 0 -1 3390
box -6 -8 66 268
use OAI21X1  _1035_
timestamp 0
transform 1 0 1830 0 -1 3390
box -6 -8 86 268
use NAND3X1  _1036_
timestamp 0
transform 1 0 2850 0 -1 3390
box -6 -8 86 268
use NAND2X1  _1037_
timestamp 0
transform 1 0 2090 0 1 2870
box -6 -8 66 268
use NAND2X1  _1038_
timestamp 0
transform -1 0 2350 0 1 3390
box -6 -8 66 268
use NAND2X1  _1039_
timestamp 0
transform 1 0 1990 0 -1 3390
box -6 -8 66 268
use NAND3X1  _1040_
timestamp 0
transform 1 0 2430 0 1 3390
box -6 -8 86 268
use NAND2X1  _1041_
timestamp 0
transform 1 0 4530 0 -1 3910
box -6 -8 66 268
use AND2X2  _1042_
timestamp 0
transform 1 0 3850 0 1 3910
box -6 -8 86 268
use OAI21X1  _1043_
timestamp 0
transform 1 0 4030 0 -1 3910
box -6 -8 86 268
use NAND3X1  _1044_
timestamp 0
transform 1 0 3410 0 1 3390
box -6 -8 86 268
use AOI21X1  _1045_
timestamp 0
transform 1 0 2590 0 1 3390
box -6 -8 86 268
use AOI22X1  _1046_
timestamp 0
transform 1 0 2550 0 -1 3390
box -6 -8 106 268
use NOR2X1  _1047_
timestamp 0
transform 1 0 3710 0 1 3910
box -6 -8 66 268
use AOI21X1  _1048_
timestamp 0
transform -1 0 3470 0 1 3910
box -6 -8 86 268
use OAI21X1  _1049_
timestamp 0
transform 1 0 2750 0 1 3390
box -6 -8 86 268
use NAND3X1  _1050_
timestamp 0
transform 1 0 3690 0 1 3390
box -6 -8 86 268
use NAND3X1  _1051_
timestamp 0
transform 1 0 3090 0 1 3390
box -6 -8 86 268
use OAI21X1  _1052_
timestamp 0
transform 1 0 2910 0 1 3390
box -6 -8 86 268
use NAND3X1  _1053_
timestamp 0
transform 1 0 3250 0 1 3390
box -6 -8 86 268
use AND2X2  _1054_
timestamp 0
transform 1 0 4590 0 1 3390
box -6 -8 86 268
use AOI21X1  _1055_
timestamp 0
transform 1 0 5890 0 1 4430
box -6 -8 86 268
use OAI21X1  _1056_
timestamp 0
transform -1 0 5990 0 -1 4430
box -6 -8 86 268
use NAND2X1  _1057_
timestamp 0
transform 1 0 3850 0 1 3390
box -6 -8 66 268
use INVX1  _1058_
timestamp 0
transform 1 0 3890 0 -1 3390
box -6 -8 46 268
use AND2X2  _1059_
timestamp 0
transform -1 0 4570 0 -1 3390
box -6 -8 86 268
use AND2X2  _1060_
timestamp 0
transform -1 0 4230 0 -1 2350
box -6 -8 86 268
use NAND2X1  _1061_
timestamp 0
transform -1 0 3830 0 1 2870
box -6 -8 66 268
use NAND2X1  _1062_
timestamp 0
transform 1 0 4310 0 1 3390
box -6 -8 66 268
use OAI21X1  _1063_
timestamp 0
transform 1 0 3730 0 -1 3390
box -6 -8 86 268
use NAND3X1  _1064_
timestamp 0
transform 1 0 4030 0 -1 3390
box -6 -8 86 268
use NAND2X1  _1065_
timestamp 0
transform 1 0 4350 0 -1 3390
box -6 -8 66 268
use OAI21X1  _1066_
timestamp 0
transform 1 0 3610 0 1 2870
box -6 -8 86 268
use NAND3X1  _1067_
timestamp 0
transform 1 0 4190 0 -1 3390
box -6 -8 86 268
use AND2X2  _1068_
timestamp 0
transform -1 0 5030 0 -1 3390
box -6 -8 86 268
use AOI21X1  _1069_
timestamp 0
transform 1 0 5630 0 -1 5470
box -6 -8 86 268
use OAI21X1  _1070_
timestamp 0
transform 1 0 5790 0 -1 5470
box -6 -8 86 268
use NAND2X1  _1071_
timestamp 0
transform -1 0 5450 0 -1 2350
box -6 -8 66 268
use INVX1  _1072_
timestamp 0
transform -1 0 5310 0 -1 2870
box -6 -8 46 268
use NAND3X1  _1073_
timestamp 0
transform -1 0 5930 0 -1 2350
box -6 -8 86 268
use INVX1  _1074_
timestamp 0
transform -1 0 5710 0 1 2350
box -6 -8 46 268
use NAND2X1  _1075_
timestamp 0
transform -1 0 5650 0 -1 270
box -6 -8 66 268
use NAND2X1  _1076_
timestamp 0
transform -1 0 5570 0 1 2350
box -6 -8 66 268
use NAND3X1  _1077_
timestamp 0
transform -1 0 5470 0 -1 2870
box -6 -8 86 268
use NAND2X1  _1078_
timestamp 0
transform 1 0 5810 0 1 2350
box -6 -8 66 268
use NAND3X1  _1079_
timestamp 0
transform 1 0 5710 0 -1 2870
box -6 -8 86 268
use NAND3X1  _1080_
timestamp 0
transform -1 0 5790 0 1 2870
box -6 -8 86 268
use NAND3X1  _1081_
timestamp 0
transform -1 0 5630 0 1 2870
box -6 -8 86 268
use INVX1  _1082_
timestamp 0
transform 1 0 5770 0 -1 3390
box -6 -8 46 268
use AOI21X1  _1083_
timestamp 0
transform 1 0 5890 0 1 2870
box -6 -8 86 268
use AOI21X1  _1084_
timestamp 0
transform 1 0 5550 0 -1 2870
box -6 -8 86 268
use OAI21X1  _1085_
timestamp 0
transform -1 0 5970 0 -1 3390
box -6 -8 86 268
use NAND3X1  _1086_
timestamp 0
transform 1 0 5110 0 -1 3390
box -6 -8 86 268
use NAND2X1  _1087_
timestamp 0
transform 1 0 5290 0 -1 3390
box -6 -8 66 268
use OAI21X1  _1088_
timestamp 0
transform -1 0 5990 0 1 3390
box -6 -8 86 268
use NAND3X1  _1089_
timestamp 0
transform 1 0 5610 0 -1 3390
box -6 -8 86 268
use NAND3X1  _1090_
timestamp 0
transform -1 0 5670 0 1 3390
box -6 -8 86 268
use NAND3X1  _1091_
timestamp 0
transform -1 0 5510 0 1 3390
box -6 -8 86 268
use INVX1  _1092_
timestamp 0
transform 1 0 5790 0 -1 4430
box -6 -8 46 268
use AOI21X1  _1093_
timestamp 0
transform 1 0 5610 0 -1 4430
box -6 -8 86 268
use AOI21X1  _1094_
timestamp 0
transform 1 0 5750 0 1 3390
box -6 -8 86 268
use AOI22X1  _1095_
timestamp 0
transform 1 0 5430 0 -1 3390
box -6 -8 106 268
use OAI21X1  _1096_
timestamp 0
transform -1 0 5870 0 -1 3910
box -6 -8 86 268
use NAND3X1  _1097_
timestamp 0
transform 1 0 4930 0 1 3390
box -6 -8 86 268
use NAND2X1  _1098_
timestamp 0
transform -1 0 4510 0 1 3390
box -6 -8 66 268
use OAI21X1  _1099_
timestamp 0
transform 1 0 5830 0 1 3910
box -6 -8 86 268
use NAND3X1  _1100_
timestamp 0
transform 1 0 5450 0 -1 3910
box -6 -8 86 268
use NAND3X1  _1101_
timestamp 0
transform -1 0 5710 0 -1 3910
box -6 -8 86 268
use NAND3X1  _1102_
timestamp 0
transform -1 0 5370 0 -1 3910
box -6 -8 86 268
use INVX1  _1103_
timestamp 0
transform -1 0 5230 0 1 4950
box -6 -8 46 268
use AOI21X1  _1104_
timestamp 0
transform 1 0 5030 0 1 4950
box -6 -8 86 268
use AOI21X1  _1105_
timestamp 0
transform -1 0 5750 0 1 3910
box -6 -8 86 268
use AOI21X1  _1106_
timestamp 0
transform 1 0 5110 0 1 3390
box -6 -8 86 268
use OAI21X1  _1107_
timestamp 0
transform -1 0 5270 0 1 3910
box -6 -8 86 268
use NAND3X1  _1108_
timestamp 0
transform -1 0 4430 0 1 3910
box -6 -8 86 268
use OAI21X1  _1109_
timestamp 0
transform -1 0 5430 0 1 3910
box -6 -8 86 268
use NAND3X1  _1110_
timestamp 0
transform -1 0 5110 0 1 3910
box -6 -8 86 268
use NAND3X1  _1111_
timestamp 0
transform -1 0 4930 0 1 3910
box -6 -8 86 268
use NAND3X1  _1112_
timestamp 0
transform -1 0 4270 0 1 3910
box -6 -8 86 268
use INVX1  _1113_
timestamp 0
transform 1 0 4730 0 1 4950
box -6 -8 46 268
use AOI21X1  _1114_
timestamp 0
transform 1 0 4570 0 1 4950
box -6 -8 86 268
use AOI21X1  _1115_
timestamp 0
transform -1 0 4770 0 1 3910
box -6 -8 86 268
use AOI21X1  _1116_
timestamp 0
transform 1 0 4510 0 1 3910
box -6 -8 86 268
use OAI21X1  _1117_
timestamp 0
transform -1 0 4630 0 -1 4430
box -6 -8 86 268
use NAND2X1  _1118_
timestamp 0
transform 1 0 4150 0 -1 4430
box -6 -8 66 268
use XNOR2X1  _1119_
timestamp 0
transform -1 0 3750 0 -1 4430
box -6 -8 126 268
use INVX1  _1120_
timestamp 0
transform -1 0 4070 0 -1 4430
box -6 -8 46 268
use AND2X2  _1121_
timestamp 0
transform -1 0 4090 0 1 4430
box -6 -8 86 268
use OAI22X1  _1122_
timestamp 0
transform -1 0 3930 0 -1 4430
box -6 -8 106 268
use INVX1  _1123_
timestamp 0
transform -1 0 4890 0 -1 3910
box -6 -8 46 268
use AOI21X1  _1124_
timestamp 0
transform 1 0 4690 0 -1 3910
box -6 -8 86 268
use NAND2X1  _1125_
timestamp 0
transform 1 0 3990 0 1 3390
box -6 -8 66 268
use INVX1  _1126_
timestamp 0
transform 1 0 4350 0 -1 2870
box -6 -8 46 268
use AOI21X1  _1127_
timestamp 0
transform -1 0 5350 0 1 3390
box -6 -8 86 268
use OAI21X1  _1128_
timestamp 0
transform 1 0 4750 0 1 3390
box -6 -8 86 268
use OAI21X1  _1129_
timestamp 0
transform 1 0 3030 0 -1 3390
box -6 -8 86 268
use NAND2X1  _1130_
timestamp 0
transform 1 0 2230 0 1 2870
box -6 -8 66 268
use INVX1  _1131_
timestamp 0
transform 1 0 2550 0 -1 2870
box -6 -8 46 268
use AND2X2  _1132_
timestamp 0
transform 1 0 2250 0 -1 2870
box -6 -8 86 268
use AND2X2  _1133_
timestamp 0
transform 1 0 2090 0 -1 2870
box -6 -8 86 268
use NAND2X1  _1134_
timestamp 0
transform 1 0 2410 0 -1 2870
box -6 -8 66 268
use INVX1  _1135_
timestamp 0
transform -1 0 1410 0 -1 2870
box -6 -8 46 268
use NAND2X1  _1136_
timestamp 0
transform -1 0 1810 0 1 2870
box -6 -8 66 268
use OAI21X1  _1137_
timestamp 0
transform 1 0 1750 0 -1 2870
box -6 -8 86 268
use NAND3X1  _1138_
timestamp 0
transform 1 0 2850 0 -1 2870
box -6 -8 86 268
use OAI21X1  _1139_
timestamp 0
transform -1 0 2450 0 1 2870
box -6 -8 86 268
use OAI21X1  _1140_
timestamp 0
transform 1 0 1910 0 -1 2870
box -6 -8 86 268
use NAND3X1  _1141_
timestamp 0
transform 1 0 2690 0 1 2870
box -6 -8 86 268
use AOI22X1  _1142_
timestamp 0
transform -1 0 4430 0 -1 3910
box -6 -8 106 268
use OAI21X1  _1143_
timestamp 0
transform -1 0 4230 0 1 3390
box -6 -8 86 268
use NAND3X1  _1144_
timestamp 0
transform 1 0 3170 0 -1 2870
box -6 -8 86 268
use AOI21X1  _1145_
timestamp 0
transform 1 0 2530 0 1 2870
box -6 -8 86 268
use AOI21X1  _1146_
timestamp 0
transform 1 0 2670 0 -1 2870
box -6 -8 86 268
use NAND2X1  _1147_
timestamp 0
transform -1 0 4530 0 -1 2350
box -6 -8 66 268
use INVX1  _1148_
timestamp 0
transform 1 0 3490 0 1 2870
box -6 -8 46 268
use AOI22X1  _1149_
timestamp 0
transform 1 0 3550 0 -1 3390
box -6 -8 106 268
use OAI21X1  _1150_
timestamp 0
transform 1 0 2850 0 1 2870
box -6 -8 86 268
use NAND3X1  _1151_
timestamp 0
transform -1 0 3090 0 -1 2870
box -6 -8 86 268
use AND2X2  _1152_
timestamp 0
transform 1 0 3210 0 -1 3390
box -6 -8 86 268
use NAND3X1  _1153_
timestamp 0
transform 1 0 3170 0 1 2870
box -6 -8 86 268
use OAI21X1  _1154_
timestamp 0
transform 1 0 3010 0 1 2870
box -6 -8 86 268
use NAND3X1  _1155_
timestamp 0
transform 1 0 3330 0 1 2870
box -6 -8 86 268
use NAND2X1  _1156_
timestamp 0
transform -1 0 3770 0 -1 2870
box -6 -8 66 268
use AOI21X1  _1157_
timestamp 0
transform -1 0 5470 0 1 2870
box -6 -8 86 268
use OAI21X1  _1158_
timestamp 0
transform -1 0 5290 0 1 2870
box -6 -8 86 268
use NAND2X1  _1159_
timestamp 0
transform -1 0 4050 0 -1 2350
box -6 -8 66 268
use INVX1  _1160_
timestamp 0
transform -1 0 3990 0 1 1830
box -6 -8 46 268
use AND2X2  _1161_
timestamp 0
transform 1 0 2970 0 1 1830
box -6 -8 86 268
use NAND2X1  _1162_
timestamp 0
transform -1 0 3710 0 1 1830
box -6 -8 66 268
use INVX1  _1163_
timestamp 0
transform -1 0 1710 0 -1 1830
box -6 -8 46 268
use OAI21X1  _1164_
timestamp 0
transform 1 0 3290 0 1 1830
box -6 -8 86 268
use NAND3X1  _1165_
timestamp 0
transform 1 0 3790 0 1 1830
box -6 -8 86 268
use NAND2X1  _1166_
timestamp 0
transform 1 0 4250 0 1 1830
box -6 -8 66 268
use NAND3X1  _1167_
timestamp 0
transform 1 0 4390 0 1 1830
box -6 -8 86 268
use NAND3X1  _1168_
timestamp 0
transform 1 0 4550 0 1 1830
box -6 -8 86 268
use NAND3X1  _1169_
timestamp 0
transform 1 0 4710 0 1 1830
box -6 -8 86 268
use NAND2X1  _1170_
timestamp 0
transform 1 0 4890 0 1 1830
box -6 -8 66 268
use AOI21X1  _1171_
timestamp 0
transform -1 0 5770 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1172_
timestamp 0
transform -1 0 5610 0 -1 2350
box -6 -8 86 268
use NAND3X1  _1173_
timestamp 0
transform -1 0 5930 0 1 1830
box -6 -8 86 268
use INVX1  _1174_
timestamp 0
transform 1 0 5870 0 -1 2870
box -6 -8 46 268
use AOI21X1  _1175_
timestamp 0
transform 1 0 5690 0 1 1830
box -6 -8 86 268
use OAI21X1  _1176_
timestamp 0
transform -1 0 5590 0 1 1830
box -6 -8 86 268
use NOR2X1  _1177_
timestamp 0
transform -1 0 5630 0 -1 5990
box -6 -8 66 268
use NAND3X1  _1178_
timestamp 0
transform -1 0 5430 0 1 1830
box -6 -8 86 268
use AOI21X1  _1179_
timestamp 0
transform -1 0 5110 0 1 1830
box -6 -8 86 268
use NAND2X1  _1180_
timestamp 0
transform 1 0 5810 0 1 1310
box -6 -8 66 268
use INVX1  _1181_
timestamp 0
transform 1 0 5850 0 -1 5990
box -6 -8 46 268
use NAND2X1  _1182_
timestamp 0
transform -1 0 5890 0 -1 1830
box -6 -8 66 268
use NAND3X1  _1183_
timestamp 0
transform -1 0 5590 0 -1 1830
box -6 -8 86 268
use AOI22X1  _1184_
timestamp 0
transform 1 0 4990 0 -1 1830
box -6 -8 106 268
use OAI21X1  _1185_
timestamp 0
transform 1 0 5070 0 -1 2350
box -6 -8 86 268
use INVX1  _1186_
timestamp 0
transform -1 0 5130 0 1 2870
box -6 -8 46 268
use AOI21X1  _1187_
timestamp 0
transform -1 0 5010 0 1 2870
box -6 -8 86 268
use AND2X2  _1188_
timestamp 0
transform 1 0 4810 0 -1 1830
box -6 -8 86 268
use NAND3X1  _1189_
timestamp 0
transform 1 0 5190 0 -1 1830
box -6 -8 86 268
use NAND3X1  _1190_
timestamp 0
transform 1 0 5190 0 1 1830
box -6 -8 86 268
use NAND3X1  _1191_
timestamp 0
transform -1 0 5090 0 1 2350
box -6 -8 86 268
use AOI21X1  _1192_
timestamp 0
transform -1 0 5030 0 -1 2870
box -6 -8 86 268
use AND2X2  _1193_
timestamp 0
transform 1 0 3870 0 -1 2870
box -6 -8 86 268
use NAND3X1  _1194_
timestamp 0
transform 1 0 5230 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1195_
timestamp 0
transform -1 0 4990 0 -1 2350
box -6 -8 86 268
use AOI21X1  _1196_
timestamp 0
transform -1 0 4770 0 1 2350
box -6 -8 86 268
use OAI21X1  _1197_
timestamp 0
transform 1 0 4630 0 -1 2870
box -6 -8 86 268
use INVX1  _1198_
timestamp 0
transform -1 0 4870 0 -1 3390
box -6 -8 46 268
use AOI21X1  _1199_
timestamp 0
transform -1 0 4730 0 -1 3390
box -6 -8 86 268
use NAND3X1  _1200_
timestamp 0
transform -1 0 4930 0 1 2350
box -6 -8 86 268
use NAND3X1  _1201_
timestamp 0
transform 1 0 5110 0 -1 2870
box -6 -8 86 268
use NAND3X1  _1202_
timestamp 0
transform -1 0 4690 0 1 2870
box -6 -8 86 268
use AOI21X1  _1203_
timestamp 0
transform -1 0 4370 0 1 2870
box -6 -8 86 268
use NAND3X1  _1204_
timestamp 0
transform -1 0 4850 0 1 2870
box -6 -8 86 268
use OAI21X1  _1205_
timestamp 0
transform -1 0 4550 0 -1 2870
box -6 -8 86 268
use AOI21X1  _1206_
timestamp 0
transform -1 0 4110 0 -1 2870
box -6 -8 86 268
use OAI21X1  _1207_
timestamp 0
transform 1 0 3930 0 1 2870
box -6 -8 86 268
use AOI21X1  _1208_
timestamp 0
transform -1 0 5210 0 -1 3910
box -6 -8 86 268
use OAI21X1  _1209_
timestamp 0
transform 1 0 4970 0 -1 3910
box -6 -8 86 268
use NAND3X1  _1210_
timestamp 0
transform -1 0 4270 0 -1 2870
box -6 -8 86 268
use NAND3X1  _1211_
timestamp 0
transform -1 0 4530 0 1 2870
box -6 -8 86 268
use NAND3X1  _1212_
timestamp 0
transform -1 0 4190 0 1 2870
box -6 -8 86 268
use NAND2X1  _1213_
timestamp 0
transform 1 0 4110 0 1 2350
box -6 -8 66 268
use XNOR2X1  _1214_
timestamp 0
transform -1 0 3370 0 1 2350
box -6 -8 126 268
use INVX1  _1215_
timestamp 0
transform 1 0 3810 0 1 2350
box -6 -8 46 268
use OAI21X1  _1216_
timestamp 0
transform 1 0 3950 0 1 2350
box -6 -8 86 268
use AOI21X1  _1217_
timestamp 0
transform -1 0 4870 0 -1 2870
box -6 -8 86 268
use OAI21X1  _1218_
timestamp 0
transform 1 0 4530 0 1 2350
box -6 -8 86 268
use NAND2X1  _1219_
timestamp 0
transform 1 0 3330 0 -1 2870
box -6 -8 66 268
use AOI21X1  _1220_
timestamp 0
transform 1 0 5170 0 1 2350
box -6 -8 86 268
use OAI21X1  _1221_
timestamp 0
transform 1 0 5350 0 1 2350
box -6 -8 86 268
use NAND2X1  _1222_
timestamp 0
transform 1 0 2070 0 1 2350
box -6 -8 66 268
use OAI21X1  _1223_
timestamp 0
transform 1 0 2930 0 1 2350
box -6 -8 86 268
use NAND2X1  _1224_
timestamp 0
transform -1 0 2410 0 1 2350
box -6 -8 66 268
use AOI22X1  _1225_
timestamp 0
transform 1 0 2110 0 -1 2350
box -6 -8 106 268
use NAND2X1  _1226_
timestamp 0
transform 1 0 1690 0 -1 2350
box -6 -8 66 268
use NOR2X1  _1227_
timestamp 0
transform -1 0 1890 0 -1 2350
box -6 -8 66 268
use OAI21X1  _1228_
timestamp 0
transform 1 0 2670 0 -1 2350
box -6 -8 86 268
use INVX1  _1229_
timestamp 0
transform 1 0 2830 0 1 1830
box -6 -8 46 268
use INVX1  _1230_
timestamp 0
transform 1 0 2310 0 -1 2350
box -6 -8 46 268
use AND2X2  _1231_
timestamp 0
transform -1 0 2570 0 1 2350
box -6 -8 86 268
use NAND2X1  _1232_
timestamp 0
transform -1 0 2710 0 1 2350
box -6 -8 66 268
use NAND3X1  _1233_
timestamp 0
transform 1 0 2990 0 -1 2350
box -6 -8 86 268
use AND2X2  _1234_
timestamp 0
transform 1 0 4070 0 1 1830
box -6 -8 86 268
use OAI21X1  _1235_
timestamp 0
transform -1 0 3910 0 -1 2350
box -6 -8 86 268
use NAND3X1  _1236_
timestamp 0
transform 1 0 3650 0 -1 2350
box -6 -8 86 268
use AOI21X1  _1237_
timestamp 0
transform 1 0 2830 0 -1 2350
box -6 -8 86 268
use NOR3X1  _1238_
timestamp 0
transform 1 0 2430 0 -1 2350
box -6 -8 166 268
use AOI22X1  _1239_
timestamp 0
transform -1 0 3570 0 1 1830
box -6 -8 106 268
use OAI21X1  _1240_
timestamp 0
transform 1 0 3150 0 -1 2350
box -6 -8 86 268
use NAND3X1  _1241_
timestamp 0
transform 1 0 3130 0 1 1830
box -6 -8 86 268
use AND2X2  _1242_
timestamp 0
transform 1 0 3090 0 1 2350
box -6 -8 86 268
use NAND3X1  _1243_
timestamp 0
transform -1 0 3570 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1244_
timestamp 0
transform 1 0 3330 0 -1 2350
box -6 -8 86 268
use NAND3X1  _1245_
timestamp 0
transform 1 0 3450 0 1 2350
box -6 -8 86 268
use AND2X2  _1246_
timestamp 0
transform 1 0 4950 0 1 790
box -6 -8 86 268
use NOR2X1  _1247_
timestamp 0
transform -1 0 5710 0 1 1310
box -6 -8 66 268
use OAI21X1  _1248_
timestamp 0
transform 1 0 5490 0 1 1310
box -6 -8 86 268
use NAND2X1  _1249_
timestamp 0
transform -1 0 3690 0 -1 1830
box -6 -8 66 268
use INVX1  _1250_
timestamp 0
transform 1 0 3170 0 -1 1310
box -6 -8 46 268
use AND2X2  _1251_
timestamp 0
transform -1 0 2910 0 -1 1830
box -6 -8 86 268
use NAND2X1  _1252_
timestamp 0
transform -1 0 3090 0 -1 1310
box -6 -8 66 268
use INVX1  _1253_
timestamp 0
transform -1 0 1150 0 -1 1830
box -6 -8 46 268
use OAI22X1  _1254_
timestamp 0
transform 1 0 2990 0 -1 1830
box -6 -8 106 268
use NAND3X1  _1255_
timestamp 0
transform 1 0 3290 0 -1 1310
box -6 -8 86 268
use OAI21X1  _1256_
timestamp 0
transform 1 0 3170 0 -1 1830
box -6 -8 86 268
use OAI21X1  _1257_
timestamp 0
transform 1 0 3330 0 -1 1830
box -6 -8 86 268
use NAND3X1  _1258_
timestamp 0
transform 1 0 3570 0 1 1310
box -6 -8 86 268
use XNOR2X1  _1259_
timestamp 0
transform -1 0 5890 0 -1 1310
box -6 -8 126 268
use NAND3X1  _1260_
timestamp 0
transform -1 0 5410 0 -1 1310
box -6 -8 86 268
use NAND2X1  _1261_
timestamp 0
transform -1 0 5550 0 -1 1310
box -6 -8 66 268
use INVX1  _1262_
timestamp 0
transform 1 0 5910 0 1 790
box -6 -8 46 268
use NAND2X1  _1263_
timestamp 0
transform -1 0 5810 0 1 790
box -6 -8 66 268
use NAND3X1  _1264_
timestamp 0
transform -1 0 5730 0 1 270
box -6 -8 86 268
use AOI21X1  _1265_
timestamp 0
transform -1 0 5750 0 -1 1830
box -6 -8 86 268
use AOI21X1  _1266_
timestamp 0
transform 1 0 5350 0 -1 1830
box -6 -8 86 268
use NAND2X1  _1267_
timestamp 0
transform -1 0 5890 0 1 270
box -6 -8 66 268
use NAND2X1  _1268_
timestamp 0
transform 1 0 5810 0 -1 790
box -6 -8 66 268
use NAND3X1  _1269_
timestamp 0
transform -1 0 5590 0 -1 790
box -6 -8 86 268
use NAND2X1  _1270_
timestamp 0
transform 1 0 5110 0 1 790
box -6 -8 66 268
use NOR2X1  _1271_
timestamp 0
transform 1 0 5730 0 -1 270
box -6 -8 66 268
use AOI21X1  _1272_
timestamp 0
transform -1 0 5570 0 1 270
box -6 -8 86 268
use OAI21X1  _1273_
timestamp 0
transform -1 0 5390 0 1 270
box -6 -8 86 268
use NAND3X1  _1274_
timestamp 0
transform -1 0 5090 0 -1 1310
box -6 -8 86 268
use INVX1  _1275_
timestamp 0
transform -1 0 4830 0 -1 2350
box -6 -8 46 268
use AOI21X1  _1276_
timestamp 0
transform 1 0 4630 0 -1 2350
box -6 -8 86 268
use NAND2X1  _1277_
timestamp 0
transform 1 0 5670 0 -1 790
box -6 -8 66 268
use NAND3X1  _1278_
timestamp 0
transform -1 0 5670 0 1 790
box -6 -8 86 268
use AOI21X1  _1279_
timestamp 0
transform -1 0 5510 0 1 790
box -6 -8 86 268
use AOI22X1  _1280_
timestamp 0
transform 1 0 5250 0 1 790
box -6 -8 106 268
use OAI21X1  _1281_
timestamp 0
transform -1 0 4910 0 1 1310
box -6 -8 86 268
use NAND3X1  _1282_
timestamp 0
transform -1 0 4730 0 -1 1830
box -6 -8 86 268
use INVX1  _1283_
timestamp 0
transform 1 0 4690 0 1 1310
box -6 -8 46 268
use OAI21X1  _1284_
timestamp 0
transform 1 0 5330 0 1 1310
box -6 -8 86 268
use NAND3X1  _1285_
timestamp 0
transform -1 0 4930 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1286_
timestamp 0
transform -1 0 5070 0 1 1310
box -6 -8 86 268
use NAND3X1  _1287_
timestamp 0
transform -1 0 4570 0 -1 1830
box -6 -8 86 268
use INVX1  _1288_
timestamp 0
transform 1 0 4250 0 1 2350
box -6 -8 46 268
use AOI21X1  _1289_
timestamp 0
transform 1 0 4370 0 1 2350
box -6 -8 86 268
use AOI21X1  _1290_
timestamp 0
transform -1 0 5250 0 1 1310
box -6 -8 86 268
use AOI21X1  _1291_
timestamp 0
transform -1 0 4610 0 1 1310
box -6 -8 86 268
use OAI21X1  _1292_
timestamp 0
transform -1 0 4450 0 1 1310
box -6 -8 86 268
use NAND2X1  _1293_
timestamp 0
transform 1 0 4210 0 -1 1830
box -6 -8 66 268
use XNOR2X1  _1294_
timestamp 0
transform -1 0 3730 0 1 2350
box -6 -8 126 268
use INVX1  _1295_
timestamp 0
transform -1 0 4410 0 -1 1830
box -6 -8 46 268
use OAI21X1  _1296_
timestamp 0
transform 1 0 4050 0 -1 1830
box -6 -8 86 268
use NOR2X1  _1297_
timestamp 0
transform -1 0 3830 0 -1 1830
box -6 -8 66 268
use AOI21X1  _1298_
timestamp 0
transform 1 0 3890 0 -1 1310
box -6 -8 86 268
use NOR3X1  _1299_
timestamp 0
transform -1 0 4590 0 -1 1310
box -6 -8 166 268
use AOI21X1  _1300_
timestamp 0
transform 1 0 4250 0 -1 1310
box -6 -8 86 268
use NAND2X1  _1301_
timestamp 0
transform 1 0 3910 0 -1 1830
box -6 -8 66 268
use INVX1  _1302_
timestamp 0
transform 1 0 4910 0 -1 790
box -6 -8 46 268
use OAI21X1  _1303_
timestamp 0
transform -1 0 5230 0 1 270
box -6 -8 86 268
use OAI21X1  _1304_
timestamp 0
transform 1 0 2670 0 1 1830
box -6 -8 86 268
use NAND2X1  _1305_
timestamp 0
transform -1 0 2030 0 -1 2350
box -6 -8 66 268
use NAND2X1  _1306_
timestamp 0
transform 1 0 1590 0 1 2350
box -6 -8 66 268
use NOR2X1  _1307_
timestamp 0
transform -1 0 1790 0 1 1830
box -6 -8 66 268
use AOI22X1  _1308_
timestamp 0
transform -1 0 1830 0 1 2350
box -6 -8 106 268
use OAI21X1  _1309_
timestamp 0
transform 1 0 2050 0 -1 1830
box -6 -8 86 268
use INVX1  _1310_
timestamp 0
transform 1 0 2190 0 1 1830
box -6 -8 46 268
use AND2X2  _1311_
timestamp 0
transform 1 0 1910 0 1 2350
box -6 -8 86 268
use NAND2X1  _1312_
timestamp 0
transform -1 0 2270 0 1 2350
box -6 -8 66 268
use INVX1  _1313_
timestamp 0
transform 1 0 2070 0 1 1830
box -6 -8 46 268
use NAND3X1  _1314_
timestamp 0
transform 1 0 2490 0 1 1830
box -6 -8 86 268
use NOR2X1  _1315_
timestamp 0
transform 1 0 2730 0 -1 1310
box -6 -8 66 268
use OAI21X1  _1316_
timestamp 0
transform 1 0 2870 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1317_
timestamp 0
transform 1 0 2730 0 1 1310
box -6 -8 86 268
use AOI21X1  _1318_
timestamp 0
transform 1 0 2330 0 1 1830
box -6 -8 86 268
use NOR3X1  _1319_
timestamp 0
transform -1 0 1950 0 -1 1830
box -6 -8 166 268
use AND2X2  _1320_
timestamp 0
transform -1 0 3470 0 1 1310
box -6 -8 86 268
use AOI21X1  _1321_
timestamp 0
transform -1 0 3310 0 1 1310
box -6 -8 86 268
use OAI21X1  _1322_
timestamp 0
transform 1 0 2410 0 1 1310
box -6 -8 86 268
use NAND3X1  _1323_
timestamp 0
transform 1 0 2890 0 1 1310
box -6 -8 86 268
use INVX1  _1324_
timestamp 0
transform 1 0 2710 0 -1 1830
box -6 -8 46 268
use NAND3X1  _1325_
timestamp 0
transform 1 0 2550 0 -1 1830
box -6 -8 86 268
use OAI21X1  _1326_
timestamp 0
transform 1 0 2570 0 1 1310
box -6 -8 86 268
use NAND3X1  _1327_
timestamp 0
transform 1 0 3070 0 1 1310
box -6 -8 86 268
use NAND2X1  _1328_
timestamp 0
transform -1 0 3670 0 1 270
box -6 -8 66 268
use NAND2X1  _1329_
timestamp 0
transform -1 0 5690 0 -1 1310
box -6 -8 66 268
use NAND2X1  _1330_
timestamp 0
transform -1 0 5510 0 -1 270
box -6 -8 66 268
use AOI22X1  _1331_
timestamp 0
transform 1 0 2370 0 -1 1830
box -6 -8 106 268
use AND2X2  _1332_
timestamp 0
transform 1 0 2230 0 -1 1310
box -6 -8 86 268
use AOI21X1  _1333_
timestamp 0
transform 1 0 2570 0 -1 1310
box -6 -8 86 268
use NAND2X1  _1334_
timestamp 0
transform -1 0 3190 0 -1 270
box -6 -8 66 268
use INVX1  _1335_
timestamp 0
transform -1 0 2610 0 1 790
box -6 -8 46 268
use AND2X2  _1336_
timestamp 0
transform -1 0 2490 0 -1 1310
box -6 -8 86 268
use OAI21X1  _1337_
timestamp 0
transform 1 0 2410 0 1 790
box -6 -8 86 268
use NAND2X1  _1338_
timestamp 0
transform 1 0 3270 0 -1 270
box -6 -8 66 268
use XOR2X1  _1339_
timestamp 0
transform -1 0 4290 0 -1 270
box -6 -8 126 268
use NOR2X1  _1340_
timestamp 0
transform 1 0 4070 0 1 270
box -6 -8 66 268
use AND2X2  _1341_
timestamp 0
transform 1 0 3450 0 1 270
box -6 -8 86 268
use NAND2X1  _1342_
timestamp 0
transform 1 0 4370 0 -1 270
box -6 -8 66 268
use AND2X2  _1343_
timestamp 0
transform 1 0 3410 0 -1 270
box -6 -8 86 268
use NAND3X1  _1344_
timestamp 0
transform -1 0 5370 0 -1 270
box -6 -8 86 268
use NAND2X1  _1345_
timestamp 0
transform 1 0 4530 0 -1 270
box -6 -8 66 268
use NOR2X1  _1346_
timestamp 0
transform -1 0 4270 0 1 270
box -6 -8 66 268
use OAI21X1  _1347_
timestamp 0
transform 1 0 4990 0 1 270
box -6 -8 86 268
use AOI21X1  _1348_
timestamp 0
transform -1 0 5430 0 -1 790
box -6 -8 86 268
use NAND3X1  _1349_
timestamp 0
transform 1 0 3750 0 1 270
box -6 -8 86 268
use NAND2X1  _1350_
timestamp 0
transform -1 0 3990 0 1 270
box -6 -8 66 268
use NAND3X1  _1351_
timestamp 0
transform 1 0 4670 0 1 270
box -6 -8 86 268
use AOI21X1  _1352_
timestamp 0
transform -1 0 5270 0 -1 790
box -6 -8 86 268
use NAND3X1  _1353_
timestamp 0
transform 1 0 4350 0 1 270
box -6 -8 86 268
use OAI21X1  _1354_
timestamp 0
transform -1 0 4910 0 1 270
box -6 -8 86 268
use AOI21X1  _1355_
timestamp 0
transform -1 0 4710 0 1 790
box -6 -8 86 268
use OAI21X1  _1356_
timestamp 0
transform -1 0 4530 0 1 790
box -6 -8 86 268
use AOI21X1  _1357_
timestamp 0
transform -1 0 5250 0 -1 1310
box -6 -8 86 268
use OAI21X1  _1358_
timestamp 0
transform -1 0 4750 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1359_
timestamp 0
transform 1 0 4750 0 -1 790
box -6 -8 86 268
use NAND3X1  _1360_
timestamp 0
transform -1 0 5110 0 -1 790
box -6 -8 86 268
use NAND3X1  _1361_
timestamp 0
transform -1 0 4870 0 1 790
box -6 -8 86 268
use NAND2X1  _1362_
timestamp 0
transform 1 0 4310 0 1 790
box -6 -8 66 268
use XOR2X1  _1363_
timestamp 0
transform 1 0 4050 0 -1 1310
box -6 -8 126 268
use OAI21X1  _1364_
timestamp 0
transform -1 0 4030 0 1 790
box -6 -8 86 268
use INVX1  _1365_
timestamp 0
transform -1 0 4470 0 -1 790
box -6 -8 46 268
use AOI21X1  _1366_
timestamp 0
transform -1 0 4350 0 -1 790
box -6 -8 86 268
use NAND2X1  _1367_
timestamp 0
transform 1 0 2850 0 1 790
box -6 -8 66 268
use INVX1  _1368_
timestamp 0
transform 1 0 3350 0 1 790
box -6 -8 46 268
use NAND2X1  _1369_
timestamp 0
transform 1 0 4030 0 -1 270
box -6 -8 66 268
use OAI21X1  _1370_
timestamp 0
transform -1 0 3950 0 -1 270
box -6 -8 86 268
use OAI21X1  _1371_
timestamp 0
transform 1 0 2210 0 -1 1830
box -6 -8 86 268
use INVX1  _1372_
timestamp 0
transform -1 0 1650 0 1 1830
box -6 -8 46 268
use NAND2X1  _1373_
timestamp 0
transform -1 0 1590 0 -1 2350
box -6 -8 66 268
use INVX1  _1374_
timestamp 0
transform 1 0 1170 0 1 2350
box -6 -8 46 268
use NAND2X1  _1375_
timestamp 0
transform 1 0 1450 0 1 2350
box -6 -8 66 268
use OAI21X1  _1376_
timestamp 0
transform 1 0 1290 0 1 2350
box -6 -8 86 268
use OAI21X1  _1377_
timestamp 0
transform -1 0 1310 0 -1 1830
box -6 -8 86 268
use OAI21X1  _1378_
timestamp 0
transform -1 0 1970 0 1 1830
box -6 -8 86 268
use NAND2X1  _1379_
timestamp 0
transform 1 0 1470 0 1 1830
box -6 -8 66 268
use INVX1  _1380_
timestamp 0
transform 1 0 1330 0 -1 1310
box -6 -8 46 268
use NOR2X1  _1381_
timestamp 0
transform 1 0 1390 0 -1 1830
box -6 -8 66 268
use INVX1  _1382_
timestamp 0
transform 1 0 1550 0 -1 1830
box -6 -8 46 268
use NAND3X1  _1383_
timestamp 0
transform 1 0 1770 0 1 1310
box -6 -8 86 268
use NAND3X1  _1384_
timestamp 0
transform -1 0 2190 0 1 1310
box -6 -8 86 268
use INVX1  _1385_
timestamp 0
transform -1 0 1810 0 -1 1310
box -6 -8 46 268
use AOI21X1  _1386_
timestamp 0
transform -1 0 1690 0 1 1310
box -6 -8 86 268
use NOR2X1  _1387_
timestamp 0
transform -1 0 1250 0 -1 1310
box -6 -8 66 268
use OAI21X1  _1388_
timestamp 0
transform 1 0 1610 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1389_
timestamp 0
transform -1 0 1990 0 1 790
box -6 -8 86 268
use INVX1  _1390_
timestamp 0
transform -1 0 2310 0 1 1310
box -6 -8 46 268
use NAND3X1  _1391_
timestamp 0
transform 1 0 1950 0 1 1310
box -6 -8 86 268
use OAI21X1  _1392_
timestamp 0
transform 1 0 1450 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1393_
timestamp 0
transform -1 0 1970 0 -1 1310
box -6 -8 86 268
use XNOR2X1  _1394_
timestamp 0
transform 1 0 2630 0 1 270
box -6 -8 126 268
use NAND2X1  _1395_
timestamp 0
transform 1 0 2990 0 -1 270
box -6 -8 66 268
use OR2X2  _1396_
timestamp 0
transform -1 0 2910 0 -1 270
box -6 -8 86 268
use NAND2X1  _1397_
timestamp 0
transform -1 0 2730 0 -1 270
box -6 -8 66 268
use INVX1  _1398_
timestamp 0
transform -1 0 2470 0 -1 790
box -6 -8 46 268
use NAND3X1  _1399_
timestamp 0
transform 1 0 2250 0 1 790
box -6 -8 86 268
use AOI21X1  _1400_
timestamp 0
transform 1 0 2050 0 -1 1310
box -6 -8 86 268
use AOI21X1  _1401_
timestamp 0
transform 1 0 2090 0 1 790
box -6 -8 86 268
use OAI21X1  _1402_
timestamp 0
transform 1 0 2550 0 -1 790
box -6 -8 86 268
use NAND2X1  _1403_
timestamp 0
transform -1 0 3050 0 1 270
box -6 -8 66 268
use NAND2X1  _1404_
timestamp 0
transform -1 0 3350 0 1 270
box -6 -8 66 268
use INVX1  _1405_
timestamp 0
transform -1 0 3790 0 -1 270
box -6 -8 46 268
use AOI21X1  _1406_
timestamp 0
transform -1 0 3650 0 -1 270
box -6 -8 86 268
use NAND3X1  _1407_
timestamp 0
transform 1 0 3030 0 -1 790
box -6 -8 86 268
use AOI21X1  _1408_
timestamp 0
transform 1 0 3670 0 -1 790
box -6 -8 86 268
use NAND3X1  _1409_
timestamp 0
transform 1 0 2870 0 -1 790
box -6 -8 86 268
use NAND2X1  _1410_
timestamp 0
transform -1 0 3210 0 1 270
box -6 -8 66 268
use AOI21X1  _1411_
timestamp 0
transform 1 0 3350 0 -1 790
box -6 -8 86 268
use OAI21X1  _1412_
timestamp 0
transform 1 0 3830 0 -1 790
box -6 -8 86 268
use AOI21X1  _1413_
timestamp 0
transform 1 0 4510 0 1 270
box -6 -8 86 268
use OAI21X1  _1414_
timestamp 0
transform -1 0 4650 0 -1 790
box -6 -8 86 268
use NAND3X1  _1415_
timestamp 0
transform -1 0 3270 0 -1 790
box -6 -8 86 268
use NAND3X1  _1416_
timestamp 0
transform 1 0 3510 0 -1 790
box -6 -8 86 268
use NAND3X1  _1417_
timestamp 0
transform -1 0 4070 0 -1 790
box -6 -8 86 268
use NAND2X1  _1418_
timestamp 0
transform 1 0 3650 0 1 790
box -6 -8 66 268
use INVX1  _1419_
timestamp 0
transform 1 0 3630 0 -1 1310
box -6 -8 46 268
use XOR2X1  _1420_
timestamp 0
transform 1 0 4110 0 1 790
box -6 -8 126 268
use NOR2X1  _1421_
timestamp 0
transform 1 0 3750 0 -1 1310
box -6 -8 66 268
use NAND3X1  _1422_
timestamp 0
transform -1 0 3530 0 -1 1310
box -6 -8 86 268
use INVX1  _1423_
timestamp 0
transform -1 0 4190 0 -1 790
box -6 -8 46 268
use NAND3X1  _1424_
timestamp 0
transform -1 0 3570 0 1 790
box -6 -8 86 268
use NAND2X1  _1425_
timestamp 0
transform 1 0 3790 0 1 790
box -6 -8 66 268
use NAND2X1  _1426_
timestamp 0
transform 1 0 2990 0 1 790
box -6 -8 66 268
use NAND3X1  _1427_
timestamp 0
transform -1 0 2770 0 1 790
box -6 -8 86 268
use NAND2X1  _1428_
timestamp 0
transform 1 0 1770 0 1 790
box -6 -8 66 268
use INVX1  _1429_
timestamp 0
transform -1 0 1270 0 -1 270
box -6 -8 46 268
use AND2X2  _1430_
timestamp 0
transform -1 0 2590 0 -1 270
box -6 -8 86 268
use OAI21X1  _1431_
timestamp 0
transform 1 0 1450 0 1 1310
box -6 -8 86 268
use NAND2X1  _1432_
timestamp 0
transform 1 0 710 0 1 2350
box -6 -8 66 268
use OAI21X1  _1433_
timestamp 0
transform -1 0 1430 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1434_
timestamp 0
transform 1 0 1170 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1435_
timestamp 0
transform 1 0 1130 0 1 1830
box -6 -8 86 268
use NAND2X1  _1436_
timestamp 0
transform 1 0 1030 0 1 2350
box -6 -8 66 268
use OR2X2  _1437_
timestamp 0
transform 1 0 1010 0 -1 2350
box -6 -8 86 268
use NAND3X1  _1438_
timestamp 0
transform -1 0 1210 0 1 1310
box -6 -8 86 268
use INVX1  _1439_
timestamp 0
transform -1 0 870 0 1 270
box -6 -8 46 268
use AOI21X1  _1440_
timestamp 0
transform 1 0 1290 0 1 1310
box -6 -8 86 268
use NOR2X1  _1441_
timestamp 0
transform -1 0 590 0 1 270
box -6 -8 66 268
use INVX1  _1442_
timestamp 0
transform 1 0 110 0 -1 270
box -6 -8 46 268
use NAND2X1  _1443_
timestamp 0
transform -1 0 2550 0 1 270
box -6 -8 66 268
use OR2X2  _1444_
timestamp 0
transform -1 0 310 0 -1 270
box -6 -8 86 268
use NAND2X1  _1445_
timestamp 0
transform 1 0 530 0 -1 270
box -6 -8 66 268
use NAND2X1  _1446_
timestamp 0
transform -1 0 450 0 -1 270
box -6 -8 66 268
use INVX1  _1447_
timestamp 0
transform -1 0 150 0 1 270
box -6 -8 46 268
use NAND2X1  _1448_
timestamp 0
transform 1 0 230 0 1 270
box -6 -8 66 268
use OAI21X1  _1449_
timestamp 0
transform -1 0 750 0 1 270
box -6 -8 86 268
use NAND2X1  _1450_
timestamp 0
transform -1 0 730 0 -1 270
box -6 -8 66 268
use NAND2X1  _1451_
timestamp 0
transform -1 0 1030 0 1 270
box -6 -8 66 268
use INVX1  _1452_
timestamp 0
transform -1 0 990 0 -1 270
box -6 -8 46 268
use NOR2X1  _1453_
timestamp 0
transform -1 0 870 0 -1 270
box -6 -8 66 268
use OAI21X1  _1454_
timestamp 0
transform 1 0 1070 0 -1 270
box -6 -8 86 268
use OR2X2  _1455_
timestamp 0
transform 1 0 1110 0 1 270
box -6 -8 86 268
use NAND3X1  _1456_
timestamp 0
transform 1 0 1290 0 1 270
box -6 -8 86 268
use NAND2X1  _1457_
timestamp 0
transform -1 0 2170 0 1 270
box -6 -8 66 268
use NAND3X1  _1458_
timestamp 0
transform -1 0 2790 0 -1 790
box -6 -8 86 268
use OAI21X1  _1459_
timestamp 0
transform -1 0 2910 0 1 270
box -6 -8 86 268
use NAND3X1  _1460_
timestamp 0
transform -1 0 2030 0 1 270
box -6 -8 86 268
use NAND2X1  _1461_
timestamp 0
transform 1 0 1850 0 -1 790
box -6 -8 66 268
use XNOR2X1  _1462_
timestamp 0
transform -1 0 2110 0 -1 790
box -6 -8 126 268
use INVX1  _1463_
timestamp 0
transform 1 0 1810 0 1 270
box -6 -8 46 268
use OAI21X1  _1464_
timestamp 0
transform -1 0 1730 0 1 270
box -6 -8 86 268
use AOI21X1  _1465_
timestamp 0
transform 1 0 1370 0 -1 270
box -6 -8 86 268
use OAI22X1  _1466_
timestamp 0
transform 1 0 850 0 1 2350
box -6 -8 106 268
use INVX1  _1467_
timestamp 0
transform -1 0 670 0 -1 2350
box -6 -8 46 268
use NOR2X1  _1468_
timestamp 0
transform 1 0 990 0 1 1830
box -6 -8 66 268
use NAND2X1  _1469_
timestamp 0
transform 1 0 690 0 1 1830
box -6 -8 66 268
use OAI21X1  _1470_
timestamp 0
transform -1 0 1390 0 1 1830
box -6 -8 86 268
use AND2X2  _1471_
timestamp 0
transform 1 0 830 0 1 1830
box -6 -8 86 268
use XOR2X1  _1472_
timestamp 0
transform -1 0 210 0 1 1830
box -6 -8 126 268
use XNOR2X1  _1473_
timestamp 0
transform -1 0 210 0 1 790
box -6 -8 126 268
use NAND3X1  _1474_
timestamp 0
transform -1 0 190 0 -1 790
box -6 -8 86 268
use INVX1  _1475_
timestamp 0
transform 1 0 590 0 -1 790
box -6 -8 46 268
use AOI21X1  _1476_
timestamp 0
transform 1 0 270 0 -1 790
box -6 -8 86 268
use OAI21X1  _1477_
timestamp 0
transform 1 0 710 0 -1 790
box -6 -8 86 268
use OAI21X1  _1478_
timestamp 0
transform 1 0 370 0 1 270
box -6 -8 86 268
use INVX1  _1479_
timestamp 0
transform 1 0 310 0 1 790
box -6 -8 46 268
use NAND2X1  _1480_
timestamp 0
transform -1 0 490 0 1 790
box -6 -8 66 268
use NAND3X1  _1481_
timestamp 0
transform 1 0 430 0 -1 790
box -6 -8 86 268
use NAND2X1  _1482_
timestamp 0
transform -1 0 930 0 -1 790
box -6 -8 66 268
use XOR2X1  _1483_
timestamp 0
transform -1 0 1570 0 1 270
box -6 -8 126 268
use XOR2X1  _1484_
timestamp 0
transform -1 0 1670 0 -1 270
box -6 -8 126 268
use NAND2X1  _1485_
timestamp 0
transform -1 0 1430 0 -1 790
box -6 -8 66 268
use NAND3X1  _1486_
timestamp 0
transform -1 0 1770 0 -1 790
box -6 -8 86 268
use INVX1  _1487_
timestamp 0
transform -1 0 1510 0 1 790
box -6 -8 46 268
use OAI21X1  _1488_
timestamp 0
transform 1 0 1530 0 -1 790
box -6 -8 86 268
use AOI22X1  _1489_
timestamp 0
transform 1 0 1290 0 1 790
box -6 -8 106 268
use INVX1  _1490_
timestamp 0
transform 1 0 570 0 1 790
box -6 -8 46 268
use NOR2X1  _1491_
timestamp 0
transform -1 0 910 0 1 790
box -6 -8 66 268
use NAND3X1  _1492_
timestamp 0
transform 1 0 690 0 -1 1830
box -6 -8 86 268
use INVX1  _1493_
timestamp 0
transform -1 0 610 0 -1 1830
box -6 -8 46 268
use INVX1  _1494_
timestamp 0
transform 1 0 270 0 -1 1830
box -6 -8 46 268
use OAI21X1  _1495_
timestamp 0
transform 1 0 390 0 -1 1830
box -6 -8 86 268
use NAND2X1  _1496_
timestamp 0
transform 1 0 790 0 1 1310
box -6 -8 66 268
use NAND2X1  _1497_
timestamp 0
transform 1 0 310 0 1 1830
box -6 -8 66 268
use NAND2X1  _1498_
timestamp 0
transform 1 0 90 0 -1 1310
box -6 -8 66 268
use NAND2X1  _1499_
timestamp 0
transform -1 0 350 0 1 1310
box -6 -8 66 268
use XNOR2X1  _1500_
timestamp 0
transform 1 0 930 0 1 1310
box -6 -8 126 268
use XNOR2X1  _1501_
timestamp 0
transform -1 0 1130 0 -1 790
box -6 -8 126 268
use INVX1  _1502_
timestamp 0
transform -1 0 1050 0 1 790
box -6 -8 46 268
use XOR2X1  _1503_
timestamp 0
transform -1 0 1090 0 -1 1310
box -6 -8 126 268
use OAI21X1  _1504_
timestamp 0
transform 1 0 690 0 1 790
box -6 -8 86 268
use OAI21X1  _1505_
timestamp 0
transform -1 0 890 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1506_
timestamp 0
transform -1 0 710 0 1 1310
box -6 -8 86 268
use OAI21X1  _1507_
timestamp 0
transform 1 0 110 0 -1 1830
box -6 -8 86 268
use XNOR2X1  _1508_
timestamp 0
transform -1 0 210 0 1 1310
box -6 -8 126 268
use XOR2X1  _1509_
timestamp 0
transform -1 0 550 0 1 1310
box -6 -8 126 268
use NAND2X1  _1510_
timestamp 0
transform 1 0 350 0 -1 1310
box -6 -8 66 268
use AOI22X1  _1511_
timestamp 0
transform 1 0 3150 0 1 790
box -6 -8 106 268
use AOI21X1  _1512_
timestamp 0
transform -1 0 1670 0 1 790
box -6 -8 86 268
use AND2X2  _1513_
timestamp 0
transform -1 0 1290 0 -1 790
box -6 -8 86 268
use OAI21X1  _1514_
timestamp 0
transform -1 0 1210 0 1 790
box -6 -8 86 268
use INVX1  _1515_
timestamp 0
transform -1 0 270 0 -1 1310
box -6 -8 46 268
use NAND3X1  _1516_
timestamp 0
transform -1 0 730 0 -1 1310
box -6 -8 86 268
use NAND2X1  _1517_
timestamp 0
transform -1 0 550 0 -1 1310
box -6 -8 66 268
use OAI21X1  _1518_
timestamp 0
transform 1 0 1350 0 -1 5470
box -6 -8 86 268
use XOR2X1  _1519_
timestamp 0
transform 1 0 2250 0 -1 5470
box -6 -8 126 268
use DFFPOSX1  _1520_
timestamp 0
transform -1 0 410 0 1 2870
box -6 -8 246 268
use DFFPOSX1  _1521_
timestamp 0
transform -1 0 650 0 1 2870
box -6 -8 246 268
use DFFPOSX1  _1522_
timestamp 0
transform -1 0 390 0 -1 4950
box -6 -8 246 268
use DFFPOSX1  _1523_
timestamp 0
transform -1 0 1270 0 -1 3910
box -6 -8 246 268
use DFFPOSX1  _1524_
timestamp 0
transform -1 0 910 0 -1 2870
box -6 -8 246 268
use DFFPOSX1  _1525_
timestamp 0
transform 1 0 3610 0 -1 5990
box -6 -8 246 268
use DFFPOSX1  _1526_
timestamp 0
transform -1 0 1330 0 -1 5990
box -6 -8 246 268
use DFFPOSX1  _1527_
timestamp 0
transform -1 0 670 0 -1 2870
box -6 -8 246 268
use DFFPOSX1  _1528_
timestamp 0
transform -1 0 390 0 1 3910
box -6 -8 246 268
use DFFPOSX1  _1529_
timestamp 0
transform -1 0 390 0 1 3390
box -6 -8 246 268
use DFFPOSX1  _1530_
timestamp 0
transform -1 0 390 0 -1 3390
box -6 -8 246 268
use DFFPOSX1  _1531_
timestamp 0
transform -1 0 690 0 -1 5990
box -6 -8 246 268
use DFFPOSX1  _1532_
timestamp 0
transform 1 0 1330 0 -1 5990
box -6 -8 246 268
use DFFPOSX1  _1533_
timestamp 0
transform 1 0 1950 0 -1 5990
box -6 -8 246 268
use DFFPOSX1  _1534_
timestamp 0
transform -1 0 3070 0 -1 5990
box -6 -8 246 268
use DFFPOSX1  _1535_
timestamp 0
transform -1 0 3410 0 1 4430
box -6 -8 246 268
use DFFPOSX1  _1536_
timestamp 0
transform -1 0 390 0 1 2350
box -6 -8 246 268
use DFFPOSX1  _1537_
timestamp 0
transform -1 0 3610 0 -1 5990
box -6 -8 246 268
use DFFPOSX1  _1538_
timestamp 0
transform -1 0 4050 0 1 1310
box -6 -8 246 268
use DFFPOSX1  _1539_
timestamp 0
transform 1 0 4830 0 -1 270
box -6 -8 246 268
use DFFPOSX1  _1540_
timestamp 0
transform 1 0 2170 0 1 270
box -6 -8 246 268
use DFFPOSX1  _1541_
timestamp 0
transform 1 0 1910 0 -1 270
box -6 -8 246 268
use DFFPOSX1  _1542_
timestamp 0
transform -1 0 910 0 -1 2350
box -6 -8 246 268
use DFFPOSX1  _1543_
timestamp 0
transform -1 0 550 0 -1 2350
box -6 -8 246 268
use DFFPOSX1  _1544_
timestamp 0
transform -1 0 390 0 -1 3910
box -6 -8 246 268
use DFFPOSX1  _1545_
timestamp 0
transform -1 0 630 0 1 3390
box -6 -8 246 268
use DFFPOSX1  _1546_
timestamp 0
transform -1 0 770 0 -1 3910
box -6 -8 246 268
use DFFPOSX1  _1547_
timestamp 0
transform -1 0 1290 0 1 5470
box -6 -8 246 268
use DFFPOSX1  _1548_
timestamp 0
transform -1 0 2350 0 1 5470
box -6 -8 246 268
use DFFPOSX1  _1549_
timestamp 0
transform -1 0 2590 0 1 5470
box -6 -8 246 268
use DFFPOSX1  _1550_
timestamp 0
transform -1 0 3490 0 1 5470
box -6 -8 246 268
use DFFPOSX1  _1551_
timestamp 0
transform -1 0 3650 0 1 4430
box -6 -8 246 268
use DFFPOSX1  _1552_
timestamp 0
transform -1 0 630 0 1 2350
box -6 -8 246 268
use DFFPOSX1  _1553_
timestamp 0
transform -1 0 3630 0 -1 2870
box -6 -8 246 268
use DFFPOSX1  _1554_
timestamp 0
transform -1 0 4290 0 1 1310
box -6 -8 246 268
use DFFPOSX1  _1555_
timestamp 0
transform 1 0 4590 0 -1 270
box -6 -8 246 268
use DFFPOSX1  _1556_
timestamp 0
transform 1 0 2110 0 -1 790
box -6 -8 246 268
use DFFPOSX1  _1557_
timestamp 0
transform 1 0 1670 0 -1 270
box -6 -8 246 268
use DFFPOSX1  _1558_
timestamp 0
transform -1 0 1010 0 -1 1830
box -6 -8 246 268
use DFFPOSX1  _1559_
timestamp 0
transform -1 0 610 0 1 1830
box -6 -8 246 268
use BUFX2  _1560_
timestamp 0
transform -1 0 170 0 1 2870
box -6 -8 66 268
use BUFX2  _1561_
timestamp 0
transform -1 0 290 0 -1 2870
box -6 -8 66 268
use BUFX2  _1562_
timestamp 0
transform -1 0 150 0 -1 4950
box -6 -8 66 268
use BUFX2  _1563_
timestamp 0
transform -1 0 150 0 -1 3910
box -6 -8 66 268
use BUFX2  _1564_
timestamp 0
transform -1 0 430 0 -1 2870
box -6 -8 66 268
use BUFX2  _1565_
timestamp 0
transform 1 0 3950 0 -1 5990
box -6 -8 66 268
use BUFX2  _1566_
timestamp 0
transform -1 0 1090 0 -1 5990
box -6 -8 66 268
use BUFX2  _1567_
timestamp 0
transform -1 0 150 0 -1 2870
box -6 -8 66 268
use BUFX2  _1568_
timestamp 0
transform -1 0 150 0 1 3910
box -6 -8 66 268
use BUFX2  _1569_
timestamp 0
transform -1 0 150 0 1 3390
box -6 -8 66 268
use BUFX2  _1570_
timestamp 0
transform -1 0 3810 0 1 1310
box -6 -8 66 268
use BUFX2  _1571_
timestamp 0
transform 1 0 5150 0 -1 270
box -6 -8 66 268
use BUFX2  _1572_
timestamp 0
transform -1 0 2430 0 -1 270
box -6 -8 66 268
use BUFX2  _1573_
timestamp 0
transform 1 0 2230 0 -1 270
box -6 -8 66 268
use BUFX2  _1574_
timestamp 0
transform -1 0 170 0 -1 2350
box -6 -8 66 268
use BUFX2  _1575_
timestamp 0
transform -1 0 310 0 -1 2350
box -6 -8 66 268
use BUFX2  _1576_
timestamp 0
transform -1 0 150 0 -1 3390
box -6 -8 66 268
use BUFX2  _1577_
timestamp 0
transform -1 0 450 0 -1 5990
box -6 -8 66 268
use BUFX2  _1578_
timestamp 0
transform 1 0 1650 0 -1 5990
box -6 -8 66 268
use BUFX2  _1579_
timestamp 0
transform 1 0 2290 0 -1 5990
box -6 -8 66 268
use BUFX2  _1580_
timestamp 0
transform -1 0 2830 0 -1 5990
box -6 -8 66 268
use BUFX2  _1581_
timestamp 0
transform -1 0 3170 0 1 4430
box -6 -8 66 268
use BUFX2  _1582_
timestamp 0
transform -1 0 150 0 1 2350
box -6 -8 66 268
use BUFX2  _1583_
timestamp 0
transform -1 0 3370 0 -1 5990
box -6 -8 66 268
use BUFX2  BUFX2_insert6
timestamp 0
transform 1 0 5130 0 -1 5990
box -6 -8 66 268
use BUFX2  BUFX2_insert7
timestamp 0
transform -1 0 3210 0 -1 5990
box -6 -8 66 268
use BUFX2  BUFX2_insert8
timestamp 0
transform -1 0 3230 0 -1 5470
box -6 -8 66 268
use BUFX2  BUFX2_insert9
timestamp 0
transform -1 0 5930 0 -1 270
box -6 -8 66 268
use BUFX2  BUFX2_insert10
timestamp 0
transform 1 0 1690 0 -1 3390
box -6 -8 66 268
use BUFX2  BUFX2_insert11
timestamp 0
transform 1 0 1810 0 1 4430
box -6 -8 66 268
use BUFX2  BUFX2_insert12
timestamp 0
transform 1 0 1570 0 1 3390
box -6 -8 66 268
use BUFX2  BUFX2_insert13
timestamp 0
transform -1 0 170 0 -1 5990
box -6 -8 66 268
use BUFX2  BUFX2_insert14
timestamp 0
transform -1 0 2850 0 1 2350
box -6 -8 66 268
use BUFX2  BUFX2_insert15
timestamp 0
transform -1 0 4150 0 -1 5990
box -6 -8 66 268
use BUFX2  BUFX2_insert16
timestamp 0
transform 1 0 4310 0 -1 2350
box -6 -8 66 268
use BUFX2  BUFX2_insert17
timestamp 0
transform 1 0 4250 0 -1 5990
box -6 -8 66 268
use CLKBUF1  CLKBUF1_insert0
timestamp 0
transform 1 0 1490 0 -1 2870
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert1
timestamp 0
transform -1 0 1490 0 1 3390
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert2
timestamp 0
transform -1 0 950 0 -1 5990
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert3
timestamp 0
transform -1 0 1290 0 -1 2870
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert4
timestamp 0
transform -1 0 1290 0 -1 3390
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert5
timestamp 0
transform 1 0 3070 0 1 5470
box -6 -8 186 268
use FILL  FILL88050x7950
timestamp 0
transform -1 0 5890 0 -1 790
box -6 -8 26 268
use FILL  FILL88050x19650
timestamp 0
transform 1 0 5870 0 1 1310
box -6 -8 26 268
use FILL  FILL88050x35250
timestamp 0
transform 1 0 5870 0 1 2350
box -6 -8 26 268
use FILL  FILL88050x54750
timestamp 0
transform -1 0 5890 0 -1 3910
box -6 -8 26 268
use FILL  FILL88050x74250
timestamp 0
transform 1 0 5870 0 1 4950
box -6 -8 26 268
use FILL  FILL88050x78150
timestamp 0
transform -1 0 5890 0 -1 5470
box -6 -8 26 268
use FILL  FILL88350x4050
timestamp 0
transform 1 0 5890 0 1 270
box -6 -8 26 268
use FILL  FILL88350x7950
timestamp 0
transform -1 0 5910 0 -1 790
box -6 -8 26 268
use FILL  FILL88350x15750
timestamp 0
transform -1 0 5910 0 -1 1310
box -6 -8 26 268
use FILL  FILL88350x19650
timestamp 0
transform 1 0 5890 0 1 1310
box -6 -8 26 268
use FILL  FILL88350x23550
timestamp 0
transform -1 0 5910 0 -1 1830
box -6 -8 26 268
use FILL  FILL88350x35250
timestamp 0
transform 1 0 5890 0 1 2350
box -6 -8 26 268
use FILL  FILL88350x54750
timestamp 0
transform -1 0 5910 0 -1 3910
box -6 -8 26 268
use FILL  FILL88350x74250
timestamp 0
transform 1 0 5890 0 1 4950
box -6 -8 26 268
use FILL  FILL88350x78150
timestamp 0
transform -1 0 5910 0 -1 5470
box -6 -8 26 268
use FILL  FILL88350x85950
timestamp 0
transform -1 0 5910 0 -1 5990
box -6 -8 26 268
use FILL  FILL88650x4050
timestamp 0
transform 1 0 5910 0 1 270
box -6 -8 26 268
use FILL  FILL88650x7950
timestamp 0
transform -1 0 5930 0 -1 790
box -6 -8 26 268
use FILL  FILL88650x15750
timestamp 0
transform -1 0 5930 0 -1 1310
box -6 -8 26 268
use FILL  FILL88650x19650
timestamp 0
transform 1 0 5910 0 1 1310
box -6 -8 26 268
use FILL  FILL88650x23550
timestamp 0
transform -1 0 5930 0 -1 1830
box -6 -8 26 268
use FILL  FILL88650x35250
timestamp 0
transform 1 0 5910 0 1 2350
box -6 -8 26 268
use FILL  FILL88650x39150
timestamp 0
transform -1 0 5930 0 -1 2870
box -6 -8 26 268
use FILL  FILL88650x54750
timestamp 0
transform -1 0 5930 0 -1 3910
box -6 -8 26 268
use FILL  FILL88650x58650
timestamp 0
transform 1 0 5910 0 1 3910
box -6 -8 26 268
use FILL  FILL88650x74250
timestamp 0
transform 1 0 5910 0 1 4950
box -6 -8 26 268
use FILL  FILL88650x78150
timestamp 0
transform -1 0 5930 0 -1 5470
box -6 -8 26 268
use FILL  FILL88650x85950
timestamp 0
transform -1 0 5930 0 -1 5990
box -6 -8 26 268
use FILL  FILL88950x150
timestamp 0
transform -1 0 5950 0 -1 270
box -6 -8 26 268
use FILL  FILL88950x4050
timestamp 0
transform 1 0 5930 0 1 270
box -6 -8 26 268
use FILL  FILL88950x7950
timestamp 0
transform -1 0 5950 0 -1 790
box -6 -8 26 268
use FILL  FILL88950x15750
timestamp 0
transform -1 0 5950 0 -1 1310
box -6 -8 26 268
use FILL  FILL88950x19650
timestamp 0
transform 1 0 5930 0 1 1310
box -6 -8 26 268
use FILL  FILL88950x23550
timestamp 0
transform -1 0 5950 0 -1 1830
box -6 -8 26 268
use FILL  FILL88950x27450
timestamp 0
transform 1 0 5930 0 1 1830
box -6 -8 26 268
use FILL  FILL88950x31350
timestamp 0
transform -1 0 5950 0 -1 2350
box -6 -8 26 268
use FILL  FILL88950x35250
timestamp 0
transform 1 0 5930 0 1 2350
box -6 -8 26 268
use FILL  FILL88950x39150
timestamp 0
transform -1 0 5950 0 -1 2870
box -6 -8 26 268
use FILL  FILL88950x54750
timestamp 0
transform -1 0 5950 0 -1 3910
box -6 -8 26 268
use FILL  FILL88950x58650
timestamp 0
transform 1 0 5930 0 1 3910
box -6 -8 26 268
use FILL  FILL88950x74250
timestamp 0
transform 1 0 5930 0 1 4950
box -6 -8 26 268
use FILL  FILL88950x78150
timestamp 0
transform -1 0 5950 0 -1 5470
box -6 -8 26 268
use FILL  FILL88950x85950
timestamp 0
transform -1 0 5950 0 -1 5990
box -6 -8 26 268
use FILL  FILL89250x150
timestamp 0
transform -1 0 5970 0 -1 270
box -6 -8 26 268
use FILL  FILL89250x4050
timestamp 0
transform 1 0 5950 0 1 270
box -6 -8 26 268
use FILL  FILL89250x7950
timestamp 0
transform -1 0 5970 0 -1 790
box -6 -8 26 268
use FILL  FILL89250x11850
timestamp 0
transform 1 0 5950 0 1 790
box -6 -8 26 268
use FILL  FILL89250x15750
timestamp 0
transform -1 0 5970 0 -1 1310
box -6 -8 26 268
use FILL  FILL89250x19650
timestamp 0
transform 1 0 5950 0 1 1310
box -6 -8 26 268
use FILL  FILL89250x23550
timestamp 0
transform -1 0 5970 0 -1 1830
box -6 -8 26 268
use FILL  FILL89250x27450
timestamp 0
transform 1 0 5950 0 1 1830
box -6 -8 26 268
use FILL  FILL89250x31350
timestamp 0
transform -1 0 5970 0 -1 2350
box -6 -8 26 268
use FILL  FILL89250x35250
timestamp 0
transform 1 0 5950 0 1 2350
box -6 -8 26 268
use FILL  FILL89250x39150
timestamp 0
transform -1 0 5970 0 -1 2870
box -6 -8 26 268
use FILL  FILL89250x54750
timestamp 0
transform -1 0 5970 0 -1 3910
box -6 -8 26 268
use FILL  FILL89250x58650
timestamp 0
transform 1 0 5950 0 1 3910
box -6 -8 26 268
use FILL  FILL89250x74250
timestamp 0
transform 1 0 5950 0 1 4950
box -6 -8 26 268
use FILL  FILL89250x78150
timestamp 0
transform -1 0 5970 0 -1 5470
box -6 -8 26 268
use FILL  FILL89250x85950
timestamp 0
transform -1 0 5970 0 -1 5990
box -6 -8 26 268
use FILL  FILL89550x150
timestamp 0
transform -1 0 5990 0 -1 270
box -6 -8 26 268
use FILL  FILL89550x4050
timestamp 0
transform 1 0 5970 0 1 270
box -6 -8 26 268
use FILL  FILL89550x7950
timestamp 0
transform -1 0 5990 0 -1 790
box -6 -8 26 268
use FILL  FILL89550x11850
timestamp 0
transform 1 0 5970 0 1 790
box -6 -8 26 268
use FILL  FILL89550x15750
timestamp 0
transform -1 0 5990 0 -1 1310
box -6 -8 26 268
use FILL  FILL89550x19650
timestamp 0
transform 1 0 5970 0 1 1310
box -6 -8 26 268
use FILL  FILL89550x23550
timestamp 0
transform -1 0 5990 0 -1 1830
box -6 -8 26 268
use FILL  FILL89550x27450
timestamp 0
transform 1 0 5970 0 1 1830
box -6 -8 26 268
use FILL  FILL89550x31350
timestamp 0
transform -1 0 5990 0 -1 2350
box -6 -8 26 268
use FILL  FILL89550x35250
timestamp 0
transform 1 0 5970 0 1 2350
box -6 -8 26 268
use FILL  FILL89550x39150
timestamp 0
transform -1 0 5990 0 -1 2870
box -6 -8 26 268
use FILL  FILL89550x43050
timestamp 0
transform 1 0 5970 0 1 2870
box -6 -8 26 268
use FILL  FILL89550x46950
timestamp 0
transform -1 0 5990 0 -1 3390
box -6 -8 26 268
use FILL  FILL89550x54750
timestamp 0
transform -1 0 5990 0 -1 3910
box -6 -8 26 268
use FILL  FILL89550x58650
timestamp 0
transform 1 0 5970 0 1 3910
box -6 -8 26 268
use FILL  FILL89550x66450
timestamp 0
transform 1 0 5970 0 1 4430
box -6 -8 26 268
use FILL  FILL89550x74250
timestamp 0
transform 1 0 5970 0 1 4950
box -6 -8 26 268
use FILL  FILL89550x78150
timestamp 0
transform -1 0 5990 0 -1 5470
box -6 -8 26 268
use FILL  FILL89550x85950
timestamp 0
transform -1 0 5990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__756_
timestamp 0
transform 1 0 1270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__757_
timestamp 0
transform 1 0 1630 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__758_
timestamp 0
transform 1 0 1390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__759_
timestamp 0
transform 1 0 530 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__760_
timestamp 0
transform 1 0 670 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__761_
timestamp 0
transform 1 0 390 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__762_
timestamp 0
transform 1 0 390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__763_
timestamp 0
transform -1 0 1130 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__764_
timestamp 0
transform 1 0 910 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__765_
timestamp 0
transform -1 0 410 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__766_
timestamp 0
transform 1 0 570 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__767_
timestamp 0
transform 1 0 730 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__768_
timestamp 0
transform -1 0 870 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__769_
timestamp 0
transform 1 0 650 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__770_
timestamp 0
transform 1 0 790 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__771_
timestamp 0
transform 1 0 950 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__772_
timestamp 0
transform -1 0 1130 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__773_
timestamp 0
transform -1 0 810 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__774_
timestamp 0
transform 1 0 630 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__775_
timestamp 0
transform -1 0 3090 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__776_
timestamp 0
transform -1 0 1430 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__777_
timestamp 0
transform -1 0 970 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__778_
timestamp 0
transform 1 0 330 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__779_
timestamp 0
transform 1 0 490 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__780_
timestamp 0
transform 1 0 10 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__781_
timestamp 0
transform 1 0 10 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__782_
timestamp 0
transform 1 0 450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__783_
timestamp 0
transform 1 0 570 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__784_
timestamp 0
transform 1 0 170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__785_
timestamp 0
transform 1 0 290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__786_
timestamp 0
transform -1 0 770 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__787_
timestamp 0
transform 1 0 910 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__788_
timestamp 0
transform 1 0 1550 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__789_
timestamp 0
transform -1 0 1150 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__790_
timestamp 0
transform -1 0 1310 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__791_
timestamp 0
transform 1 0 1250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__792_
timestamp 0
transform -1 0 1390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__793_
timestamp 0
transform -1 0 990 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__794_
timestamp 0
transform 1 0 910 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__795_
timestamp 0
transform -1 0 830 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__796_
timestamp 0
transform 1 0 770 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__797_
timestamp 0
transform 1 0 1070 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__798_
timestamp 0
transform -1 0 870 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__799_
timestamp 0
transform -1 0 3430 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__800_
timestamp 0
transform 1 0 2190 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__801_
timestamp 0
transform 1 0 2270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__802_
timestamp 0
transform 1 0 1850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__803_
timestamp 0
transform -1 0 1550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__804_
timestamp 0
transform -1 0 1250 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__805_
timestamp 0
transform -1 0 190 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__806_
timestamp 0
transform -1 0 730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__807_
timestamp 0
transform 1 0 830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__808_
timestamp 0
transform 1 0 430 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__809_
timestamp 0
transform 1 0 10 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__810_
timestamp 0
transform -1 0 190 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__811_
timestamp 0
transform 1 0 130 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__812_
timestamp 0
transform -1 0 690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__813_
timestamp 0
transform -1 0 310 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__814_
timestamp 0
transform -1 0 30 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__815_
timestamp 0
transform 1 0 330 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__816_
timestamp 0
transform 1 0 390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__817_
timestamp 0
transform -1 0 30 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__818_
timestamp 0
transform -1 0 190 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__819_
timestamp 0
transform -1 0 530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__820_
timestamp 0
transform -1 0 150 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__821_
timestamp 0
transform 1 0 870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__822_
timestamp 0
transform 1 0 1990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__823_
timestamp 0
transform -1 0 1710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__824_
timestamp 0
transform 1 0 610 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__825_
timestamp 0
transform 1 0 550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__826_
timestamp 0
transform 1 0 910 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__827_
timestamp 0
transform -1 0 1230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__828_
timestamp 0
transform 1 0 710 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__829_
timestamp 0
transform -1 0 1050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__830_
timestamp 0
transform 1 0 310 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__831_
timestamp 0
transform -1 0 1450 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__832_
timestamp 0
transform 1 0 550 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__833_
timestamp 0
transform -1 0 1130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__834_
timestamp 0
transform 1 0 2050 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__835_
timestamp 0
transform 1 0 1070 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__836_
timestamp 0
transform 1 0 590 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__837_
timestamp 0
transform 1 0 950 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__838_
timestamp 0
transform -1 0 2370 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__839_
timestamp 0
transform -1 0 2550 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__840_
timestamp 0
transform -1 0 1730 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__841_
timestamp 0
transform -1 0 2530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__842_
timestamp 0
transform 1 0 2050 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__843_
timestamp 0
transform -1 0 1790 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__844_
timestamp 0
transform 1 0 1830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__845_
timestamp 0
transform -1 0 1910 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__846_
timestamp 0
transform -1 0 1570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__847_
timestamp 0
transform -1 0 950 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__848_
timestamp 0
transform 1 0 750 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__849_
timestamp 0
transform -1 0 1970 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__850_
timestamp 0
transform -1 0 1630 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__851_
timestamp 0
transform -1 0 1310 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__852_
timestamp 0
transform 1 0 2310 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__853_
timestamp 0
transform 1 0 2750 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__854_
timestamp 0
transform 1 0 2010 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__855_
timestamp 0
transform -1 0 1570 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__856_
timestamp 0
transform 1 0 1550 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__857_
timestamp 0
transform -1 0 1890 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__858_
timestamp 0
transform -1 0 2230 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__859_
timestamp 0
transform 1 0 2630 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__860_
timestamp 0
transform -1 0 2490 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__861_
timestamp 0
transform 1 0 1670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__862_
timestamp 0
transform -1 0 1730 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__863_
timestamp 0
transform 1 0 1850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__864_
timestamp 0
transform -1 0 990 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__865_
timestamp 0
transform 1 0 1450 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__866_
timestamp 0
transform -1 0 1730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__867_
timestamp 0
transform 1 0 2050 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__868_
timestamp 0
transform 1 0 2150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__869_
timestamp 0
transform 1 0 2130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__870_
timestamp 0
transform 1 0 1530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__871_
timestamp 0
transform 1 0 1390 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__872_
timestamp 0
transform -1 0 770 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__873_
timestamp 0
transform 1 0 1690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__874_
timestamp 0
transform 1 0 1130 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__875_
timestamp 0
transform 1 0 2010 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__876_
timestamp 0
transform -1 0 2210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__877_
timestamp 0
transform 1 0 1350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__878_
timestamp 0
transform 1 0 1570 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__879_
timestamp 0
transform 1 0 1850 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__880_
timestamp 0
transform -1 0 1630 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__881_
timestamp 0
transform 1 0 2370 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__882_
timestamp 0
transform 1 0 1790 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__883_
timestamp 0
transform 1 0 1950 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__884_
timestamp 0
transform -1 0 1890 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__885_
timestamp 0
transform 1 0 1250 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__886_
timestamp 0
transform 1 0 1750 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__887_
timestamp 0
transform -1 0 2350 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__888_
timestamp 0
transform 1 0 2450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__889_
timestamp 0
transform 1 0 2670 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__890_
timestamp 0
transform 1 0 1450 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__891_
timestamp 0
transform 1 0 2630 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__892_
timestamp 0
transform 1 0 2770 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__893_
timestamp 0
transform 1 0 3190 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__894_
timestamp 0
transform 1 0 2910 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__895_
timestamp 0
transform 1 0 3350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__896_
timestamp 0
transform 1 0 2470 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__897_
timestamp 0
transform 1 0 2890 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__898_
timestamp 0
transform 1 0 2610 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__899_
timestamp 0
transform -1 0 3130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__900_
timestamp 0
transform -1 0 2970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__901_
timestamp 0
transform 1 0 2790 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__902_
timestamp 0
transform 1 0 3550 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__903_
timestamp 0
transform 1 0 2590 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__904_
timestamp 0
transform -1 0 4510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__905_
timestamp 0
transform -1 0 4810 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__906_
timestamp 0
transform -1 0 5270 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__907_
timestamp 0
transform -1 0 4510 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__908_
timestamp 0
transform -1 0 4930 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__909_
timestamp 0
transform 1 0 4630 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__910_
timestamp 0
transform -1 0 4650 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__911_
timestamp 0
transform -1 0 4790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__912_
timestamp 0
transform 1 0 4310 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__913_
timestamp 0
transform -1 0 4770 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__914_
timestamp 0
transform 1 0 4330 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__915_
timestamp 0
transform 1 0 4310 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__916_
timestamp 0
transform -1 0 4610 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__917_
timestamp 0
transform -1 0 4930 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__918_
timestamp 0
transform 1 0 4150 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__919_
timestamp 0
transform -1 0 3730 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__920_
timestamp 0
transform 1 0 3550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__921_
timestamp 0
transform -1 0 3990 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__922_
timestamp 0
transform -1 0 4450 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__923_
timestamp 0
transform -1 0 3830 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__924_
timestamp 0
transform 1 0 2910 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__925_
timestamp 0
transform 1 0 1290 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__926_
timestamp 0
transform -1 0 3650 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__927_
timestamp 0
transform 1 0 3690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__928_
timestamp 0
transform 1 0 3390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__929_
timestamp 0
transform -1 0 3030 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__930_
timestamp 0
transform 1 0 2330 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__931_
timestamp 0
transform -1 0 2490 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__932_
timestamp 0
transform -1 0 3250 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__933_
timestamp 0
transform -1 0 2770 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__934_
timestamp 0
transform 1 0 2590 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__935_
timestamp 0
transform -1 0 2690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__936_
timestamp 0
transform 1 0 2350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__937_
timestamp 0
transform 1 0 2430 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__938_
timestamp 0
transform -1 0 2870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__939_
timestamp 0
transform -1 0 2530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__940_
timestamp 0
transform 1 0 2250 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__941_
timestamp 0
transform -1 0 2090 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__942_
timestamp 0
transform 1 0 2950 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__943_
timestamp 0
transform 1 0 2810 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__944_
timestamp 0
transform -1 0 2790 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__945_
timestamp 0
transform 1 0 2650 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__946_
timestamp 0
transform -1 0 2910 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__947_
timestamp 0
transform 1 0 3070 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__948_
timestamp 0
transform 1 0 3170 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__949_
timestamp 0
transform 1 0 1290 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__950_
timestamp 0
transform 1 0 1370 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__951_
timestamp 0
transform 1 0 1890 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__952_
timestamp 0
transform 1 0 3250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__953_
timestamp 0
transform 1 0 4830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__954_
timestamp 0
transform -1 0 4190 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__955_
timestamp 0
transform 1 0 3870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__956_
timestamp 0
transform 1 0 3050 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__957_
timestamp 0
transform 1 0 3190 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__958_
timestamp 0
transform 1 0 3290 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__959_
timestamp 0
transform -1 0 4130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__960_
timestamp 0
transform 1 0 2050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__961_
timestamp 0
transform 1 0 3410 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__962_
timestamp 0
transform 1 0 3470 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__963_
timestamp 0
transform 1 0 3930 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__964_
timestamp 0
transform 1 0 3630 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__965_
timestamp 0
transform 1 0 3470 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__966_
timestamp 0
transform 1 0 3790 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__967_
timestamp 0
transform 1 0 5210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__968_
timestamp 0
transform -1 0 5110 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__969_
timestamp 0
transform 1 0 4910 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__970_
timestamp 0
transform 1 0 5070 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__971_
timestamp 0
transform -1 0 5210 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__972_
timestamp 0
transform -1 0 5350 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__973_
timestamp 0
transform -1 0 5890 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__974_
timestamp 0
transform -1 0 5430 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__975_
timestamp 0
transform -1 0 5230 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__976_
timestamp 0
transform -1 0 5650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__977_
timestamp 0
transform 1 0 5570 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__978_
timestamp 0
transform -1 0 5750 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__979_
timestamp 0
transform -1 0 5570 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__980_
timestamp 0
transform -1 0 5410 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__981_
timestamp 0
transform -1 0 5870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__982_
timestamp 0
transform 1 0 5710 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__983_
timestamp 0
transform 1 0 5370 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__984_
timestamp 0
transform -1 0 5710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__985_
timestamp 0
transform -1 0 5230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__986_
timestamp 0
transform -1 0 5630 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__987_
timestamp 0
transform 1 0 5530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__988_
timestamp 0
transform 1 0 5430 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__989_
timestamp 0
transform -1 0 5130 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__990_
timestamp 0
transform 1 0 4030 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__991_
timestamp 0
transform 1 0 4150 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__992_
timestamp 0
transform -1 0 5450 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__993_
timestamp 0
transform -1 0 5390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__994_
timestamp 0
transform -1 0 5390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__995_
timestamp 0
transform -1 0 4870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__996_
timestamp 0
transform -1 0 4790 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__997_
timestamp 0
transform 1 0 4630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__998_
timestamp 0
transform -1 0 5250 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__999_
timestamp 0
transform -1 0 5050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1000_
timestamp 0
transform -1 0 4790 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1001_
timestamp 0
transform -1 0 4550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1002_
timestamp 0
transform -1 0 3350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1003_
timestamp 0
transform 1 0 3450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1004_
timestamp 0
transform -1 0 4710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1005_
timestamp 0
transform -1 0 4950 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1006_
timestamp 0
transform -1 0 4290 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1007_
timestamp 0
transform -1 0 3790 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1008_
timestamp 0
transform 1 0 4090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1009_
timestamp 0
transform -1 0 4610 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1010_
timestamp 0
transform -1 0 4390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1011_
timestamp 0
transform -1 0 4230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1012_
timestamp 0
transform -1 0 3630 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1013_
timestamp 0
transform 1 0 3870 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1014_
timestamp 0
transform -1 0 4330 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1015_
timestamp 0
transform 1 0 3930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1016_
timestamp 0
transform -1 0 4010 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1017_
timestamp 0
transform 1 0 3390 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1018_
timestamp 0
transform -1 0 3670 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1019_
timestamp 0
transform -1 0 3250 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1020_
timestamp 0
transform 1 0 3490 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1021_
timestamp 0
transform -1 0 3810 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1022_
timestamp 0
transform -1 0 4450 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1023_
timestamp 0
transform 1 0 4090 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1024_
timestamp 0
transform 1 0 4210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1025_
timestamp 0
transform 1 0 4350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1026_
timestamp 0
transform -1 0 5290 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1027_
timestamp 0
transform 1 0 5050 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1028_
timestamp 0
transform -1 0 2070 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1029_
timestamp 0
transform 1 0 3490 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1030_
timestamp 0
transform 1 0 2310 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1031_
timestamp 0
transform 1 0 2650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1032_
timestamp 0
transform -1 0 1830 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1033_
timestamp 0
transform -1 0 2190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1034_
timestamp 0
transform -1 0 1490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1035_
timestamp 0
transform 1 0 1750 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1036_
timestamp 0
transform 1 0 2770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1037_
timestamp 0
transform 1 0 1990 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1038_
timestamp 0
transform -1 0 2230 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1039_
timestamp 0
transform 1 0 1910 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1040_
timestamp 0
transform 1 0 2350 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1041_
timestamp 0
transform 1 0 4430 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1042_
timestamp 0
transform 1 0 3770 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1043_
timestamp 0
transform 1 0 3950 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1044_
timestamp 0
transform 1 0 3330 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1045_
timestamp 0
transform 1 0 2510 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1046_
timestamp 0
transform 1 0 2450 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1047_
timestamp 0
transform 1 0 3630 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1048_
timestamp 0
transform -1 0 3330 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1049_
timestamp 0
transform 1 0 2670 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1050_
timestamp 0
transform 1 0 3610 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1051_
timestamp 0
transform 1 0 2990 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1052_
timestamp 0
transform 1 0 2830 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1053_
timestamp 0
transform 1 0 3170 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1054_
timestamp 0
transform 1 0 4510 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1055_
timestamp 0
transform 1 0 5790 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1056_
timestamp 0
transform -1 0 5850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1057_
timestamp 0
transform 1 0 3770 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1058_
timestamp 0
transform 1 0 3810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1059_
timestamp 0
transform -1 0 4430 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1060_
timestamp 0
transform -1 0 4070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1061_
timestamp 0
transform -1 0 3710 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1062_
timestamp 0
transform 1 0 4230 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1063_
timestamp 0
transform 1 0 3650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1064_
timestamp 0
transform 1 0 3930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1065_
timestamp 0
transform 1 0 4270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1066_
timestamp 0
transform 1 0 3530 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1067_
timestamp 0
transform 1 0 4110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1068_
timestamp 0
transform -1 0 4890 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1069_
timestamp 0
transform 1 0 5530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1070_
timestamp 0
transform 1 0 5710 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1071_
timestamp 0
transform -1 0 5330 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1072_
timestamp 0
transform -1 0 5210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1073_
timestamp 0
transform -1 0 5790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1074_
timestamp 0
transform -1 0 5590 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1075_
timestamp 0
transform -1 0 5530 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1076_
timestamp 0
transform -1 0 5450 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1077_
timestamp 0
transform -1 0 5330 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1078_
timestamp 0
transform 1 0 5710 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1079_
timestamp 0
transform 1 0 5630 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1080_
timestamp 0
transform -1 0 5650 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1081_
timestamp 0
transform -1 0 5490 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1082_
timestamp 0
transform 1 0 5690 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1083_
timestamp 0
transform 1 0 5790 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1084_
timestamp 0
transform 1 0 5470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1085_
timestamp 0
transform -1 0 5830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1086_
timestamp 0
transform 1 0 5030 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1087_
timestamp 0
transform 1 0 5190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1088_
timestamp 0
transform -1 0 5850 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1089_
timestamp 0
transform 1 0 5530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1090_
timestamp 0
transform -1 0 5530 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1091_
timestamp 0
transform -1 0 5370 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1092_
timestamp 0
transform 1 0 5690 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1093_
timestamp 0
transform 1 0 5530 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1094_
timestamp 0
transform 1 0 5670 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1095_
timestamp 0
transform 1 0 5350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1096_
timestamp 0
transform -1 0 5730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1097_
timestamp 0
transform 1 0 4830 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1098_
timestamp 0
transform -1 0 4390 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1099_
timestamp 0
transform 1 0 5750 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1100_
timestamp 0
transform 1 0 5370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1101_
timestamp 0
transform -1 0 5550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1102_
timestamp 0
transform -1 0 5230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1103_
timestamp 0
transform -1 0 5130 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1104_
timestamp 0
transform 1 0 4950 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1105_
timestamp 0
transform -1 0 5610 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1106_
timestamp 0
transform 1 0 5010 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1107_
timestamp 0
transform -1 0 5130 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1108_
timestamp 0
transform -1 0 4290 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1109_
timestamp 0
transform -1 0 5290 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1110_
timestamp 0
transform -1 0 4950 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1111_
timestamp 0
transform -1 0 4790 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1112_
timestamp 0
transform -1 0 4130 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1113_
timestamp 0
transform 1 0 4650 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1114_
timestamp 0
transform 1 0 4490 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1115_
timestamp 0
transform -1 0 4610 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1116_
timestamp 0
transform 1 0 4430 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1117_
timestamp 0
transform -1 0 4490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1118_
timestamp 0
transform 1 0 4070 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1119_
timestamp 0
transform -1 0 3570 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1120_
timestamp 0
transform -1 0 3950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1121_
timestamp 0
transform -1 0 3950 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1122_
timestamp 0
transform -1 0 3770 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1123_
timestamp 0
transform -1 0 4790 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1124_
timestamp 0
transform 1 0 4590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1125_
timestamp 0
transform 1 0 3910 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1126_
timestamp 0
transform 1 0 4270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1127_
timestamp 0
transform -1 0 5210 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1128_
timestamp 0
transform 1 0 4670 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1129_
timestamp 0
transform 1 0 2930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1130_
timestamp 0
transform 1 0 2150 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1131_
timestamp 0
transform 1 0 2470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1132_
timestamp 0
transform 1 0 2170 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1133_
timestamp 0
transform 1 0 1990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1134_
timestamp 0
transform 1 0 2330 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1135_
timestamp 0
transform -1 0 1310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1136_
timestamp 0
transform -1 0 1690 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1137_
timestamp 0
transform 1 0 1670 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1138_
timestamp 0
transform 1 0 2750 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1139_
timestamp 0
transform -1 0 2310 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1140_
timestamp 0
transform 1 0 1830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1141_
timestamp 0
transform 1 0 2610 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1142_
timestamp 0
transform -1 0 4270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1143_
timestamp 0
transform -1 0 4070 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1144_
timestamp 0
transform 1 0 3090 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1145_
timestamp 0
transform 1 0 2450 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1146_
timestamp 0
transform 1 0 2590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1147_
timestamp 0
transform -1 0 4390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1148_
timestamp 0
transform 1 0 3410 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1149_
timestamp 0
transform 1 0 3470 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1150_
timestamp 0
transform 1 0 2770 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1151_
timestamp 0
transform -1 0 2950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1152_
timestamp 0
transform 1 0 3110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1153_
timestamp 0
transform 1 0 3090 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1154_
timestamp 0
transform 1 0 2930 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1155_
timestamp 0
transform 1 0 3250 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1156_
timestamp 0
transform -1 0 3650 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1157_
timestamp 0
transform -1 0 5310 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1158_
timestamp 0
transform -1 0 5150 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1159_
timestamp 0
transform -1 0 3930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1160_
timestamp 0
transform -1 0 3890 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1161_
timestamp 0
transform 1 0 2870 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1162_
timestamp 0
transform -1 0 3590 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1163_
timestamp 0
transform -1 0 1610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1164_
timestamp 0
transform 1 0 3210 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1165_
timestamp 0
transform 1 0 3710 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1166_
timestamp 0
transform 1 0 4150 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1167_
timestamp 0
transform 1 0 4310 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1168_
timestamp 0
transform 1 0 4470 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1169_
timestamp 0
transform 1 0 4630 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1170_
timestamp 0
transform 1 0 4790 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1171_
timestamp 0
transform -1 0 5630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1172_
timestamp 0
transform -1 0 5470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1173_
timestamp 0
transform -1 0 5790 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1174_
timestamp 0
transform 1 0 5790 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1175_
timestamp 0
transform 1 0 5590 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1176_
timestamp 0
transform -1 0 5450 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1177_
timestamp 0
transform -1 0 5510 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1178_
timestamp 0
transform -1 0 5290 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1179_
timestamp 0
transform -1 0 4970 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1180_
timestamp 0
transform 1 0 5710 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1181_
timestamp 0
transform 1 0 5770 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1182_
timestamp 0
transform -1 0 5770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1183_
timestamp 0
transform -1 0 5450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1184_
timestamp 0
transform 1 0 4890 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1185_
timestamp 0
transform 1 0 4990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1186_
timestamp 0
transform -1 0 5030 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1187_
timestamp 0
transform -1 0 4870 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1188_
timestamp 0
transform 1 0 4730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1189_
timestamp 0
transform 1 0 5090 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1190_
timestamp 0
transform 1 0 5110 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1191_
timestamp 0
transform -1 0 4950 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1192_
timestamp 0
transform -1 0 4890 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1193_
timestamp 0
transform 1 0 3770 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1194_
timestamp 0
transform 1 0 5150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1195_
timestamp 0
transform -1 0 4850 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1196_
timestamp 0
transform -1 0 4630 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1197_
timestamp 0
transform 1 0 4550 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1198_
timestamp 0
transform -1 0 4750 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1199_
timestamp 0
transform -1 0 4590 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1200_
timestamp 0
transform -1 0 4790 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1201_
timestamp 0
transform 1 0 5030 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1202_
timestamp 0
transform -1 0 4550 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1203_
timestamp 0
transform -1 0 4210 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1204_
timestamp 0
transform -1 0 4710 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1205_
timestamp 0
transform -1 0 4410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1206_
timestamp 0
transform -1 0 3970 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1207_
timestamp 0
transform 1 0 3830 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1208_
timestamp 0
transform -1 0 5070 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1209_
timestamp 0
transform 1 0 4890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1210_
timestamp 0
transform -1 0 4130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1211_
timestamp 0
transform -1 0 4390 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1212_
timestamp 0
transform -1 0 4030 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1213_
timestamp 0
transform 1 0 4030 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1214_
timestamp 0
transform -1 0 3190 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1215_
timestamp 0
transform 1 0 3730 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1216_
timestamp 0
transform 1 0 3850 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1217_
timestamp 0
transform -1 0 4730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1218_
timestamp 0
transform 1 0 4450 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1219_
timestamp 0
transform 1 0 3250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1220_
timestamp 0
transform 1 0 5090 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1221_
timestamp 0
transform 1 0 5250 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1222_
timestamp 0
transform 1 0 1990 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1223_
timestamp 0
transform 1 0 2850 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1224_
timestamp 0
transform -1 0 2290 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1225_
timestamp 0
transform 1 0 2030 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1226_
timestamp 0
transform 1 0 1590 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1227_
timestamp 0
transform -1 0 1770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1228_
timestamp 0
transform 1 0 2590 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1229_
timestamp 0
transform 1 0 2750 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1230_
timestamp 0
transform 1 0 2210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1231_
timestamp 0
transform -1 0 2430 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1232_
timestamp 0
transform -1 0 2590 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1233_
timestamp 0
transform 1 0 2910 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1234_
timestamp 0
transform 1 0 3990 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1235_
timestamp 0
transform -1 0 3750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1236_
timestamp 0
transform 1 0 3570 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1237_
timestamp 0
transform 1 0 2750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1238_
timestamp 0
transform 1 0 2350 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1239_
timestamp 0
transform -1 0 3390 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1240_
timestamp 0
transform 1 0 3070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1241_
timestamp 0
transform 1 0 3050 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1242_
timestamp 0
transform 1 0 3010 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1243_
timestamp 0
transform -1 0 3430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1244_
timestamp 0
transform 1 0 3230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1245_
timestamp 0
transform 1 0 3370 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1246_
timestamp 0
transform 1 0 4870 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1247_
timestamp 0
transform -1 0 5590 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1248_
timestamp 0
transform 1 0 5410 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1249_
timestamp 0
transform -1 0 3550 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1250_
timestamp 0
transform 1 0 3090 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1251_
timestamp 0
transform -1 0 2770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1252_
timestamp 0
transform -1 0 2970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1253_
timestamp 0
transform -1 0 1030 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1254_
timestamp 0
transform 1 0 2910 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1255_
timestamp 0
transform 1 0 3210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1256_
timestamp 0
transform 1 0 3090 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1257_
timestamp 0
transform 1 0 3250 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1258_
timestamp 0
transform 1 0 3470 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1259_
timestamp 0
transform -1 0 5710 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1260_
timestamp 0
transform -1 0 5270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1261_
timestamp 0
transform -1 0 5430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1262_
timestamp 0
transform 1 0 5810 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1263_
timestamp 0
transform -1 0 5690 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1264_
timestamp 0
transform -1 0 5590 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1265_
timestamp 0
transform -1 0 5610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1266_
timestamp 0
transform 1 0 5270 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1267_
timestamp 0
transform -1 0 5750 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1268_
timestamp 0
transform 1 0 5730 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1269_
timestamp 0
transform -1 0 5450 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1270_
timestamp 0
transform 1 0 5030 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1271_
timestamp 0
transform 1 0 5650 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1272_
timestamp 0
transform -1 0 5410 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1273_
timestamp 0
transform -1 0 5250 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1274_
timestamp 0
transform -1 0 4950 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1275_
timestamp 0
transform -1 0 4730 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1276_
timestamp 0
transform 1 0 4530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1277_
timestamp 0
transform 1 0 5590 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1278_
timestamp 0
transform -1 0 5530 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1279_
timestamp 0
transform -1 0 5370 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1280_
timestamp 0
transform 1 0 5170 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1281_
timestamp 0
transform -1 0 4750 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1282_
timestamp 0
transform -1 0 4590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1283_
timestamp 0
transform 1 0 4610 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1284_
timestamp 0
transform 1 0 5250 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1285_
timestamp 0
transform -1 0 4770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1286_
timestamp 0
transform -1 0 4930 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1287_
timestamp 0
transform -1 0 4430 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1288_
timestamp 0
transform 1 0 4170 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1289_
timestamp 0
transform 1 0 4290 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1290_
timestamp 0
transform -1 0 5090 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1291_
timestamp 0
transform -1 0 4470 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1292_
timestamp 0
transform -1 0 4310 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1293_
timestamp 0
transform 1 0 4130 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1294_
timestamp 0
transform -1 0 3550 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1295_
timestamp 0
transform -1 0 4290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1296_
timestamp 0
transform 1 0 3970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1297_
timestamp 0
transform -1 0 3710 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1298_
timestamp 0
transform 1 0 3810 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1299_
timestamp 0
transform -1 0 4350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1300_
timestamp 0
transform 1 0 4170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1301_
timestamp 0
transform 1 0 3830 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1302_
timestamp 0
transform 1 0 4830 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1303_
timestamp 0
transform -1 0 5090 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1304_
timestamp 0
transform 1 0 2570 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1305_
timestamp 0
transform -1 0 1910 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1306_
timestamp 0
transform 1 0 1510 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1307_
timestamp 0
transform -1 0 1670 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1308_
timestamp 0
transform -1 0 1670 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1309_
timestamp 0
transform 1 0 1950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1310_
timestamp 0
transform 1 0 2110 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1311_
timestamp 0
transform 1 0 1830 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1312_
timestamp 0
transform -1 0 2150 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1313_
timestamp 0
transform 1 0 1970 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1314_
timestamp 0
transform 1 0 2410 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1315_
timestamp 0
transform 1 0 2650 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1316_
timestamp 0
transform 1 0 2790 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1317_
timestamp 0
transform 1 0 2650 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1318_
timestamp 0
transform 1 0 2230 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1319_
timestamp 0
transform -1 0 1730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1320_
timestamp 0
transform -1 0 3330 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1321_
timestamp 0
transform -1 0 3170 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1322_
timestamp 0
transform 1 0 2310 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1323_
timestamp 0
transform 1 0 2810 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1324_
timestamp 0
transform 1 0 2630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1325_
timestamp 0
transform 1 0 2470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1326_
timestamp 0
transform 1 0 2490 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1327_
timestamp 0
transform 1 0 2970 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1328_
timestamp 0
transform -1 0 3550 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1329_
timestamp 0
transform -1 0 5570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1330_
timestamp 0
transform -1 0 5390 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1331_
timestamp 0
transform 1 0 2290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1332_
timestamp 0
transform 1 0 2130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1333_
timestamp 0
transform 1 0 2490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1334_
timestamp 0
transform -1 0 3070 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1335_
timestamp 0
transform -1 0 2510 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1336_
timestamp 0
transform -1 0 2330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1337_
timestamp 0
transform 1 0 2330 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1338_
timestamp 0
transform 1 0 3190 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1339_
timestamp 0
transform -1 0 4110 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1340_
timestamp 0
transform 1 0 3990 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1341_
timestamp 0
transform 1 0 3350 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1342_
timestamp 0
transform 1 0 4290 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1343_
timestamp 0
transform 1 0 3330 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1344_
timestamp 0
transform -1 0 5230 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1345_
timestamp 0
transform 1 0 4430 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1346_
timestamp 0
transform -1 0 4150 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1347_
timestamp 0
transform 1 0 4910 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1348_
timestamp 0
transform -1 0 5290 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1349_
timestamp 0
transform 1 0 3670 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1350_
timestamp 0
transform -1 0 3850 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1351_
timestamp 0
transform 1 0 4590 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1352_
timestamp 0
transform -1 0 5130 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1353_
timestamp 0
transform 1 0 4270 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1354_
timestamp 0
transform -1 0 4770 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1355_
timestamp 0
transform -1 0 4550 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1356_
timestamp 0
transform -1 0 4390 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1357_
timestamp 0
transform -1 0 5110 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1358_
timestamp 0
transform -1 0 4610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1359_
timestamp 0
transform 1 0 4650 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1360_
timestamp 0
transform -1 0 4970 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1361_
timestamp 0
transform -1 0 4730 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1362_
timestamp 0
transform 1 0 4230 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1363_
timestamp 0
transform 1 0 3970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1364_
timestamp 0
transform -1 0 3870 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1365_
timestamp 0
transform -1 0 4370 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1366_
timestamp 0
transform -1 0 4210 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1367_
timestamp 0
transform 1 0 2770 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1368_
timestamp 0
transform 1 0 3250 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1369_
timestamp 0
transform 1 0 3950 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1370_
timestamp 0
transform -1 0 3810 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1371_
timestamp 0
transform 1 0 2130 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1372_
timestamp 0
transform -1 0 1550 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1373_
timestamp 0
transform -1 0 1450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1374_
timestamp 0
transform 1 0 1090 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1375_
timestamp 0
transform 1 0 1370 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1376_
timestamp 0
transform 1 0 1210 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1377_
timestamp 0
transform -1 0 1170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1378_
timestamp 0
transform -1 0 1810 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1379_
timestamp 0
transform 1 0 1390 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1380_
timestamp 0
transform 1 0 1250 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1381_
timestamp 0
transform 1 0 1310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1382_
timestamp 0
transform 1 0 1450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1383_
timestamp 0
transform 1 0 1690 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1384_
timestamp 0
transform -1 0 2050 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1385_
timestamp 0
transform -1 0 1710 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1386_
timestamp 0
transform -1 0 1550 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1387_
timestamp 0
transform -1 0 1110 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1388_
timestamp 0
transform 1 0 1530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1389_
timestamp 0
transform -1 0 1850 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1390_
timestamp 0
transform -1 0 2210 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1391_
timestamp 0
transform 1 0 1850 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1392_
timestamp 0
transform 1 0 1370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1393_
timestamp 0
transform -1 0 1830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1394_
timestamp 0
transform 1 0 2550 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1395_
timestamp 0
transform 1 0 2910 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1396_
timestamp 0
transform -1 0 2750 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1397_
timestamp 0
transform -1 0 2610 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1398_
timestamp 0
transform -1 0 2370 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1399_
timestamp 0
transform 1 0 2170 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1400_
timestamp 0
transform 1 0 1970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1401_
timestamp 0
transform 1 0 1990 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1402_
timestamp 0
transform 1 0 2470 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1403_
timestamp 0
transform -1 0 2930 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1404_
timestamp 0
transform -1 0 3230 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1405_
timestamp 0
transform -1 0 3670 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1406_
timestamp 0
transform -1 0 3510 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1407_
timestamp 0
transform 1 0 2950 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1408_
timestamp 0
transform 1 0 3590 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1409_
timestamp 0
transform 1 0 2790 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1410_
timestamp 0
transform -1 0 3070 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1411_
timestamp 0
transform 1 0 3270 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1412_
timestamp 0
transform 1 0 3750 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1413_
timestamp 0
transform 1 0 4430 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1414_
timestamp 0
transform -1 0 4490 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1415_
timestamp 0
transform -1 0 3130 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1416_
timestamp 0
transform 1 0 3430 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1417_
timestamp 0
transform -1 0 3930 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1418_
timestamp 0
transform 1 0 3570 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1419_
timestamp 0
transform 1 0 3530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1420_
timestamp 0
transform 1 0 4030 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1421_
timestamp 0
transform 1 0 3670 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1422_
timestamp 0
transform -1 0 3390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1423_
timestamp 0
transform -1 0 4090 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1424_
timestamp 0
transform -1 0 3410 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1425_
timestamp 0
transform 1 0 3710 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1426_
timestamp 0
transform 1 0 2910 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1427_
timestamp 0
transform -1 0 2630 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1428_
timestamp 0
transform 1 0 1670 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1429_
timestamp 0
transform -1 0 1170 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1430_
timestamp 0
transform -1 0 2450 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1431_
timestamp 0
transform 1 0 1370 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1432_
timestamp 0
transform 1 0 630 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1433_
timestamp 0
transform -1 0 1270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1434_
timestamp 0
transform 1 0 1090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1435_
timestamp 0
transform 1 0 1050 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1436_
timestamp 0
transform 1 0 950 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1437_
timestamp 0
transform 1 0 910 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1438_
timestamp 0
transform -1 0 1070 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1439_
timestamp 0
transform -1 0 770 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1440_
timestamp 0
transform 1 0 1210 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1441_
timestamp 0
transform -1 0 470 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1442_
timestamp 0
transform 1 0 10 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1443_
timestamp 0
transform -1 0 2430 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1444_
timestamp 0
transform -1 0 170 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1445_
timestamp 0
transform 1 0 450 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1446_
timestamp 0
transform -1 0 330 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1447_
timestamp 0
transform -1 0 30 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1448_
timestamp 0
transform 1 0 150 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1449_
timestamp 0
transform -1 0 610 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1450_
timestamp 0
transform -1 0 610 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1451_
timestamp 0
transform -1 0 890 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1452_
timestamp 0
transform -1 0 890 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1453_
timestamp 0
transform -1 0 750 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1454_
timestamp 0
transform 1 0 990 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1455_
timestamp 0
transform 1 0 1030 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1456_
timestamp 0
transform 1 0 1190 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1457_
timestamp 0
transform -1 0 2050 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1458_
timestamp 0
transform -1 0 2650 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1459_
timestamp 0
transform -1 0 2770 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1460_
timestamp 0
transform -1 0 1870 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1461_
timestamp 0
transform 1 0 1770 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1462_
timestamp 0
transform -1 0 1930 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1463_
timestamp 0
transform 1 0 1730 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1464_
timestamp 0
transform -1 0 1590 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1465_
timestamp 0
transform 1 0 1270 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1466_
timestamp 0
transform 1 0 770 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1467_
timestamp 0
transform -1 0 570 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1468_
timestamp 0
transform 1 0 910 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1469_
timestamp 0
transform 1 0 610 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1470_
timestamp 0
transform -1 0 1230 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1471_
timestamp 0
transform 1 0 750 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1472_
timestamp 0
transform -1 0 30 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1473_
timestamp 0
transform -1 0 30 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1474_
timestamp 0
transform -1 0 30 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1475_
timestamp 0
transform 1 0 510 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1476_
timestamp 0
transform 1 0 190 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1477_
timestamp 0
transform 1 0 630 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1478_
timestamp 0
transform 1 0 290 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1479_
timestamp 0
transform 1 0 210 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1480_
timestamp 0
transform -1 0 370 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1481_
timestamp 0
transform 1 0 350 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1482_
timestamp 0
transform -1 0 810 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1483_
timestamp 0
transform -1 0 1390 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1484_
timestamp 0
transform -1 0 1470 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1485_
timestamp 0
transform -1 0 1310 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1486_
timestamp 0
transform -1 0 1630 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1487_
timestamp 0
transform -1 0 1410 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1488_
timestamp 0
transform 1 0 1430 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1489_
timestamp 0
transform 1 0 1210 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1490_
timestamp 0
transform 1 0 490 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1491_
timestamp 0
transform -1 0 790 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1492_
timestamp 0
transform 1 0 610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1493_
timestamp 0
transform -1 0 490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1494_
timestamp 0
transform 1 0 190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1495_
timestamp 0
transform 1 0 310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1496_
timestamp 0
transform 1 0 710 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1497_
timestamp 0
transform 1 0 210 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1498_
timestamp 0
transform 1 0 10 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1499_
timestamp 0
transform -1 0 230 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1500_
timestamp 0
transform 1 0 850 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1501_
timestamp 0
transform -1 0 950 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1502_
timestamp 0
transform -1 0 930 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1503_
timestamp 0
transform -1 0 910 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1504_
timestamp 0
transform 1 0 610 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1505_
timestamp 0
transform -1 0 750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1506_
timestamp 0
transform -1 0 570 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1507_
timestamp 0
transform 1 0 10 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1508_
timestamp 0
transform -1 0 30 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1509_
timestamp 0
transform -1 0 370 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1510_
timestamp 0
transform 1 0 270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1511_
timestamp 0
transform 1 0 3050 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1512_
timestamp 0
transform -1 0 1530 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1513_
timestamp 0
transform -1 0 1150 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1514_
timestamp 0
transform -1 0 1070 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1515_
timestamp 0
transform -1 0 170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1516_
timestamp 0
transform -1 0 570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1517_
timestamp 0
transform -1 0 430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1518_
timestamp 0
transform 1 0 1270 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1519_
timestamp 0
transform 1 0 2170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1560_
timestamp 0
transform -1 0 30 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1561_
timestamp 0
transform -1 0 170 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1562_
timestamp 0
transform -1 0 30 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1563_
timestamp 0
transform -1 0 30 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1564_
timestamp 0
transform -1 0 310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1565_
timestamp 0
transform 1 0 3850 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1566_
timestamp 0
transform -1 0 970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1567_
timestamp 0
transform -1 0 30 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1568_
timestamp 0
transform -1 0 30 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1569_
timestamp 0
transform -1 0 30 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1570_
timestamp 0
transform -1 0 3670 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1571_
timestamp 0
transform 1 0 5070 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1572_
timestamp 0
transform -1 0 2310 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1573_
timestamp 0
transform 1 0 2150 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1574_
timestamp 0
transform -1 0 30 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1575_
timestamp 0
transform -1 0 190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1576_
timestamp 0
transform -1 0 30 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1577_
timestamp 0
transform -1 0 330 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1578_
timestamp 0
transform 1 0 1570 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1579_
timestamp 0
transform 1 0 2190 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1580_
timestamp 0
transform -1 0 2710 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1581_
timestamp 0
transform -1 0 3050 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1582_
timestamp 0
transform -1 0 30 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1583_
timestamp 0
transform -1 0 3230 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert6
timestamp 0
transform 1 0 5050 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert7
timestamp 0
transform -1 0 3090 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert8
timestamp 0
transform -1 0 3090 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert9
timestamp 0
transform -1 0 5810 0 -1 270
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert10
timestamp 0
transform 1 0 1610 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert11
timestamp 0
transform 1 0 1730 0 1 4430
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert12
timestamp 0
transform 1 0 1490 0 1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert13
timestamp 0
transform -1 0 30 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert14
timestamp 0
transform -1 0 2730 0 1 2350
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert15
timestamp 0
transform -1 0 4030 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert16
timestamp 0
transform 1 0 4230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert17
timestamp 0
transform 1 0 4150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert0
timestamp 0
transform 1 0 1410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert1
timestamp 0
transform -1 0 1250 0 1 3390
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert2
timestamp 0
transform -1 0 710 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert3
timestamp 0
transform -1 0 1050 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert4
timestamp 0
transform -1 0 1030 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert5
timestamp 0
transform 1 0 2990 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__756_
timestamp 0
transform 1 0 1290 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__757_
timestamp 0
transform 1 0 1650 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__758_
timestamp 0
transform 1 0 1410 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__759_
timestamp 0
transform 1 0 550 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__760_
timestamp 0
transform 1 0 690 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__761_
timestamp 0
transform 1 0 410 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__762_
timestamp 0
transform 1 0 410 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__763_
timestamp 0
transform -1 0 1150 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__764_
timestamp 0
transform 1 0 930 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__765_
timestamp 0
transform -1 0 430 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__766_
timestamp 0
transform 1 0 590 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__767_
timestamp 0
transform 1 0 750 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__768_
timestamp 0
transform -1 0 890 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__769_
timestamp 0
transform 1 0 670 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__770_
timestamp 0
transform 1 0 810 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__771_
timestamp 0
transform 1 0 970 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__772_
timestamp 0
transform -1 0 1150 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__773_
timestamp 0
transform -1 0 830 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__774_
timestamp 0
transform 1 0 650 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__775_
timestamp 0
transform -1 0 3110 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__776_
timestamp 0
transform -1 0 1450 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__777_
timestamp 0
transform -1 0 990 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__778_
timestamp 0
transform 1 0 350 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__779_
timestamp 0
transform 1 0 510 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__780_
timestamp 0
transform 1 0 30 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__781_
timestamp 0
transform 1 0 30 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__782_
timestamp 0
transform 1 0 470 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__783_
timestamp 0
transform 1 0 590 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__784_
timestamp 0
transform 1 0 190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__785_
timestamp 0
transform 1 0 310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__786_
timestamp 0
transform -1 0 790 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__787_
timestamp 0
transform 1 0 930 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__788_
timestamp 0
transform 1 0 1570 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__789_
timestamp 0
transform -1 0 1170 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__790_
timestamp 0
transform -1 0 1330 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__791_
timestamp 0
transform 1 0 1270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__792_
timestamp 0
transform -1 0 1410 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__793_
timestamp 0
transform -1 0 1010 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__794_
timestamp 0
transform 1 0 930 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__795_
timestamp 0
transform -1 0 850 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__796_
timestamp 0
transform 1 0 790 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__797_
timestamp 0
transform 1 0 1090 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__798_
timestamp 0
transform -1 0 890 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__799_
timestamp 0
transform -1 0 3450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__800_
timestamp 0
transform 1 0 2210 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__801_
timestamp 0
transform 1 0 2290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__802_
timestamp 0
transform 1 0 1870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__803_
timestamp 0
transform -1 0 1570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__804_
timestamp 0
transform -1 0 1270 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__805_
timestamp 0
transform -1 0 210 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__806_
timestamp 0
transform -1 0 750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__807_
timestamp 0
transform 1 0 850 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__808_
timestamp 0
transform 1 0 450 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__809_
timestamp 0
transform 1 0 30 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__810_
timestamp 0
transform -1 0 210 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__811_
timestamp 0
transform 1 0 150 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__812_
timestamp 0
transform -1 0 710 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__813_
timestamp 0
transform -1 0 330 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__814_
timestamp 0
transform -1 0 50 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__815_
timestamp 0
transform 1 0 350 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__816_
timestamp 0
transform 1 0 410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__817_
timestamp 0
transform -1 0 50 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__818_
timestamp 0
transform -1 0 210 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__819_
timestamp 0
transform -1 0 550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__820_
timestamp 0
transform -1 0 170 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__821_
timestamp 0
transform 1 0 890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__822_
timestamp 0
transform 1 0 2010 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__823_
timestamp 0
transform -1 0 1730 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__824_
timestamp 0
transform 1 0 630 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__825_
timestamp 0
transform 1 0 570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__826_
timestamp 0
transform 1 0 930 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__827_
timestamp 0
transform -1 0 1250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__828_
timestamp 0
transform 1 0 730 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__829_
timestamp 0
transform -1 0 1070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__830_
timestamp 0
transform 1 0 330 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__831_
timestamp 0
transform -1 0 1470 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__832_
timestamp 0
transform 1 0 570 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__833_
timestamp 0
transform -1 0 1150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__834_
timestamp 0
transform 1 0 2070 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__835_
timestamp 0
transform 1 0 1090 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__836_
timestamp 0
transform 1 0 610 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__837_
timestamp 0
transform 1 0 970 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__838_
timestamp 0
transform -1 0 2390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__839_
timestamp 0
transform -1 0 2570 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__840_
timestamp 0
transform -1 0 1750 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__841_
timestamp 0
transform -1 0 2550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__842_
timestamp 0
transform 1 0 2070 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__843_
timestamp 0
transform -1 0 1810 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__844_
timestamp 0
transform 1 0 1850 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__845_
timestamp 0
transform -1 0 1930 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__846_
timestamp 0
transform -1 0 1590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__847_
timestamp 0
transform -1 0 970 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__848_
timestamp 0
transform 1 0 770 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__849_
timestamp 0
transform -1 0 1990 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__850_
timestamp 0
transform -1 0 1650 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__851_
timestamp 0
transform -1 0 1330 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__852_
timestamp 0
transform 1 0 2330 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__853_
timestamp 0
transform 1 0 2770 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__854_
timestamp 0
transform 1 0 2030 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__855_
timestamp 0
transform -1 0 1590 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__856_
timestamp 0
transform 1 0 1570 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__857_
timestamp 0
transform -1 0 1910 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__858_
timestamp 0
transform -1 0 2250 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__859_
timestamp 0
transform 1 0 2650 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__860_
timestamp 0
transform -1 0 2510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__861_
timestamp 0
transform 1 0 1690 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__862_
timestamp 0
transform -1 0 1750 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__863_
timestamp 0
transform 1 0 1870 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__864_
timestamp 0
transform -1 0 1010 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__865_
timestamp 0
transform 1 0 1470 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__866_
timestamp 0
transform -1 0 1750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__867_
timestamp 0
transform 1 0 2070 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__868_
timestamp 0
transform 1 0 2170 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__869_
timestamp 0
transform 1 0 2150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__870_
timestamp 0
transform 1 0 1550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__871_
timestamp 0
transform 1 0 1410 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__872_
timestamp 0
transform -1 0 790 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__873_
timestamp 0
transform 1 0 1710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__874_
timestamp 0
transform 1 0 1150 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__875_
timestamp 0
transform 1 0 2030 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__876_
timestamp 0
transform -1 0 2230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__877_
timestamp 0
transform 1 0 1370 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__878_
timestamp 0
transform 1 0 1590 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__879_
timestamp 0
transform 1 0 1870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__880_
timestamp 0
transform -1 0 1650 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__881_
timestamp 0
transform 1 0 2390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__882_
timestamp 0
transform 1 0 1810 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__883_
timestamp 0
transform 1 0 1970 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__884_
timestamp 0
transform -1 0 1910 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__885_
timestamp 0
transform 1 0 1270 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__886_
timestamp 0
transform 1 0 1770 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__887_
timestamp 0
transform -1 0 2370 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__888_
timestamp 0
transform 1 0 2470 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__889_
timestamp 0
transform 1 0 2690 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__890_
timestamp 0
transform 1 0 1470 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__891_
timestamp 0
transform 1 0 2650 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__892_
timestamp 0
transform 1 0 2790 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__893_
timestamp 0
transform 1 0 3210 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__894_
timestamp 0
transform 1 0 2930 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__895_
timestamp 0
transform 1 0 3370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__896_
timestamp 0
transform 1 0 2490 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__897_
timestamp 0
transform 1 0 2910 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__898_
timestamp 0
transform 1 0 2630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__899_
timestamp 0
transform -1 0 3150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__900_
timestamp 0
transform -1 0 2990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__901_
timestamp 0
transform 1 0 2810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__902_
timestamp 0
transform 1 0 3570 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__903_
timestamp 0
transform 1 0 2610 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__904_
timestamp 0
transform -1 0 4530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__905_
timestamp 0
transform -1 0 4830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__906_
timestamp 0
transform -1 0 5290 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__907_
timestamp 0
transform -1 0 4530 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__908_
timestamp 0
transform -1 0 4950 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__909_
timestamp 0
transform 1 0 4650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__910_
timestamp 0
transform -1 0 4670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__911_
timestamp 0
transform -1 0 4810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__912_
timestamp 0
transform 1 0 4330 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__913_
timestamp 0
transform -1 0 4790 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__914_
timestamp 0
transform 1 0 4350 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__915_
timestamp 0
transform 1 0 4330 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__916_
timestamp 0
transform -1 0 4630 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__917_
timestamp 0
transform -1 0 4950 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__918_
timestamp 0
transform 1 0 4170 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__919_
timestamp 0
transform -1 0 3750 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__920_
timestamp 0
transform 1 0 3570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__921_
timestamp 0
transform -1 0 4010 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__922_
timestamp 0
transform -1 0 4470 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__923_
timestamp 0
transform -1 0 3850 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__924_
timestamp 0
transform 1 0 2930 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__925_
timestamp 0
transform 1 0 1310 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__926_
timestamp 0
transform -1 0 3670 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__927_
timestamp 0
transform 1 0 3710 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__928_
timestamp 0
transform 1 0 3410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__929_
timestamp 0
transform -1 0 3050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__930_
timestamp 0
transform 1 0 2350 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__931_
timestamp 0
transform -1 0 2510 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__932_
timestamp 0
transform -1 0 3270 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__933_
timestamp 0
transform -1 0 2790 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__934_
timestamp 0
transform 1 0 2610 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__935_
timestamp 0
transform -1 0 2710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__936_
timestamp 0
transform 1 0 2370 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__937_
timestamp 0
transform 1 0 2450 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__938_
timestamp 0
transform -1 0 2890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__939_
timestamp 0
transform -1 0 2550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__940_
timestamp 0
transform 1 0 2270 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__941_
timestamp 0
transform -1 0 2110 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__942_
timestamp 0
transform 1 0 2970 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__943_
timestamp 0
transform 1 0 2830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__944_
timestamp 0
transform -1 0 2810 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__945_
timestamp 0
transform 1 0 2670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__946_
timestamp 0
transform -1 0 2930 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__947_
timestamp 0
transform 1 0 3090 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__948_
timestamp 0
transform 1 0 3190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__949_
timestamp 0
transform 1 0 1310 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__950_
timestamp 0
transform 1 0 1390 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__951_
timestamp 0
transform 1 0 1910 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__952_
timestamp 0
transform 1 0 3270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__953_
timestamp 0
transform 1 0 4850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__954_
timestamp 0
transform -1 0 4210 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__955_
timestamp 0
transform 1 0 3890 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__956_
timestamp 0
transform 1 0 3070 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__957_
timestamp 0
transform 1 0 3210 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__958_
timestamp 0
transform 1 0 3310 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__959_
timestamp 0
transform -1 0 4150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__960_
timestamp 0
transform 1 0 2070 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__961_
timestamp 0
transform 1 0 3430 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__962_
timestamp 0
transform 1 0 3490 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__963_
timestamp 0
transform 1 0 3950 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__964_
timestamp 0
transform 1 0 3650 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__965_
timestamp 0
transform 1 0 3490 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__966_
timestamp 0
transform 1 0 3810 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__967_
timestamp 0
transform 1 0 5230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__968_
timestamp 0
transform -1 0 5130 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__969_
timestamp 0
transform 1 0 4930 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__970_
timestamp 0
transform 1 0 5090 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__971_
timestamp 0
transform -1 0 5230 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__972_
timestamp 0
transform -1 0 5370 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__973_
timestamp 0
transform -1 0 5910 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__974_
timestamp 0
transform -1 0 5450 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__975_
timestamp 0
transform -1 0 5250 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__976_
timestamp 0
transform -1 0 5670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__977_
timestamp 0
transform 1 0 5590 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__978_
timestamp 0
transform -1 0 5770 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__979_
timestamp 0
transform -1 0 5590 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__980_
timestamp 0
transform -1 0 5430 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__981_
timestamp 0
transform -1 0 5890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__982_
timestamp 0
transform 1 0 5730 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__983_
timestamp 0
transform 1 0 5390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__984_
timestamp 0
transform -1 0 5730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__985_
timestamp 0
transform -1 0 5250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__986_
timestamp 0
transform -1 0 5650 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__987_
timestamp 0
transform 1 0 5550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__988_
timestamp 0
transform 1 0 5450 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__989_
timestamp 0
transform -1 0 5150 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__990_
timestamp 0
transform 1 0 4050 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__991_
timestamp 0
transform 1 0 4170 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__992_
timestamp 0
transform -1 0 5470 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__993_
timestamp 0
transform -1 0 5410 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__994_
timestamp 0
transform -1 0 5410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__995_
timestamp 0
transform -1 0 4890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__996_
timestamp 0
transform -1 0 4810 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__997_
timestamp 0
transform 1 0 4650 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__998_
timestamp 0
transform -1 0 5270 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__999_
timestamp 0
transform -1 0 5070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1000_
timestamp 0
transform -1 0 4810 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1001_
timestamp 0
transform -1 0 4570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1002_
timestamp 0
transform -1 0 3370 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1003_
timestamp 0
transform 1 0 3470 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1004_
timestamp 0
transform -1 0 4730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1005_
timestamp 0
transform -1 0 4970 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1006_
timestamp 0
transform -1 0 4310 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1007_
timestamp 0
transform -1 0 3810 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1008_
timestamp 0
transform 1 0 4110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1009_
timestamp 0
transform -1 0 4630 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1010_
timestamp 0
transform -1 0 4410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1011_
timestamp 0
transform -1 0 4250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1012_
timestamp 0
transform -1 0 3650 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1013_
timestamp 0
transform 1 0 3890 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1014_
timestamp 0
transform -1 0 4350 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1015_
timestamp 0
transform 1 0 3950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1016_
timestamp 0
transform -1 0 4030 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1017_
timestamp 0
transform 1 0 3410 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1018_
timestamp 0
transform -1 0 3690 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1019_
timestamp 0
transform -1 0 3270 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1020_
timestamp 0
transform 1 0 3510 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1021_
timestamp 0
transform -1 0 3830 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1022_
timestamp 0
transform -1 0 4470 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1023_
timestamp 0
transform 1 0 4110 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1024_
timestamp 0
transform 1 0 4230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1025_
timestamp 0
transform 1 0 4370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1026_
timestamp 0
transform -1 0 5310 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1027_
timestamp 0
transform 1 0 5070 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1028_
timestamp 0
transform -1 0 2090 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1029_
timestamp 0
transform 1 0 3510 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1030_
timestamp 0
transform 1 0 2330 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1031_
timestamp 0
transform 1 0 2670 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1032_
timestamp 0
transform -1 0 1850 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1033_
timestamp 0
transform -1 0 2210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1034_
timestamp 0
transform -1 0 1510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1035_
timestamp 0
transform 1 0 1770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1036_
timestamp 0
transform 1 0 2790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1037_
timestamp 0
transform 1 0 2010 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1038_
timestamp 0
transform -1 0 2250 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1039_
timestamp 0
transform 1 0 1930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1040_
timestamp 0
transform 1 0 2370 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1041_
timestamp 0
transform 1 0 4450 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1042_
timestamp 0
transform 1 0 3790 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1043_
timestamp 0
transform 1 0 3970 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1044_
timestamp 0
transform 1 0 3350 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1045_
timestamp 0
transform 1 0 2530 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1046_
timestamp 0
transform 1 0 2470 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1047_
timestamp 0
transform 1 0 3650 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1048_
timestamp 0
transform -1 0 3350 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1049_
timestamp 0
transform 1 0 2690 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1050_
timestamp 0
transform 1 0 3630 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1051_
timestamp 0
transform 1 0 3010 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1052_
timestamp 0
transform 1 0 2850 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1053_
timestamp 0
transform 1 0 3190 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1054_
timestamp 0
transform 1 0 4530 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1055_
timestamp 0
transform 1 0 5810 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1056_
timestamp 0
transform -1 0 5870 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1057_
timestamp 0
transform 1 0 3790 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1058_
timestamp 0
transform 1 0 3830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1059_
timestamp 0
transform -1 0 4450 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1060_
timestamp 0
transform -1 0 4090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1061_
timestamp 0
transform -1 0 3730 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1062_
timestamp 0
transform 1 0 4250 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1063_
timestamp 0
transform 1 0 3670 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1064_
timestamp 0
transform 1 0 3950 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1065_
timestamp 0
transform 1 0 4290 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1066_
timestamp 0
transform 1 0 3550 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1067_
timestamp 0
transform 1 0 4130 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1068_
timestamp 0
transform -1 0 4910 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1069_
timestamp 0
transform 1 0 5550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1070_
timestamp 0
transform 1 0 5730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1071_
timestamp 0
transform -1 0 5350 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1072_
timestamp 0
transform -1 0 5230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1073_
timestamp 0
transform -1 0 5810 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1074_
timestamp 0
transform -1 0 5610 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1075_
timestamp 0
transform -1 0 5550 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1076_
timestamp 0
transform -1 0 5470 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1077_
timestamp 0
transform -1 0 5350 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1078_
timestamp 0
transform 1 0 5730 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1079_
timestamp 0
transform 1 0 5650 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1080_
timestamp 0
transform -1 0 5670 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1081_
timestamp 0
transform -1 0 5510 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1082_
timestamp 0
transform 1 0 5710 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1083_
timestamp 0
transform 1 0 5810 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1084_
timestamp 0
transform 1 0 5490 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1085_
timestamp 0
transform -1 0 5850 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1086_
timestamp 0
transform 1 0 5050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1087_
timestamp 0
transform 1 0 5210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1088_
timestamp 0
transform -1 0 5870 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1089_
timestamp 0
transform 1 0 5550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1090_
timestamp 0
transform -1 0 5550 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1091_
timestamp 0
transform -1 0 5390 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1092_
timestamp 0
transform 1 0 5710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1093_
timestamp 0
transform 1 0 5550 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1094_
timestamp 0
transform 1 0 5690 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1095_
timestamp 0
transform 1 0 5370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1096_
timestamp 0
transform -1 0 5750 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1097_
timestamp 0
transform 1 0 4850 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1098_
timestamp 0
transform -1 0 4410 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1099_
timestamp 0
transform 1 0 5770 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1100_
timestamp 0
transform 1 0 5390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1101_
timestamp 0
transform -1 0 5570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1102_
timestamp 0
transform -1 0 5250 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1103_
timestamp 0
transform -1 0 5150 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1104_
timestamp 0
transform 1 0 4970 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1105_
timestamp 0
transform -1 0 5630 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1106_
timestamp 0
transform 1 0 5030 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1107_
timestamp 0
transform -1 0 5150 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1108_
timestamp 0
transform -1 0 4310 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1109_
timestamp 0
transform -1 0 5310 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1110_
timestamp 0
transform -1 0 4970 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1111_
timestamp 0
transform -1 0 4810 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1112_
timestamp 0
transform -1 0 4150 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1113_
timestamp 0
transform 1 0 4670 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1114_
timestamp 0
transform 1 0 4510 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1115_
timestamp 0
transform -1 0 4630 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1116_
timestamp 0
transform 1 0 4450 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1117_
timestamp 0
transform -1 0 4510 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1118_
timestamp 0
transform 1 0 4090 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1119_
timestamp 0
transform -1 0 3590 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1120_
timestamp 0
transform -1 0 3970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1121_
timestamp 0
transform -1 0 3970 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1122_
timestamp 0
transform -1 0 3790 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1123_
timestamp 0
transform -1 0 4810 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1124_
timestamp 0
transform 1 0 4610 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1125_
timestamp 0
transform 1 0 3930 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1126_
timestamp 0
transform 1 0 4290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1127_
timestamp 0
transform -1 0 5230 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1128_
timestamp 0
transform 1 0 4690 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1129_
timestamp 0
transform 1 0 2950 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1130_
timestamp 0
transform 1 0 2170 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1131_
timestamp 0
transform 1 0 2490 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1132_
timestamp 0
transform 1 0 2190 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1133_
timestamp 0
transform 1 0 2010 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1134_
timestamp 0
transform 1 0 2350 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1135_
timestamp 0
transform -1 0 1330 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1136_
timestamp 0
transform -1 0 1710 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1137_
timestamp 0
transform 1 0 1690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1138_
timestamp 0
transform 1 0 2770 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1139_
timestamp 0
transform -1 0 2330 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1140_
timestamp 0
transform 1 0 1850 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1141_
timestamp 0
transform 1 0 2630 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1142_
timestamp 0
transform -1 0 4290 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1143_
timestamp 0
transform -1 0 4090 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1144_
timestamp 0
transform 1 0 3110 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1145_
timestamp 0
transform 1 0 2470 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1146_
timestamp 0
transform 1 0 2610 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1147_
timestamp 0
transform -1 0 4410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1148_
timestamp 0
transform 1 0 3430 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1149_
timestamp 0
transform 1 0 3490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1150_
timestamp 0
transform 1 0 2790 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1151_
timestamp 0
transform -1 0 2970 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1152_
timestamp 0
transform 1 0 3130 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1153_
timestamp 0
transform 1 0 3110 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1154_
timestamp 0
transform 1 0 2950 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1155_
timestamp 0
transform 1 0 3270 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1156_
timestamp 0
transform -1 0 3670 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1157_
timestamp 0
transform -1 0 5330 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1158_
timestamp 0
transform -1 0 5170 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1159_
timestamp 0
transform -1 0 3950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1160_
timestamp 0
transform -1 0 3910 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1161_
timestamp 0
transform 1 0 2890 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1162_
timestamp 0
transform -1 0 3610 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1163_
timestamp 0
transform -1 0 1630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1164_
timestamp 0
transform 1 0 3230 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1165_
timestamp 0
transform 1 0 3730 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1166_
timestamp 0
transform 1 0 4170 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1167_
timestamp 0
transform 1 0 4330 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1168_
timestamp 0
transform 1 0 4490 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1169_
timestamp 0
transform 1 0 4650 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1170_
timestamp 0
transform 1 0 4810 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1171_
timestamp 0
transform -1 0 5650 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1172_
timestamp 0
transform -1 0 5490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1173_
timestamp 0
transform -1 0 5810 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1174_
timestamp 0
transform 1 0 5810 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1175_
timestamp 0
transform 1 0 5610 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1176_
timestamp 0
transform -1 0 5470 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1177_
timestamp 0
transform -1 0 5530 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1178_
timestamp 0
transform -1 0 5310 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1179_
timestamp 0
transform -1 0 4990 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1180_
timestamp 0
transform 1 0 5730 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1181_
timestamp 0
transform 1 0 5790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1182_
timestamp 0
transform -1 0 5790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1183_
timestamp 0
transform -1 0 5470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1184_
timestamp 0
transform 1 0 4910 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1185_
timestamp 0
transform 1 0 5010 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1186_
timestamp 0
transform -1 0 5050 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1187_
timestamp 0
transform -1 0 4890 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1188_
timestamp 0
transform 1 0 4750 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1189_
timestamp 0
transform 1 0 5110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1190_
timestamp 0
transform 1 0 5130 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1191_
timestamp 0
transform -1 0 4970 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1192_
timestamp 0
transform -1 0 4910 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1193_
timestamp 0
transform 1 0 3790 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1194_
timestamp 0
transform 1 0 5170 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1195_
timestamp 0
transform -1 0 4870 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1196_
timestamp 0
transform -1 0 4650 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1197_
timestamp 0
transform 1 0 4570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1198_
timestamp 0
transform -1 0 4770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1199_
timestamp 0
transform -1 0 4610 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1200_
timestamp 0
transform -1 0 4810 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1201_
timestamp 0
transform 1 0 5050 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1202_
timestamp 0
transform -1 0 4570 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1203_
timestamp 0
transform -1 0 4230 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1204_
timestamp 0
transform -1 0 4730 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1205_
timestamp 0
transform -1 0 4430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1206_
timestamp 0
transform -1 0 3990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1207_
timestamp 0
transform 1 0 3850 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1208_
timestamp 0
transform -1 0 5090 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1209_
timestamp 0
transform 1 0 4910 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1210_
timestamp 0
transform -1 0 4150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1211_
timestamp 0
transform -1 0 4410 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1212_
timestamp 0
transform -1 0 4050 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1213_
timestamp 0
transform 1 0 4050 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1214_
timestamp 0
transform -1 0 3210 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1215_
timestamp 0
transform 1 0 3750 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1216_
timestamp 0
transform 1 0 3870 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1217_
timestamp 0
transform -1 0 4750 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1218_
timestamp 0
transform 1 0 4470 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1219_
timestamp 0
transform 1 0 3270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1220_
timestamp 0
transform 1 0 5110 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1221_
timestamp 0
transform 1 0 5270 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1222_
timestamp 0
transform 1 0 2010 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1223_
timestamp 0
transform 1 0 2870 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1224_
timestamp 0
transform -1 0 2310 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1225_
timestamp 0
transform 1 0 2050 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1226_
timestamp 0
transform 1 0 1610 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1227_
timestamp 0
transform -1 0 1790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1228_
timestamp 0
transform 1 0 2610 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1229_
timestamp 0
transform 1 0 2770 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1230_
timestamp 0
transform 1 0 2230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1231_
timestamp 0
transform -1 0 2450 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1232_
timestamp 0
transform -1 0 2610 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1233_
timestamp 0
transform 1 0 2930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1234_
timestamp 0
transform 1 0 4010 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1235_
timestamp 0
transform -1 0 3770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1236_
timestamp 0
transform 1 0 3590 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1237_
timestamp 0
transform 1 0 2770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1238_
timestamp 0
transform 1 0 2370 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1239_
timestamp 0
transform -1 0 3410 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1240_
timestamp 0
transform 1 0 3090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1241_
timestamp 0
transform 1 0 3070 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1242_
timestamp 0
transform 1 0 3030 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1243_
timestamp 0
transform -1 0 3450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1244_
timestamp 0
transform 1 0 3250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1245_
timestamp 0
transform 1 0 3390 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1246_
timestamp 0
transform 1 0 4890 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1247_
timestamp 0
transform -1 0 5610 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1248_
timestamp 0
transform 1 0 5430 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1249_
timestamp 0
transform -1 0 3570 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1250_
timestamp 0
transform 1 0 3110 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1251_
timestamp 0
transform -1 0 2790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1252_
timestamp 0
transform -1 0 2990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1253_
timestamp 0
transform -1 0 1050 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1254_
timestamp 0
transform 1 0 2930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1255_
timestamp 0
transform 1 0 3230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1256_
timestamp 0
transform 1 0 3110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1257_
timestamp 0
transform 1 0 3270 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1258_
timestamp 0
transform 1 0 3490 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1259_
timestamp 0
transform -1 0 5730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1260_
timestamp 0
transform -1 0 5290 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1261_
timestamp 0
transform -1 0 5450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1262_
timestamp 0
transform 1 0 5830 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1263_
timestamp 0
transform -1 0 5710 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1264_
timestamp 0
transform -1 0 5610 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1265_
timestamp 0
transform -1 0 5630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1266_
timestamp 0
transform 1 0 5290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1267_
timestamp 0
transform -1 0 5770 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1268_
timestamp 0
transform 1 0 5750 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1269_
timestamp 0
transform -1 0 5470 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1270_
timestamp 0
transform 1 0 5050 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1271_
timestamp 0
transform 1 0 5670 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1272_
timestamp 0
transform -1 0 5430 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1273_
timestamp 0
transform -1 0 5270 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1274_
timestamp 0
transform -1 0 4970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1275_
timestamp 0
transform -1 0 4750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1276_
timestamp 0
transform 1 0 4550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1277_
timestamp 0
transform 1 0 5610 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1278_
timestamp 0
transform -1 0 5550 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1279_
timestamp 0
transform -1 0 5390 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1280_
timestamp 0
transform 1 0 5190 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1281_
timestamp 0
transform -1 0 4770 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1282_
timestamp 0
transform -1 0 4610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1283_
timestamp 0
transform 1 0 4630 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1284_
timestamp 0
transform 1 0 5270 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1285_
timestamp 0
transform -1 0 4790 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1286_
timestamp 0
transform -1 0 4950 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1287_
timestamp 0
transform -1 0 4450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1288_
timestamp 0
transform 1 0 4190 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1289_
timestamp 0
transform 1 0 4310 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1290_
timestamp 0
transform -1 0 5110 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1291_
timestamp 0
transform -1 0 4490 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1292_
timestamp 0
transform -1 0 4330 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1293_
timestamp 0
transform 1 0 4150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1294_
timestamp 0
transform -1 0 3570 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1295_
timestamp 0
transform -1 0 4310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1296_
timestamp 0
transform 1 0 3990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1297_
timestamp 0
transform -1 0 3730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1298_
timestamp 0
transform 1 0 3830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1299_
timestamp 0
transform -1 0 4370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1300_
timestamp 0
transform 1 0 4190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1301_
timestamp 0
transform 1 0 3850 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1302_
timestamp 0
transform 1 0 4850 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1303_
timestamp 0
transform -1 0 5110 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1304_
timestamp 0
transform 1 0 2590 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1305_
timestamp 0
transform -1 0 1930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1306_
timestamp 0
transform 1 0 1530 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1307_
timestamp 0
transform -1 0 1690 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1308_
timestamp 0
transform -1 0 1690 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1309_
timestamp 0
transform 1 0 1970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1310_
timestamp 0
transform 1 0 2130 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1311_
timestamp 0
transform 1 0 1850 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1312_
timestamp 0
transform -1 0 2170 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1313_
timestamp 0
transform 1 0 1990 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1314_
timestamp 0
transform 1 0 2430 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1315_
timestamp 0
transform 1 0 2670 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1316_
timestamp 0
transform 1 0 2810 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1317_
timestamp 0
transform 1 0 2670 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1318_
timestamp 0
transform 1 0 2250 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1319_
timestamp 0
transform -1 0 1750 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1320_
timestamp 0
transform -1 0 3350 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1321_
timestamp 0
transform -1 0 3190 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1322_
timestamp 0
transform 1 0 2330 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1323_
timestamp 0
transform 1 0 2830 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1324_
timestamp 0
transform 1 0 2650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1325_
timestamp 0
transform 1 0 2490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1326_
timestamp 0
transform 1 0 2510 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1327_
timestamp 0
transform 1 0 2990 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1328_
timestamp 0
transform -1 0 3570 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1329_
timestamp 0
transform -1 0 5590 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1330_
timestamp 0
transform -1 0 5410 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1331_
timestamp 0
transform 1 0 2310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1332_
timestamp 0
transform 1 0 2150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1333_
timestamp 0
transform 1 0 2510 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1334_
timestamp 0
transform -1 0 3090 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1335_
timestamp 0
transform -1 0 2530 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1336_
timestamp 0
transform -1 0 2350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1337_
timestamp 0
transform 1 0 2350 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1338_
timestamp 0
transform 1 0 3210 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1339_
timestamp 0
transform -1 0 4130 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1340_
timestamp 0
transform 1 0 4010 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1341_
timestamp 0
transform 1 0 3370 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1342_
timestamp 0
transform 1 0 4310 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1343_
timestamp 0
transform 1 0 3350 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1344_
timestamp 0
transform -1 0 5250 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1345_
timestamp 0
transform 1 0 4450 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1346_
timestamp 0
transform -1 0 4170 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1347_
timestamp 0
transform 1 0 4930 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1348_
timestamp 0
transform -1 0 5310 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1349_
timestamp 0
transform 1 0 3690 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1350_
timestamp 0
transform -1 0 3870 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1351_
timestamp 0
transform 1 0 4610 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1352_
timestamp 0
transform -1 0 5150 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1353_
timestamp 0
transform 1 0 4290 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1354_
timestamp 0
transform -1 0 4790 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1355_
timestamp 0
transform -1 0 4570 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1356_
timestamp 0
transform -1 0 4410 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1357_
timestamp 0
transform -1 0 5130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1358_
timestamp 0
transform -1 0 4630 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1359_
timestamp 0
transform 1 0 4670 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1360_
timestamp 0
transform -1 0 4990 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1361_
timestamp 0
transform -1 0 4750 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1362_
timestamp 0
transform 1 0 4250 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1363_
timestamp 0
transform 1 0 3990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1364_
timestamp 0
transform -1 0 3890 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1365_
timestamp 0
transform -1 0 4390 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1366_
timestamp 0
transform -1 0 4230 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1367_
timestamp 0
transform 1 0 2790 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1368_
timestamp 0
transform 1 0 3270 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1369_
timestamp 0
transform 1 0 3970 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1370_
timestamp 0
transform -1 0 3830 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1371_
timestamp 0
transform 1 0 2150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1372_
timestamp 0
transform -1 0 1570 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1373_
timestamp 0
transform -1 0 1470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1374_
timestamp 0
transform 1 0 1110 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1375_
timestamp 0
transform 1 0 1390 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1376_
timestamp 0
transform 1 0 1230 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1377_
timestamp 0
transform -1 0 1190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1378_
timestamp 0
transform -1 0 1830 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1379_
timestamp 0
transform 1 0 1410 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1380_
timestamp 0
transform 1 0 1270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1381_
timestamp 0
transform 1 0 1330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1382_
timestamp 0
transform 1 0 1470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1383_
timestamp 0
transform 1 0 1710 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1384_
timestamp 0
transform -1 0 2070 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1385_
timestamp 0
transform -1 0 1730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1386_
timestamp 0
transform -1 0 1570 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1387_
timestamp 0
transform -1 0 1130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1388_
timestamp 0
transform 1 0 1550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1389_
timestamp 0
transform -1 0 1870 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1390_
timestamp 0
transform -1 0 2230 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1391_
timestamp 0
transform 1 0 1870 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1392_
timestamp 0
transform 1 0 1390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1393_
timestamp 0
transform -1 0 1850 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1394_
timestamp 0
transform 1 0 2570 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1395_
timestamp 0
transform 1 0 2930 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1396_
timestamp 0
transform -1 0 2770 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1397_
timestamp 0
transform -1 0 2630 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1398_
timestamp 0
transform -1 0 2390 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1399_
timestamp 0
transform 1 0 2190 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1400_
timestamp 0
transform 1 0 1990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1401_
timestamp 0
transform 1 0 2010 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1402_
timestamp 0
transform 1 0 2490 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1403_
timestamp 0
transform -1 0 2950 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1404_
timestamp 0
transform -1 0 3250 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1405_
timestamp 0
transform -1 0 3690 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1406_
timestamp 0
transform -1 0 3530 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1407_
timestamp 0
transform 1 0 2970 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1408_
timestamp 0
transform 1 0 3610 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1409_
timestamp 0
transform 1 0 2810 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1410_
timestamp 0
transform -1 0 3090 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1411_
timestamp 0
transform 1 0 3290 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1412_
timestamp 0
transform 1 0 3770 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1413_
timestamp 0
transform 1 0 4450 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1414_
timestamp 0
transform -1 0 4510 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1415_
timestamp 0
transform -1 0 3150 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1416_
timestamp 0
transform 1 0 3450 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1417_
timestamp 0
transform -1 0 3950 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1418_
timestamp 0
transform 1 0 3590 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1419_
timestamp 0
transform 1 0 3550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1420_
timestamp 0
transform 1 0 4050 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1421_
timestamp 0
transform 1 0 3690 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1422_
timestamp 0
transform -1 0 3410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1423_
timestamp 0
transform -1 0 4110 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1424_
timestamp 0
transform -1 0 3430 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1425_
timestamp 0
transform 1 0 3730 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1426_
timestamp 0
transform 1 0 2930 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1427_
timestamp 0
transform -1 0 2650 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1428_
timestamp 0
transform 1 0 1690 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1429_
timestamp 0
transform -1 0 1190 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1430_
timestamp 0
transform -1 0 2470 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1431_
timestamp 0
transform 1 0 1390 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1432_
timestamp 0
transform 1 0 650 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1433_
timestamp 0
transform -1 0 1290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1434_
timestamp 0
transform 1 0 1110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1435_
timestamp 0
transform 1 0 1070 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1436_
timestamp 0
transform 1 0 970 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1437_
timestamp 0
transform 1 0 930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1438_
timestamp 0
transform -1 0 1090 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1439_
timestamp 0
transform -1 0 790 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1440_
timestamp 0
transform 1 0 1230 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1441_
timestamp 0
transform -1 0 490 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1442_
timestamp 0
transform 1 0 30 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1443_
timestamp 0
transform -1 0 2450 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1444_
timestamp 0
transform -1 0 190 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1445_
timestamp 0
transform 1 0 470 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1446_
timestamp 0
transform -1 0 350 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1447_
timestamp 0
transform -1 0 50 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1448_
timestamp 0
transform 1 0 170 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1449_
timestamp 0
transform -1 0 630 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1450_
timestamp 0
transform -1 0 630 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1451_
timestamp 0
transform -1 0 910 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1452_
timestamp 0
transform -1 0 910 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1453_
timestamp 0
transform -1 0 770 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1454_
timestamp 0
transform 1 0 1010 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1455_
timestamp 0
transform 1 0 1050 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1456_
timestamp 0
transform 1 0 1210 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1457_
timestamp 0
transform -1 0 2070 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1458_
timestamp 0
transform -1 0 2670 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1459_
timestamp 0
transform -1 0 2790 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1460_
timestamp 0
transform -1 0 1890 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1461_
timestamp 0
transform 1 0 1790 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1462_
timestamp 0
transform -1 0 1950 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1463_
timestamp 0
transform 1 0 1750 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1464_
timestamp 0
transform -1 0 1610 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1465_
timestamp 0
transform 1 0 1290 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1466_
timestamp 0
transform 1 0 790 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1467_
timestamp 0
transform -1 0 590 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1468_
timestamp 0
transform 1 0 930 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1469_
timestamp 0
transform 1 0 630 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1470_
timestamp 0
transform -1 0 1250 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1471_
timestamp 0
transform 1 0 770 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1472_
timestamp 0
transform -1 0 50 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1473_
timestamp 0
transform -1 0 50 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1474_
timestamp 0
transform -1 0 50 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1475_
timestamp 0
transform 1 0 530 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1476_
timestamp 0
transform 1 0 210 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1477_
timestamp 0
transform 1 0 650 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1478_
timestamp 0
transform 1 0 310 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1479_
timestamp 0
transform 1 0 230 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1480_
timestamp 0
transform -1 0 390 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1481_
timestamp 0
transform 1 0 370 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1482_
timestamp 0
transform -1 0 830 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1483_
timestamp 0
transform -1 0 1410 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1484_
timestamp 0
transform -1 0 1490 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1485_
timestamp 0
transform -1 0 1330 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1486_
timestamp 0
transform -1 0 1650 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1487_
timestamp 0
transform -1 0 1430 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1488_
timestamp 0
transform 1 0 1450 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1489_
timestamp 0
transform 1 0 1230 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1490_
timestamp 0
transform 1 0 510 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1491_
timestamp 0
transform -1 0 810 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1492_
timestamp 0
transform 1 0 630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1493_
timestamp 0
transform -1 0 510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1494_
timestamp 0
transform 1 0 210 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1495_
timestamp 0
transform 1 0 330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1496_
timestamp 0
transform 1 0 730 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1497_
timestamp 0
transform 1 0 230 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1498_
timestamp 0
transform 1 0 30 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1499_
timestamp 0
transform -1 0 250 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1500_
timestamp 0
transform 1 0 870 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1501_
timestamp 0
transform -1 0 970 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1502_
timestamp 0
transform -1 0 950 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1503_
timestamp 0
transform -1 0 930 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1504_
timestamp 0
transform 1 0 630 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1505_
timestamp 0
transform -1 0 770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1506_
timestamp 0
transform -1 0 590 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1507_
timestamp 0
transform 1 0 30 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1508_
timestamp 0
transform -1 0 50 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1509_
timestamp 0
transform -1 0 390 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1510_
timestamp 0
transform 1 0 290 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1511_
timestamp 0
transform 1 0 3070 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1512_
timestamp 0
transform -1 0 1550 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1513_
timestamp 0
transform -1 0 1170 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1514_
timestamp 0
transform -1 0 1090 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1515_
timestamp 0
transform -1 0 190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1516_
timestamp 0
transform -1 0 590 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1517_
timestamp 0
transform -1 0 450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1518_
timestamp 0
transform 1 0 1290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1519_
timestamp 0
transform 1 0 2190 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1560_
timestamp 0
transform -1 0 50 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1561_
timestamp 0
transform -1 0 190 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1562_
timestamp 0
transform -1 0 50 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1563_
timestamp 0
transform -1 0 50 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1564_
timestamp 0
transform -1 0 330 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1565_
timestamp 0
transform 1 0 3870 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1566_
timestamp 0
transform -1 0 990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1567_
timestamp 0
transform -1 0 50 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1568_
timestamp 0
transform -1 0 50 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1569_
timestamp 0
transform -1 0 50 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1570_
timestamp 0
transform -1 0 3690 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1571_
timestamp 0
transform 1 0 5090 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1572_
timestamp 0
transform -1 0 2330 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1573_
timestamp 0
transform 1 0 2170 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1574_
timestamp 0
transform -1 0 50 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1575_
timestamp 0
transform -1 0 210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1576_
timestamp 0
transform -1 0 50 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1577_
timestamp 0
transform -1 0 350 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1578_
timestamp 0
transform 1 0 1590 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1579_
timestamp 0
transform 1 0 2210 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1580_
timestamp 0
transform -1 0 2730 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1581_
timestamp 0
transform -1 0 3070 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1582_
timestamp 0
transform -1 0 50 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1583_
timestamp 0
transform -1 0 3250 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert6
timestamp 0
transform 1 0 5070 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert7
timestamp 0
transform -1 0 3110 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert8
timestamp 0
transform -1 0 3110 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert9
timestamp 0
transform -1 0 5830 0 -1 270
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert10
timestamp 0
transform 1 0 1630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert11
timestamp 0
transform 1 0 1750 0 1 4430
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert12
timestamp 0
transform 1 0 1510 0 1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert13
timestamp 0
transform -1 0 50 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert14
timestamp 0
transform -1 0 2750 0 1 2350
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert15
timestamp 0
transform -1 0 4050 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert16
timestamp 0
transform 1 0 4250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert17
timestamp 0
transform 1 0 4170 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert0
timestamp 0
transform 1 0 1430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert1
timestamp 0
transform -1 0 1270 0 1 3390
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert2
timestamp 0
transform -1 0 730 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert3
timestamp 0
transform -1 0 1070 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert4
timestamp 0
transform -1 0 1050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert5
timestamp 0
transform 1 0 3010 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__756_
timestamp 0
transform 1 0 1310 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__757_
timestamp 0
transform 1 0 1670 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__758_
timestamp 0
transform 1 0 1430 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__759_
timestamp 0
transform 1 0 570 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__760_
timestamp 0
transform 1 0 710 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__761_
timestamp 0
transform 1 0 430 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__762_
timestamp 0
transform 1 0 430 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__763_
timestamp 0
transform -1 0 1170 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__764_
timestamp 0
transform 1 0 950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__765_
timestamp 0
transform -1 0 450 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__766_
timestamp 0
transform 1 0 610 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__767_
timestamp 0
transform 1 0 770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__768_
timestamp 0
transform -1 0 910 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__769_
timestamp 0
transform 1 0 690 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__770_
timestamp 0
transform 1 0 830 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__771_
timestamp 0
transform 1 0 990 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__772_
timestamp 0
transform -1 0 1170 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__773_
timestamp 0
transform -1 0 850 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__774_
timestamp 0
transform 1 0 670 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__775_
timestamp 0
transform -1 0 3130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__776_
timestamp 0
transform -1 0 1470 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__777_
timestamp 0
transform -1 0 1010 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__778_
timestamp 0
transform 1 0 370 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__779_
timestamp 0
transform 1 0 530 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__780_
timestamp 0
transform 1 0 50 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__781_
timestamp 0
transform 1 0 50 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__782_
timestamp 0
transform 1 0 490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__783_
timestamp 0
transform 1 0 610 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__784_
timestamp 0
transform 1 0 210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__785_
timestamp 0
transform 1 0 330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__786_
timestamp 0
transform -1 0 810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__787_
timestamp 0
transform 1 0 950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__788_
timestamp 0
transform 1 0 1590 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__789_
timestamp 0
transform -1 0 1190 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__790_
timestamp 0
transform -1 0 1350 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__791_
timestamp 0
transform 1 0 1290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__792_
timestamp 0
transform -1 0 1430 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__793_
timestamp 0
transform -1 0 1030 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__794_
timestamp 0
transform 1 0 950 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__795_
timestamp 0
transform -1 0 870 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__796_
timestamp 0
transform 1 0 810 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__797_
timestamp 0
transform 1 0 1110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__798_
timestamp 0
transform -1 0 910 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__799_
timestamp 0
transform -1 0 3470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__800_
timestamp 0
transform 1 0 2230 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__801_
timestamp 0
transform 1 0 2310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__802_
timestamp 0
transform 1 0 1890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__803_
timestamp 0
transform -1 0 1590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__804_
timestamp 0
transform -1 0 1290 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__805_
timestamp 0
transform -1 0 230 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__806_
timestamp 0
transform -1 0 770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__807_
timestamp 0
transform 1 0 870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__808_
timestamp 0
transform 1 0 470 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__809_
timestamp 0
transform 1 0 50 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__810_
timestamp 0
transform -1 0 230 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__811_
timestamp 0
transform 1 0 170 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__812_
timestamp 0
transform -1 0 730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__813_
timestamp 0
transform -1 0 350 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__814_
timestamp 0
transform -1 0 70 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__815_
timestamp 0
transform 1 0 370 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__816_
timestamp 0
transform 1 0 430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__817_
timestamp 0
transform -1 0 70 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__818_
timestamp 0
transform -1 0 230 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__819_
timestamp 0
transform -1 0 570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__820_
timestamp 0
transform -1 0 190 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__821_
timestamp 0
transform 1 0 910 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__822_
timestamp 0
transform 1 0 2030 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__823_
timestamp 0
transform -1 0 1750 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__824_
timestamp 0
transform 1 0 650 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__825_
timestamp 0
transform 1 0 590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__826_
timestamp 0
transform 1 0 950 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__827_
timestamp 0
transform -1 0 1270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__828_
timestamp 0
transform 1 0 750 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__829_
timestamp 0
transform -1 0 1090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__830_
timestamp 0
transform 1 0 350 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__831_
timestamp 0
transform -1 0 1490 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__832_
timestamp 0
transform 1 0 590 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__833_
timestamp 0
transform -1 0 1170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__834_
timestamp 0
transform 1 0 2090 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__835_
timestamp 0
transform 1 0 1110 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__836_
timestamp 0
transform 1 0 630 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__837_
timestamp 0
transform 1 0 990 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__838_
timestamp 0
transform -1 0 2410 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__839_
timestamp 0
transform -1 0 2590 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__840_
timestamp 0
transform -1 0 1770 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__841_
timestamp 0
transform -1 0 2570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__842_
timestamp 0
transform 1 0 2090 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__843_
timestamp 0
transform -1 0 1830 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__844_
timestamp 0
transform 1 0 1870 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__845_
timestamp 0
transform -1 0 1950 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__846_
timestamp 0
transform -1 0 1610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__847_
timestamp 0
transform -1 0 990 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__848_
timestamp 0
transform 1 0 790 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__849_
timestamp 0
transform -1 0 2010 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__850_
timestamp 0
transform -1 0 1670 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__851_
timestamp 0
transform -1 0 1350 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__852_
timestamp 0
transform 1 0 2350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__853_
timestamp 0
transform 1 0 2790 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__854_
timestamp 0
transform 1 0 2050 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__855_
timestamp 0
transform -1 0 1610 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__856_
timestamp 0
transform 1 0 1590 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__857_
timestamp 0
transform -1 0 1930 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__858_
timestamp 0
transform -1 0 2270 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__859_
timestamp 0
transform 1 0 2670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__860_
timestamp 0
transform -1 0 2530 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__861_
timestamp 0
transform 1 0 1710 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__862_
timestamp 0
transform -1 0 1770 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__863_
timestamp 0
transform 1 0 1890 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__864_
timestamp 0
transform -1 0 1030 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__865_
timestamp 0
transform 1 0 1490 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__866_
timestamp 0
transform -1 0 1770 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__867_
timestamp 0
transform 1 0 2090 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__868_
timestamp 0
transform 1 0 2190 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__869_
timestamp 0
transform 1 0 2170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__870_
timestamp 0
transform 1 0 1570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__871_
timestamp 0
transform 1 0 1430 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__872_
timestamp 0
transform -1 0 810 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__873_
timestamp 0
transform 1 0 1730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__874_
timestamp 0
transform 1 0 1170 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__875_
timestamp 0
transform 1 0 2050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__876_
timestamp 0
transform -1 0 2250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__877_
timestamp 0
transform 1 0 1390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__878_
timestamp 0
transform 1 0 1610 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__879_
timestamp 0
transform 1 0 1890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__880_
timestamp 0
transform -1 0 1670 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__881_
timestamp 0
transform 1 0 2410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__882_
timestamp 0
transform 1 0 1830 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__883_
timestamp 0
transform 1 0 1990 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__884_
timestamp 0
transform -1 0 1930 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__885_
timestamp 0
transform 1 0 1290 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__886_
timestamp 0
transform 1 0 1790 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__887_
timestamp 0
transform -1 0 2390 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__888_
timestamp 0
transform 1 0 2490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__889_
timestamp 0
transform 1 0 2710 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__890_
timestamp 0
transform 1 0 1490 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__891_
timestamp 0
transform 1 0 2670 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__892_
timestamp 0
transform 1 0 2810 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__893_
timestamp 0
transform 1 0 3230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__894_
timestamp 0
transform 1 0 2950 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__895_
timestamp 0
transform 1 0 3390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__896_
timestamp 0
transform 1 0 2510 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__897_
timestamp 0
transform 1 0 2930 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__898_
timestamp 0
transform 1 0 2650 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__899_
timestamp 0
transform -1 0 3170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__900_
timestamp 0
transform -1 0 3010 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__901_
timestamp 0
transform 1 0 2830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__902_
timestamp 0
transform 1 0 3590 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__903_
timestamp 0
transform 1 0 2630 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__904_
timestamp 0
transform -1 0 4550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__905_
timestamp 0
transform -1 0 4850 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__906_
timestamp 0
transform -1 0 5310 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__907_
timestamp 0
transform -1 0 4550 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__908_
timestamp 0
transform -1 0 4970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__909_
timestamp 0
transform 1 0 4670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__910_
timestamp 0
transform -1 0 4690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__911_
timestamp 0
transform -1 0 4830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__912_
timestamp 0
transform 1 0 4350 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__913_
timestamp 0
transform -1 0 4810 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__914_
timestamp 0
transform 1 0 4370 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__915_
timestamp 0
transform 1 0 4350 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__916_
timestamp 0
transform -1 0 4650 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__917_
timestamp 0
transform -1 0 4970 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__918_
timestamp 0
transform 1 0 4190 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__919_
timestamp 0
transform -1 0 3770 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__920_
timestamp 0
transform 1 0 3590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__921_
timestamp 0
transform -1 0 4030 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__922_
timestamp 0
transform -1 0 4490 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__923_
timestamp 0
transform -1 0 3870 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__924_
timestamp 0
transform 1 0 2950 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__925_
timestamp 0
transform 1 0 1330 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__926_
timestamp 0
transform -1 0 3690 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__927_
timestamp 0
transform 1 0 3730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__928_
timestamp 0
transform 1 0 3430 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__929_
timestamp 0
transform -1 0 3070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__930_
timestamp 0
transform 1 0 2370 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__931_
timestamp 0
transform -1 0 2530 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__932_
timestamp 0
transform -1 0 3290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__933_
timestamp 0
transform -1 0 2810 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__934_
timestamp 0
transform 1 0 2630 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__935_
timestamp 0
transform -1 0 2730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__936_
timestamp 0
transform 1 0 2390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__937_
timestamp 0
transform 1 0 2470 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__938_
timestamp 0
transform -1 0 2910 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__939_
timestamp 0
transform -1 0 2570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__940_
timestamp 0
transform 1 0 2290 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__941_
timestamp 0
transform -1 0 2130 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__942_
timestamp 0
transform 1 0 2990 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__943_
timestamp 0
transform 1 0 2850 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__944_
timestamp 0
transform -1 0 2830 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__945_
timestamp 0
transform 1 0 2690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__946_
timestamp 0
transform -1 0 2950 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__947_
timestamp 0
transform 1 0 3110 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__948_
timestamp 0
transform 1 0 3210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__949_
timestamp 0
transform 1 0 1330 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__950_
timestamp 0
transform 1 0 1410 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__951_
timestamp 0
transform 1 0 1930 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__952_
timestamp 0
transform 1 0 3290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__953_
timestamp 0
transform 1 0 4870 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__954_
timestamp 0
transform -1 0 4230 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__955_
timestamp 0
transform 1 0 3910 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__956_
timestamp 0
transform 1 0 3090 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__957_
timestamp 0
transform 1 0 3230 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__958_
timestamp 0
transform 1 0 3330 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__959_
timestamp 0
transform -1 0 4170 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__960_
timestamp 0
transform 1 0 2090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__961_
timestamp 0
transform 1 0 3450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__962_
timestamp 0
transform 1 0 3510 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__963_
timestamp 0
transform 1 0 3970 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__964_
timestamp 0
transform 1 0 3670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__965_
timestamp 0
transform 1 0 3510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__966_
timestamp 0
transform 1 0 3830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__967_
timestamp 0
transform 1 0 5250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__968_
timestamp 0
transform -1 0 5150 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__969_
timestamp 0
transform 1 0 4950 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__970_
timestamp 0
transform 1 0 5110 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__971_
timestamp 0
transform -1 0 5250 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__972_
timestamp 0
transform -1 0 5390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__973_
timestamp 0
transform -1 0 5930 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__974_
timestamp 0
transform -1 0 5470 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__975_
timestamp 0
transform -1 0 5270 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__976_
timestamp 0
transform -1 0 5690 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__977_
timestamp 0
transform 1 0 5610 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__978_
timestamp 0
transform -1 0 5790 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__979_
timestamp 0
transform -1 0 5610 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__980_
timestamp 0
transform -1 0 5450 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__981_
timestamp 0
transform -1 0 5910 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__982_
timestamp 0
transform 1 0 5750 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__983_
timestamp 0
transform 1 0 5410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__984_
timestamp 0
transform -1 0 5750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__985_
timestamp 0
transform -1 0 5270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__986_
timestamp 0
transform -1 0 5670 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__987_
timestamp 0
transform 1 0 5570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__988_
timestamp 0
transform 1 0 5470 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__989_
timestamp 0
transform -1 0 5170 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__990_
timestamp 0
transform 1 0 4070 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__991_
timestamp 0
transform 1 0 4190 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__992_
timestamp 0
transform -1 0 5490 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__993_
timestamp 0
transform -1 0 5430 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__994_
timestamp 0
transform -1 0 5430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__995_
timestamp 0
transform -1 0 4910 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__996_
timestamp 0
transform -1 0 4830 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__997_
timestamp 0
transform 1 0 4670 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__998_
timestamp 0
transform -1 0 5290 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__999_
timestamp 0
transform -1 0 5090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1000_
timestamp 0
transform -1 0 4830 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1001_
timestamp 0
transform -1 0 4590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1002_
timestamp 0
transform -1 0 3390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1003_
timestamp 0
transform 1 0 3490 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1004_
timestamp 0
transform -1 0 4750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1005_
timestamp 0
transform -1 0 4990 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1006_
timestamp 0
transform -1 0 4330 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1007_
timestamp 0
transform -1 0 3830 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1008_
timestamp 0
transform 1 0 4130 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1009_
timestamp 0
transform -1 0 4650 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1010_
timestamp 0
transform -1 0 4430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1011_
timestamp 0
transform -1 0 4270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1012_
timestamp 0
transform -1 0 3670 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1013_
timestamp 0
transform 1 0 3910 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1014_
timestamp 0
transform -1 0 4370 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1015_
timestamp 0
transform 1 0 3970 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1016_
timestamp 0
transform -1 0 4050 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1017_
timestamp 0
transform 1 0 3430 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1018_
timestamp 0
transform -1 0 3710 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1019_
timestamp 0
transform -1 0 3290 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1020_
timestamp 0
transform 1 0 3530 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1021_
timestamp 0
transform -1 0 3850 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1022_
timestamp 0
transform -1 0 4490 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1023_
timestamp 0
transform 1 0 4130 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1024_
timestamp 0
transform 1 0 4250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1025_
timestamp 0
transform 1 0 4390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1026_
timestamp 0
transform -1 0 5330 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1027_
timestamp 0
transform 1 0 5090 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1028_
timestamp 0
transform -1 0 2110 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1029_
timestamp 0
transform 1 0 3530 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1030_
timestamp 0
transform 1 0 2350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1031_
timestamp 0
transform 1 0 2690 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1032_
timestamp 0
transform -1 0 1870 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1033_
timestamp 0
transform -1 0 2230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1034_
timestamp 0
transform -1 0 1530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1035_
timestamp 0
transform 1 0 1790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1036_
timestamp 0
transform 1 0 2810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1037_
timestamp 0
transform 1 0 2030 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1038_
timestamp 0
transform -1 0 2270 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1039_
timestamp 0
transform 1 0 1950 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1040_
timestamp 0
transform 1 0 2390 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1041_
timestamp 0
transform 1 0 4470 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1042_
timestamp 0
transform 1 0 3810 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1043_
timestamp 0
transform 1 0 3990 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1044_
timestamp 0
transform 1 0 3370 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1045_
timestamp 0
transform 1 0 2550 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1046_
timestamp 0
transform 1 0 2490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1047_
timestamp 0
transform 1 0 3670 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1048_
timestamp 0
transform -1 0 3370 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1049_
timestamp 0
transform 1 0 2710 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1050_
timestamp 0
transform 1 0 3650 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1051_
timestamp 0
transform 1 0 3030 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1052_
timestamp 0
transform 1 0 2870 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1053_
timestamp 0
transform 1 0 3210 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1054_
timestamp 0
transform 1 0 4550 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1055_
timestamp 0
transform 1 0 5830 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1056_
timestamp 0
transform -1 0 5890 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1057_
timestamp 0
transform 1 0 3810 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1058_
timestamp 0
transform 1 0 3850 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1059_
timestamp 0
transform -1 0 4470 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1060_
timestamp 0
transform -1 0 4110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1061_
timestamp 0
transform -1 0 3750 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1062_
timestamp 0
transform 1 0 4270 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1063_
timestamp 0
transform 1 0 3690 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1064_
timestamp 0
transform 1 0 3970 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1065_
timestamp 0
transform 1 0 4310 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1066_
timestamp 0
transform 1 0 3570 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1067_
timestamp 0
transform 1 0 4150 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1068_
timestamp 0
transform -1 0 4930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1069_
timestamp 0
transform 1 0 5570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1070_
timestamp 0
transform 1 0 5750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1071_
timestamp 0
transform -1 0 5370 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1072_
timestamp 0
transform -1 0 5250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1073_
timestamp 0
transform -1 0 5830 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1074_
timestamp 0
transform -1 0 5630 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1075_
timestamp 0
transform -1 0 5570 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1076_
timestamp 0
transform -1 0 5490 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1077_
timestamp 0
transform -1 0 5370 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1078_
timestamp 0
transform 1 0 5750 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1079_
timestamp 0
transform 1 0 5670 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1080_
timestamp 0
transform -1 0 5690 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1081_
timestamp 0
transform -1 0 5530 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1082_
timestamp 0
transform 1 0 5730 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1083_
timestamp 0
transform 1 0 5830 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1084_
timestamp 0
transform 1 0 5510 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1085_
timestamp 0
transform -1 0 5870 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1086_
timestamp 0
transform 1 0 5070 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1087_
timestamp 0
transform 1 0 5230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1088_
timestamp 0
transform -1 0 5890 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1089_
timestamp 0
transform 1 0 5570 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1090_
timestamp 0
transform -1 0 5570 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1091_
timestamp 0
transform -1 0 5410 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1092_
timestamp 0
transform 1 0 5730 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1093_
timestamp 0
transform 1 0 5570 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1094_
timestamp 0
transform 1 0 5710 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1095_
timestamp 0
transform 1 0 5390 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1096_
timestamp 0
transform -1 0 5770 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1097_
timestamp 0
transform 1 0 4870 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1098_
timestamp 0
transform -1 0 4430 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1099_
timestamp 0
transform 1 0 5790 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1100_
timestamp 0
transform 1 0 5410 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1101_
timestamp 0
transform -1 0 5590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1102_
timestamp 0
transform -1 0 5270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1103_
timestamp 0
transform -1 0 5170 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1104_
timestamp 0
transform 1 0 4990 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1105_
timestamp 0
transform -1 0 5650 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1106_
timestamp 0
transform 1 0 5050 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1107_
timestamp 0
transform -1 0 5170 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1108_
timestamp 0
transform -1 0 4330 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1109_
timestamp 0
transform -1 0 5330 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1110_
timestamp 0
transform -1 0 4990 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1111_
timestamp 0
transform -1 0 4830 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1112_
timestamp 0
transform -1 0 4170 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1113_
timestamp 0
transform 1 0 4690 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1114_
timestamp 0
transform 1 0 4530 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1115_
timestamp 0
transform -1 0 4650 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1116_
timestamp 0
transform 1 0 4470 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1117_
timestamp 0
transform -1 0 4530 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1118_
timestamp 0
transform 1 0 4110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1119_
timestamp 0
transform -1 0 3610 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1120_
timestamp 0
transform -1 0 3990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1121_
timestamp 0
transform -1 0 3990 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1122_
timestamp 0
transform -1 0 3810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1123_
timestamp 0
transform -1 0 4830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1124_
timestamp 0
transform 1 0 4630 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1125_
timestamp 0
transform 1 0 3950 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1126_
timestamp 0
transform 1 0 4310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1127_
timestamp 0
transform -1 0 5250 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1128_
timestamp 0
transform 1 0 4710 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1129_
timestamp 0
transform 1 0 2970 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1130_
timestamp 0
transform 1 0 2190 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1131_
timestamp 0
transform 1 0 2510 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1132_
timestamp 0
transform 1 0 2210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1133_
timestamp 0
transform 1 0 2030 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1134_
timestamp 0
transform 1 0 2370 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1135_
timestamp 0
transform -1 0 1350 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1136_
timestamp 0
transform -1 0 1730 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1137_
timestamp 0
transform 1 0 1710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1138_
timestamp 0
transform 1 0 2790 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1139_
timestamp 0
transform -1 0 2350 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1140_
timestamp 0
transform 1 0 1870 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1141_
timestamp 0
transform 1 0 2650 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1142_
timestamp 0
transform -1 0 4310 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1143_
timestamp 0
transform -1 0 4110 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1144_
timestamp 0
transform 1 0 3130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1145_
timestamp 0
transform 1 0 2490 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1146_
timestamp 0
transform 1 0 2630 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1147_
timestamp 0
transform -1 0 4430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1148_
timestamp 0
transform 1 0 3450 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1149_
timestamp 0
transform 1 0 3510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1150_
timestamp 0
transform 1 0 2810 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1151_
timestamp 0
transform -1 0 2990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1152_
timestamp 0
transform 1 0 3150 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1153_
timestamp 0
transform 1 0 3130 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1154_
timestamp 0
transform 1 0 2970 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1155_
timestamp 0
transform 1 0 3290 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1156_
timestamp 0
transform -1 0 3690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1157_
timestamp 0
transform -1 0 5350 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1158_
timestamp 0
transform -1 0 5190 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1159_
timestamp 0
transform -1 0 3970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1160_
timestamp 0
transform -1 0 3930 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1161_
timestamp 0
transform 1 0 2910 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1162_
timestamp 0
transform -1 0 3630 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1163_
timestamp 0
transform -1 0 1650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1164_
timestamp 0
transform 1 0 3250 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1165_
timestamp 0
transform 1 0 3750 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1166_
timestamp 0
transform 1 0 4190 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1167_
timestamp 0
transform 1 0 4350 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1168_
timestamp 0
transform 1 0 4510 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1169_
timestamp 0
transform 1 0 4670 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1170_
timestamp 0
transform 1 0 4830 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1171_
timestamp 0
transform -1 0 5670 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1172_
timestamp 0
transform -1 0 5510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1173_
timestamp 0
transform -1 0 5830 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1174_
timestamp 0
transform 1 0 5830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1175_
timestamp 0
transform 1 0 5630 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1176_
timestamp 0
transform -1 0 5490 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1177_
timestamp 0
transform -1 0 5550 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1178_
timestamp 0
transform -1 0 5330 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1179_
timestamp 0
transform -1 0 5010 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1180_
timestamp 0
transform 1 0 5750 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1181_
timestamp 0
transform 1 0 5810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1182_
timestamp 0
transform -1 0 5810 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1183_
timestamp 0
transform -1 0 5490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1184_
timestamp 0
transform 1 0 4930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1185_
timestamp 0
transform 1 0 5030 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1186_
timestamp 0
transform -1 0 5070 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1187_
timestamp 0
transform -1 0 4910 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1188_
timestamp 0
transform 1 0 4770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1189_
timestamp 0
transform 1 0 5130 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1190_
timestamp 0
transform 1 0 5150 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1191_
timestamp 0
transform -1 0 4990 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1192_
timestamp 0
transform -1 0 4930 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1193_
timestamp 0
transform 1 0 3810 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1194_
timestamp 0
transform 1 0 5190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1195_
timestamp 0
transform -1 0 4890 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1196_
timestamp 0
transform -1 0 4670 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1197_
timestamp 0
transform 1 0 4590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1198_
timestamp 0
transform -1 0 4790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1199_
timestamp 0
transform -1 0 4630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1200_
timestamp 0
transform -1 0 4830 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1201_
timestamp 0
transform 1 0 5070 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1202_
timestamp 0
transform -1 0 4590 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1203_
timestamp 0
transform -1 0 4250 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1204_
timestamp 0
transform -1 0 4750 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1205_
timestamp 0
transform -1 0 4450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1206_
timestamp 0
transform -1 0 4010 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1207_
timestamp 0
transform 1 0 3870 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1208_
timestamp 0
transform -1 0 5110 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1209_
timestamp 0
transform 1 0 4930 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1210_
timestamp 0
transform -1 0 4170 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1211_
timestamp 0
transform -1 0 4430 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1212_
timestamp 0
transform -1 0 4070 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1213_
timestamp 0
transform 1 0 4070 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1214_
timestamp 0
transform -1 0 3230 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1215_
timestamp 0
transform 1 0 3770 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1216_
timestamp 0
transform 1 0 3890 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1217_
timestamp 0
transform -1 0 4770 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1218_
timestamp 0
transform 1 0 4490 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1219_
timestamp 0
transform 1 0 3290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1220_
timestamp 0
transform 1 0 5130 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1221_
timestamp 0
transform 1 0 5290 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1222_
timestamp 0
transform 1 0 2030 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1223_
timestamp 0
transform 1 0 2890 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1224_
timestamp 0
transform -1 0 2330 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1225_
timestamp 0
transform 1 0 2070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1226_
timestamp 0
transform 1 0 1630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1227_
timestamp 0
transform -1 0 1810 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1228_
timestamp 0
transform 1 0 2630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1229_
timestamp 0
transform 1 0 2790 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1230_
timestamp 0
transform 1 0 2250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1231_
timestamp 0
transform -1 0 2470 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1232_
timestamp 0
transform -1 0 2630 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1233_
timestamp 0
transform 1 0 2950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1234_
timestamp 0
transform 1 0 4030 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1235_
timestamp 0
transform -1 0 3790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1236_
timestamp 0
transform 1 0 3610 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1237_
timestamp 0
transform 1 0 2790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1238_
timestamp 0
transform 1 0 2390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1239_
timestamp 0
transform -1 0 3430 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1240_
timestamp 0
transform 1 0 3110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1241_
timestamp 0
transform 1 0 3090 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1242_
timestamp 0
transform 1 0 3050 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1243_
timestamp 0
transform -1 0 3470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1244_
timestamp 0
transform 1 0 3270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1245_
timestamp 0
transform 1 0 3410 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1246_
timestamp 0
transform 1 0 4910 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1247_
timestamp 0
transform -1 0 5630 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1248_
timestamp 0
transform 1 0 5450 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1249_
timestamp 0
transform -1 0 3590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1250_
timestamp 0
transform 1 0 3130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1251_
timestamp 0
transform -1 0 2810 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1252_
timestamp 0
transform -1 0 3010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1253_
timestamp 0
transform -1 0 1070 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1254_
timestamp 0
transform 1 0 2950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1255_
timestamp 0
transform 1 0 3250 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1256_
timestamp 0
transform 1 0 3130 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1257_
timestamp 0
transform 1 0 3290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1258_
timestamp 0
transform 1 0 3510 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1259_
timestamp 0
transform -1 0 5750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1260_
timestamp 0
transform -1 0 5310 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1261_
timestamp 0
transform -1 0 5470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1262_
timestamp 0
transform 1 0 5850 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1263_
timestamp 0
transform -1 0 5730 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1264_
timestamp 0
transform -1 0 5630 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1265_
timestamp 0
transform -1 0 5650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1266_
timestamp 0
transform 1 0 5310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1267_
timestamp 0
transform -1 0 5790 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1268_
timestamp 0
transform 1 0 5770 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1269_
timestamp 0
transform -1 0 5490 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1270_
timestamp 0
transform 1 0 5070 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1271_
timestamp 0
transform 1 0 5690 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1272_
timestamp 0
transform -1 0 5450 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1273_
timestamp 0
transform -1 0 5290 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1274_
timestamp 0
transform -1 0 4990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1275_
timestamp 0
transform -1 0 4770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1276_
timestamp 0
transform 1 0 4570 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1277_
timestamp 0
transform 1 0 5630 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1278_
timestamp 0
transform -1 0 5570 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1279_
timestamp 0
transform -1 0 5410 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1280_
timestamp 0
transform 1 0 5210 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1281_
timestamp 0
transform -1 0 4790 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1282_
timestamp 0
transform -1 0 4630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1283_
timestamp 0
transform 1 0 4650 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1284_
timestamp 0
transform 1 0 5290 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1285_
timestamp 0
transform -1 0 4810 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1286_
timestamp 0
transform -1 0 4970 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1287_
timestamp 0
transform -1 0 4470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1288_
timestamp 0
transform 1 0 4210 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1289_
timestamp 0
transform 1 0 4330 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1290_
timestamp 0
transform -1 0 5130 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1291_
timestamp 0
transform -1 0 4510 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1292_
timestamp 0
transform -1 0 4350 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1293_
timestamp 0
transform 1 0 4170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1294_
timestamp 0
transform -1 0 3590 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1295_
timestamp 0
transform -1 0 4330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1296_
timestamp 0
transform 1 0 4010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1297_
timestamp 0
transform -1 0 3750 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1298_
timestamp 0
transform 1 0 3850 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1299_
timestamp 0
transform -1 0 4390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1300_
timestamp 0
transform 1 0 4210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1301_
timestamp 0
transform 1 0 3870 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1302_
timestamp 0
transform 1 0 4870 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1303_
timestamp 0
transform -1 0 5130 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1304_
timestamp 0
transform 1 0 2610 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1305_
timestamp 0
transform -1 0 1950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1306_
timestamp 0
transform 1 0 1550 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1307_
timestamp 0
transform -1 0 1710 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1308_
timestamp 0
transform -1 0 1710 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1309_
timestamp 0
transform 1 0 1990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1310_
timestamp 0
transform 1 0 2150 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1311_
timestamp 0
transform 1 0 1870 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1312_
timestamp 0
transform -1 0 2190 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1313_
timestamp 0
transform 1 0 2010 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1314_
timestamp 0
transform 1 0 2450 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1315_
timestamp 0
transform 1 0 2690 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1316_
timestamp 0
transform 1 0 2830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1317_
timestamp 0
transform 1 0 2690 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1318_
timestamp 0
transform 1 0 2270 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1319_
timestamp 0
transform -1 0 1770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1320_
timestamp 0
transform -1 0 3370 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1321_
timestamp 0
transform -1 0 3210 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1322_
timestamp 0
transform 1 0 2350 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1323_
timestamp 0
transform 1 0 2850 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1324_
timestamp 0
transform 1 0 2670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1325_
timestamp 0
transform 1 0 2510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1326_
timestamp 0
transform 1 0 2530 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1327_
timestamp 0
transform 1 0 3010 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1328_
timestamp 0
transform -1 0 3590 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1329_
timestamp 0
transform -1 0 5610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1330_
timestamp 0
transform -1 0 5430 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1331_
timestamp 0
transform 1 0 2330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1332_
timestamp 0
transform 1 0 2170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1333_
timestamp 0
transform 1 0 2530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1334_
timestamp 0
transform -1 0 3110 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1335_
timestamp 0
transform -1 0 2550 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1336_
timestamp 0
transform -1 0 2370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1337_
timestamp 0
transform 1 0 2370 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1338_
timestamp 0
transform 1 0 3230 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1339_
timestamp 0
transform -1 0 4150 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1340_
timestamp 0
transform 1 0 4030 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1341_
timestamp 0
transform 1 0 3390 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1342_
timestamp 0
transform 1 0 4330 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1343_
timestamp 0
transform 1 0 3370 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1344_
timestamp 0
transform -1 0 5270 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1345_
timestamp 0
transform 1 0 4470 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1346_
timestamp 0
transform -1 0 4190 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1347_
timestamp 0
transform 1 0 4950 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1348_
timestamp 0
transform -1 0 5330 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1349_
timestamp 0
transform 1 0 3710 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1350_
timestamp 0
transform -1 0 3890 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1351_
timestamp 0
transform 1 0 4630 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1352_
timestamp 0
transform -1 0 5170 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1353_
timestamp 0
transform 1 0 4310 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1354_
timestamp 0
transform -1 0 4810 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1355_
timestamp 0
transform -1 0 4590 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1356_
timestamp 0
transform -1 0 4430 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1357_
timestamp 0
transform -1 0 5150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1358_
timestamp 0
transform -1 0 4650 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1359_
timestamp 0
transform 1 0 4690 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1360_
timestamp 0
transform -1 0 5010 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1361_
timestamp 0
transform -1 0 4770 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1362_
timestamp 0
transform 1 0 4270 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1363_
timestamp 0
transform 1 0 4010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1364_
timestamp 0
transform -1 0 3910 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1365_
timestamp 0
transform -1 0 4410 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1366_
timestamp 0
transform -1 0 4250 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1367_
timestamp 0
transform 1 0 2810 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1368_
timestamp 0
transform 1 0 3290 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1369_
timestamp 0
transform 1 0 3990 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1370_
timestamp 0
transform -1 0 3850 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1371_
timestamp 0
transform 1 0 2170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1372_
timestamp 0
transform -1 0 1590 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1373_
timestamp 0
transform -1 0 1490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1374_
timestamp 0
transform 1 0 1130 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1375_
timestamp 0
transform 1 0 1410 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1376_
timestamp 0
transform 1 0 1250 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1377_
timestamp 0
transform -1 0 1210 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1378_
timestamp 0
transform -1 0 1850 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1379_
timestamp 0
transform 1 0 1430 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1380_
timestamp 0
transform 1 0 1290 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1381_
timestamp 0
transform 1 0 1350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1382_
timestamp 0
transform 1 0 1490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1383_
timestamp 0
transform 1 0 1730 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1384_
timestamp 0
transform -1 0 2090 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1385_
timestamp 0
transform -1 0 1750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1386_
timestamp 0
transform -1 0 1590 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1387_
timestamp 0
transform -1 0 1150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1388_
timestamp 0
transform 1 0 1570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1389_
timestamp 0
transform -1 0 1890 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1390_
timestamp 0
transform -1 0 2250 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1391_
timestamp 0
transform 1 0 1890 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1392_
timestamp 0
transform 1 0 1410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1393_
timestamp 0
transform -1 0 1870 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1394_
timestamp 0
transform 1 0 2590 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1395_
timestamp 0
transform 1 0 2950 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1396_
timestamp 0
transform -1 0 2790 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1397_
timestamp 0
transform -1 0 2650 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1398_
timestamp 0
transform -1 0 2410 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1399_
timestamp 0
transform 1 0 2210 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1400_
timestamp 0
transform 1 0 2010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1401_
timestamp 0
transform 1 0 2030 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1402_
timestamp 0
transform 1 0 2510 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1403_
timestamp 0
transform -1 0 2970 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1404_
timestamp 0
transform -1 0 3270 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1405_
timestamp 0
transform -1 0 3710 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1406_
timestamp 0
transform -1 0 3550 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1407_
timestamp 0
transform 1 0 2990 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1408_
timestamp 0
transform 1 0 3630 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1409_
timestamp 0
transform 1 0 2830 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1410_
timestamp 0
transform -1 0 3110 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1411_
timestamp 0
transform 1 0 3310 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1412_
timestamp 0
transform 1 0 3790 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1413_
timestamp 0
transform 1 0 4470 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1414_
timestamp 0
transform -1 0 4530 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1415_
timestamp 0
transform -1 0 3170 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1416_
timestamp 0
transform 1 0 3470 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1417_
timestamp 0
transform -1 0 3970 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1418_
timestamp 0
transform 1 0 3610 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1419_
timestamp 0
transform 1 0 3570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1420_
timestamp 0
transform 1 0 4070 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1421_
timestamp 0
transform 1 0 3710 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1422_
timestamp 0
transform -1 0 3430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1423_
timestamp 0
transform -1 0 4130 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1424_
timestamp 0
transform -1 0 3450 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1425_
timestamp 0
transform 1 0 3750 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1426_
timestamp 0
transform 1 0 2950 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1427_
timestamp 0
transform -1 0 2670 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1428_
timestamp 0
transform 1 0 1710 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1429_
timestamp 0
transform -1 0 1210 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1430_
timestamp 0
transform -1 0 2490 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1431_
timestamp 0
transform 1 0 1410 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1432_
timestamp 0
transform 1 0 670 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1433_
timestamp 0
transform -1 0 1310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1434_
timestamp 0
transform 1 0 1130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1435_
timestamp 0
transform 1 0 1090 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1436_
timestamp 0
transform 1 0 990 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1437_
timestamp 0
transform 1 0 950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1438_
timestamp 0
transform -1 0 1110 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1439_
timestamp 0
transform -1 0 810 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1440_
timestamp 0
transform 1 0 1250 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1441_
timestamp 0
transform -1 0 510 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1442_
timestamp 0
transform 1 0 50 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1443_
timestamp 0
transform -1 0 2470 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1444_
timestamp 0
transform -1 0 210 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1445_
timestamp 0
transform 1 0 490 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1446_
timestamp 0
transform -1 0 370 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1447_
timestamp 0
transform -1 0 70 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1448_
timestamp 0
transform 1 0 190 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1449_
timestamp 0
transform -1 0 650 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1450_
timestamp 0
transform -1 0 650 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1451_
timestamp 0
transform -1 0 930 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1452_
timestamp 0
transform -1 0 930 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1453_
timestamp 0
transform -1 0 790 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1454_
timestamp 0
transform 1 0 1030 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1455_
timestamp 0
transform 1 0 1070 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1456_
timestamp 0
transform 1 0 1230 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1457_
timestamp 0
transform -1 0 2090 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1458_
timestamp 0
transform -1 0 2690 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1459_
timestamp 0
transform -1 0 2810 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1460_
timestamp 0
transform -1 0 1910 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1461_
timestamp 0
transform 1 0 1810 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1462_
timestamp 0
transform -1 0 1970 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1463_
timestamp 0
transform 1 0 1770 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1464_
timestamp 0
transform -1 0 1630 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1465_
timestamp 0
transform 1 0 1310 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1466_
timestamp 0
transform 1 0 810 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1467_
timestamp 0
transform -1 0 610 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1468_
timestamp 0
transform 1 0 950 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1469_
timestamp 0
transform 1 0 650 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1470_
timestamp 0
transform -1 0 1270 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1471_
timestamp 0
transform 1 0 790 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1472_
timestamp 0
transform -1 0 70 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1473_
timestamp 0
transform -1 0 70 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1474_
timestamp 0
transform -1 0 70 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1475_
timestamp 0
transform 1 0 550 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1476_
timestamp 0
transform 1 0 230 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1477_
timestamp 0
transform 1 0 670 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1478_
timestamp 0
transform 1 0 330 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1479_
timestamp 0
transform 1 0 250 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1480_
timestamp 0
transform -1 0 410 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1481_
timestamp 0
transform 1 0 390 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1482_
timestamp 0
transform -1 0 850 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1483_
timestamp 0
transform -1 0 1430 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1484_
timestamp 0
transform -1 0 1510 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1485_
timestamp 0
transform -1 0 1350 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1486_
timestamp 0
transform -1 0 1670 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1487_
timestamp 0
transform -1 0 1450 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1488_
timestamp 0
transform 1 0 1470 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1489_
timestamp 0
transform 1 0 1250 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1490_
timestamp 0
transform 1 0 530 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1491_
timestamp 0
transform -1 0 830 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1492_
timestamp 0
transform 1 0 650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1493_
timestamp 0
transform -1 0 530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1494_
timestamp 0
transform 1 0 230 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1495_
timestamp 0
transform 1 0 350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1496_
timestamp 0
transform 1 0 750 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1497_
timestamp 0
transform 1 0 250 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1498_
timestamp 0
transform 1 0 50 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1499_
timestamp 0
transform -1 0 270 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1500_
timestamp 0
transform 1 0 890 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1501_
timestamp 0
transform -1 0 990 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1502_
timestamp 0
transform -1 0 970 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1503_
timestamp 0
transform -1 0 950 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1504_
timestamp 0
transform 1 0 650 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1505_
timestamp 0
transform -1 0 790 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1506_
timestamp 0
transform -1 0 610 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1507_
timestamp 0
transform 1 0 50 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1508_
timestamp 0
transform -1 0 70 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1509_
timestamp 0
transform -1 0 410 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1510_
timestamp 0
transform 1 0 310 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1511_
timestamp 0
transform 1 0 3090 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1512_
timestamp 0
transform -1 0 1570 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1513_
timestamp 0
transform -1 0 1190 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1514_
timestamp 0
transform -1 0 1110 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1515_
timestamp 0
transform -1 0 210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1516_
timestamp 0
transform -1 0 610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1517_
timestamp 0
transform -1 0 470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1518_
timestamp 0
transform 1 0 1310 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1519_
timestamp 0
transform 1 0 2210 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1560_
timestamp 0
transform -1 0 70 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1561_
timestamp 0
transform -1 0 210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1562_
timestamp 0
transform -1 0 70 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1563_
timestamp 0
transform -1 0 70 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1564_
timestamp 0
transform -1 0 350 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1565_
timestamp 0
transform 1 0 3890 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1566_
timestamp 0
transform -1 0 1010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1567_
timestamp 0
transform -1 0 70 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1568_
timestamp 0
transform -1 0 70 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1569_
timestamp 0
transform -1 0 70 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1570_
timestamp 0
transform -1 0 3710 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1571_
timestamp 0
transform 1 0 5110 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1572_
timestamp 0
transform -1 0 2350 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1573_
timestamp 0
transform 1 0 2190 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1574_
timestamp 0
transform -1 0 70 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1575_
timestamp 0
transform -1 0 230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1576_
timestamp 0
transform -1 0 70 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1577_
timestamp 0
transform -1 0 370 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1578_
timestamp 0
transform 1 0 1610 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1579_
timestamp 0
transform 1 0 2230 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1580_
timestamp 0
transform -1 0 2750 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1581_
timestamp 0
transform -1 0 3090 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1582_
timestamp 0
transform -1 0 70 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1583_
timestamp 0
transform -1 0 3270 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert6
timestamp 0
transform 1 0 5090 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert7
timestamp 0
transform -1 0 3130 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert8
timestamp 0
transform -1 0 3130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert9
timestamp 0
transform -1 0 5850 0 -1 270
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert10
timestamp 0
transform 1 0 1650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert11
timestamp 0
transform 1 0 1770 0 1 4430
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert12
timestamp 0
transform 1 0 1530 0 1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert13
timestamp 0
transform -1 0 70 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert14
timestamp 0
transform -1 0 2770 0 1 2350
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert15
timestamp 0
transform -1 0 4070 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert16
timestamp 0
transform 1 0 4270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert17
timestamp 0
transform 1 0 4190 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert0
timestamp 0
transform 1 0 1450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert1
timestamp 0
transform -1 0 1290 0 1 3390
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert2
timestamp 0
transform -1 0 750 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert3
timestamp 0
transform -1 0 1090 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert4
timestamp 0
transform -1 0 1070 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert5
timestamp 0
transform 1 0 3030 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__756_
timestamp 0
transform 1 0 1330 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__757_
timestamp 0
transform 1 0 1690 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__758_
timestamp 0
transform 1 0 1450 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__759_
timestamp 0
transform 1 0 590 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__760_
timestamp 0
transform 1 0 730 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__761_
timestamp 0
transform 1 0 450 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__762_
timestamp 0
transform 1 0 450 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__763_
timestamp 0
transform -1 0 1190 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__764_
timestamp 0
transform 1 0 970 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__765_
timestamp 0
transform -1 0 470 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__766_
timestamp 0
transform 1 0 630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__767_
timestamp 0
transform 1 0 790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__768_
timestamp 0
transform -1 0 930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__769_
timestamp 0
transform 1 0 710 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__770_
timestamp 0
transform 1 0 850 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__771_
timestamp 0
transform 1 0 1010 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__772_
timestamp 0
transform -1 0 1190 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__773_
timestamp 0
transform -1 0 870 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__774_
timestamp 0
transform 1 0 690 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__775_
timestamp 0
transform -1 0 3150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__776_
timestamp 0
transform -1 0 1490 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__777_
timestamp 0
transform -1 0 1030 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__778_
timestamp 0
transform 1 0 390 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__779_
timestamp 0
transform 1 0 550 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__780_
timestamp 0
transform 1 0 70 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__781_
timestamp 0
transform 1 0 70 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__782_
timestamp 0
transform 1 0 510 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__783_
timestamp 0
transform 1 0 630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__784_
timestamp 0
transform 1 0 230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__785_
timestamp 0
transform 1 0 350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__786_
timestamp 0
transform -1 0 830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__787_
timestamp 0
transform 1 0 970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__788_
timestamp 0
transform 1 0 1610 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__789_
timestamp 0
transform -1 0 1210 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__790_
timestamp 0
transform -1 0 1370 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__791_
timestamp 0
transform 1 0 1310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__792_
timestamp 0
transform -1 0 1450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__793_
timestamp 0
transform -1 0 1050 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__794_
timestamp 0
transform 1 0 970 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__795_
timestamp 0
transform -1 0 890 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__796_
timestamp 0
transform 1 0 830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__797_
timestamp 0
transform 1 0 1130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__798_
timestamp 0
transform -1 0 930 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__799_
timestamp 0
transform -1 0 3490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__800_
timestamp 0
transform 1 0 2250 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__801_
timestamp 0
transform 1 0 2330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__802_
timestamp 0
transform 1 0 1910 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__803_
timestamp 0
transform -1 0 1610 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__804_
timestamp 0
transform -1 0 1310 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__805_
timestamp 0
transform -1 0 250 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__806_
timestamp 0
transform -1 0 790 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__807_
timestamp 0
transform 1 0 890 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__808_
timestamp 0
transform 1 0 490 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__809_
timestamp 0
transform 1 0 70 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__810_
timestamp 0
transform -1 0 250 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__811_
timestamp 0
transform 1 0 190 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__812_
timestamp 0
transform -1 0 750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__813_
timestamp 0
transform -1 0 370 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__814_
timestamp 0
transform -1 0 90 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__815_
timestamp 0
transform 1 0 390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__816_
timestamp 0
transform 1 0 450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__817_
timestamp 0
transform -1 0 90 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__818_
timestamp 0
transform -1 0 250 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__819_
timestamp 0
transform -1 0 590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__820_
timestamp 0
transform -1 0 210 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__821_
timestamp 0
transform 1 0 930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__822_
timestamp 0
transform 1 0 2050 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__823_
timestamp 0
transform -1 0 1770 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__824_
timestamp 0
transform 1 0 670 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__825_
timestamp 0
transform 1 0 610 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__826_
timestamp 0
transform 1 0 970 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__827_
timestamp 0
transform -1 0 1290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__828_
timestamp 0
transform 1 0 770 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__829_
timestamp 0
transform -1 0 1110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__830_
timestamp 0
transform 1 0 370 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__831_
timestamp 0
transform -1 0 1510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__832_
timestamp 0
transform 1 0 610 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__833_
timestamp 0
transform -1 0 1190 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__834_
timestamp 0
transform 1 0 2110 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__835_
timestamp 0
transform 1 0 1130 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__836_
timestamp 0
transform 1 0 650 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__837_
timestamp 0
transform 1 0 1010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__838_
timestamp 0
transform -1 0 2430 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__839_
timestamp 0
transform -1 0 2610 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__840_
timestamp 0
transform -1 0 1790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__841_
timestamp 0
transform -1 0 2590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__842_
timestamp 0
transform 1 0 2110 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__843_
timestamp 0
transform -1 0 1850 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__844_
timestamp 0
transform 1 0 1890 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__845_
timestamp 0
transform -1 0 1970 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__846_
timestamp 0
transform -1 0 1630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__847_
timestamp 0
transform -1 0 1010 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__848_
timestamp 0
transform 1 0 810 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__849_
timestamp 0
transform -1 0 2030 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__850_
timestamp 0
transform -1 0 1690 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__851_
timestamp 0
transform -1 0 1370 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__852_
timestamp 0
transform 1 0 2370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__853_
timestamp 0
transform 1 0 2810 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__854_
timestamp 0
transform 1 0 2070 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__855_
timestamp 0
transform -1 0 1630 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__856_
timestamp 0
transform 1 0 1610 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__857_
timestamp 0
transform -1 0 1950 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__858_
timestamp 0
transform -1 0 2290 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__859_
timestamp 0
transform 1 0 2690 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__860_
timestamp 0
transform -1 0 2550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__861_
timestamp 0
transform 1 0 1730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__862_
timestamp 0
transform -1 0 1790 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__863_
timestamp 0
transform 1 0 1910 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__864_
timestamp 0
transform -1 0 1050 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__865_
timestamp 0
transform 1 0 1510 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__866_
timestamp 0
transform -1 0 1790 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__867_
timestamp 0
transform 1 0 2110 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__868_
timestamp 0
transform 1 0 2210 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__869_
timestamp 0
transform 1 0 2190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__870_
timestamp 0
transform 1 0 1590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__871_
timestamp 0
transform 1 0 1450 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__872_
timestamp 0
transform -1 0 830 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__873_
timestamp 0
transform 1 0 1750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__874_
timestamp 0
transform 1 0 1190 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__875_
timestamp 0
transform 1 0 2070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__876_
timestamp 0
transform -1 0 2270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__877_
timestamp 0
transform 1 0 1410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__878_
timestamp 0
transform 1 0 1630 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__879_
timestamp 0
transform 1 0 1910 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__880_
timestamp 0
transform -1 0 1690 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__881_
timestamp 0
transform 1 0 2430 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__882_
timestamp 0
transform 1 0 1850 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__883_
timestamp 0
transform 1 0 2010 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__884_
timestamp 0
transform -1 0 1950 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__885_
timestamp 0
transform 1 0 1310 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__886_
timestamp 0
transform 1 0 1810 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__887_
timestamp 0
transform -1 0 2410 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__888_
timestamp 0
transform 1 0 2510 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__889_
timestamp 0
transform 1 0 2730 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__890_
timestamp 0
transform 1 0 1510 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__891_
timestamp 0
transform 1 0 2690 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__892_
timestamp 0
transform 1 0 2830 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__893_
timestamp 0
transform 1 0 3250 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__894_
timestamp 0
transform 1 0 2970 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__895_
timestamp 0
transform 1 0 3410 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__896_
timestamp 0
transform 1 0 2530 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__897_
timestamp 0
transform 1 0 2950 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__898_
timestamp 0
transform 1 0 2670 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__899_
timestamp 0
transform -1 0 3190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__900_
timestamp 0
transform -1 0 3030 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__901_
timestamp 0
transform 1 0 2850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__902_
timestamp 0
transform 1 0 3610 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__903_
timestamp 0
transform 1 0 2650 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__904_
timestamp 0
transform -1 0 4570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__905_
timestamp 0
transform -1 0 4870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__906_
timestamp 0
transform -1 0 5330 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__907_
timestamp 0
transform -1 0 4570 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__908_
timestamp 0
transform -1 0 4990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__909_
timestamp 0
transform 1 0 4690 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__910_
timestamp 0
transform -1 0 4710 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__911_
timestamp 0
transform -1 0 4850 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__912_
timestamp 0
transform 1 0 4370 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__913_
timestamp 0
transform -1 0 4830 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__914_
timestamp 0
transform 1 0 4390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__915_
timestamp 0
transform 1 0 4370 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__916_
timestamp 0
transform -1 0 4670 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__917_
timestamp 0
transform -1 0 4990 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__918_
timestamp 0
transform 1 0 4210 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__919_
timestamp 0
transform -1 0 3790 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__920_
timestamp 0
transform 1 0 3610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__921_
timestamp 0
transform -1 0 4050 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__922_
timestamp 0
transform -1 0 4510 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__923_
timestamp 0
transform -1 0 3890 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__924_
timestamp 0
transform 1 0 2970 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__925_
timestamp 0
transform 1 0 1350 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__926_
timestamp 0
transform -1 0 3710 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__927_
timestamp 0
transform 1 0 3750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__928_
timestamp 0
transform 1 0 3450 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__929_
timestamp 0
transform -1 0 3090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__930_
timestamp 0
transform 1 0 2390 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__931_
timestamp 0
transform -1 0 2550 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__932_
timestamp 0
transform -1 0 3310 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__933_
timestamp 0
transform -1 0 2830 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__934_
timestamp 0
transform 1 0 2650 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__935_
timestamp 0
transform -1 0 2750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__936_
timestamp 0
transform 1 0 2410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__937_
timestamp 0
transform 1 0 2490 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__938_
timestamp 0
transform -1 0 2930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__939_
timestamp 0
transform -1 0 2590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__940_
timestamp 0
transform 1 0 2310 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__941_
timestamp 0
transform -1 0 2150 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__942_
timestamp 0
transform 1 0 3010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__943_
timestamp 0
transform 1 0 2870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__944_
timestamp 0
transform -1 0 2850 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__945_
timestamp 0
transform 1 0 2710 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__946_
timestamp 0
transform -1 0 2970 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__947_
timestamp 0
transform 1 0 3130 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__948_
timestamp 0
transform 1 0 3230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__949_
timestamp 0
transform 1 0 1350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__950_
timestamp 0
transform 1 0 1430 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__951_
timestamp 0
transform 1 0 1950 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__952_
timestamp 0
transform 1 0 3310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__953_
timestamp 0
transform 1 0 4890 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__954_
timestamp 0
transform -1 0 4250 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__955_
timestamp 0
transform 1 0 3930 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__956_
timestamp 0
transform 1 0 3110 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__957_
timestamp 0
transform 1 0 3250 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__958_
timestamp 0
transform 1 0 3350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__959_
timestamp 0
transform -1 0 4190 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__960_
timestamp 0
transform 1 0 2110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__961_
timestamp 0
transform 1 0 3470 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__962_
timestamp 0
transform 1 0 3530 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__963_
timestamp 0
transform 1 0 3990 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__964_
timestamp 0
transform 1 0 3690 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__965_
timestamp 0
transform 1 0 3530 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__966_
timestamp 0
transform 1 0 3850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__967_
timestamp 0
transform 1 0 5270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__968_
timestamp 0
transform -1 0 5170 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__969_
timestamp 0
transform 1 0 4970 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__970_
timestamp 0
transform 1 0 5130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__971_
timestamp 0
transform -1 0 5270 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__972_
timestamp 0
transform -1 0 5410 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__973_
timestamp 0
transform -1 0 5950 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__974_
timestamp 0
transform -1 0 5490 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__975_
timestamp 0
transform -1 0 5290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__976_
timestamp 0
transform -1 0 5710 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__977_
timestamp 0
transform 1 0 5630 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__978_
timestamp 0
transform -1 0 5810 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__979_
timestamp 0
transform -1 0 5630 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__980_
timestamp 0
transform -1 0 5470 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__981_
timestamp 0
transform -1 0 5930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__982_
timestamp 0
transform 1 0 5770 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__983_
timestamp 0
transform 1 0 5430 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__984_
timestamp 0
transform -1 0 5770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__985_
timestamp 0
transform -1 0 5290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__986_
timestamp 0
transform -1 0 5690 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__987_
timestamp 0
transform 1 0 5590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__988_
timestamp 0
transform 1 0 5490 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__989_
timestamp 0
transform -1 0 5190 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__990_
timestamp 0
transform 1 0 4090 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__991_
timestamp 0
transform 1 0 4210 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__992_
timestamp 0
transform -1 0 5510 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__993_
timestamp 0
transform -1 0 5450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__994_
timestamp 0
transform -1 0 5450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__995_
timestamp 0
transform -1 0 4930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__996_
timestamp 0
transform -1 0 4850 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__997_
timestamp 0
transform 1 0 4690 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__998_
timestamp 0
transform -1 0 5310 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__999_
timestamp 0
transform -1 0 5110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1000_
timestamp 0
transform -1 0 4850 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1001_
timestamp 0
transform -1 0 4610 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1002_
timestamp 0
transform -1 0 3410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1003_
timestamp 0
transform 1 0 3510 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1004_
timestamp 0
transform -1 0 4770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1005_
timestamp 0
transform -1 0 5010 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1006_
timestamp 0
transform -1 0 4350 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1007_
timestamp 0
transform -1 0 3850 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1008_
timestamp 0
transform 1 0 4150 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1009_
timestamp 0
transform -1 0 4670 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1010_
timestamp 0
transform -1 0 4450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1011_
timestamp 0
transform -1 0 4290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1012_
timestamp 0
transform -1 0 3690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1013_
timestamp 0
transform 1 0 3930 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1014_
timestamp 0
transform -1 0 4390 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1015_
timestamp 0
transform 1 0 3990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1016_
timestamp 0
transform -1 0 4070 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1017_
timestamp 0
transform 1 0 3450 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1018_
timestamp 0
transform -1 0 3730 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1019_
timestamp 0
transform -1 0 3310 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1020_
timestamp 0
transform 1 0 3550 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1021_
timestamp 0
transform -1 0 3870 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1022_
timestamp 0
transform -1 0 4510 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1023_
timestamp 0
transform 1 0 4150 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1024_
timestamp 0
transform 1 0 4270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1025_
timestamp 0
transform 1 0 4410 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1026_
timestamp 0
transform -1 0 5350 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1027_
timestamp 0
transform 1 0 5110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1028_
timestamp 0
transform -1 0 2130 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1029_
timestamp 0
transform 1 0 3550 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1030_
timestamp 0
transform 1 0 2370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1031_
timestamp 0
transform 1 0 2710 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1032_
timestamp 0
transform -1 0 1890 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1033_
timestamp 0
transform -1 0 2250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1034_
timestamp 0
transform -1 0 1550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1035_
timestamp 0
transform 1 0 1810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1036_
timestamp 0
transform 1 0 2830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1037_
timestamp 0
transform 1 0 2050 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1038_
timestamp 0
transform -1 0 2290 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1039_
timestamp 0
transform 1 0 1970 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1040_
timestamp 0
transform 1 0 2410 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1041_
timestamp 0
transform 1 0 4490 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1042_
timestamp 0
transform 1 0 3830 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1043_
timestamp 0
transform 1 0 4010 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1044_
timestamp 0
transform 1 0 3390 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1045_
timestamp 0
transform 1 0 2570 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1046_
timestamp 0
transform 1 0 2510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1047_
timestamp 0
transform 1 0 3690 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1048_
timestamp 0
transform -1 0 3390 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1049_
timestamp 0
transform 1 0 2730 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1050_
timestamp 0
transform 1 0 3670 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1051_
timestamp 0
transform 1 0 3050 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1052_
timestamp 0
transform 1 0 2890 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1053_
timestamp 0
transform 1 0 3230 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1054_
timestamp 0
transform 1 0 4570 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1055_
timestamp 0
transform 1 0 5850 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1056_
timestamp 0
transform -1 0 5910 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1057_
timestamp 0
transform 1 0 3830 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1058_
timestamp 0
transform 1 0 3870 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1059_
timestamp 0
transform -1 0 4490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1060_
timestamp 0
transform -1 0 4130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1061_
timestamp 0
transform -1 0 3770 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1062_
timestamp 0
transform 1 0 4290 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1063_
timestamp 0
transform 1 0 3710 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1064_
timestamp 0
transform 1 0 3990 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1065_
timestamp 0
transform 1 0 4330 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1066_
timestamp 0
transform 1 0 3590 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1067_
timestamp 0
transform 1 0 4170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1068_
timestamp 0
transform -1 0 4950 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1069_
timestamp 0
transform 1 0 5590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1070_
timestamp 0
transform 1 0 5770 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1071_
timestamp 0
transform -1 0 5390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1072_
timestamp 0
transform -1 0 5270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1073_
timestamp 0
transform -1 0 5850 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1074_
timestamp 0
transform -1 0 5650 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1075_
timestamp 0
transform -1 0 5590 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1076_
timestamp 0
transform -1 0 5510 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1077_
timestamp 0
transform -1 0 5390 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1078_
timestamp 0
transform 1 0 5770 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1079_
timestamp 0
transform 1 0 5690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1080_
timestamp 0
transform -1 0 5710 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1081_
timestamp 0
transform -1 0 5550 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1082_
timestamp 0
transform 1 0 5750 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1083_
timestamp 0
transform 1 0 5850 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1084_
timestamp 0
transform 1 0 5530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1085_
timestamp 0
transform -1 0 5890 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1086_
timestamp 0
transform 1 0 5090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1087_
timestamp 0
transform 1 0 5250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1088_
timestamp 0
transform -1 0 5910 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1089_
timestamp 0
transform 1 0 5590 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1090_
timestamp 0
transform -1 0 5590 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1091_
timestamp 0
transform -1 0 5430 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1092_
timestamp 0
transform 1 0 5750 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1093_
timestamp 0
transform 1 0 5590 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1094_
timestamp 0
transform 1 0 5730 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1095_
timestamp 0
transform 1 0 5410 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1096_
timestamp 0
transform -1 0 5790 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1097_
timestamp 0
transform 1 0 4890 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1098_
timestamp 0
transform -1 0 4450 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1099_
timestamp 0
transform 1 0 5810 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1100_
timestamp 0
transform 1 0 5430 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1101_
timestamp 0
transform -1 0 5610 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1102_
timestamp 0
transform -1 0 5290 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1103_
timestamp 0
transform -1 0 5190 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1104_
timestamp 0
transform 1 0 5010 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1105_
timestamp 0
transform -1 0 5670 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1106_
timestamp 0
transform 1 0 5070 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1107_
timestamp 0
transform -1 0 5190 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1108_
timestamp 0
transform -1 0 4350 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1109_
timestamp 0
transform -1 0 5350 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1110_
timestamp 0
transform -1 0 5010 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1111_
timestamp 0
transform -1 0 4850 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1112_
timestamp 0
transform -1 0 4190 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1113_
timestamp 0
transform 1 0 4710 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1114_
timestamp 0
transform 1 0 4550 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1115_
timestamp 0
transform -1 0 4670 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1116_
timestamp 0
transform 1 0 4490 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1117_
timestamp 0
transform -1 0 4550 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1118_
timestamp 0
transform 1 0 4130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1119_
timestamp 0
transform -1 0 3630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1120_
timestamp 0
transform -1 0 4010 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1121_
timestamp 0
transform -1 0 4010 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1122_
timestamp 0
transform -1 0 3830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1123_
timestamp 0
transform -1 0 4850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1124_
timestamp 0
transform 1 0 4650 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1125_
timestamp 0
transform 1 0 3970 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1126_
timestamp 0
transform 1 0 4330 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1127_
timestamp 0
transform -1 0 5270 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1128_
timestamp 0
transform 1 0 4730 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1129_
timestamp 0
transform 1 0 2990 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1130_
timestamp 0
transform 1 0 2210 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1131_
timestamp 0
transform 1 0 2530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1132_
timestamp 0
transform 1 0 2230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1133_
timestamp 0
transform 1 0 2050 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1134_
timestamp 0
transform 1 0 2390 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1135_
timestamp 0
transform -1 0 1370 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1136_
timestamp 0
transform -1 0 1750 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1137_
timestamp 0
transform 1 0 1730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1138_
timestamp 0
transform 1 0 2810 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1139_
timestamp 0
transform -1 0 2370 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1140_
timestamp 0
transform 1 0 1890 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1141_
timestamp 0
transform 1 0 2670 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1142_
timestamp 0
transform -1 0 4330 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1143_
timestamp 0
transform -1 0 4130 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1144_
timestamp 0
transform 1 0 3150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1145_
timestamp 0
transform 1 0 2510 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1146_
timestamp 0
transform 1 0 2650 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1147_
timestamp 0
transform -1 0 4450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1148_
timestamp 0
transform 1 0 3470 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1149_
timestamp 0
transform 1 0 3530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1150_
timestamp 0
transform 1 0 2830 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1151_
timestamp 0
transform -1 0 3010 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1152_
timestamp 0
transform 1 0 3170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1153_
timestamp 0
transform 1 0 3150 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1154_
timestamp 0
transform 1 0 2990 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1155_
timestamp 0
transform 1 0 3310 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1156_
timestamp 0
transform -1 0 3710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1157_
timestamp 0
transform -1 0 5370 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1158_
timestamp 0
transform -1 0 5210 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1159_
timestamp 0
transform -1 0 3990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1160_
timestamp 0
transform -1 0 3950 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1161_
timestamp 0
transform 1 0 2930 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1162_
timestamp 0
transform -1 0 3650 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1163_
timestamp 0
transform -1 0 1670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1164_
timestamp 0
transform 1 0 3270 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1165_
timestamp 0
transform 1 0 3770 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1166_
timestamp 0
transform 1 0 4210 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1167_
timestamp 0
transform 1 0 4370 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1168_
timestamp 0
transform 1 0 4530 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1169_
timestamp 0
transform 1 0 4690 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1170_
timestamp 0
transform 1 0 4850 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1171_
timestamp 0
transform -1 0 5690 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1172_
timestamp 0
transform -1 0 5530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1173_
timestamp 0
transform -1 0 5850 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1174_
timestamp 0
transform 1 0 5850 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1175_
timestamp 0
transform 1 0 5650 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1176_
timestamp 0
transform -1 0 5510 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1177_
timestamp 0
transform -1 0 5570 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1178_
timestamp 0
transform -1 0 5350 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1179_
timestamp 0
transform -1 0 5030 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1180_
timestamp 0
transform 1 0 5770 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1181_
timestamp 0
transform 1 0 5830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1182_
timestamp 0
transform -1 0 5830 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1183_
timestamp 0
transform -1 0 5510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1184_
timestamp 0
transform 1 0 4950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1185_
timestamp 0
transform 1 0 5050 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1186_
timestamp 0
transform -1 0 5090 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1187_
timestamp 0
transform -1 0 4930 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1188_
timestamp 0
transform 1 0 4790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1189_
timestamp 0
transform 1 0 5150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1190_
timestamp 0
transform 1 0 5170 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1191_
timestamp 0
transform -1 0 5010 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1192_
timestamp 0
transform -1 0 4950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1193_
timestamp 0
transform 1 0 3830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1194_
timestamp 0
transform 1 0 5210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1195_
timestamp 0
transform -1 0 4910 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1196_
timestamp 0
transform -1 0 4690 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1197_
timestamp 0
transform 1 0 4610 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1198_
timestamp 0
transform -1 0 4810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1199_
timestamp 0
transform -1 0 4650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1200_
timestamp 0
transform -1 0 4850 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1201_
timestamp 0
transform 1 0 5090 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1202_
timestamp 0
transform -1 0 4610 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1203_
timestamp 0
transform -1 0 4270 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1204_
timestamp 0
transform -1 0 4770 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1205_
timestamp 0
transform -1 0 4470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1206_
timestamp 0
transform -1 0 4030 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1207_
timestamp 0
transform 1 0 3890 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1208_
timestamp 0
transform -1 0 5130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1209_
timestamp 0
transform 1 0 4950 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1210_
timestamp 0
transform -1 0 4190 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1211_
timestamp 0
transform -1 0 4450 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1212_
timestamp 0
transform -1 0 4090 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1213_
timestamp 0
transform 1 0 4090 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1214_
timestamp 0
transform -1 0 3250 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1215_
timestamp 0
transform 1 0 3790 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1216_
timestamp 0
transform 1 0 3910 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1217_
timestamp 0
transform -1 0 4790 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1218_
timestamp 0
transform 1 0 4510 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1219_
timestamp 0
transform 1 0 3310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1220_
timestamp 0
transform 1 0 5150 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1221_
timestamp 0
transform 1 0 5310 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1222_
timestamp 0
transform 1 0 2050 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1223_
timestamp 0
transform 1 0 2910 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1224_
timestamp 0
transform -1 0 2350 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1225_
timestamp 0
transform 1 0 2090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1226_
timestamp 0
transform 1 0 1650 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1227_
timestamp 0
transform -1 0 1830 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1228_
timestamp 0
transform 1 0 2650 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1229_
timestamp 0
transform 1 0 2810 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1230_
timestamp 0
transform 1 0 2270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1231_
timestamp 0
transform -1 0 2490 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1232_
timestamp 0
transform -1 0 2650 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1233_
timestamp 0
transform 1 0 2970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1234_
timestamp 0
transform 1 0 4050 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1235_
timestamp 0
transform -1 0 3810 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1236_
timestamp 0
transform 1 0 3630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1237_
timestamp 0
transform 1 0 2810 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1238_
timestamp 0
transform 1 0 2410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1239_
timestamp 0
transform -1 0 3450 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1240_
timestamp 0
transform 1 0 3130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1241_
timestamp 0
transform 1 0 3110 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1242_
timestamp 0
transform 1 0 3070 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1243_
timestamp 0
transform -1 0 3490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1244_
timestamp 0
transform 1 0 3290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1245_
timestamp 0
transform 1 0 3430 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1246_
timestamp 0
transform 1 0 4930 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1247_
timestamp 0
transform -1 0 5650 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1248_
timestamp 0
transform 1 0 5470 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1249_
timestamp 0
transform -1 0 3610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1250_
timestamp 0
transform 1 0 3150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1251_
timestamp 0
transform -1 0 2830 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1252_
timestamp 0
transform -1 0 3030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1253_
timestamp 0
transform -1 0 1090 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1254_
timestamp 0
transform 1 0 2970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1255_
timestamp 0
transform 1 0 3270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1256_
timestamp 0
transform 1 0 3150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1257_
timestamp 0
transform 1 0 3310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1258_
timestamp 0
transform 1 0 3530 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1259_
timestamp 0
transform -1 0 5770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1260_
timestamp 0
transform -1 0 5330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1261_
timestamp 0
transform -1 0 5490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1262_
timestamp 0
transform 1 0 5870 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1263_
timestamp 0
transform -1 0 5750 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1264_
timestamp 0
transform -1 0 5650 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1265_
timestamp 0
transform -1 0 5670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1266_
timestamp 0
transform 1 0 5330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1267_
timestamp 0
transform -1 0 5810 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1268_
timestamp 0
transform 1 0 5790 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1269_
timestamp 0
transform -1 0 5510 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1270_
timestamp 0
transform 1 0 5090 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1271_
timestamp 0
transform 1 0 5710 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1272_
timestamp 0
transform -1 0 5470 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1273_
timestamp 0
transform -1 0 5310 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1274_
timestamp 0
transform -1 0 5010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1275_
timestamp 0
transform -1 0 4790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1276_
timestamp 0
transform 1 0 4590 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1277_
timestamp 0
transform 1 0 5650 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1278_
timestamp 0
transform -1 0 5590 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1279_
timestamp 0
transform -1 0 5430 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1280_
timestamp 0
transform 1 0 5230 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1281_
timestamp 0
transform -1 0 4810 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1282_
timestamp 0
transform -1 0 4650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1283_
timestamp 0
transform 1 0 4670 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1284_
timestamp 0
transform 1 0 5310 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1285_
timestamp 0
transform -1 0 4830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1286_
timestamp 0
transform -1 0 4990 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1287_
timestamp 0
transform -1 0 4490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1288_
timestamp 0
transform 1 0 4230 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1289_
timestamp 0
transform 1 0 4350 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1290_
timestamp 0
transform -1 0 5150 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1291_
timestamp 0
transform -1 0 4530 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1292_
timestamp 0
transform -1 0 4370 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1293_
timestamp 0
transform 1 0 4190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1294_
timestamp 0
transform -1 0 3610 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1295_
timestamp 0
transform -1 0 4350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1296_
timestamp 0
transform 1 0 4030 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1297_
timestamp 0
transform -1 0 3770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1298_
timestamp 0
transform 1 0 3870 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1299_
timestamp 0
transform -1 0 4410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1300_
timestamp 0
transform 1 0 4230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1301_
timestamp 0
transform 1 0 3890 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1302_
timestamp 0
transform 1 0 4890 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1303_
timestamp 0
transform -1 0 5150 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1304_
timestamp 0
transform 1 0 2630 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1305_
timestamp 0
transform -1 0 1970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1306_
timestamp 0
transform 1 0 1570 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1307_
timestamp 0
transform -1 0 1730 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1308_
timestamp 0
transform -1 0 1730 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1309_
timestamp 0
transform 1 0 2010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1310_
timestamp 0
transform 1 0 2170 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1311_
timestamp 0
transform 1 0 1890 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1312_
timestamp 0
transform -1 0 2210 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1313_
timestamp 0
transform 1 0 2030 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1314_
timestamp 0
transform 1 0 2470 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1315_
timestamp 0
transform 1 0 2710 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1316_
timestamp 0
transform 1 0 2850 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1317_
timestamp 0
transform 1 0 2710 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1318_
timestamp 0
transform 1 0 2290 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1319_
timestamp 0
transform -1 0 1790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1320_
timestamp 0
transform -1 0 3390 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1321_
timestamp 0
transform -1 0 3230 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1322_
timestamp 0
transform 1 0 2370 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1323_
timestamp 0
transform 1 0 2870 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1324_
timestamp 0
transform 1 0 2690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1325_
timestamp 0
transform 1 0 2530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1326_
timestamp 0
transform 1 0 2550 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1327_
timestamp 0
transform 1 0 3030 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1328_
timestamp 0
transform -1 0 3610 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1329_
timestamp 0
transform -1 0 5630 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1330_
timestamp 0
transform -1 0 5450 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1331_
timestamp 0
transform 1 0 2350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1332_
timestamp 0
transform 1 0 2190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1333_
timestamp 0
transform 1 0 2550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1334_
timestamp 0
transform -1 0 3130 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1335_
timestamp 0
transform -1 0 2570 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1336_
timestamp 0
transform -1 0 2390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1337_
timestamp 0
transform 1 0 2390 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1338_
timestamp 0
transform 1 0 3250 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1339_
timestamp 0
transform -1 0 4170 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1340_
timestamp 0
transform 1 0 4050 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1341_
timestamp 0
transform 1 0 3410 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1342_
timestamp 0
transform 1 0 4350 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1343_
timestamp 0
transform 1 0 3390 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1344_
timestamp 0
transform -1 0 5290 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1345_
timestamp 0
transform 1 0 4490 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1346_
timestamp 0
transform -1 0 4210 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1347_
timestamp 0
transform 1 0 4970 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1348_
timestamp 0
transform -1 0 5350 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1349_
timestamp 0
transform 1 0 3730 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1350_
timestamp 0
transform -1 0 3910 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1351_
timestamp 0
transform 1 0 4650 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1352_
timestamp 0
transform -1 0 5190 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1353_
timestamp 0
transform 1 0 4330 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1354_
timestamp 0
transform -1 0 4830 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1355_
timestamp 0
transform -1 0 4610 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1356_
timestamp 0
transform -1 0 4450 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1357_
timestamp 0
transform -1 0 5170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1358_
timestamp 0
transform -1 0 4670 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1359_
timestamp 0
transform 1 0 4710 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1360_
timestamp 0
transform -1 0 5030 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1361_
timestamp 0
transform -1 0 4790 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1362_
timestamp 0
transform 1 0 4290 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1363_
timestamp 0
transform 1 0 4030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1364_
timestamp 0
transform -1 0 3930 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1365_
timestamp 0
transform -1 0 4430 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1366_
timestamp 0
transform -1 0 4270 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1367_
timestamp 0
transform 1 0 2830 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1368_
timestamp 0
transform 1 0 3310 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1369_
timestamp 0
transform 1 0 4010 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1370_
timestamp 0
transform -1 0 3870 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1371_
timestamp 0
transform 1 0 2190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1372_
timestamp 0
transform -1 0 1610 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1373_
timestamp 0
transform -1 0 1510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1374_
timestamp 0
transform 1 0 1150 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1375_
timestamp 0
transform 1 0 1430 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1376_
timestamp 0
transform 1 0 1270 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1377_
timestamp 0
transform -1 0 1230 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1378_
timestamp 0
transform -1 0 1870 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1379_
timestamp 0
transform 1 0 1450 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1380_
timestamp 0
transform 1 0 1310 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1381_
timestamp 0
transform 1 0 1370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1382_
timestamp 0
transform 1 0 1510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1383_
timestamp 0
transform 1 0 1750 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1384_
timestamp 0
transform -1 0 2110 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1385_
timestamp 0
transform -1 0 1770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1386_
timestamp 0
transform -1 0 1610 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1387_
timestamp 0
transform -1 0 1170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1388_
timestamp 0
transform 1 0 1590 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1389_
timestamp 0
transform -1 0 1910 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1390_
timestamp 0
transform -1 0 2270 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1391_
timestamp 0
transform 1 0 1910 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1392_
timestamp 0
transform 1 0 1430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1393_
timestamp 0
transform -1 0 1890 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1394_
timestamp 0
transform 1 0 2610 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1395_
timestamp 0
transform 1 0 2970 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1396_
timestamp 0
transform -1 0 2810 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1397_
timestamp 0
transform -1 0 2670 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1398_
timestamp 0
transform -1 0 2430 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1399_
timestamp 0
transform 1 0 2230 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1400_
timestamp 0
transform 1 0 2030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1401_
timestamp 0
transform 1 0 2050 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1402_
timestamp 0
transform 1 0 2530 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1403_
timestamp 0
transform -1 0 2990 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1404_
timestamp 0
transform -1 0 3290 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1405_
timestamp 0
transform -1 0 3730 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1406_
timestamp 0
transform -1 0 3570 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1407_
timestamp 0
transform 1 0 3010 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1408_
timestamp 0
transform 1 0 3650 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1409_
timestamp 0
transform 1 0 2850 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1410_
timestamp 0
transform -1 0 3130 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1411_
timestamp 0
transform 1 0 3330 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1412_
timestamp 0
transform 1 0 3810 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1413_
timestamp 0
transform 1 0 4490 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1414_
timestamp 0
transform -1 0 4550 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1415_
timestamp 0
transform -1 0 3190 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1416_
timestamp 0
transform 1 0 3490 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1417_
timestamp 0
transform -1 0 3990 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1418_
timestamp 0
transform 1 0 3630 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1419_
timestamp 0
transform 1 0 3590 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1420_
timestamp 0
transform 1 0 4090 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1421_
timestamp 0
transform 1 0 3730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1422_
timestamp 0
transform -1 0 3450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1423_
timestamp 0
transform -1 0 4150 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1424_
timestamp 0
transform -1 0 3470 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1425_
timestamp 0
transform 1 0 3770 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1426_
timestamp 0
transform 1 0 2970 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1427_
timestamp 0
transform -1 0 2690 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1428_
timestamp 0
transform 1 0 1730 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1429_
timestamp 0
transform -1 0 1230 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1430_
timestamp 0
transform -1 0 2510 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1431_
timestamp 0
transform 1 0 1430 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1432_
timestamp 0
transform 1 0 690 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1433_
timestamp 0
transform -1 0 1330 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1434_
timestamp 0
transform 1 0 1150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1435_
timestamp 0
transform 1 0 1110 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1436_
timestamp 0
transform 1 0 1010 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1437_
timestamp 0
transform 1 0 970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1438_
timestamp 0
transform -1 0 1130 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1439_
timestamp 0
transform -1 0 830 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1440_
timestamp 0
transform 1 0 1270 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1441_
timestamp 0
transform -1 0 530 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1442_
timestamp 0
transform 1 0 70 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1443_
timestamp 0
transform -1 0 2490 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1444_
timestamp 0
transform -1 0 230 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1445_
timestamp 0
transform 1 0 510 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1446_
timestamp 0
transform -1 0 390 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1447_
timestamp 0
transform -1 0 90 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1448_
timestamp 0
transform 1 0 210 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1449_
timestamp 0
transform -1 0 670 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1450_
timestamp 0
transform -1 0 670 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1451_
timestamp 0
transform -1 0 950 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1452_
timestamp 0
transform -1 0 950 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1453_
timestamp 0
transform -1 0 810 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1454_
timestamp 0
transform 1 0 1050 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1455_
timestamp 0
transform 1 0 1090 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1456_
timestamp 0
transform 1 0 1250 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1457_
timestamp 0
transform -1 0 2110 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1458_
timestamp 0
transform -1 0 2710 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1459_
timestamp 0
transform -1 0 2830 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1460_
timestamp 0
transform -1 0 1930 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1461_
timestamp 0
transform 1 0 1830 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1462_
timestamp 0
transform -1 0 1990 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1463_
timestamp 0
transform 1 0 1790 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1464_
timestamp 0
transform -1 0 1650 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1465_
timestamp 0
transform 1 0 1330 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1466_
timestamp 0
transform 1 0 830 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1467_
timestamp 0
transform -1 0 630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1468_
timestamp 0
transform 1 0 970 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1469_
timestamp 0
transform 1 0 670 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1470_
timestamp 0
transform -1 0 1290 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1471_
timestamp 0
transform 1 0 810 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1472_
timestamp 0
transform -1 0 90 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1473_
timestamp 0
transform -1 0 90 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1474_
timestamp 0
transform -1 0 90 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1475_
timestamp 0
transform 1 0 570 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1476_
timestamp 0
transform 1 0 250 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1477_
timestamp 0
transform 1 0 690 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1478_
timestamp 0
transform 1 0 350 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1479_
timestamp 0
transform 1 0 270 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1480_
timestamp 0
transform -1 0 430 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1481_
timestamp 0
transform 1 0 410 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1482_
timestamp 0
transform -1 0 870 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1483_
timestamp 0
transform -1 0 1450 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1484_
timestamp 0
transform -1 0 1530 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1485_
timestamp 0
transform -1 0 1370 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1486_
timestamp 0
transform -1 0 1690 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1487_
timestamp 0
transform -1 0 1470 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1488_
timestamp 0
transform 1 0 1490 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1489_
timestamp 0
transform 1 0 1270 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1490_
timestamp 0
transform 1 0 550 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1491_
timestamp 0
transform -1 0 850 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1492_
timestamp 0
transform 1 0 670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1493_
timestamp 0
transform -1 0 550 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1494_
timestamp 0
transform 1 0 250 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1495_
timestamp 0
transform 1 0 370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1496_
timestamp 0
transform 1 0 770 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1497_
timestamp 0
transform 1 0 270 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1498_
timestamp 0
transform 1 0 70 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1499_
timestamp 0
transform -1 0 290 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1500_
timestamp 0
transform 1 0 910 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1501_
timestamp 0
transform -1 0 1010 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1502_
timestamp 0
transform -1 0 990 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1503_
timestamp 0
transform -1 0 970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1504_
timestamp 0
transform 1 0 670 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1505_
timestamp 0
transform -1 0 810 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1506_
timestamp 0
transform -1 0 630 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1507_
timestamp 0
transform 1 0 70 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1508_
timestamp 0
transform -1 0 90 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1509_
timestamp 0
transform -1 0 430 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1510_
timestamp 0
transform 1 0 330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1511_
timestamp 0
transform 1 0 3110 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1512_
timestamp 0
transform -1 0 1590 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1513_
timestamp 0
transform -1 0 1210 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1514_
timestamp 0
transform -1 0 1130 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1515_
timestamp 0
transform -1 0 230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1516_
timestamp 0
transform -1 0 630 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1517_
timestamp 0
transform -1 0 490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1518_
timestamp 0
transform 1 0 1330 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1519_
timestamp 0
transform 1 0 2230 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1560_
timestamp 0
transform -1 0 90 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1561_
timestamp 0
transform -1 0 230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1562_
timestamp 0
transform -1 0 90 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1563_
timestamp 0
transform -1 0 90 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1564_
timestamp 0
transform -1 0 370 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1565_
timestamp 0
transform 1 0 3910 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1566_
timestamp 0
transform -1 0 1030 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1567_
timestamp 0
transform -1 0 90 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1568_
timestamp 0
transform -1 0 90 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1569_
timestamp 0
transform -1 0 90 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1570_
timestamp 0
transform -1 0 3730 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1571_
timestamp 0
transform 1 0 5130 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1572_
timestamp 0
transform -1 0 2370 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1573_
timestamp 0
transform 1 0 2210 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1574_
timestamp 0
transform -1 0 90 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1575_
timestamp 0
transform -1 0 250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1576_
timestamp 0
transform -1 0 90 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1577_
timestamp 0
transform -1 0 390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1578_
timestamp 0
transform 1 0 1630 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1579_
timestamp 0
transform 1 0 2250 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1580_
timestamp 0
transform -1 0 2770 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1581_
timestamp 0
transform -1 0 3110 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1582_
timestamp 0
transform -1 0 90 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1583_
timestamp 0
transform -1 0 3290 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert6
timestamp 0
transform 1 0 5110 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert7
timestamp 0
transform -1 0 3150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert8
timestamp 0
transform -1 0 3150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert9
timestamp 0
transform -1 0 5870 0 -1 270
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert10
timestamp 0
transform 1 0 1670 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert11
timestamp 0
transform 1 0 1790 0 1 4430
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert12
timestamp 0
transform 1 0 1550 0 1 3390
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert13
timestamp 0
transform -1 0 90 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert14
timestamp 0
transform -1 0 2790 0 1 2350
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert15
timestamp 0
transform -1 0 4090 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert16
timestamp 0
transform 1 0 4290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert17
timestamp 0
transform 1 0 4210 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert0
timestamp 0
transform 1 0 1470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert1
timestamp 0
transform -1 0 1310 0 1 3390
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert2
timestamp 0
transform -1 0 770 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert3
timestamp 0
transform -1 0 1110 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert4
timestamp 0
transform -1 0 1090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert5
timestamp 0
transform 1 0 3050 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__760_
timestamp 0
transform 1 0 750 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__765_
timestamp 0
transform -1 0 490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__769_
timestamp 0
transform 1 0 730 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__774_
timestamp 0
transform 1 0 710 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__778_
timestamp 0
transform 1 0 410 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__783_
timestamp 0
transform 1 0 650 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__788_
timestamp 0
transform 1 0 1630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__792_
timestamp 0
transform -1 0 1470 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__797_
timestamp 0
transform 1 0 1150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__801_
timestamp 0
transform 1 0 2350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__806_
timestamp 0
transform -1 0 810 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__811_
timestamp 0
transform 1 0 210 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__815_
timestamp 0
transform 1 0 410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__820_
timestamp 0
transform -1 0 230 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__824_
timestamp 0
transform 1 0 690 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__829_
timestamp 0
transform -1 0 1130 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__834_
timestamp 0
transform 1 0 2130 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__838_
timestamp 0
transform -1 0 2450 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__843_
timestamp 0
transform -1 0 1870 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__848_
timestamp 0
transform 1 0 830 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__852_
timestamp 0
transform 1 0 2390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__857_
timestamp 0
transform -1 0 1970 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__861_
timestamp 0
transform 1 0 1750 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__866_
timestamp 0
transform -1 0 1810 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__871_
timestamp 0
transform 1 0 1470 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__875_
timestamp 0
transform 1 0 2090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__880_
timestamp 0
transform -1 0 1710 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__884_
timestamp 0
transform -1 0 1970 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__889_
timestamp 0
transform 1 0 2750 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__894_
timestamp 0
transform 1 0 2990 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__898_
timestamp 0
transform 1 0 2690 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__903_
timestamp 0
transform 1 0 2670 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__907_
timestamp 0
transform -1 0 4590 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__912_
timestamp 0
transform 1 0 4390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__917_
timestamp 0
transform -1 0 5010 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__921_
timestamp 0
transform -1 0 4070 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__926_
timestamp 0
transform -1 0 3730 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__930_
timestamp 0
transform 1 0 2410 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__935_
timestamp 0
transform -1 0 2770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__940_
timestamp 0
transform 1 0 2330 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__944_
timestamp 0
transform -1 0 2870 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__949_
timestamp 0
transform 1 0 1370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__953_
timestamp 0
transform 1 0 4910 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__958_
timestamp 0
transform 1 0 3370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__963_
timestamp 0
transform 1 0 4010 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__967_
timestamp 0
transform 1 0 5290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__972_
timestamp 0
transform -1 0 5430 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__976_
timestamp 0
transform -1 0 5730 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__981_
timestamp 0
transform -1 0 5950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__986_
timestamp 0
transform -1 0 5710 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__990_
timestamp 0
transform 1 0 4110 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__995_
timestamp 0
transform -1 0 4950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__999_
timestamp 0
transform -1 0 5130 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1000_
timestamp 0
transform -1 0 4870 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1005_
timestamp 0
transform -1 0 5030 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1009_
timestamp 0
transform -1 0 4690 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1014_
timestamp 0
transform -1 0 4410 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1018_
timestamp 0
transform -1 0 3750 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1023_
timestamp 0
transform 1 0 4170 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1028_
timestamp 0
transform -1 0 2150 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1032_
timestamp 0
transform -1 0 1910 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1037_
timestamp 0
transform 1 0 2070 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1041_
timestamp 0
transform 1 0 4510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1046_
timestamp 0
transform 1 0 2530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1051_
timestamp 0
transform 1 0 3070 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1055_
timestamp 0
transform 1 0 5870 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1060_
timestamp 0
transform -1 0 4150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1064_
timestamp 0
transform 1 0 4010 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1069_
timestamp 0
transform 1 0 5610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1074_
timestamp 0
transform -1 0 5670 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1078_
timestamp 0
transform 1 0 5790 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1083_
timestamp 0
transform 1 0 5870 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1087_
timestamp 0
transform 1 0 5270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1092_
timestamp 0
transform 1 0 5770 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1097_
timestamp 0
transform 1 0 4910 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1101_
timestamp 0
transform -1 0 5630 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1106_
timestamp 0
transform 1 0 5090 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1110_
timestamp 0
transform -1 0 5030 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1115_
timestamp 0
transform -1 0 4690 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1120_
timestamp 0
transform -1 0 4030 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1124_
timestamp 0
transform 1 0 4670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1129_
timestamp 0
transform 1 0 3010 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1133_
timestamp 0
transform 1 0 2070 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1138_
timestamp 0
transform 1 0 2830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1143_
timestamp 0
transform -1 0 4150 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1147_
timestamp 0
transform -1 0 4470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1152_
timestamp 0
transform 1 0 3190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1157_
timestamp 0
transform -1 0 5390 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1161_
timestamp 0
transform 1 0 2950 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1166_
timestamp 0
transform 1 0 4230 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1170_
timestamp 0
transform 1 0 4870 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1175_
timestamp 0
transform 1 0 5670 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1180_
timestamp 0
transform 1 0 5790 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1184_
timestamp 0
transform 1 0 4970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1189_
timestamp 0
transform 1 0 5170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1193_
timestamp 0
transform 1 0 3850 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1198_
timestamp 0
transform -1 0 4830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1203_
timestamp 0
transform -1 0 4290 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1207_
timestamp 0
transform 1 0 3910 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1212_
timestamp 0
transform -1 0 4110 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1216_
timestamp 0
transform 1 0 3930 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1221_
timestamp 0
transform 1 0 5330 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1226_
timestamp 0
transform 1 0 1670 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1230_
timestamp 0
transform 1 0 2290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1235_
timestamp 0
transform -1 0 3830 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1239_
timestamp 0
transform -1 0 3470 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1244_
timestamp 0
transform 1 0 3310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1249_
timestamp 0
transform -1 0 3630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1253_
timestamp 0
transform -1 0 1110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1258_
timestamp 0
transform 1 0 3550 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1262_
timestamp 0
transform 1 0 5890 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1267_
timestamp 0
transform -1 0 5830 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1272_
timestamp 0
transform -1 0 5490 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1276_
timestamp 0
transform 1 0 4610 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1281_
timestamp 0
transform -1 0 4830 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1285_
timestamp 0
transform -1 0 4850 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1290_
timestamp 0
transform -1 0 5170 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1295_
timestamp 0
transform -1 0 4370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1299_
timestamp 0
transform -1 0 4430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1304_
timestamp 0
transform 1 0 2650 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1309_
timestamp 0
transform 1 0 2030 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1313_
timestamp 0
transform 1 0 2050 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1318_
timestamp 0
transform 1 0 2310 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1322_
timestamp 0
transform 1 0 2390 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1327_
timestamp 0
transform 1 0 3050 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1332_
timestamp 0
transform 1 0 2210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1336_
timestamp 0
transform -1 0 2410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1341_
timestamp 0
transform 1 0 3430 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1345_
timestamp 0
transform 1 0 4510 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1350_
timestamp 0
transform -1 0 3930 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1355_
timestamp 0
transform -1 0 4630 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1359_
timestamp 0
transform 1 0 4730 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1364_
timestamp 0
transform -1 0 3950 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1368_
timestamp 0
transform 1 0 3330 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1373_
timestamp 0
transform -1 0 1530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1378_
timestamp 0
transform -1 0 1890 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1382_
timestamp 0
transform 1 0 1530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1387_
timestamp 0
transform -1 0 1190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1391_
timestamp 0
transform 1 0 1930 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1396_
timestamp 0
transform -1 0 2830 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1401_
timestamp 0
transform 1 0 2070 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1405_
timestamp 0
transform -1 0 3750 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1410_
timestamp 0
transform -1 0 3150 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1414_
timestamp 0
transform -1 0 4570 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1419_
timestamp 0
transform 1 0 3610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1424_
timestamp 0
transform -1 0 3490 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1428_
timestamp 0
transform 1 0 1750 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1433_
timestamp 0
transform -1 0 1350 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1437_
timestamp 0
transform 1 0 990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1442_
timestamp 0
transform 1 0 90 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1447_
timestamp 0
transform -1 0 110 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1451_
timestamp 0
transform -1 0 970 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1456_
timestamp 0
transform 1 0 1270 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1460_
timestamp 0
transform -1 0 1950 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1465_
timestamp 0
transform 1 0 1350 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1470_
timestamp 0
transform -1 0 1310 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1474_
timestamp 0
transform -1 0 110 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1479_
timestamp 0
transform 1 0 290 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1484_
timestamp 0
transform -1 0 1550 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1488_
timestamp 0
transform 1 0 1510 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1493_
timestamp 0
transform -1 0 570 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1497_
timestamp 0
transform 1 0 290 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1502_
timestamp 0
transform -1 0 1010 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1507_
timestamp 0
transform 1 0 90 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1511_
timestamp 0
transform 1 0 3130 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1516_
timestamp 0
transform -1 0 650 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1560_
timestamp 0
transform -1 0 110 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1565_
timestamp 0
transform 1 0 3930 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1570_
timestamp 0
transform -1 0 3750 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1574_
timestamp 0
transform -1 0 110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1579_
timestamp 0
transform 1 0 2270 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1583_
timestamp 0
transform -1 0 3310 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert8
timestamp 0
transform -1 0 3170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert13
timestamp 0
transform -1 0 110 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert17
timestamp 0
transform 1 0 4230 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4_CLKBUF1_insert4
timestamp 0
transform -1 0 1110 0 -1 3390
box -6 -8 26 268
<< labels >>
flabel metal1 s 6003 2 6063 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -63 2 -3 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal3 s -24 2556 -16 2564 7 FreeSans 16 0 0 0 Cin[7]
port 2 nsew
flabel metal3 s -24 2476 -16 2484 7 FreeSans 16 0 0 0 Cin[6]
port 3 nsew
flabel metal3 s -24 2956 -16 2964 7 FreeSans 16 0 0 0 Cin[5]
port 4 nsew
flabel metal2 s 2217 -23 2223 -17 7 FreeSans 16 270 0 0 Cin[4]
port 5 nsew
flabel metal3 s 6036 3516 6044 3524 3 FreeSans 16 0 0 0 Cin[3]
port 6 nsew
flabel metal2 s 2297 6037 2303 6043 3 FreeSans 16 90 0 0 Cin[2]
port 7 nsew
flabel metal3 s 6036 1956 6044 1964 3 FreeSans 16 0 0 0 Cin[1]
port 8 nsew
flabel metal3 s 6036 176 6044 184 3 FreeSans 16 0 0 0 Cin[0]
port 9 nsew
flabel metal3 s 6036 2036 6044 2044 3 FreeSans 16 0 0 0 Xin[7]
port 10 nsew
flabel metal2 s 5237 6037 5243 6043 3 FreeSans 16 90 0 0 Xin[6]
port 11 nsew
flabel metal2 s 4097 6037 4103 6043 3 FreeSans 16 90 0 0 Xin[5]
port 12 nsew
flabel metal2 s 2637 6037 2643 6043 3 FreeSans 16 90 0 0 Xin[4]
port 13 nsew
flabel metal2 s 137 6037 143 6043 3 FreeSans 16 90 0 0 Xin[3]
port 14 nsew
flabel metal3 s -24 4516 -16 4524 7 FreeSans 16 0 0 0 Xin[2]
port 15 nsew
flabel metal3 s -24 4096 -16 4104 7 FreeSans 16 0 0 0 Xin[1]
port 16 nsew
flabel metal3 s -24 3056 -16 3064 7 FreeSans 16 0 0 0 Xin[0]
port 17 nsew
flabel metal3 s -24 2776 -16 2784 7 FreeSans 16 0 0 0 Xout[7]
port 18 nsew
flabel metal2 s 1057 6037 1063 6043 3 FreeSans 16 90 0 0 Xout[6]
port 19 nsew
flabel metal2 s 3977 6037 3983 6043 3 FreeSans 16 90 0 0 Xout[5]
port 20 nsew
flabel metal3 s -24 2816 -16 2824 7 FreeSans 16 0 0 0 Xout[4]
port 21 nsew
flabel metal3 s -24 3776 -16 3784 7 FreeSans 16 0 0 0 Xout[3]
port 22 nsew
flabel metal3 s -24 4816 -16 4824 7 FreeSans 16 0 0 0 Xout[2]
port 23 nsew
flabel metal3 s -24 2736 -16 2744 7 FreeSans 16 0 0 0 Xout[1]
port 24 nsew
flabel metal3 s -24 2996 -16 3004 7 FreeSans 16 0 0 0 Xout[0]
port 25 nsew
flabel metal3 s -24 1436 -16 1444 7 FreeSans 16 0 0 0 Yin[15]
port 26 nsew
flabel metal3 s -24 1696 -16 1704 7 FreeSans 16 0 0 0 Yin[14]
port 27 nsew
flabel metal3 s -24 916 -16 924 7 FreeSans 16 0 0 0 Yin[13]
port 28 nsew
flabel metal3 s -24 136 -16 144 7 FreeSans 16 0 0 0 Yin[12]
port 29 nsew
flabel metal2 s 2657 -23 2663 -17 7 FreeSans 16 270 0 0 Yin[11]
port 30 nsew
flabel metal2 s 3117 -23 3123 -17 7 FreeSans 16 270 0 0 Yin[10]
port 31 nsew
flabel metal3 s 6036 1176 6044 1184 3 FreeSans 16 0 0 0 Yin[9]
port 32 nsew
flabel metal3 s 6036 1996 6044 2004 3 FreeSans 16 0 0 0 Yin[8]
port 33 nsew
flabel metal3 s 6036 2216 6044 2224 3 FreeSans 16 0 0 0 Yin[7]
port 34 nsew
flabel metal3 s 6036 5556 6044 5564 3 FreeSans 16 0 0 0 Yin[6]
port 35 nsew
flabel metal2 s 4597 6037 4603 6043 3 FreeSans 16 90 0 0 Yin[5]
port 36 nsew
flabel metal2 s 2597 6037 2603 6043 3 FreeSans 16 90 0 0 Yin[4]
port 37 nsew
flabel metal3 s -24 5596 -16 5604 7 FreeSans 16 0 0 0 Yin[3]
port 38 nsew
flabel metal3 s -24 4556 -16 4564 7 FreeSans 16 0 0 0 Yin[2]
port 39 nsew
flabel metal3 s -24 3256 -16 3264 7 FreeSans 16 0 0 0 Yin[1]
port 40 nsew
flabel metal3 s -24 3996 -16 4004 7 FreeSans 16 0 0 0 Yin[0]
port 41 nsew
flabel metal3 s -24 2256 -16 2264 7 FreeSans 16 0 0 0 Yout[15]
port 42 nsew
flabel metal3 s -24 2216 -16 2224 7 FreeSans 16 0 0 0 Yout[14]
port 43 nsew
flabel metal2 s 2257 -23 2263 -17 7 FreeSans 16 270 0 0 Yout[13]
port 44 nsew
flabel metal2 s 2397 -23 2403 -17 7 FreeSans 16 270 0 0 Yout[12]
port 45 nsew
flabel metal2 s 5177 -23 5183 -17 7 FreeSans 16 270 0 0 Yout[11]
port 46 nsew
flabel metal2 s 3777 -23 3783 -17 7 FreeSans 16 270 0 0 Yout[10]
port 47 nsew
flabel metal2 s 3337 6037 3343 6043 3 FreeSans 16 90 0 0 Yout[9]
port 48 nsew
flabel metal3 s -24 2516 -16 2524 7 FreeSans 16 0 0 0 Yout[8]
port 49 nsew
flabel metal2 s 3137 6037 3143 6043 3 FreeSans 16 90 0 0 Yout[7]
port 50 nsew
flabel metal2 s 2797 6037 2803 6043 3 FreeSans 16 90 0 0 Yout[6]
port 51 nsew
flabel metal2 s 2337 6037 2343 6043 3 FreeSans 16 90 0 0 Yout[5]
port 52 nsew
flabel metal2 s 1677 6037 1683 6043 3 FreeSans 16 90 0 0 Yout[4]
port 53 nsew
flabel metal2 s 417 6037 423 6043 3 FreeSans 16 90 0 0 Yout[3]
port 54 nsew
flabel metal3 s -24 3296 -16 3304 7 FreeSans 16 0 0 0 Yout[2]
port 55 nsew
flabel metal3 s -24 3516 -16 3524 7 FreeSans 16 0 0 0 Yout[1]
port 56 nsew
flabel metal3 s -24 4036 -16 4044 7 FreeSans 16 0 0 0 Yout[0]
port 57 nsew
flabel metal2 s 877 6037 883 6043 3 FreeSans 16 90 0 0 clk
port 58 nsew
<< properties >>
string FIXED_BBOX -40 -40 6040 6040
<< end >>

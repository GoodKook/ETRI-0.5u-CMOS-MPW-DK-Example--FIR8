/* Verilog module written by vlog2Verilog (qflow) */
/* With explicit power connections */

module fir_pe(
    inout vdd,
    inout gnd,
    input [7:0] Cin,
    input Rdy,
    output Vld,
    input [3:0] Xin,
    output [3:0] Xout,
    input [3:0] Yin,
    output [3:0] Yout,
    input clk
);

wire [15:0] y ;
wire _588_ ;
wire _168_ ;
wire _800_ ;
wire _60_ ;
wire _397_ ;
wire _703_ ;
wire _19_ ;
wire _512_ ;
wire [4:0] LoadCtl ;
wire _741_ ;
wire _321_ ;
wire _57_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _835_ ;
wire _415_ ;
wire _95_ ;
wire _148__bF$buf0 ;
wire _148__bF$buf1 ;
wire _148__bF$buf2 ;
wire _148__bF$buf3 ;
wire _148__bF$buf4 ;
wire _644_ ;
wire _224_ ;
wire _873_ ;
wire _453_ ;
wire _509_ ;
wire _682_ ;
wire _262_ ;
wire _738_ ;
wire _318_ ;
wire _491_ ;
wire _547_ ;
wire _127_ ;
wire _776_ ;
wire _356_ ;
wire _585_ ;
wire _165_ ;
wire _394_ ;
wire _679_ ;
wire _259_ ;
wire _488_ ;
wire _700_ ;
wire _297_ ;
wire _16_ ;
wire _54_ ;
wire _603_ ;
wire _832_ ;
wire _412_ ;
wire _92_ ;
wire _641_ ;
wire _221_ ;
wire _870_ ;
wire _450_ ;
wire _506_ ;
wire _735_ ;
wire _315_ ;
wire _544_ ;
wire _124_ ;
wire _773_ ;
wire _353_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _582_ ;
wire _162_ ;
wire _638_ ;
wire _218_ ;
wire _391_ ;
wire _867_ ;
wire _447_ ;
wire _676_ ;
wire _256_ ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire _388_ ;
wire _600_ ;
wire Rdy ;
wire _197_ ;
wire _7_ ;
wire _503_ ;
wire _732_ ;
wire _312_ ;
wire _48_ ;
wire _541_ ;
wire _121_ ;
wire _770_ ;
wire _350_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _635_ ;
wire _215_ ;
wire _864_ ;
wire _444_ ;
wire _673_ ;
wire _253_ ;
wire _729_ ;
wire _309_ ;
wire _482_ ;
wire _538_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _767_ ;
wire _347_ ;
wire _576_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire [3:0] XinHL ;
wire _899_ ;
wire _479_ ;
wire _288_ ;
wire _4_ ;
wire [3:0] _920_ ;
wire _500_ ;
wire _45_ ;
wire _823_ ;
wire _403_ ;
wire _83_ ;
wire _632_ ;
wire _212_ ;
wire _861_ ;
wire _441_ ;
wire _917_ ;
wire _670_ ;
wire _250_ ;
wire _726_ ;
wire _306_ ;
wire _535_ ;
wire _115_ ;
wire _764_ ;
wire _344_ ;
wire _573_ ;
wire _153_ ;
wire _629_ ;
wire _209_ ;
wire _382_ ;
wire _858_ ;
wire _438_ ;
wire _191_ ;
wire _667_ ;
wire _247_ ;
wire _896_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire _285_ ;
wire _1_ ;
wire _42_ ;
wire _799_ ;
wire _379_ ;
wire _188_ ;
wire _820_ ;
wire _400_ ;
wire _80_ ;
wire _914_ ;
wire _723_ ;
wire _303_ ;
wire _39_ ;
wire _532_ ;
wire _112_ ;
wire _761_ ;
wire _341_ ;
wire clk ;
wire _817_ ;
wire _77_ ;
wire _570_ ;
wire _150_ ;
wire _626_ ;
wire _206_ ;
wire _855_ ;
wire _435_ ;
wire _664_ ;
wire _244_ ;
wire _893_ ;
wire _473_ ;
wire _529_ ;
wire _109_ ;
wire _282_ ;
wire _758_ ;
wire _338_ ;
wire _567_ ;
wire _147_ ;
wire _796_ ;
wire _376_ ;
wire _185_ ;
wire _699_ ;
wire _279_ ;
wire _911_ ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire _814_ ;
wire _74_ ;
wire _623_ ;
wire _203_ ;
wire _852_ ;
wire _432_ ;
wire _908_ ;
wire _661_ ;
wire _241_ ;
wire _717_ ;
wire _890_ ;
wire _470_ ;
wire _526_ ;
wire _106_ ;
wire _755_ ;
wire _335_ ;
wire _564_ ;
wire _144_ ;
wire _793_ ;
wire _373_ ;
wire _849_ ;
wire _429_ ;
wire _182_ ;
wire LoadCtl_0_bF$buf0 ;
wire LoadCtl_0_bF$buf1 ;
wire LoadCtl_0_bF$buf2 ;
wire LoadCtl_0_bF$buf3 ;
wire LoadCtl_0_bF$buf4 ;
wire _658_ ;
wire _238_ ;
wire _887_ ;
wire _467_ ;
wire _696_ ;
wire _276_ ;
wire _33_ ;
wire _599_ ;
wire _179_ ;
wire _811_ ;
wire _71_ ;
wire _620_ ;
wire _200_ ;
wire _905_ ;
wire _714_ ;
wire _523_ ;
wire _103_ ;
wire _752_ ;
wire _332_ ;
wire _808_ ;
wire _68_ ;
wire _561_ ;
wire _141_ ;
wire _617_ ;
wire _790_ ;
wire _370_ ;
wire _846_ ;
wire _426_ ;
wire _655_ ;
wire _235_ ;
wire _884_ ;
wire _464_ ;
wire _693_ ;
wire _273_ ;
wire _749_ ;
wire _329_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _787_ ;
wire _367_ ;
wire _596_ ;
wire _176_ ;
wire _902_ ;
wire _499_ ;
wire _711_ ;
wire _27_ ;
wire _520_ ;
wire _100_ ;
wire _805_ ;
wire _65_ ;
wire _614_ ;
wire _843_ ;
wire _423_ ;
wire _652_ ;
wire _232_ ;
wire _708_ ;
wire _881_ ;
wire _461_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _746_ ;
wire _326_ ;
wire _555_ ;
wire _135_ ;
wire _784_ ;
wire _364_ ;
wire _593_ ;
wire _173_ ;
wire _649_ ;
wire _229_ ;
wire _878_ ;
wire _458_ ;
wire _687_ ;
wire _267_ ;
wire _496_ ;
wire _24_ ;
wire _802_ ;
wire _62_ ;
wire _399_ ;
wire _611_ ;
wire _840_ ;
wire _420_ ;
wire _705_ ;
wire [15:0] _y ;
wire _514_ ;
wire _743_ ;
wire _323_ ;
wire _59_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _781_ ;
wire _361_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _646_ ;
wire _226_ ;
wire _875_ ;
wire _455_ ;
wire _684_ ;
wire _264_ ;
wire _493_ ;
wire _549_ ;
wire _129_ ;
wire _21_ ;
wire _778_ ;
wire _358_ ;
wire _587_ ;
wire _167_ ;
wire _396_ ;
wire _702_ ;
wire _299_ ;
wire _18_ ;
wire _511_ ;
wire _740_ ;
wire _320_ ;
wire _56_ ;
wire _605_ ;
wire _834_ ;
wire _414_ ;
wire _94_ ;
wire _643_ ;
wire _223_ ;
wire _872_ ;
wire _452_ ;
wire _508_ ;
wire _681_ ;
wire _261_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _546_ ;
wire _126_ ;
wire _775_ ;
wire _355_ ;
wire _584_ ;
wire _164_ ;
wire _393_ ;
wire _869_ ;
wire _449_ ;
wire _678_ ;
wire _258_ ;
wire _487_ ;
wire _296_ ;
wire _15_ ;
wire _53_ ;
wire _602_ ;
wire _199_ ;
wire _831_ ;
wire _411_ ;
wire _91_ ;
wire _640_ ;
wire _220_ ;
wire _9_ ;
wire _505_ ;
wire _734_ ;
wire _314_ ;
wire _543_ ;
wire _123_ ;
wire _772_ ;
wire _352_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _581_ ;
wire _161_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _866_ ;
wire _446_ ;
wire [3:0] Yin ;
wire _675_ ;
wire _255_ ;
wire _484_ ;
wire _293_ ;
wire _12_ ;
wire _769_ ;
wire _349_ ;
wire _578_ ;
wire _158_ ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire _6_ ;
wire _502_ ;
wire _731_ ;
wire _311_ ;
wire _47_ ;
wire _540_ ;
wire _120_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire [3:0] Yin0 ;
wire [3:0] Yin1 ;
wire [3:0] Yin2 ;
wire [3:0] Yin3 ;
wire _634_ ;
wire _214_ ;
wire _863_ ;
wire _443_ ;
wire _919_ ;
wire _672_ ;
wire _252_ ;
wire _728_ ;
wire _308_ ;
wire _481_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _766_ ;
wire _346_ ;
wire _575_ ;
wire _155_ ;
wire _384_ ;
wire _193_ ;
wire _669_ ;
wire _249_ ;
wire _898_ ;
wire _478_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _822_ ;
wire _402_ ;
wire _82_ ;
wire _631_ ;
wire _211_ ;
wire _860_ ;
wire _440_ ;
wire _916_ ;
wire _725_ ;
wire _305_ ;
wire [3:0] XinH ;
wire _534_ ;
wire _114_ ;
wire _763_ ;
wire _343_ ;
wire _819_ ;
wire _79_ ;
wire _572_ ;
wire _152_ ;
wire _628_ ;
wire _208_ ;
wire _381_ ;
wire _857_ ;
wire _437_ ;
wire _190_ ;
wire _666_ ;
wire _246_ ;
wire _895_ ;
wire _475_ ;
wire _284_ ;
wire _0_ ;
wire _569_ ;
wire _149_ ;
wire _41_ ;
wire _798_ ;
wire _378_ ;
wire _187_ ;
wire [3:0] Yout ;
wire _913_ ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _531_ ;
wire _111_ ;
wire _760_ ;
wire _340_ ;
wire _816_ ;
wire _76_ ;
wire _625_ ;
wire _205_ ;
wire _854_ ;
wire _434_ ;
wire _663_ ;
wire _243_ ;
wire _719_ ;
wire _892_ ;
wire _472_ ;
wire _528_ ;
wire _108_ ;
wire _281_ ;
wire _757_ ;
wire _337_ ;
wire _566_ ;
wire _146_ ;
wire _795_ ;
wire _375_ ;
wire _184_ ;
wire _889_ ;
wire _469_ ;
wire _698_ ;
wire _278_ ;
wire _910_ ;
wire _35_ ;
wire [3:0] Xout ;
wire _813_ ;
wire _73_ ;
wire _622_ ;
wire _202_ ;
wire _851_ ;
wire _431_ ;
wire _907_ ;
wire _660_ ;
wire _240_ ;
wire _716_ ;
wire _525_ ;
wire _105_ ;
wire _754_ ;
wire _334_ ;
wire _563_ ;
wire _143_ ;
wire _619_ ;
wire _792_ ;
wire _372_ ;
wire _848_ ;
wire _428_ ;
wire _181_ ;
wire _657_ ;
wire _237_ ;
wire _886_ ;
wire _466_ ;
wire _695_ ;
wire _275_ ;
wire _32_ ;
wire _789_ ;
wire _369_ ;
wire _598_ ;
wire _178_ ;
wire _810_ ;
wire _70_ ;
wire LoadCtl_4_bF$buf0 ;
wire LoadCtl_4_bF$buf1 ;
wire LoadCtl_4_bF$buf2 ;
wire LoadCtl_4_bF$buf3 ;
wire LoadCtl_4_bF$buf4 ;
wire _904_ ;
wire _713_ ;
wire _29_ ;
wire _522_ ;
wire _102_ ;
wire _751_ ;
wire _331_ ;
wire _807_ ;
wire _67_ ;
wire _560_ ;
wire _140_ ;
wire _616_ ;
wire _845_ ;
wire _425_ ;
wire _654_ ;
wire _234_ ;
wire _883_ ;
wire _463_ ;
wire _519_ ;
wire _692_ ;
wire _272_ ;
wire _748_ ;
wire _328_ ;
wire _557_ ;
wire _137_ ;
wire _786_ ;
wire _366_ ;
wire _595_ ;
wire _175_ ;
wire _689_ ;
wire _269_ ;
wire _901_ ;
wire _498_ ;
wire _710_ ;
wire _26_ ;
wire Cin_0_bF$buf0 ;
wire Cin_0_bF$buf1 ;
wire Cin_0_bF$buf2 ;
wire Cin_0_bF$buf3 ;
wire _804_ ;
wire _64_ ;
wire _613_ ;
wire _842_ ;
wire _422_ ;
wire _651_ ;
wire _231_ ;
wire _707_ ;
wire _880_ ;
wire _460_ ;
wire _516_ ;
wire _745_ ;
wire _325_ ;
wire _554_ ;
wire _134_ ;
wire _783_ ;
wire _363_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _592_ ;
wire _172_ ;
wire Vld ;
wire _648_ ;
wire _228_ ;
wire _877_ ;
wire _457_ ;
wire _686_ ;
wire _266_ ;
wire _495_ ;
wire _23_ ;
wire _589_ ;
wire _169_ ;
wire _801_ ;
wire _61_ ;
wire _398_ ;
wire _610_ ;
wire _704_ ;
wire _513_ ;
wire _742_ ;
wire _322_ ;
wire _58_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _780_ ;
wire _360_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire [7:0] Cin ;
wire _645_ ;
wire _225_ ;
wire _874_ ;
wire _454_ ;
wire _683_ ;
wire _263_ ;
wire _739_ ;
wire _319_ ;
wire _492_ ;
wire _548_ ;
wire _128_ ;
wire _20_ ;
wire _777_ ;
wire _357_ ;
wire _586_ ;
wire _166_ ;
wire _395_ ;
wire _489_ ;
wire _701_ ;
wire _298_ ;
wire _17_ ;
wire _510_ ;
wire _55_ ;
wire _604_ ;
wire _833_ ;
wire _413_ ;
wire _93_ ;
wire _642_ ;
wire _222_ ;
wire _871_ ;
wire _451_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _736_ ;
wire _316_ ;
wire _545_ ;
wire _125_ ;
wire _774_ ;
wire _354_ ;
wire _583_ ;
wire _163_ ;
wire _639_ ;
wire _219_ ;
wire _392_ ;
wire _868_ ;
wire _448_ ;
wire _677_ ;
wire _257_ ;
wire _486_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _601_ ;
wire _198_ ;
wire _830_ ;
wire _410_ ;
wire _90_ ;
wire _8_ ;
wire _504_ ;
wire _733_ ;
wire _313_ ;
wire _49_ ;
wire _542_ ;
wire _122_ ;
wire _771_ ;
wire _351_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _636_ ;
wire _216_ ;
wire _865_ ;
wire _445_ ;
wire _674_ ;
wire _254_ ;
wire _483_ ;
wire _539_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _768_ ;
wire _348_ ;
wire _577_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire _289_ ;
wire _5_ ;
wire [3:0] _921_ ;
wire _501_ ;
wire _730_ ;
wire _310_ ;
wire _46_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _633_ ;
wire _213_ ;
wire _862_ ;
wire _442_ ;
wire _918_ ;
wire _671_ ;
wire _251_ ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire _536_ ;
wire _116_ ;
wire _765_ ;
wire _345_ ;
wire _574_ ;
wire _154_ ;
wire _383_ ;
wire _859_ ;
wire _439_ ;
wire _192_ ;
wire _668_ ;
wire _248_ ;
wire _897_ ;
wire _477_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire _189_ ;
wire _821_ ;
wire _401_ ;
wire _81_ ;
wire _630_ ;
wire _210_ ;
wire _915_ ;
wire _724_ ;
wire _304_ ;
wire _533_ ;
wire _113_ ;
wire _762_ ;
wire _342_ ;
wire _818_ ;
wire _78_ ;
wire _571_ ;
wire _151_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _856_ ;
wire _436_ ;
wire [3:0] Xin ;
wire _665_ ;
wire _245_ ;
wire _894_ ;
wire _474_ ;
wire _283_ ;
wire _759_ ;
wire _339_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire _797_ ;
wire _377_ ;
wire _186_ ;
wire _912_ ;
wire _721_ ;
wire _301_ ;
wire _37_ ;
wire _530_ ;
wire _110_ ;
wire _815_ ;
wire _75_ ;
wire _624_ ;
wire _204_ ;
wire _853_ ;
wire _433_ ;
wire _909_ ;
wire _662_ ;
wire _242_ ;
wire _718_ ;
wire _891_ ;
wire _471_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _756_ ;
wire _336_ ;
wire _565_ ;
wire _145_ ;
wire _794_ ;
wire _374_ ;
wire _183_ ;
wire _659_ ;
wire _239_ ;
wire _888_ ;
wire _468_ ;
wire _697_ ;
wire _277_ ;
wire _34_ ;
wire _812_ ;
wire _72_ ;
wire _621_ ;
wire _201_ ;
wire _850_ ;
wire _430_ ;
wire _906_ ;
wire _715_ ;
wire _524_ ;
wire _104_ ;
wire _753_ ;
wire _333_ ;
wire _809_ ;
wire _69_ ;
wire _562_ ;
wire _142_ ;
wire _618_ ;
wire _791_ ;
wire _371_ ;
wire _847_ ;
wire _427_ ;
wire _180_ ;
wire _656_ ;
wire _236_ ;
wire _885_ ;
wire _465_ ;
wire _694_ ;
wire _274_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _788_ ;
wire _368_ ;
wire _597_ ;
wire _177_ ;
wire _903_ ;
wire _712_ ;
wire _28_ ;
wire _521_ ;
wire _101_ ;
wire _750_ ;
wire _330_ ;
wire _806_ ;
wire _66_ ;
wire _615_ ;
wire _844_ ;
wire _424_ ;
wire _653_ ;
wire _233_ ;
wire _709_ ;
wire _882_ ;
wire _462_ ;
wire _518_ ;
wire _691_ ;
wire _271_ ;
wire _747_ ;
wire _327_ ;
wire _556_ ;
wire _136_ ;
wire _785_ ;
wire _365_ ;
wire _594_ ;
wire _174_ ;
wire _879_ ;
wire _459_ ;
wire _688_ ;
wire _268_ ;
wire _900_ ;
wire _497_ ;
wire _25_ ;
wire _803_ ;
wire _63_ ;
wire _612_ ;
wire _841_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire _706_ ;
wire _515_ ;
wire _744_ ;
wire _324_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _782_ ;
wire _362_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _591_ ;
wire _171_ ;
wire _647_ ;
wire _227_ ;
wire _876_ ;
wire _456_ ;
wire _685_ ;
wire _265_ ;
wire _494_ ;
wire _22_ ;
wire _779_ ;
wire _359_ ;

FILL FILL_2__1679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1259_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1328_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_819_),
    .B(_818_),
    .Y(_820_)
);

OAI21X1 _1257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_128_),
    .B(_167_),
    .C(Yin1[2]),
    .Y(_405_)
);

FILL FILL_3__1081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1137_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_618_),
    .B(_623_),
    .C(_546_),
    .Y(_632_)
);

AOI22X1 _1066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[0]),
    .B(Cin[3]),
    .C(XinHL[1]),
    .D(Cin[2]),
    .Y(_217_)
);

FILL FILL_2__1700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100950x93750 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_435_),
    .Y(_442_)
);

FILL FILL_4__1015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1114_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_442_),
    .B(_443_),
    .Y(_536_)
);

FILL FILL_2__1603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1182_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_729_),
    .B(_734_),
    .C(_741_),
    .Y(_745_)
);

NAND2X1 _932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[2]),
    .B(_112_),
    .Y(_113_)
);

FILL FILL_1__1763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1269_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_338_),
    .B(_332_),
    .C(_321_),
    .Y(_347_)
);

FILL FILL_2__1832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1819_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf4),
    .B(_109_),
    .C(Yin1[2]),
    .Y(_94_)
);

OAI21X1 _1410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_271_),
    .B(_456_),
    .C(_555_),
    .Y(_556_)
);

FILL FILL_1__1572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1208_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf1),
    .B(_y[1]),
    .Y(_139_)
);

FILL FILL_1__1381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1085_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _1504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_645_),
    .B(_648_),
    .C(_647_),
    .Y(_649_)
);

FILL FILL_3__976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1804_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_818_),
    .B(_825_),
    .C(_874_),
    .Y(_875_)
);

OAI21X1 _1313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_380_),
    .B(_383_),
    .C(_387_),
    .Y(_460_)
);

FILL FILL_1__1475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1613_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_596_),
    .B(_593_),
    .Y(_687_)
);

OAI21X1 _1122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_271_),
    .B(_187_),
    .C(_215_),
    .Y(_272_)
);

FILL FILL_1__1284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1002_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf4),
    .B(y[0]),
    .C(_110_),
    .D(y[4]),
    .Y(_111_)
);

NAND3X1 _1771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_881_),
    .B(_905_),
    .C(_884_),
    .Y(_911_)
);

AOI21X1 _1351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_495_),
    .B(_494_),
    .C(_493_),
    .Y(_498_)
);

FILL FILL100650x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1162_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_76_),
    .B(_91_),
    .C(_92_),
    .Y(_44_)
);

AND2X2 _1407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[3]),
    .B(Cin[5]),
    .Y(_553_)
);

FILL FILL100050x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1149_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_723_),
    .Y(_724_)
);

XOR2X1 _1160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_308_),
    .B(_306_),
    .Y(_309_)
);

FILL FILL_1__942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1707_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_775_),
    .B(_774_),
    .C(_720_),
    .Y(_780_)
);

OAI21X1 _1216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148__bF$buf3),
    .B(_364_),
    .C(_301_),
    .Y(_25_)
);

FILL FILL_0__964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1040_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_y[0]),
    .B(LoadCtl_4_bF$buf3),
    .Y(_137_)
);

FILL FILL_1__1798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1516_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1865_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_15_),
    .CLK(clk_bF$buf6),
    .Q(y[11])
);

NAND3X1 _1445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[3]),
    .B(Cin[1]),
    .C(Yin2[0]),
    .Y(_591_)
);

INVX1 _1025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_175_),
    .Y(_178_)
);

FILL FILL100950x58650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1325_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_751_),
    .B(_816_),
    .Y(_817_)
);

AOI21X1 _1254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_399_),
    .B(_394_),
    .C(_398_),
    .Y(_402_)
);

FILL FILL_4__1814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1134_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_525_),
    .Y(_629_)
);

OAI21X1 _1063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_206_),
    .B(_213_),
    .C(_203_),
    .Y(_214_)
);

FILL FILL_4__1623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1294_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_681_),
    .B(_679_),
    .C(_675_),
    .Y(_684_)
);

AND2X2 _1119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[2]),
    .B(Cin[2]),
    .Y(_269_)
);

FILL FILL_3__1783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1363_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_435_),
    .B(_365_),
    .C(_438_),
    .Y(_440_)
);

FILL FILL_4__1012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1419_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_908_),
    .B(_905_),
    .C(_148__bF$buf0),
    .Y(_909_)
);

NAND2X1 _1348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_488_),
    .B(_490_),
    .Y(_495_)
);

FILL FILL_3__1592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1228_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_720_),
    .Y(_721_)
);

INVX1 _1157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_305_),
    .Y(_306_)
);

FILL FILL_1__939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1037_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_530_),
    .B(_531_),
    .C(_532_),
    .Y(_533_)
);

FILL FILL_2__1600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1266_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_339_),
    .B(_343_),
    .C(_310_),
    .Y(_344_)
);

FILL FILL_1__977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100950x46950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1014_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_424_),
    .B(_429_),
    .C(_367_),
    .Y(_437_)
);

FILL FILL_2__1503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1082_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[0]),
    .B(Cin[6]),
    .Y(_646_)
);

FILL FILL_3__973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1169_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148__bF$buf3),
    .B(_248_),
    .C(_212_),
    .Y(_23_)
);

FILL FILL_2__1732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1719_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_862_),
    .B(_871_),
    .C(_870_),
    .Y(_872_)
);

OAI21X1 _1310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_190_),
    .B(_456_),
    .C(_451_),
    .Y(_457_)
);

FILL FILL_1__1472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL101250x78150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__923_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[2]),
    .B(y[12]),
    .C(_107_),
    .Y(_108_)
);

FILL FILL_1__1757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1406_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_816_),
    .B(_86_),
    .C(_90_),
    .Y(_43_)
);

NAND2X1 _1404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[1]),
    .B(Cin[7]),
    .Y(_550_)
);

FILL FILL_1__1566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1635_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1704_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_773_),
    .B(_776_),
    .C(_719_),
    .Y(_777_)
);

AOI22X1 _1213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_361_),
    .B(_244_),
    .C(_354_),
    .D(_358_),
    .Y(_362_)
);

FILL FILL_0__961_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[3]),
    .B(_110_),
    .Y(_135_)
);

FILL FILL_1__1795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1513_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1862_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_12_),
    .CLK(clk_bF$buf5),
    .Q(y[8])
);

NAND3X1 _1442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_584_),
    .B(_587_),
    .C(_586_),
    .Y(_588_)
);

NAND2X1 _1022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[0]),
    .B(Cin[1]),
    .Y(_175_)
);

FILL FILL_1__1184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1079_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_921_[2]),
    .Y(Yout[2])
);

FILL FILL_3__1742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1322_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_805_),
    .B(_807_),
    .C(_802_),
    .Y(_814_)
);

INVX1 _1251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_396_),
    .Y(_399_)
);

FILL FILL_4__1811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1062_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_861_),
    .B(_863_),
    .C(_868_),
    .Y(_869_)
);

OAI21X1 _1307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_271_),
    .B(_304_),
    .C(_453_),
    .Y(_454_)
);

FILL FILL_3__1551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1049_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_621_),
    .B(_622_),
    .C(_548_),
    .Y(_626_)
);

OAI21X1 _1060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_209_),
    .B(_211_),
    .C(_185_),
    .Y(_22_)
);

FILL FILL_4__1620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1607_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _1536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_591_),
    .B(Yin2[1]),
    .Y(_681_)
);

NAND2X1 _1116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[0]),
    .B(Cin[4]),
    .Y(_266_)
);

FILL FILL_3__1780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1416_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_905_),
    .Y(_906_)
);

NAND3X1 _1345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_),
    .B(_491_),
    .C(_489_),
    .Y(_492_)
);

FILL FILL_1__1087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL101250x66450 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_690_),
    .B(_694_),
    .C(_697_),
    .Y(_718_)
);

OAI21X1 _1154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_250_),
    .B(_284_),
    .C(_292_),
    .Y(_303_)
);

FILL FILL_1__936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1034_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_367_),
    .B(_529_),
    .C(_432_),
    .Y(_530_)
);

FILL FILL_0__1843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1194_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1859_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_9_),
    .CLK(clk_bF$buf1),
    .Q(y[5])
);

AND2X2 _1439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[2]),
    .B(Cin[3]),
    .Y(_585_)
);

AOI21X1 _1019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[1]),
    .B(Cin_0_bF$buf1),
    .C(Yin0[1]),
    .Y(_172_)
);

FILL FILL_3__1683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1263_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_322_),
    .B(_331_),
    .C(_328_),
    .Y(_341_)
);

FILL FILL_1__974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1319_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_810_),
    .B(_806_),
    .C(_795_),
    .Y(_811_)
);

AOI21X1 _1248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[2]),
    .B(Cin_0_bF$buf3),
    .C(Yin1[2]),
    .Y(_396_)
);

FILL FILL_0__996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1072_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[12]),
    .Y(_157_)
);

FILL FILL_4__1808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1128_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1897_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_47_),
    .CLK(clk_bF$buf3),
    .Q(Yin1[3])
);

OAI21X1 _1477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_622_),
    .B(_621_),
    .C(_620_),
    .Y(_623_)
);

AOI21X1 _1057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_205_),
    .B(_208_),
    .C(_186_),
    .Y(_209_)
);

FILL FILL_4__1617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1357_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_431_),
    .B(_432_),
    .C(_433_),
    .Y(_434_)
);

FILL FILL_2__1500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1166_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _1095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_244_),
    .B(_210_),
    .C(_243_),
    .Y(_246_)
);

FILL FILL_0__1555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL101250x54750 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_104_),
    .Y(_105_)
);

FILL FILL_1__1754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1334_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_333_),
    .B(_337_),
    .C(_322_),
    .Y(_338_)
);

FILL FILL_2__1823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1229_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[2]),
    .B(_86_),
    .Y(_89_)
);

INVX1 _1401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_514_),
    .Y(_547_)
);

FILL FILL_1__1563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1619_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_763_),
    .B(_767_),
    .C(_769_),
    .Y(_774_)
);

NAND3X1 _1210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_354_),
    .B(_358_),
    .C(_302_),
    .Y(_359_)
);

OAI21X1 _961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_126_),
    .B(_110_),
    .C(_133_),
    .Y(_1_)
);

FILL FILL_1__1792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1076_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_920_[3]),
    .Y(Xout[3])
);

FILL FILL_1_BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1657_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1306_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_864_),
    .B(_865_),
    .Y(_866_)
);

AND2X2 _1304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[2]),
    .B(Cin[5]),
    .Y(_451_)
);

FILL FILL_1__1466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL99750x15750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1604_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _1533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_128_),
    .B(_275_),
    .C(_130_),
    .D(_187_),
    .Y(_678_)
);

NAND3X1 _1113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_256_),
    .B(_260_),
    .C(_255_),
    .Y(_263_)
);

FILL FILL_1__1695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1413_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_898_),
    .B(_902_),
    .C(_862_),
    .Y(_903_)
);

NAND3X1 _1342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[3]),
    .B(Cin_0_bF$buf0),
    .C(_488_),
    .Y(_489_)
);

FILL FILL_1__1084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1399_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_76_),
    .B(_86_),
    .C(_87_),
    .Y(_40_)
);

FILL FILL_3__1642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_628_),
    .B(_711_),
    .C(_710_),
    .Y(_715_)
);

OAI21X1 _1151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_298_),
    .B(_300_),
    .C(_249_),
    .Y(_24_)
);

FILL FILL_1__933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1382_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_747_),
    .B(_762_),
    .Y(_771_)
);

AOI21X1 _1207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_352_),
    .B(_351_),
    .C(_350_),
    .Y(_356_)
);

FILL FILL_0__955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1031_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[0]),
    .B(_110_),
    .Y(_132_)
);

FILL FILL_1__1789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1369_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_526_),
    .B(_525_),
    .C(_524_),
    .Y(_527_)
);

FILL FILL_0__1840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1507_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1856_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6_),
    .CLK(clk_bF$buf0),
    .Q(y[2])
);

NAND3X1 _1436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[1]),
    .B(Cin[3]),
    .C(_581_),
    .Y(_582_)
);

NAND2X1 _1016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_165_),
    .B(_169_),
    .Y(_170_)
);

FILL FILL_3__1680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1316_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _1665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_796_),
    .B(_798_),
    .C(_804_),
    .Y(_808_)
);

NAND2X1 _1245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[1]),
    .B(Cin[1]),
    .Y(_393_)
);

FILL FILL_0__993_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf1),
    .B(_116_),
    .C(_155_),
    .Y(_14_)
);

FILL FILL_4__1805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1125_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1894_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_44_),
    .CLK(clk_bF$buf2),
    .Q(Yin1[0])
);

OAI21X1 _1474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_470_),
    .B(_619_),
    .C(_514_),
    .Y(_620_)
);

NAND2X1 _1054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[0]),
    .B(Cin[2]),
    .Y(_206_)
);

FILL FILL_0__1514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1354_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_367_),
    .Y(_431_)
);

FILL FILL_4__1003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL101250x19650 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_867_),
    .B(_897_),
    .C(_872_),
    .Y(_900_)
);

INVX1 _1339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_485_),
    .Y(_486_)
);

FILL FILL_3__1583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1163_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_214_),
    .B(_242_),
    .Y(_243_)
);

FILL FILL_0__1552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1219_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_y[9]),
    .B(_148__bF$buf2),
    .Y(_713_)
);

AOI21X1 _1148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297_),
    .B(_294_),
    .C(_246_),
    .Y(_298_)
);

FILL FILL_3__1392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1028_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_71_),
    .Y(_72_)
);

INVX1 _1377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_446_),
    .Y(_524_)
);

FILL FILL100050x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1257_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[1]),
    .B(Cin_0_bF$buf3),
    .C(_334_),
    .Y(_335_)
);

FILL FILL_1__968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1073_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_920_[0]),
    .Y(Xout[0])
);

FILL FILL_3__964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1234_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_234_),
    .B(_239_),
    .C(_233_),
    .Y(_240_)
);

FILL FILL_2__1723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1129_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_862_),
    .Y(_863_)
);

AOI21X1 _1301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_420_),
    .B(_422_),
    .C(_447_),
    .Y(_448_)
);

FILL FILL_1__1463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1519_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_671_),
    .B(_673_),
    .C(_674_),
    .Y(_675_)
);

INVX1 _1110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_257_),
    .Y(_260_)
);

FILL FILL_1__1692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1396_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_84_),
    .B(_78_),
    .C(_85_),
    .Y(_39_)
);

FILL FILL_1__1557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1206_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_763_),
    .B(_767_),
    .C(_722_),
    .Y(_768_)
);

NAND3X1 _1204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_351_),
    .B(_350_),
    .C(_352_),
    .Y(_353_)
);

FILL FILL_0__952_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[3]),
    .Y(_130_)
);

FILL FILL_1__1786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1504_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1853_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3_),
    .CLK(clk_bF$buf4),
    .Q(XinH[3])
);

NAND2X1 _1433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[1]),
    .B(Cin[3]),
    .Y(_579_)
);

INVX1 _1013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf3),
    .Y(_167_)
);

FILL FILL_1__1595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1244_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1909_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(LoadCtl[2]),
    .CLK(clk_bF$buf4),
    .Q(LoadCtl[3])
);

FILL FILL_3__1733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1313_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_798_),
    .B(_804_),
    .C(_796_),
    .Y(_805_)
);

NAND2X1 _1242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_389_),
    .B(_384_),
    .Y(_390_)
);

FILL FILL_0__990_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf1),
    .B(_y[9]),
    .Y(_154_)
);

FILL FILL_4__1802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1299_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _1718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_859_),
    .B(_854_),
    .Y(_860_)
);

FILL FILL_3__1542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1122_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1891_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_41_),
    .CLK(clk_bF$buf3),
    .Q(Yin2[1])
);

NAND3X1 _1471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_615_),
    .B(_616_),
    .C(_614_),
    .Y(_617_)
);

NAND3X1 _1051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_188_),
    .B(_202_),
    .C(_201_),
    .Y(_203_)
);

FILL FILL_0__1511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1282_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[3]),
    .B(Cin[2]),
    .Y(_672_)
);

NAND2X1 _1107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[3]),
    .B(Cin[1]),
    .Y(_257_)
);

FILL FILL_3__999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1269_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_418_),
    .B(_413_),
    .C(_377_),
    .Y(_428_)
);

FILL FILL_4__1000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1407_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _1756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_896_),
    .B(Yin3[1]),
    .Y(_897_)
);

NAND3X1 _1336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_479_),
    .B(_482_),
    .C(_481_),
    .Y(_483_)
);

FILL FILL_3__1580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1216_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _1565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_708_),
    .B(_709_),
    .C(_638_),
    .D(_632_),
    .Y(_710_)
);

INVX1 _1145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_244_),
    .Y(_295_)
);

FILL FILL_1__927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin3[2]),
    .B(_800_),
    .C(_893_),
    .Y(_69_)
);

AOI21X1 _1374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_506_),
    .B(_511_),
    .C(_470_),
    .Y(_521_)
);

FILL FILL_0__1834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1254_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_331_),
    .B(_328_),
    .C(_323_),
    .Y(_332_)
);

FILL FILL_1__965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1804_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_799_),
    .B(_797_),
    .C(_801_),
    .Y(_802_)
);

NAND2X1 _1239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_314_),
    .B(_386_),
    .Y(_387_)
);

FILL FILL_0__987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1119_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1888_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_38_),
    .CLK(clk_bF$buf3),
    .Q(Yin3[2])
);

AND2X2 _1468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_569_),
    .B(_574_),
    .Y(_614_)
);

NAND3X1 _1048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_189_),
    .B(_199_),
    .C(_196_),
    .Y(_200_)
);

FILL FILL_3__1292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1348_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_834_),
    .B(_839_),
    .Y(_840_)
);

AOI21X1 _1277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_343_),
    .B(_339_),
    .C(_345_),
    .Y(_425_)
);

FILL FILL_2__1911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1157_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _1086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[3]),
    .Y(_237_)
);

FILL FILL_2__1720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1393_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_82_),
    .B(_78_),
    .C(_83_),
    .Y(_38_)
);

FILL FILL_1__1554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__978_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_760_),
    .B(_749_),
    .Y(_765_)
);

INVX1 _1201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_309_),
    .Y(_350_)
);

INVX2 _952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[2]),
    .Y(_128_)
);

FILL FILL_1__1783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1419_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1850_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_0_),
    .CLK(clk_bF$buf0),
    .Q(XinH[0])
);

INVX1 _1430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_503_),
    .Y(_576_)
);

OAI21X1 _1010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148__bF$buf1),
    .B(_163_),
    .C(_164_),
    .Y(_19_)
);

FILL FILL_1__1592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1067_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1906_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(Rdy),
    .CLK(clk_bF$buf2),
    .Q(LoadCtl[0])
);

FILL FILL_3__958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1228_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148__bF$buf4),
    .B(_151_),
    .C(_152_),
    .Y(_11_)
);

FILL FILL_2__1717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1296_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[3]),
    .B(Cin[6]),
    .Y(_857_)
);

FILL FILL_1__1457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1106_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_494_),
    .B(_496_),
    .C(_601_),
    .Y(_669_)
);

AOI21X1 _1104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[0]),
    .B(Cin_0_bF$buf2),
    .C(Yin1[0]),
    .Y(_254_)
);

FILL FILL_3__996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1404_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_800_),
    .B(_893_),
    .Y(_894_)
);

AND2X2 _1333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[1]),
    .B(Cin[2]),
    .Y(_480_)
);

FILL FILL_1__1495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1144_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_80_),
    .B(_78_),
    .C(_81_),
    .Y(_37_)
);

FILL FILL_3__1633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1213_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_703_),
    .B(_706_),
    .C(_639_),
    .Y(_707_)
);

NAND3X1 _1142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_251_),
    .B(_279_),
    .C(_283_),
    .Y(_292_)
);

FILL FILL_1__924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1199_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_761_),
    .B(_758_),
    .Y(_762_)
);

FILL FILL_0__946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1022_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[1]),
    .Y(_126_)
);

OAI21X1 _1791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_914_),
    .B(_912_),
    .C(_64_),
    .Y(_66_)
);

AOI21X1 _1371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_412_),
    .B(_408_),
    .C(_415_),
    .Y(_518_)
);

FILL FILL_0__1831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1918_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf1),
    .B(_271_),
    .C(_102_),
    .Y(_54_)
);

OAI21X1 _1427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_557_),
    .B(_560_),
    .C(_567_),
    .Y(_573_)
);

OAI21X1 _1007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf0),
    .B(_161_),
    .C(_162_),
    .Y(_18_)
);

FILL FILL_3__1671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1169_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_324_),
    .Y(_329_)
);

FILL FILL_1__962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100650x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1307_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_798_),
    .Y(_799_)
);

OAI21X1 _1236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_382_),
    .B(_383_),
    .C(_380_),
    .Y(_384_)
);

FILL FILL_0__984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1060_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148__bF$buf4),
    .B(_149_),
    .C(_150_),
    .Y(_10_)
);

FILL FILL_1__1398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1885_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_35_),
    .CLK(clk_bF$buf6),
    .Q(_y[15])
);

AOI21X1 _1465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_594_),
    .B(_597_),
    .C(_589_),
    .Y(_611_)
);

NAND2X1 _1045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[1]),
    .B(Cin[1]),
    .Y(_197_)
);

FILL FILL_0__1505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1345_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_832_),
    .B(_831_),
    .C(_790_),
    .Y(_837_)
);

OAI21X1 _1274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_417_),
    .B(_416_),
    .C(_379_),
    .Y(_422_)
);

FILL FILL100050x39150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100950x82050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1154_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_226_),
    .B(_221_),
    .C(_225_),
    .Y(_234_)
);

FILL FILL_0__1543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1704_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_697_),
    .B(_694_),
    .C(_690_),
    .Y(_704_)
);

OAI21X1 _1139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_288_),
    .B(_284_),
    .C(_250_),
    .Y(_289_)
);

FILL FILL_3__1383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1019_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_62_),
    .B(_63_),
    .Y(_64_)
);

OAI21X1 _1368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_510_),
    .B(_509_),
    .C(_472_),
    .Y(_515_)
);

FILL FILL_3__1192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1248_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_676_),
    .B(_678_),
    .C(_740_),
    .Y(_741_)
);

INVX1 _1177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_325_),
    .Y(_326_)
);

FILL FILL_1__959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100650x31350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1064_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1903_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_53_),
    .CLK(clk_bF$buf0),
    .Q(XinHL[1])
);

FILL FILL_3__955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1293_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[1]),
    .B(Cin[7]),
    .Y(_854_)
);

FILL FILL_1__1454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100950x70350 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_654_),
    .B(_649_),
    .C(_660_),
    .Y(_666_)
);

OAI21X1 _1101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_232_),
    .B(_230_),
    .C(_228_),
    .Y(_251_)
);

FILL FILL_3__993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1319_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[7]),
    .Y(_891_)
);

NAND2X1 _1330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_476_),
    .B(_386_),
    .Y(_477_)
);

FILL FILL_1__1492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1387_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_76_),
    .B(_78_),
    .C(_79_),
    .Y(_36_)
);

FILL FILL_3__1630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100350x66450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1196_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin2[1]),
    .B(_592_),
    .Y(_759_)
);

FILL FILL_0__943_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[0]),
    .Y(_124_)
);

FILL FILL_1__1777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1915_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf1),
    .B(Xin[1]),
    .Y(_101_)
);

INVX1 _1424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_451_),
    .Y(_570_)
);

OAI21X1 _1004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148__bF$buf1),
    .B(_159_),
    .C(_160_),
    .Y(_17_)
);

FILL FILL_1__1586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1304_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[0]),
    .B(Cin[7]),
    .Y(_796_)
);

NAND2X1 _1233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[0]),
    .B(Cin[2]),
    .Y(_381_)
);

FILL FILL_0__981_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf2),
    .Y(_148_)
);

FILL FILL_1__1395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1044_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_806_),
    .B(_823_),
    .Y(_851_)
);

FILL FILL_3__1533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1113_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1882_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_32_),
    .CLK(clk_bF$buf6),
    .Q(_y[12])
);

NAND2X1 _1462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_596_),
    .B(_593_),
    .Y(_608_)
);

INVX1 _1042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_193_),
    .Y(_194_)
);

FILL FILL_0__1502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1099_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[3]),
    .B(Cin[6]),
    .Y(_663_)
);

FILL FILL_3__1762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1342_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_833_),
    .B(_789_),
    .C(_829_),
    .Y(_834_)
);

NAND3X1 _1271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_377_),
    .B(_413_),
    .C(_418_),
    .Y(_419_)
);

FILL FILL_0__1731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1818_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_849_),
    .B(_885_),
    .Y(_888_)
);

NAND2X1 _1327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[0]),
    .B(Cin[3]),
    .Y(_474_)
);

FILL FILL_3__1571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100050x15750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1069_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_230_),
    .B(_229_),
    .C(_218_),
    .Y(_231_)
);

FILL FILL_0__1540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1207_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_700_),
    .B(_699_),
    .C(_668_),
    .Y(_701_)
);

NAND3X1 _1136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_265_),
    .B(_282_),
    .C(_262_),
    .Y(_286_)
);

FILL FILL_3__1380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1016_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_917_),
    .B(_919_),
    .C(_60_),
    .Y(_61_)
);

NAND3X1 _1365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_470_),
    .B(_511_),
    .C(_506_),
    .Y(_512_)
);

FILL FILL_0__1825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1245_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_731_),
    .B(_730_),
    .C(_733_),
    .Y(_738_)
);

INVX1 _1174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_322_),
    .Y(_323_)
);

FILL FILL_1__956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1604_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1879_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_29_),
    .CLK(clk_bF$buf5),
    .Q(_y[9])
);

NAND3X1 _1459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_598_),
    .B(_604_),
    .C(_577_),
    .Y(_605_)
);

INVX1 _1039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[1]),
    .Y(_191_)
);

FILL FILL_3__1283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100950x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1339_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_821_),
    .B(_825_),
    .C(_830_),
    .Y(_831_)
);

AOI21X1 _1268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_410_),
    .B(_411_),
    .C(_409_),
    .Y(_416_)
);

FILL FILL_3__1092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1079_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1900_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_50_),
    .CLK(clk_bF$buf2),
    .Q(Yin0[2])
);

FILL FILL_3__952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1148_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_615_),
    .Y(_642_)
);

NAND3X1 _1077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_219_),
    .B(_227_),
    .C(_224_),
    .Y(_228_)
);

FILL FILL_2__1711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1384_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[2]),
    .Y(_77_)
);

FILL FILL_1__1545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1193_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin2[2]),
    .B(_755_),
    .Y(_756_)
);

FILL FILL_0__940_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[2]),
    .B(y[15]),
    .C(_121_),
    .Y(_122_)
);

FILL FILL_1__1774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1912_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf2),
    .B(_235_),
    .C(_99_),
    .Y(_51_)
);

AOI21X1 _1421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_479_),
    .B(_482_),
    .C(_566_),
    .Y(_567_)
);

OAI21X1 _1001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf2),
    .B(_157_),
    .C(_158_),
    .Y(_16_)
);

FILL FILL_1__1583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1219_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_758_),
    .Y(_793_)
);

INVX1 _1230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_341_),
    .Y(_378_)
);

INVX1 _981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[5]),
    .Y(_146_)
);

FILL FILL_1__1392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100950x23550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1287_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_839_),
    .B(_847_),
    .C(_845_),
    .D(_715_),
    .Y(_848_)
);

FILL FILL_3__1530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1096_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_480_),
    .B(_585_),
    .C(_587_),
    .D(_584_),
    .Y(_660_)
);

FILL FILL_3__987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1815_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _1744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_849_),
    .B(_885_),
    .Y(_886_)
);

INVX1 _1324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_410_),
    .Y(_471_)
);

FILL FILL_1__1486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1204_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_662_),
    .B(_667_),
    .C(_693_),
    .D(_692_),
    .Y(_698_)
);

OAI21X1 _1133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_280_),
    .B(_281_),
    .C(_282_),
    .Y(_283_)
);

FILL FILL_1__1295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[2]),
    .B(Cin[4]),
    .C(XinH[3]),
    .D(Cin[3]),
    .Y(_753_)
);

FILL FILL_0__937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1013_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_919_),
    .B(_56_),
    .Y(_58_)
);

AOI21X1 _1362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_503_),
    .B(_504_),
    .C(_502_),
    .Y(_509_)
);

FILL FILL_0__1822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1099_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf2),
    .B(Yin0[2]),
    .Y(_98_)
);

NAND3X1 _1418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_550_),
    .B(_558_),
    .C(_559_),
    .Y(_564_)
);

FILL FILL_3__1662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100650x58650 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_585_),
    .B(_672_),
    .Y(_735_)
);

NAND3X1 _1171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_317_),
    .B(_319_),
    .C(_318_),
    .Y(_320_)
);

FILL FILL_1__953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1718_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_744_),
    .B(_746_),
    .Y(_790_)
);

NAND2X1 _1227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[3]),
    .B(Cin[3]),
    .Y(_375_)
);

FILL FILL_0__975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1051_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[4]),
    .Y(_144_)
);

FILL FILL_1__1389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1107_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1876_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_26_),
    .CLK(clk_bF$buf1),
    .Q(_y[6])
);

NOR2X1 _1456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_596_),
    .B(_601_),
    .Y(_602_)
);

OAI21X1 _1036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_175_),
    .B(_172_),
    .C(_173_),
    .Y(_188_)
);

FILL FILL_3__1280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1336_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_793_),
    .B(_771_),
    .C(_827_),
    .Y(_828_)
);

NAND3X1 _1265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_408_),
    .B(_412_),
    .C(_379_),
    .Y(_413_)
);

FILL FILL_0__1725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100950x11850 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1145_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_545_),
    .B(_626_),
    .C(_638_),
    .Y(_639_)
);

INVX1 _1074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_220_),
    .Y(_225_)
);

FILL FILL_0__1534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1374_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf4)
);

BUFX2 BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf3)
);

BUFX2 BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf2)
);

BUFX2 BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf1)
);

BUFX2 BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf0)
);

FILL FILL_0__1763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1504_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918_),
    .B(Yin3[2]),
    .Y(_919_)
);

NAND3X1 _1359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_501_),
    .B(_505_),
    .C(_472_),
    .Y(_506_)
);

FILL FILL_3__1183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1239_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_727_),
    .Y(_732_)
);

INVX1 _1168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_311_),
    .Y(_317_)
);

FILL FILL_2__1802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL101250x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1381_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_74_),
    .B(LoadCtl_4_bF$buf0),
    .Y(_75_)
);

FILL FILL_1__1542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1048_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_512_),
    .B(_516_),
    .C(_519_),
    .Y(_543_)
);

FILL FILL_2__1611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100650x46950 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_105_),
    .B(_118_),
    .C(_119_),
    .Y(_921_[2])
);

FILL FILL_1__1771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1284_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_840_),
    .B(_783_),
    .Y(_845_)
);

FILL FILL100950x85950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1093_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_654_),
    .B(_649_),
    .C(_656_),
    .Y(_657_)
);

FILL FILL_3__984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1812_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_876_),
    .B(_880_),
    .Y(_883_)
);

OAI21X1 _1321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_455_),
    .B(_459_),
    .C(_464_),
    .Y(_468_)
);

FILL FILL_1__1483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1119_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_694_),
    .B(_690_),
    .C(_643_),
    .Y(_695_)
);

AOI21X1 _1130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_264_),
    .B(_263_),
    .C(_252_),
    .Y(_280_)
);

FILL FILL_1__1292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1187_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin2[2]),
    .Y(_750_)
);

FILL FILL_0__934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1010_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[2]),
    .B(_116_),
    .Y(_117_)
);

FILL FILL_1__1768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL101250x31350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1096_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf3),
    .B(_168_),
    .C(_96_),
    .Y(_48_)
);

AND2X2 _1415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_474_),
    .B(_476_),
    .Y(_561_)
);

FILL FILL_4_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1715_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_783_),
    .B(_717_),
    .C(_777_),
    .Y(_787_)
);

NAND2X1 _1224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_371_),
    .B(_305_),
    .Y(_372_)
);

FILL FILL_0__972_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[3]),
    .Y(_142_)
);

FILL FILL_1__1386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1104_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1873_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_23_),
    .CLK(clk_bF$buf0),
    .Q(_y[3])
);

AND2X2 _1453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_588_),
    .B(_583_),
    .Y(_599_)
);

NAND2X1 _1033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_y[2]),
    .B(_148__bF$buf3),
    .Y(_185_)
);

FILL FILL_1__1195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1264_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_652_),
    .B(_653_),
    .C(_650_),
    .Y(_654_)
);

FILL FILL_3__1753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1333_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_822_),
    .B(_823_),
    .C(_824_),
    .Y(_825_)
);

NAND3X1 _1262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_391_),
    .B(_400_),
    .C(_397_),
    .Y(_410_)
);

FILL FILL_0__1722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1809_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_878_),
    .B(_879_),
    .C(_877_),
    .Y(_880_)
);

NAND3X1 _1318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_463_),
    .B(_462_),
    .C(_464_),
    .Y(_465_)
);

FILL FILL_3__1562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1142_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_628_),
    .Y(_636_)
);

INVX1 _1071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_221_),
    .Y(_222_)
);

FILL FILL_4__997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL99750x150 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_683_),
    .B(_684_),
    .C(_688_),
    .Y(_692_)
);

NAND3X1 _1127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_266_),
    .B(_274_),
    .C(_276_),
    .Y(_277_)
);

FILL FILL_3__1791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1007_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_863_),
    .B(_900_),
    .C(_898_),
    .Y(_916_)
);

NAND3X1 _1356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_485_),
    .B(_496_),
    .C(_492_),
    .Y(_503_)
);

FILL FILL_3__1180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1236_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _1585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_725_),
    .B(_726_),
    .C(_728_),
    .Y(_729_)
);

AND2X2 _1165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[3]),
    .B(Cin[2]),
    .Y(_314_)
);

FILL FILL_1__947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1045_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_528_),
    .Y(_540_)
);

FILL FILL_4__1534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1404_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_812_),
    .B(_814_),
    .C(_813_),
    .Y(_822_)
);

OAI21X1 _1259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_402_),
    .B(_406_),
    .C(_391_),
    .Y(_407_)
);

FILL FILL_3__1083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1139_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_628_),
    .B(_633_),
    .Y(_634_)
);

OAI21X1 _1068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_197_),
    .B(_192_),
    .C(_193_),
    .Y(_219_)
);

FILL FILL_2__1702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1281_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_842_),
    .B(_841_),
    .C(LoadCtl_4_bF$buf2),
    .Y(_843_)
);

FILL FILL_1__1442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1368_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_432_),
    .Y(_444_)
);

FILL FILL_2__1511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL99750x66450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1184_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_746_),
    .B(_743_),
    .Y(_747_)
);

FILL FILL_0__931_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf4),
    .B(y[1]),
    .C(_110_),
    .D(y[5]),
    .Y(_115_)
);

FILL FILL_1__1765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL101250x93750 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf0),
    .B(_109_),
    .C(Yin1[3]),
    .Y(_95_)
);

OAI21X1 _1412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_271_),
    .B(_456_),
    .C(_553_),
    .Y(_558_)
);

FILL FILL_1__1574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1712_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_783_),
    .B(_717_),
    .C(LoadCtl_4_bF$buf2),
    .Y(_785_)
);

AOI21X1 _1221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_350_),
    .B(_352_),
    .C(_368_),
    .Y(_369_)
);

INVX1 _972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[2]),
    .Y(_140_)
);

FILL FILL_1__1383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1019_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1870_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_20_),
    .CLK(clk_bF$buf0),
    .Q(_y[0])
);

OAI21X1 _1450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_),
    .B(_595_),
    .C(_494_),
    .Y(_596_)
);

NAND2X1 _1030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_182_),
    .B(_181_),
    .Y(_183_)
);

FILL FILL_1__1192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL99450x15750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1087_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[0]),
    .B(Cin[6]),
    .Y(_651_)
);

FILL FILL_3__978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1806_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_851_),
    .Y(_877_)
);

NAND3X1 _1315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_449_),
    .B(_457_),
    .C(_458_),
    .Y(_462_)
);

FILL FILL_1__1477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1615_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_683_),
    .B(_684_),
    .C(_688_),
    .Y(_689_)
);

OAI21X1 _1124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_271_),
    .B(_187_),
    .C(_268_),
    .Y(_274_)
);

FILL FILL_1__1286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1004_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_905_),
    .B(_887_),
    .Y(_913_)
);

OAI21X1 _1353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_498_),
    .B(_499_),
    .C(_485_),
    .Y(_500_)
);

FILL FILL_1__1095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1164_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_80_),
    .B(_91_),
    .C(_93_),
    .Y(_45_)
);

NAND2X1 _1409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[3]),
    .B(Cin[5]),
    .Y(_555_)
);

FILL FILL_3__1653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1233_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[0]),
    .B(Cin[6]),
    .C(XinH[1]),
    .D(Cin[5]),
    .Y(_726_)
);

NAND2X1 _1162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[1]),
    .B(Cin[4]),
    .Y(_311_)
);

FILL FILL_1__944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL99750x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1709_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_780_),
    .B(_781_),
    .C(_779_),
    .Y(_782_)
);

INVX1 _1218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_354_),
    .Y(_366_)
);

FILL FILL_0__966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1042_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[1]),
    .Y(_138_)
);

AOI21X1 _1391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_536_),
    .B(_537_),
    .C(_148__bF$buf4),
    .Y(_538_)
);

FILL FILL_4__1531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1518_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1867_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_17_),
    .CLK(clk_bF$buf6),
    .Q(y[13])
);

NOR2X1 _1447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_590_),
    .B(_592_),
    .Y(_593_)
);

NAND2X1 _1027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_179_),
    .B(_176_),
    .Y(_180_)
);

FILL FILL_3__1691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1327_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_817_),
    .B(_756_),
    .Y(_819_)
);

NAND3X1 _1256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[2]),
    .B(Cin_0_bF$buf0),
    .C(_403_),
    .Y(_404_)
);

FILL FILL_3__1080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1136_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_626_),
    .B(_625_),
    .C(_545_),
    .Y(_631_)
);

NOR2X1 _1065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_206_),
    .B(_215_),
    .Y(_216_)
);

FILL FILL_0__1525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1365_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _1294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf4),
    .B(_149_),
    .C(_439_),
    .D(_441_),
    .Y(_26_)
);

FILL FILL_0__1754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL101250x58650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_645_),
    .B(_648_),
    .C(_652_),
    .Y(_723_)
);

FILL FILL_0_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_215_),
    .B(_307_),
    .C(_273_),
    .Y(_308_)
);

FILL FILL_0_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1039_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_442_),
    .B(_443_),
    .C(_534_),
    .Y(_535_)
);

FILL FILL_2__1602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1199_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_738_),
    .B(_739_),
    .C(_736_),
    .Y(_744_)
);

INVX1 _931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[9]),
    .Y(_112_)
);

FILL FILL_1__1762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1268_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_341_),
    .B(_342_),
    .C(_340_),
    .Y(_346_)
);

FILL FILL_1__979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1657_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1077_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf0)
);

BUFX2 BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148_),
    .Y(_148__bF$buf4)
);

BUFX2 BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148_),
    .Y(_148__bF$buf3)
);

BUFX2 BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148_),
    .Y(_148__bF$buf2)
);

BUFX2 BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148_),
    .Y(_148__bF$buf1)
);

BUFX2 BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148_),
    .Y(_148__bF$buf0)
);

FILL FILL_2__1640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1084_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[0]),
    .B(Cin[5]),
    .C(XinHL[3]),
    .D(Cin[6]),
    .Y(_648_)
);

FILL FILL_3__975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1803_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_872_),
    .B(_869_),
    .Y(_874_)
);

AOI21X1 _1312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_457_),
    .B(_458_),
    .C(_449_),
    .Y(_459_)
);

FILL FILL_1__1474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1612_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_670_),
    .B(_685_),
    .Y(_686_)
);

INVX2 _1121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[2]),
    .Y(_271_)
);

FILL FILL_1__1283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL101250x46950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1001_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf4),
    .B(_109_),
    .Y(_110_)
);

FILL FILL_1__1759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1339_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_y[14]),
    .B(_148__bF$buf0),
    .Y(_910_)
);

NAND3X1 _1350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_492_),
    .B(_496_),
    .C(_486_),
    .Y(_497_)
);

FILL FILL_1__1092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1087_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf3),
    .B(_109_),
    .C(Yin1[0]),
    .Y(_92_)
);

AND2X2 _1406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[2]),
    .B(Cin[6]),
    .Y(_552_)
);

FILL FILL_3__1650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1706_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_640_),
    .B(_705_),
    .C(_778_),
    .Y(_779_)
);

XOR2X1 _1215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_363_),
    .B(_299_),
    .Y(_364_)
);

FILL FILL_0__963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[0]),
    .Y(_136_)
);

FILL FILL_2_CLKBUF1_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1515_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1864_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_14_),
    .CLK(clk_bF$buf5),
    .Q(y[10])
);

AOI21X1 _1444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[3]),
    .B(Cin[1]),
    .C(Yin2[0]),
    .Y(_590_)
);

INVX1 _1024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172_),
    .Y(_177_)
);

FILL FILL_1__1186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1324_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin2[3]),
    .Y(_816_)
);

NAND3X1 _1253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_400_),
    .B(_397_),
    .C(_392_),
    .Y(_401_)
);

FILL FILL_0__1713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1064_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_868_),
    .Y(_871_)
);

INVX1 _1309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[6]),
    .Y(_456_)
);

FILL FILL_3__1553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1133_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_627_),
    .B(_624_),
    .C(_544_),
    .Y(_628_)
);

AOI21X1 _1062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_201_),
    .B(_202_),
    .C(_188_),
    .Y(_213_)
);

FILL FILL_4__988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1609_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_682_),
    .B(_680_),
    .Y(_683_)
);

AND2X2 _1118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[1]),
    .B(Cin[3]),
    .Y(_268_)
);

FILL FILL_3__1782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1362_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_438_),
    .B(_435_),
    .C(_365_),
    .Y(_439_)
);

FILL FILL_2__1769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1418_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887_),
    .B(_888_),
    .Y(_908_)
);

NAND3X1 _1347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[3]),
    .B(Cin_0_bF$buf0),
    .C(Yin1[3]),
    .Y(_494_)
);

FILL FILL_3__1591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1227_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_665_),
    .B(_667_),
    .Y(_720_)
);

NOR2X1 _1156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_166_),
    .B(_304_),
    .Y(_305_)
);

FILL FILL_1__938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1036_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_446_),
    .B(_522_),
    .C(_517_),
    .Y(_532_)
);

FILL FILL_4__1525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1265_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_341_),
    .B(_342_),
    .C(_340_),
    .Y(_343_)
);

FILL FILL_1__976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1204_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1899_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_49_),
    .CLK(clk_bF$buf2),
    .Q(Yin0[1])
);

NAND3X1 _1479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_613_),
    .B(_617_),
    .C(_620_),
    .Y(_625_)
);

NAND2X1 _1059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf3),
    .B(_210_),
    .Y(_211_)
);

FILL FILL_0__1519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1359_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_433_),
    .B(_432_),
    .C(_431_),
    .Y(_436_)
);

FILL FILL_2__1502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1081_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[2]),
    .B(Cin[7]),
    .Y(_645_)
);

FILL FILL_3__972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1168_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_245_),
    .B(_247_),
    .Y(_248_)
);

FILL FILL_2__1731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__922_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[2]),
    .B(_106_),
    .Y(_107_)
);

FILL FILL_1__1756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1084_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[3]),
    .B(_86_),
    .Y(_90_)
);

AND2X2 _1403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_463_),
    .B(_452_),
    .Y(_549_)
);

FILL FILL_1__1565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1703_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_774_),
    .B(_720_),
    .C(_775_),
    .Y(_776_)
);

AND2X2 _1212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_293_),
    .B(_289_),
    .Y(_361_)
);

FILL FILL_0__960_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_128_),
    .B(_110_),
    .C(_134_),
    .Y(_2_)
);

FILL FILL_1__1794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1512_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1861_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_11_),
    .CLK(clk_bF$buf0),
    .Q(y[7])
);

OAI21X1 _1441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_128_),
    .B(_187_),
    .C(_579_),
    .Y(_587_)
);

INVX1 _1021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_173_),
    .Y(_174_)
);

FILL FILL_1__1183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1078_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_921_[1]),
    .Y(Yout[1])
);

FILL FILL_3__969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1239_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_808_),
    .B(_809_),
    .C(_752_),
    .Y(_813_)
);

INVX1 _1250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_393_),
    .Y(_398_)
);

FILL FILL_0__1710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1061_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_866_),
    .B(_867_),
    .Y(_868_)
);

NAND2X1 _1306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[1]),
    .B(Cin[6]),
    .Y(_453_)
);

FILL FILL_3__1550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1606_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_679_),
    .B(_675_),
    .Y(_680_)
);

NAND3X1 _1115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_252_),
    .B(_263_),
    .C(_264_),
    .Y(_265_)
);

FILL FILL_1__1697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1415_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_904_),
    .B(_889_),
    .Y(_905_)
);

NAND2X1 _1344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin1[3]),
    .B(_490_),
    .Y(_491_)
);

FILL FILL_1__1086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1224_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_542_),
    .B(_716_),
    .C(_715_),
    .Y(_717_)
);

INVX1 _1153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_294_),
    .Y(_302_)
);

FILL FILL_1__935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100350x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1384_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_721_),
    .B(_772_),
    .C(_768_),
    .Y(_773_)
);

OAI21X1 _1209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_356_),
    .B(_357_),
    .C(_355_),
    .Y(_358_)
);

FILL FILL_0__957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1033_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_419_),
    .B(_423_),
    .C(_426_),
    .Y(_529_)
);

FILL FILL_4__1522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1509_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1858_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_8_),
    .CLK(clk_bF$buf5),
    .Q(y[4])
);

INVX1 _1438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_578_),
    .Y(_584_)
);

OAI21X1 _1018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148__bF$buf3),
    .B(_170_),
    .C(_171_),
    .Y(_20_)
);

FILL FILL_3__1682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1262_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_316_),
    .B(_320_),
    .Y(_340_)
);

FILL FILL_1__973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1318_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_808_),
    .B(_809_),
    .C(_807_),
    .Y(_810_)
);

INVX1 _1247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_394_),
    .Y(_395_)
);

FILL FILL_0__995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1071_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf0),
    .B(_120_),
    .C(_156_),
    .Y(_15_)
);

FILL FILL_0__1707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1127_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1896_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_46_),
    .CLK(clk_bF$buf4),
    .Q(Yin1[2])
);

AOI21X1 _1476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_612_),
    .B(_605_),
    .C(_575_),
    .Y(_622_)
);

NAND3X1 _1056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_207_),
    .B(_203_),
    .C(_200_),
    .Y(_208_)
);

FILL FILL_0__1516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1356_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_427_),
    .B(_428_),
    .C(_369_),
    .Y(_433_)
);

FILL FILL_0__1745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1165_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_244_),
    .B(_243_),
    .C(_210_),
    .Y(_245_)
);

FILL FILL_0__1554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1104_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_62_),
    .B(_71_),
    .C(_66_),
    .Y(_74_)
);

OAI21X1 _1379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_520_),
    .B(_521_),
    .C(_448_),
    .Y(_526_)
);

FILL FILL_4__1519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1172_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[1]),
    .B(LoadCtl_0_bF$buf0),
    .Y(_104_)
);

FILL FILL_1__1753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1259_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_336_),
    .B(_335_),
    .C(_324_),
    .Y(_337_)
);

FILL FILL_2__1822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100350x31350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1809_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_748_),
    .B(_86_),
    .C(_88_),
    .Y(_41_)
);

INVX1 _1400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_545_),
    .Y(_546_)
);

FILL FILL_1__1562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1618_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[1]),
    .B(_110_),
    .Y(_133_)
);

FILL FILL_1__1791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100650x70350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1075_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_920_[2]),
    .Y(Xout[2])
);

FILL FILL_3__966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1305_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin2[3]),
    .B(_751_),
    .Y(_865_)
);

INVX1 _1303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_449_),
    .Y(_450_)
);

FILL FILL_1__1465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1603_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_585_),
    .B(_672_),
    .Y(_677_)
);

NAND3X1 _1112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_258_),
    .B(_261_),
    .C(_253_),
    .Y(_262_)
);

FILL FILL100050x66450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1412_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_900_),
    .Y(_902_)
);

INVX1 _1341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin1[3]),
    .Y(_488_)
);

FILL FILL_1__1083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1398_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin2[0]),
    .B(_86_),
    .Y(_87_)
);

FILL FILL_3__1641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1139_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_y[10]),
    .B(_148__bF$buf2),
    .Y(_714_)
);

NAND2X1 _1150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf4),
    .B(_299_),
    .Y(_300_)
);

FILL FILL_1__932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1381_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_743_),
    .B(_746_),
    .C(_766_),
    .Y(_770_)
);

AOI21X1 _1206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_291_),
    .B(_216_),
    .C(_288_),
    .Y(_355_)
);

FILL FILL_0__954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1030_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf0),
    .B(_130_),
    .C(_131_),
    .Y(_920_[3])
);

FILL FILL_1__1788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1506_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1855_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5_),
    .CLK(clk_bF$buf5),
    .Q(y[1])
);

NAND2X1 _1435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[2]),
    .B(Cin[2]),
    .Y(_581_)
);

OAI21X1 _1015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_166_),
    .B(_167_),
    .C(_168_),
    .Y(_169_)
);

FILL FILL_1__1597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1315_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_752_),
    .Y(_807_)
);

INVX1 _1244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_391_),
    .Y(_392_)
);

FILL FILL_0__992_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf1),
    .B(_y[10]),
    .Y(_155_)
);

FILL FILL_0__1704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1124_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1893_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_43_),
    .CLK(clk_bF$buf3),
    .Q(Yin2[3])
);

AOI21X1 _1473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_505_),
    .B(_501_),
    .C(_508_),
    .Y(_619_)
);

OAI21X1 _1053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_166_),
    .B(_187_),
    .C(_204_),
    .Y(_205_)
);

FILL FILL_4__979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1284_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_130_),
    .B(_187_),
    .C(_585_),
    .Y(_674_)
);

INVX1 _1109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_256_),
    .Y(_259_)
);

FILL FILL_3__1773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1353_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_367_),
    .B(_429_),
    .C(_424_),
    .Y(_430_)
);

FILL FILL_0__1742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1409_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_898_),
    .Y(_899_)
);

OAI21X1 _1338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_393_),
    .B(_396_),
    .C(_394_),
    .Y(_485_)
);

FILL FILL_3__1582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1162_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_241_),
    .B(_231_),
    .Y(_242_)
);

FILL FILL_0__1551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1218_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _1567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_637_),
    .B(_711_),
    .Y(_712_)
);

NAND2X1 _1147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_295_),
    .B(_296_),
    .Y(_297_)
);

FILL FILL_1__929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1027_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _1796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_68_),
    .B(_70_),
    .Y(_71_)
);

AOI21X1 _1376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_517_),
    .B(_522_),
    .C(_446_),
    .Y(_523_)
);

FILL FILL_4__1516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1256_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin1[1]),
    .Y(_334_)
);

FILL FILL_1__967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100650x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1004_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_840_),
    .B(_787_),
    .Y(_842_)
);

AOI21X1 _1279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_422_),
    .B(_421_),
    .C(_420_),
    .Y(_427_)
);

FILL FILL_2__1913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100950x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1072_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf4),
    .Y(Vld)
);

FILL FILL_3__963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1159_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_238_),
    .B(_236_),
    .C(_220_),
    .Y(_239_)
);

FILL FILL_2__1722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1709_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_804_),
    .B(_808_),
    .C(_860_),
    .Y(_862_)
);

INVX1 _1300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_421_),
    .Y(_447_)
);

FILL FILL_1__1462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1395_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin3[3]),
    .B(_78_),
    .Y(_85_)
);

FILL FILL_1__1556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1205_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_743_),
    .B(_746_),
    .C(_766_),
    .Y(_767_)
);

OAI21X1 _1203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_347_),
    .B(_346_),
    .C(_310_),
    .Y(_352_)
);

FILL FILL_0__951_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf0),
    .B(_128_),
    .C(_129_),
    .Y(_920_[2])
);

FILL FILL_1__1785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100650x23550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1503_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1852_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2_),
    .CLK(clk_bF$buf1),
    .Q(XinH[2])
);

NAND2X1 _1432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[0]),
    .B(Cin[4]),
    .Y(_578_)
);

INVX1 _1012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[0]),
    .Y(_166_)
);

FILL FILL_1__1594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1069_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1908_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(LoadCtl[1]),
    .CLK(clk_bF$buf2),
    .Q(LoadCtl[2])
);

FILL FILL_3__1732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1312_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_727_),
    .B(_803_),
    .Y(_804_)
);

NAND3X1 _1241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_388_),
    .B(_385_),
    .C(_387_),
    .Y(_389_)
);

OAI21X1 _992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf2),
    .B(_106_),
    .C(_153_),
    .Y(_12_)
);

FILL FILL_2__1719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1298_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_858_),
    .B(_855_),
    .Y(_859_)
);

FILL FILL_3__1541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1039_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1890_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_40_),
    .CLK(clk_bF$buf3),
    .Q(Yin2[0])
);

OAI21X1 _1470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_611_),
    .B(_610_),
    .C(_577_),
    .Y(_616_)
);

OAI21X1 _1050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_192_),
    .B(_194_),
    .C(_197_),
    .Y(_202_)
);

FILL FILL_4__976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1281_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[1]),
    .B(Cin[4]),
    .Y(_671_)
);

NAND3X1 _1106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[0]),
    .B(Cin_0_bF$buf1),
    .C(Yin1[0]),
    .Y(_256_)
);

FILL FILL_3__998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1268_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1406_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_895_),
    .B(_890_),
    .Y(_896_)
);

OAI21X1 _1335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_126_),
    .B(_187_),
    .C(_474_),
    .Y(_482_)
);

FILL FILL_1__1497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1635_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100350x58650 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_695_),
    .B(_702_),
    .C(_640_),
    .Y(_709_)
);

NAND3X1 _1144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_244_),
    .B(_289_),
    .C(_293_),
    .Y(_294_)
);

FILL FILL_1__926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_917_),
    .B(_919_),
    .C(_57_),
    .Y(_68_)
);

AOI21X1 _1373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_515_),
    .B(_514_),
    .C(_513_),
    .Y(_520_)
);

FILL FILL_4__1513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1184_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf2),
    .B(_237_),
    .C(_103_),
    .Y(_55_)
);

NAND2X1 _1429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_569_),
    .B(_574_),
    .Y(_575_)
);

NAND2X1 _1009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[15]),
    .B(_148__bF$buf1),
    .Y(_164_)
);

FILL FILL_3__1673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1253_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_329_),
    .B(_325_),
    .C(_330_),
    .Y(_331_)
);

FILL FILL_1__964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100950x39150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1309_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_800_),
    .B(_732_),
    .Y(_801_)
);

AND2X2 _1238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[0]),
    .B(Cin[3]),
    .Y(_386_)
);

FILL FILL_0__986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1062_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[7]),
    .B(_148__bF$buf4),
    .Y(_152_)
);

FILL FILL100650x11850 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1118_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1887_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_37_),
    .CLK(clk_bF$buf3),
    .Q(Yin3[1])
);

NAND3X1 _1467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_575_),
    .B(_605_),
    .C(_612_),
    .Y(_613_)
);

OAI21X1 _1047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_192_),
    .B(_194_),
    .C(_198_),
    .Y(_199_)
);

FILL FILL_3__1291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1347_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_837_),
    .B(_838_),
    .C(_836_),
    .Y(_839_)
);

NAND3X1 _1276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_419_),
    .B(_423_),
    .C(_369_),
    .Y(_424_)
);

FILL FILL_0__1736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1156_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[3]),
    .B(Cin_0_bF$buf2),
    .C(_235_),
    .Y(_236_)
);

FILL FILL_0__1545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100350x46950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1324_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_724_),
    .B(_742_),
    .C(_737_),
    .Y(_743_)
);

OAI21X1 _1179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_327_),
    .B(_326_),
    .C(_324_),
    .Y(_328_)
);

FILL FILL_2__1813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1392_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin3[2]),
    .B(_78_),
    .Y(_83_)
);

FILL FILL_1__1553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL101250x82050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1609_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_759_),
    .B(_684_),
    .C(_757_),
    .Y(_764_)
);

NAND3X1 _1200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_309_),
    .B(_344_),
    .C(_348_),
    .Y(_349_)
);

OAI21X1 _951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf1),
    .B(_126_),
    .C(_127_),
    .Y(_920_[1])
);

FILL FILL_1__1782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100950x27450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100650x85950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1066_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1905_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_55_),
    .CLK(clk_bF$buf2),
    .Q(XinHL[3])
);

FILL FILL_3__957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1295_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[2]),
    .B(Cin[5]),
    .Y(_856_)
);

FILL FILL_1__1456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1105_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_662_),
    .B(_667_),
    .Y(_668_)
);

INVX1 _1103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_252_),
    .Y(_253_)
);

FILL FILL_3__995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1403_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_130_),
    .B(_891_),
    .Y(_893_)
);

INVX1 _1332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_473_),
    .Y(_479_)
);

FILL FILL_1__1494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1389_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin3[1]),
    .B(_78_),
    .Y(_81_)
);

FILL FILL_3__1632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1212_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_705_),
    .B(_704_),
    .C(_640_),
    .Y(_706_)
);

NAND3X1 _1141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_286_),
    .B(_287_),
    .C(_290_),
    .Y(_291_)
);

FILL FILL_1__923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1198_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_759_),
    .B(_684_),
    .C(_760_),
    .Y(_761_)
);

FILL FILL_0__945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1021_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf2),
    .B(_124_),
    .C(_125_),
    .Y(_920_[0])
);

FILL FILL_1__1779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1359_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148__bF$buf0),
    .B(_65_),
    .C(_910_),
    .Y(_34_)
);

NAND3X1 _1370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_512_),
    .B(_516_),
    .C(_448_),
    .Y(_517_)
);

FILL FILL_4__1510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1917_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf1),
    .B(Xin[2]),
    .Y(_102_)
);

NAND3X1 _1426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_565_),
    .B(_564_),
    .C(_562_),
    .Y(_572_)
);

NAND2X1 _1006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf0),
    .B(_y[14]),
    .Y(_162_)
);

FILL FILL_3__1670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL101250x70350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1657_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1306_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[1]),
    .B(Cin[6]),
    .C(XinH[2]),
    .D(Cin[5]),
    .Y(_798_)
);

AND2X2 _1235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_375_),
    .B(_381_),
    .Y(_383_)
);

FILL FILL_0__983_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[6]),
    .B(_148__bF$buf4),
    .Y(_150_)
);

FILL FILL_1__1397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100950x15750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1115_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1884_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_34_),
    .CLK(clk_bF$buf6),
    .Q(_y[14])
);

AOI21X1 _1464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_608_),
    .B(_609_),
    .C(_599_),
    .Y(_610_)
);

OAI21X1 _1044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_190_),
    .B(_191_),
    .C(_195_),
    .Y(_196_)
);

FILL FILL_0__1504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1344_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_720_),
    .B(_775_),
    .C(_835_),
    .Y(_836_)
);

NAND3X1 _1273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_408_),
    .B(_415_),
    .C(_412_),
    .Y(_421_)
);

FILL FILL_0__1733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1084_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _1749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_856_),
    .B(_857_),
    .C(_854_),
    .D(_855_),
    .Y(_890_)
);

NAND2X1 _1329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[1]),
    .B(Cin[2]),
    .Y(_476_)
);

FILL FILL_3__1573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1153_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_219_),
    .Y(_233_)
);

FILL FILL_0__1542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1209_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_695_),
    .B(_702_),
    .C(_641_),
    .Y(_703_)
);

AOI22X1 _1138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_228_),
    .B(_285_),
    .C(_287_),
    .D(_286_),
    .Y(_288_)
);

FILL FILL_3__1382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100950x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1018_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_916_),
    .B(_61_),
    .Y(_63_)
);

NAND3X1 _1367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_501_),
    .B(_505_),
    .C(_508_),
    .Y(_514_)
);

FILL FILL99750x31350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1247_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_585_),
    .B(_672_),
    .Y(_740_)
);

NAND3X1 _1176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[1]),
    .B(Cin_0_bF$buf3),
    .C(Yin1[1]),
    .Y(_325_)
);

FILL FILL_1__958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1063_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1902_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_52_),
    .CLK(clk_bF$buf4),
    .Q(XinHL[0])
);

FILL FILL_3__954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1224_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_565_),
    .B(_554_),
    .Y(_644_)
);

AOI21X1 _1079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_224_),
    .B(_227_),
    .C(_219_),
    .Y(_230_)
);

FILL FILL_2__1713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL99450x66450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1292_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_796_),
    .B(_798_),
    .C(_801_),
    .Y(_853_)
);

FILL FILL_1__1453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1509_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_658_),
    .B(_659_),
    .C(_656_),
    .Y(_665_)
);

INVX1 _1100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_216_),
    .Y(_250_)
);

FILL FILL_3__992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL101250x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1386_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin3[0]),
    .B(_78_),
    .Y(_79_)
);

FILL FILL_1__1547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1195_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_757_),
    .B(_749_),
    .Y(_758_)
);

FILL FILL_0__942_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_105_),
    .B(_122_),
    .C(_123_),
    .Y(_921_[3])
);

FILL FILL_1__1776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1914_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf3),
    .B(_166_),
    .C(_100_),
    .Y(_52_)
);

NAND3X1 _1423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549_),
    .B(_568_),
    .C(_563_),
    .Y(_569_)
);

NAND2X1 _1003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[13]),
    .B(_148__bF$buf0),
    .Y(_160_)
);

FILL FILL_1__1585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1303_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_725_),
    .B(_726_),
    .C(_733_),
    .Y(_795_)
);

NAND2X1 _1232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[2]),
    .B(Cin[4]),
    .Y(_380_)
);

FILL FILL_0__980_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf4),
    .B(_146_),
    .C(_147_),
    .Y(_9_)
);

FILL FILL_1__1394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1289_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_794_),
    .B(_827_),
    .C(_833_),
    .Y(_850_)
);

FILL FILL_3__1532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1112_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1881_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_31_),
    .CLK(clk_bF$buf6),
    .Q(_y[11])
);

OAI21X1 _1461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_484_),
    .B(_606_),
    .C(_503_),
    .Y(_607_)
);

NAND3X1 _1041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[2]),
    .B(Cin_0_bF$buf2),
    .C(Yin0[2]),
    .Y(_193_)
);

FILL FILL_4__967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1098_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_644_),
    .B(_661_),
    .C(_657_),
    .Y(_662_)
);

FILL FILL_3__989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1259_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_790_),
    .B(_831_),
    .C(_832_),
    .Y(_833_)
);

OAI21X1 _1270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_417_),
    .B(_416_),
    .C(_415_),
    .Y(_418_)
);

FILL FILL_2__1748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1817_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_881_),
    .Y(_887_)
);

NAND2X1 _1326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[3]),
    .B(Cin[4]),
    .Y(_473_)
);

FILL FILL_3__1570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1206_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_669_),
    .B(_611_),
    .C(_685_),
    .Y(_700_)
);

NAND3X1 _1135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_218_),
    .B(_228_),
    .C(_240_),
    .Y(_285_)
);

FILL FILL_1__1297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1015_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_917_),
    .B(_59_),
    .Y(_60_)
);

OAI21X1 _1364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_510_),
    .B(_509_),
    .C(_508_),
    .Y(_511_)
);

FILL FILL101250x23550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1244_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_729_),
    .B(_734_),
    .C(_736_),
    .Y(_737_)
);

OAI21X1 _1173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_257_),
    .B(_254_),
    .C(_256_),
    .Y(_322_)
);

FILL FILL_1__955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1213_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_743_),
    .B(_746_),
    .Y(_792_)
);

XNOR2X1 _1229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_374_),
    .B(_376_),
    .Y(_377_)
);

FILL FILL_0__977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1109_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1878_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_28_),
    .CLK(clk_bF$buf5),
    .Q(_y[8])
);

OAI21X1 _1458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_602_),
    .B(_603_),
    .C(_599_),
    .Y(_604_)
);

INVX1 _1038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[1]),
    .Y(_190_)
);

FILL FILL_3__1282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1338_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_747_),
    .B(_762_),
    .C(_758_),
    .Y(_830_)
);

OAI21X1 _1267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_321_),
    .B(_414_),
    .C(_341_),
    .Y(_415_)
);

FILL FILL_3__1091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1147_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_640_),
    .Y(_641_)
);

NAND3X1 _1076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_225_),
    .B(_221_),
    .C(_226_),
    .Y(_227_)
);

FILL FILL_2__1710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1383_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[0]),
    .Y(_76_)
);

FILL FILL_1__1544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL101250x11850 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_467_),
    .B(_469_),
    .Y(_545_)
);

FILL FILL_2__1613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1192_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_585_),
    .B(_751_),
    .C(_753_),
    .Y(_755_)
);

NAND2X1 _942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[2]),
    .B(_120_),
    .Y(_121_)
);

FILL FILL_1__1773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1911_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert10 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf1)
);

FILL FILL_1__1829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1409_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert11 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf0)
);

NAND2X1 _1840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf2),
    .B(Yin[3]),
    .Y(_99_)
);

NOR2X1 _1420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_474_),
    .B(_476_),
    .Y(_566_)
);

NAND2X1 _1000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf2),
    .B(_y[12]),
    .Y(_158_)
);

FILL FILL_1__1582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1218_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf1),
    .B(_144_),
    .C(_145_),
    .Y(_8_)
);

FILL FILL_1__1391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1286_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_834_),
    .B(_777_),
    .Y(_847_)
);

FILL FILL_1__1447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1095_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_648_),
    .B(_647_),
    .C(_645_),
    .Y(_659_)
);

FILL FILL_3__986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1814_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_884_),
    .B(_881_),
    .Y(_885_)
);

NAND2X1 _1323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_466_),
    .B(_469_),
    .Y(_470_)
);

FILL FILL_1__1485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1203_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_575_),
    .B(_696_),
    .C(_615_),
    .Y(_697_)
);

NAND2X1 _1132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_273_),
    .B(_277_),
    .Y(_282_)
);

FILL FILL_1__1294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1189_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_585_),
    .B(_751_),
    .Y(_752_)
);

FILL FILL_0__936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1012_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf4),
    .B(y[2]),
    .C(_110_),
    .D(y[6]),
    .Y(_119_)
);

OR2X2 _1781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_56_),
    .B(_919_),
    .Y(_57_)
);

OAI21X1 _1361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_390_),
    .B(_507_),
    .C(_410_),
    .Y(_508_)
);

FILL FILL_4__1501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL101250x85950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1172_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf3),
    .B(_80_),
    .C(_97_),
    .Y(_49_)
);

OAI21X1 _1417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_557_),
    .B(_560_),
    .C(_562_),
    .Y(_563_)
);

FILL FILL_3__1661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1159_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_733_),
    .B(_731_),
    .C(_730_),
    .Y(_734_)
);

OAI22X1 _1170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_271_),
    .B(_275_),
    .C(_237_),
    .D(_187_),
    .Y(_319_)
);

FILL FILL_1__952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1717_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_721_),
    .B(_788_),
    .C(_774_),
    .Y(_789_)
);

NOR2X1 _1226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_370_),
    .B(_373_),
    .Y(_374_)
);

FILL FILL_0__974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1050_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf3),
    .B(_142_),
    .C(_143_),
    .Y(_7_)
);

FILL FILL_1__1388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1106_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1875_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_25_),
    .CLK(clk_bF$buf0),
    .Q(_y[5])
);

NAND2X1 _1455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_591_),
    .B(_600_),
    .Y(_601_)
);

INVX4 _1035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[2]),
    .Y(_187_)
);

FILL FILL_1__1197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1335_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_821_),
    .B(_825_),
    .Y(_827_)
);

NAND3X1 _1264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_410_),
    .B(_411_),
    .C(_409_),
    .Y(_412_)
);

FILL FILL100050x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1144_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_625_),
    .Y(_638_)
);

OAI21X1 _1073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_223_),
    .B(_222_),
    .C(_220_),
    .Y(_224_)
);

FILL FILL_0__1533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1113_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_692_),
    .B(_693_),
    .C(_691_),
    .Y(_694_)
);

NAND3X1 _1129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_262_),
    .B(_265_),
    .C(_278_),
    .Y(_279_)
);

FILL FILL_3__1793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL99750x46950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1009_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_128_),
    .B(_456_),
    .C(_893_),
    .Y(_918_)
);

NAND3X1 _1358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_503_),
    .B(_504_),
    .C(_502_),
    .Y(_505_)
);

FILL FILL_3__1182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1238_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_726_),
    .Y(_731_)
);

NAND3X1 _1167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_311_),
    .B(_313_),
    .C(_315_),
    .Y(_316_)
);

FILL FILL_1__949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1047_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _1396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_540_),
    .B(_541_),
    .C(_534_),
    .D(_440_),
    .Y(_542_)
);

FILL FILL_2__1610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1635_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1283_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_y[12]),
    .B(_148__bF$buf2),
    .Y(_844_)
);

FILL FILL_1__1444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__961_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_376_),
    .B(_374_),
    .Y(_446_)
);

FILL FILL_2__1513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1092_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_578_),
    .B(_655_),
    .C(_586_),
    .Y(_656_)
);

FILL FILL_3__983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100950x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1309_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_850_),
    .Y(_882_)
);

NAND3X1 _1320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_463_),
    .B(_462_),
    .C(_460_),
    .Y(_467_)
);

FILL FILL_1__1482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100350x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1186_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_748_),
    .B(_591_),
    .C(_684_),
    .Y(_749_)
);

FILL FILL_0__933_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[10]),
    .Y(_116_)
);

FILL FILL_1__1767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1416_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf2),
    .B(Yin[0]),
    .Y(_96_)
);

AOI21X1 _1414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_558_),
    .B(_559_),
    .C(_550_),
    .Y(_560_)
);

FILL FILL_4_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1714_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_y[11]),
    .Y(_786_)
);

AND2X2 _1223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[1]),
    .B(Cin[6]),
    .Y(_371_)
);

FILL FILL_0__971_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf3),
    .B(_140_),
    .C(_141_),
    .Y(_6_)
);

FILL FILL_1__1385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1103_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1872_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_22_),
    .CLK(clk_bF$buf0),
    .Q(_y[2])
);

NAND3X1 _1452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_597_),
    .B(_589_),
    .C(_594_),
    .Y(_598_)
);

OAI21X1 _1032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148__bF$buf1),
    .B(_183_),
    .C(_184_),
    .Y(_21_)
);

FILL FILL_4__958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1089_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_648_),
    .Y(_653_)
);

FILL FILL_3__1752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1332_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_820_),
    .Y(_824_)
);

AND2X2 _1261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_384_),
    .B(_389_),
    .Y(_409_)
);

FILL FILL_2__1739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1808_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_875_),
    .Y(_879_)
);

AOI21X1 _1317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_385_),
    .B(_388_),
    .C(_382_),
    .Y(_464_)
);

FILL FILL_3__1561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1059_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148__bF$buf2),
    .B(_635_),
    .C(_539_),
    .Y(_28_)
);

NAND3X1 _1070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[3]),
    .B(Cin_0_bF$buf2),
    .C(Yin0[3]),
    .Y(_221_)
);

FILL FILL_2__1548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1617_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_662_),
    .B(_667_),
    .Y(_691_)
);

OAI21X1 _1126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_190_),
    .B(_275_),
    .C(_269_),
    .Y(_276_)
);

FILL FILL_3__1790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1006_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_914_),
    .B(_912_),
    .Y(_915_)
);

AND2X2 _1355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_483_),
    .B(_478_),
    .Y(_502_)
);

FILL FILL_1__1097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1235_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_646_),
    .B(_727_),
    .Y(_728_)
);

OAI21X1 _1164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237_),
    .B(_187_),
    .C(_312_),
    .Y(_313_)
);

FILL FILL_1__946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1044_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_y[8]),
    .B(_148__bF$buf2),
    .Y(_539_)
);

FILL FILL_0__1433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__962_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1869_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_19_),
    .CLK(clk_bF$buf6),
    .Q(y[15])
);

AOI21X1 _1449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[3]),
    .B(Cin_0_bF$buf0),
    .C(Yin1[3]),
    .Y(_595_)
);

NAND2X1 _1029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_165_),
    .B(_180_),
    .Y(_182_)
);

FILL FILL_3__1693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1329_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_811_),
    .B(_815_),
    .C(_820_),
    .Y(_821_)
);

AOI21X1 _1258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_405_),
    .B(_404_),
    .C(_393_),
    .Y(_406_)
);

FILL FILL_3__1082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1138_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_631_),
    .B(_632_),
    .C(_630_),
    .Y(_633_)
);

NOR2X1 _1067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_217_),
    .B(_216_),
    .Y(_218_)
);

FILL FILL_2__1701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1367_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_440_),
    .Y(_443_)
);

FILL FILL_2__1510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100050x31350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1183_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_723_),
    .B(_744_),
    .C(_745_),
    .Y(_746_)
);

FILL FILL_0__930_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[2]),
    .B(y[13]),
    .C(_113_),
    .Y(_114_)
);

FILL FILL_1__1764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1344_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_347_),
    .B(_346_),
    .C(_345_),
    .Y(_348_)
);

FILL FILL_2__1833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1239_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_82_),
    .B(_91_),
    .C(_94_),
    .Y(_46_)
);

AOI21X1 _1411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_554_),
    .B(_556_),
    .C(_551_),
    .Y(_557_)
);

FILL FILL_1__1573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100350x70350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1209_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_717_),
    .B(_783_),
    .Y(_784_)
);

INVX1 _1220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_351_),
    .Y(_368_)
);

OAI21X1 _971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf1),
    .B(_138_),
    .C(_139_),
    .Y(_5_)
);

FILL FILL_1__1382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1086_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_645_),
    .Y(_650_)
);

FILL FILL_3__977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1805_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_851_),
    .B(_873_),
    .C(_875_),
    .Y(_876_)
);

OAI21X1 _1314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_455_),
    .B(_459_),
    .C(_460_),
    .Y(_461_)
);

FILL FILL_1__1476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1614_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_589_),
    .B(_687_),
    .C(_608_),
    .Y(_688_)
);

NAND3X1 _1123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_),
    .B(_267_),
    .C(_270_),
    .Y(_273_)
);

FILL FILL_1__1285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1003_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_848_),
    .B(_846_),
    .C(_911_),
    .Y(_912_)
);

AOI21X1 _1352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_489_),
    .B(_491_),
    .C(_487_),
    .Y(_499_)
);

FILL FILL_1__1094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1163_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf4),
    .B(_109_),
    .C(Yin1[1]),
    .Y(_93_)
);

NAND2X1 _1408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_552_),
    .B(_553_),
    .Y(_554_)
);

FILL FILL_3__1652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1232_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[3]),
    .B(Cin[7]),
    .Y(_725_)
);

AOI21X1 _1161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_278_),
    .B(_262_),
    .C(_281_),
    .Y(_310_)
);

FILL FILL_1__943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1708_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_768_),
    .B(_772_),
    .C(_721_),
    .Y(_781_)
);

OAI21X1 _1217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_362_),
    .B(_299_),
    .C(_359_),
    .Y(_365_)
);

FILL FILL_0__965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1041_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf3),
    .B(_136_),
    .C(_137_),
    .Y(_4_)
);

FILL FILL_1__1799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1379_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_534_),
    .Y(_537_)
);

FILL FILL_2__1448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1517_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1866_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_16_),
    .CLK(clk_bF$buf6),
    .Q(y[12])
);

INVX1 _1446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_591_),
    .Y(_592_)
);

NAND3X1 _1026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_173_),
    .B(_178_),
    .C(_177_),
    .Y(_179_)
);

FILL FILL_3__1690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1326_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_756_),
    .B(_817_),
    .Y(_818_)
);

INVX1 _1255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin1[2]),
    .Y(_403_)
);

FILL FILL_0__1715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1135_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_524_),
    .B(_526_),
    .C(_629_),
    .Y(_630_)
);

NAND2X1 _1064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[1]),
    .B(Cin[3]),
    .Y(_215_)
);

FILL FILL_0__1524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1364_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf4),
    .B(_440_),
    .Y(_441_)
);

FILL FILL_4__1433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1914_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148__bF$buf0),
    .B(_159_),
    .C(_909_),
    .D(_907_),
    .Y(_33_)
);

NAND3X1 _1349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_494_),
    .B(_493_),
    .C(_495_),
    .Y(_496_)
);

FILL FILL_3__1593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1229_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691_),
    .B(_693_),
    .C(_686_),
    .Y(_722_)
);

INVX1 _1158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_269_),
    .Y(_307_)
);

FILL FILL_0__1618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100350x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1038_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_533_),
    .B(_528_),
    .Y(_534_)
);

FILL FILL_2__1601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1198_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_105_),
    .B(_108_),
    .C(_111_),
    .Y(_921_[0])
);

FILL FILL_1__1761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1267_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_282_),
    .B(_280_),
    .C(_265_),
    .Y(_345_)
);

FILL FILL_1__978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1076_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[0]),
    .Y(Cin_0_bF$buf3)
);

BUFX2 BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[0]),
    .Y(Cin_0_bF$buf2)
);

BUFX2 BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[0]),
    .Y(Cin_0_bF$buf1)
);

BUFX2 BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[0]),
    .Y(Cin_0_bF$buf0)
);

BUFX2 BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf4)
);

BUFX2 BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf3)
);

BUFX2 BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf2)
);

BUFX2 BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf1)
);

FILL FILL100650x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1083_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_555_),
    .B(_646_),
    .Y(_647_)
);

FILL FILL_3__974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1244_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_y[4]),
    .B(_148__bF$buf3),
    .Y(_249_)
);

FILL FILL_2__1733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1802_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_872_),
    .B(_852_),
    .C(_869_),
    .Y(_873_)
);

OAI21X1 _1311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_271_),
    .B(_304_),
    .C(_371_),
    .Y(_458_)
);

FILL FILL_1__1473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1109_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_684_),
    .B(_683_),
    .Y(_685_)
);

NAND2X1 _1120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_268_),
    .B(_269_),
    .Y(_270_)
);

FILL FILL_1__1282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100350x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1000_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[1]),
    .Y(_109_)
);

FILL FILL_1__1758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100350x23550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1160_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_110_),
    .Y(_91_)
);

INVX1 _1405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_550_),
    .Y(_551_)
);

FILL FILL_1__1567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1705_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _1634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_698_),
    .B(_701_),
    .C(_643_),
    .Y(_778_)
);

NOR2X1 _1214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_362_),
    .B(_360_),
    .Y(_363_)
);

FILL FILL_0__962_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_130_),
    .B(_110_),
    .C(_135_),
    .Y(_3_)
);

FILL FILL_1__1796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1514_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1863_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_13_),
    .CLK(clk_bF$buf5),
    .Q(y[9])
);

NAND2X1 _1443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_583_),
    .B(_588_),
    .Y(_589_)
);

OAI21X1 _1023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172_),
    .B(_174_),
    .C(_175_),
    .Y(_176_)
);

FILL FILL_4__949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1254_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_921_[3]),
    .Y(Yout[3])
);

FILL FILL_3__1743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1323_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_813_),
    .B(_814_),
    .C(_812_),
    .Y(_815_)
);

NAND3X1 _1252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_398_),
    .B(_394_),
    .C(_399_),
    .Y(_400_)
);

FILL FILL_0__1712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1063_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_860_),
    .B(_853_),
    .Y(_870_)
);

AOI21X1 _1308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_452_),
    .B(_454_),
    .C(_450_),
    .Y(_455_)
);

FILL FILL_3__1552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1132_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_545_),
    .B(_625_),
    .C(_626_),
    .Y(_627_)
);

NAND2X1 _1061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_y[3]),
    .B(_148__bF$buf3),
    .Y(_212_)
);

FILL FILL_0__1521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1608_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_681_),
    .Y(_682_)
);

INVX1 _1117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_266_),
    .Y(_267_)
);

FILL FILL_3__1781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1279_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_436_),
    .B(_437_),
    .C(_354_),
    .Y(_438_)
);

FILL FILL_4__1430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100350x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1417_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887_),
    .B(_888_),
    .C(_906_),
    .Y(_907_)
);

INVX1 _1346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_),
    .Y(_493_)
);

FILL FILL_3__1590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1226_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_641_),
    .B(_718_),
    .C(_704_),
    .Y(_719_)
);

INVX1 _1155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[5]),
    .Y(_304_)
);

FILL FILL_1__937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100650x39150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1035_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_524_),
    .B(_525_),
    .C(_526_),
    .Y(_531_)
);

FILL FILL100350x11850 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1264_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_333_),
    .B(_337_),
    .C(_323_),
    .Y(_342_)
);

FILL FILL_1__975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1814_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_795_),
    .Y(_812_)
);

OAI21X1 _1249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_396_),
    .B(_395_),
    .C(_393_),
    .Y(_397_)
);

FILL FILL_0__997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100950x78150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1129_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1898_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_48_),
    .CLK(clk_bF$buf2),
    .Q(Yin0[0])
);

NAND3X1 _1478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_546_),
    .B(_623_),
    .C(_618_),
    .Y(_624_)
);

NAND3X1 _1058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_186_),
    .B(_208_),
    .C(_205_),
    .Y(_210_)
);

FILL FILL_0__1518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1358_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_366_),
    .B(_434_),
    .C(_430_),
    .Y(_435_)
);

FILL FILL_2__1501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1167_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_246_),
    .Y(_247_)
);

FILL FILL_2__1730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100050x46950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1174_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[8]),
    .Y(_106_)
);

FILL FILL_1__1755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100650x27450 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_750_),
    .B(_86_),
    .C(_89_),
    .Y(_42_)
);

AOI21X1 _1402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_513_),
    .B(_515_),
    .C(_547_),
    .Y(_548_)
);

FILL FILL_1__1564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1702_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_771_),
    .B(_770_),
    .C(_722_),
    .Y(_775_)
);

INVX1 _1211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_359_),
    .Y(_360_)
);

NAND2X1 _962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[2]),
    .B(_110_),
    .Y(_134_)
);

FILL FILL_1__1793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1268_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1009_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1860_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_10_),
    .CLK(clk_bF$buf5),
    .Q(y[6])
);

NAND2X1 _1440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_480_),
    .B(_585_),
    .Y(_586_)
);

NAND3X1 _1020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[1]),
    .B(Cin_0_bF$buf1),
    .C(Yin0[1]),
    .Y(_173_)
);

FILL FILL_4__946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100950x66450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1077_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_921_[0]),
    .Y(Yout[0])
);

FILL FILL_3__968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1060_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_865_),
    .B(_864_),
    .Y(_867_)
);

NAND2X1 _1305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_371_),
    .B(_451_),
    .Y(_452_)
);

FILL FILL_1__1467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1605_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_676_),
    .B(_678_),
    .C(_677_),
    .Y(_679_)
);

OAI21X1 _1114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254_),
    .B(_259_),
    .C(_257_),
    .Y(_264_)
);

FILL FILL_1__1696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1414_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_901_),
    .B(_903_),
    .Y(_904_)
);

NAND2X1 _1343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[3]),
    .B(Cin_0_bF$buf0),
    .Y(_490_)
);

FILL FILL_1__1085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1154_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[1]),
    .B(_86_),
    .Y(_88_)
);

FILL FILL_3__1643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1223_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_711_),
    .B(_634_),
    .Y(_716_)
);

NAND2X1 _1152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_y[5]),
    .B(_148__bF$buf3),
    .Y(_301_)
);

FILL FILL_1__934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1383_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_771_),
    .B(_770_),
    .C(_769_),
    .Y(_772_)
);

AOI21X1 _1208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_348_),
    .B(_344_),
    .C(_309_),
    .Y(_357_)
);

FILL FILL_0__956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1032_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_124_),
    .B(_110_),
    .C(_132_),
    .Y(_0_)
);

OAI21X1 _1381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_527_),
    .B(_523_),
    .C(_445_),
    .Y(_528_)
);

FILL FILL100650x15750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1508_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1857_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_7_),
    .CLK(clk_bF$buf4),
    .Q(y[3])
);

NAND3X1 _1437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_578_),
    .B(_580_),
    .C(_582_),
    .Y(_583_)
);

NAND2X1 _1017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_y[0]),
    .B(_148__bF$buf4),
    .Y(_171_)
);

FILL FILL_3__1681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1179_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_321_),
    .B(_332_),
    .C(_338_),
    .Y(_339_)
);

FILL FILL_1__972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1317_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_801_),
    .B(_799_),
    .C(_797_),
    .Y(_809_)
);

NAND3X1 _1246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[2]),
    .B(Cin_0_bF$buf3),
    .C(Yin1[2]),
    .Y(_394_)
);

FILL FILL_0__994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1070_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf0),
    .B(_y[11]),
    .Y(_156_)
);

FILL FILL_0__1706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1126_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1895_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_45_),
    .CLK(clk_bF$buf4),
    .Q(Yin1[1])
);

AOI21X1 _1475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_615_),
    .B(_616_),
    .C(_614_),
    .Y(_621_)
);

INVX1 _1055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_206_),
    .Y(_207_)
);

FILL FILL_4__1615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1355_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_426_),
    .B(_423_),
    .C(_419_),
    .Y(_432_)
);

FILL FILL_4__1844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1164_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_208_),
    .B(_203_),
    .C(_231_),
    .D(_241_),
    .Y(_244_)
);

FILL FILL_4__1653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1714_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148__bF$buf2),
    .B(_712_),
    .C(_713_),
    .Y(_29_)
);

NAND3X1 _1149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_294_),
    .B(_246_),
    .C(_297_),
    .Y(_299_)
);

FILL FILL_3__1393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1029_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_72_),
    .B(_67_),
    .Y(_73_)
);

NAND3X1 _1378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_516_),
    .B(_512_),
    .C(_519_),
    .Y(_525_)
);

FILL FILL_0__1838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL99750x70350 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_126_),
    .B(_167_),
    .C(Yin1[1]),
    .Y(_336_)
);

FILL FILL_1__969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1074_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_920_[1]),
    .Y(Xout[1])
);

FILL FILL_3__965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1304_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin3[0]),
    .Y(_864_)
);

NAND2X1 _1302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[0]),
    .B(Cin[7]),
    .Y(_449_)
);

FILL FILL_1__1464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1602_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_671_),
    .Y(_676_)
);

OAI21X1 _1111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254_),
    .B(_259_),
    .C(_260_),
    .Y(_261_)
);

FILL FILL_1__1693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL101250x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1329_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_863_),
    .B(_900_),
    .C(_899_),
    .Y(_901_)
);

NAND2X1 _1340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[2]),
    .B(Cin[1]),
    .Y(_487_)
);

FILL FILL_1__1082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1397_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_77_),
    .B(_105_),
    .Y(_86_)
);

FILL FILL_3__1640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL101250x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1380_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_689_),
    .B(_668_),
    .C(_692_),
    .Y(_769_)
);

NAND3X1 _1205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_349_),
    .B(_353_),
    .C(_303_),
    .Y(_354_)
);

FILL FILL_0__953_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf0),
    .B(XinHL[3]),
    .Y(_131_)
);

FILL FILL_1__1787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100950x19650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1505_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1854_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4_),
    .CLK(clk_bF$buf1),
    .Q(y[0])
);

NAND3X1 _1434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[2]),
    .B(Cin[2]),
    .C(_579_),
    .Y(_580_)
);

INVX1 _1014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin0[0]),
    .Y(_168_)
);

FILL FILL_1__1596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1314_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_752_),
    .B(_805_),
    .C(_802_),
    .Y(_806_)
);

OAI21X1 _1243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_324_),
    .B(_327_),
    .C(_325_),
    .Y(_391_)
);

FILL FILL_0__991_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf1),
    .B(_112_),
    .C(_154_),
    .Y(_13_)
);

FILL FILL_0__1703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1054_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853_),
    .B(_860_),
    .Y(_861_)
);

FILL FILL_3__1543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1123_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1892_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_42_),
    .CLK(clk_bF$buf3),
    .Q(Yin2[2])
);

NAND3X1 _1472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_613_),
    .B(_617_),
    .C(_548_),
    .Y(_618_)
);

NAND2X1 _1052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_203_),
    .B(_200_),
    .Y(_204_)
);

FILL FILL_4__1612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1283_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_128_),
    .B(_275_),
    .C(_672_),
    .Y(_673_)
);

NAND3X1 _1108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_256_),
    .B(_257_),
    .C(_255_),
    .Y(_258_)
);

FILL FILL_3__1772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1352_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_427_),
    .B(_428_),
    .C(_426_),
    .Y(_429_)
);

FILL FILL_4__1841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1408_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_872_),
    .B(_867_),
    .C(_897_),
    .Y(_898_)
);

NAND2X1 _1337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_478_),
    .B(_483_),
    .Y(_484_)
);

FILL FILL_3__1581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1079_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_232_),
    .B(_228_),
    .C(_240_),
    .Y(_241_)
);

FILL FILL_4__1650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1217_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_707_),
    .B(_710_),
    .Y(_711_)
);

NAND2X1 _1146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_289_),
    .B(_293_),
    .Y(_296_)
);

FILL FILL_1__928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1026_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_69_),
    .B(Yin3[3]),
    .Y(_70_)
);

OAI21X1 _1375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_520_),
    .B(_521_),
    .C(_519_),
    .Y(_522_)
);

FILL FILL_0__1835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1255_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_330_),
    .B(_325_),
    .C(_329_),
    .Y(_333_)
);

FILL FILL_1__966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100650x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1614_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1889_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_39_),
    .CLK(clk_bF$buf3),
    .Q(Yin3[3])
);

NAND3X1 _1469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_598_),
    .B(_607_),
    .C(_604_),
    .Y(_615_)
);

NAND2X1 _1049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_198_),
    .B(_195_),
    .Y(_201_)
);

FILL FILL_3__1293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__940_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_787_),
    .B(_840_),
    .Y(_841_)
);

OAI21X1 _1278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_309_),
    .B(_425_),
    .C(_351_),
    .Y(_426_)
);

FILL FILL_2__1912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1071_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1910_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(LoadCtl[3]),
    .CLK(clk_bF$buf4),
    .Q(LoadCtl[4])
);

FILL FILL_3__962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1158_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237_),
    .B(_167_),
    .C(Yin0[3]),
    .Y(_238_)
);

FILL FILL_2__1721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL101250x39150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL99750x23550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1394_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[3]),
    .Y(_84_)
);

FILL FILL_1__1555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__979_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_764_),
    .B(_765_),
    .Y(_766_)
);

NAND3X1 _1202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_339_),
    .B(_345_),
    .C(_343_),
    .Y(_351_)
);

FILL FILL_0__950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL101250x50850 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf0),
    .B(XinHL[2]),
    .Y(_129_)
);

FILL FILL_1__1784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1259_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1502_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1851_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1_),
    .CLK(clk_bF$buf1),
    .Q(XinH[1])
);

AOI21X1 _1431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_502_),
    .B(_504_),
    .C(_576_),
    .Y(_577_)
);

NAND3X1 _1011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[0]),
    .B(Cin_0_bF$buf1),
    .C(Yin0[0]),
    .Y(_165_)
);

FILL FILL_4__937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1068_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1907_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(LoadCtl_0_bF$buf0),
    .CLK(clk_bF$buf2),
    .Q(LoadCtl[1])
);

FILL FILL_3__959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1229_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[2]),
    .B(Cin[6]),
    .Y(_803_)
);

OAI21X1 _1240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_124_),
    .B(_187_),
    .C(_375_),
    .Y(_388_)
);

NAND2X1 _991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf2),
    .B(_y[8]),
    .Y(_153_)
);

FILL FILL_2__1718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1297_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_856_),
    .B(_857_),
    .Y(_858_)
);

FILL FILL_3__1540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1280_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_599_),
    .B(_609_),
    .C(_669_),
    .Y(_670_)
);

INVX1 _1105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254_),
    .Y(_255_)
);

FILL FILL_3__997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1405_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_894_),
    .B(_892_),
    .Y(_895_)
);

NAND2X1 _1334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_386_),
    .B(_480_),
    .Y(_481_)
);

FILL FILL101250x27450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1214_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_705_),
    .B(_704_),
    .C(_641_),
    .Y(_708_)
);

NAND3X1 _1143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_216_),
    .B(_292_),
    .C(_291_),
    .Y(_293_)
);

FILL FILL_1__925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1374_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_747_),
    .B(_762_),
    .Y(_763_)
);

FILL FILL_0__947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1023_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_916_),
    .B(_61_),
    .C(_66_),
    .Y(_67_)
);

OAI21X1 _1372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_518_),
    .B(_377_),
    .C(_421_),
    .Y(_519_)
);

FILL FILL_0__1832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1919_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf3),
    .B(Xin[3]),
    .Y(_103_)
);

NAND3X1 _1428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_571_),
    .B(_572_),
    .C(_573_),
    .Y(_574_)
);

INVX1 _1008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_y[15]),
    .Y(_163_)
);

FILL FILL_3__1672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1252_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_327_),
    .Y(_330_)
);

FILL FILL_1__963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1308_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[2]),
    .B(Cin[6]),
    .Y(_800_)
);

INVX1 _1237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_380_),
    .Y(_385_)
);

FILL FILL_0__985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1061_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_y[7]),
    .Y(_151_)
);

FILL FILL_1__1399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1117_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1886_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_36_),
    .CLK(clk_bF$buf3),
    .Q(Yin3[0])
);

OAI21X1 _1466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_611_),
    .B(_610_),
    .C(_607_),
    .Y(_612_)
);

INVX1 _1046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_197_),
    .Y(_198_)
);

FILL FILL_3__1290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1346_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_826_),
    .B(_828_),
    .C(_791_),
    .Y(_838_)
);

NAND3X1 _1275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_420_),
    .B(_421_),
    .C(_422_),
    .Y(_423_)
);

FILL FILL_4__1835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1155_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin0[3]),
    .Y(_235_)
);

FILL FILL_4__1644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL101250x15750 (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_915_),
    .B(_64_),
    .Y(_65_)
);

NAND3X1 _1369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_514_),
    .B(_513_),
    .C(_515_),
    .Y(_516_)
);

FILL FILL_3__1193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1249_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_738_),
    .B(_739_),
    .C(_741_),
    .Y(_742_)
);

AOI21X1 _1178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[1]),
    .B(Cin_0_bF$buf3),
    .C(Yin1[1]),
    .Y(_327_)
);

FILL FILL_2__1812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1391_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[2]),
    .Y(_82_)
);

FILL FILL_1__1552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1608_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf1),
    .B(XinHL[1]),
    .Y(_127_)
);

FILL FILL_1__1781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1065_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1904_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_54_),
    .CLK(clk_bF$buf1),
    .Q(XinHL[2])
);

FILL FILL_3__956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1294_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[3]),
    .B(Cin[5]),
    .C(_800_),
    .Y(_855_)
);

FILL FILL_1__1455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1104_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_664_),
    .B(_665_),
    .C(_666_),
    .Y(_667_)
);

OAI21X1 _1102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_220_),
    .B(_223_),
    .C(_221_),
    .Y(_252_)
);

FILL FILL_3__994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1402_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_128_),
    .B(_891_),
    .C(_857_),
    .Y(_892_)
);

NAND3X1 _1331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_473_),
    .B(_475_),
    .C(_477_),
    .Y(_478_)
);

FILL FILL_1__1493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL101250x89850 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1388_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[1]),
    .Y(_80_)
);

FILL FILL_3__1631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1129_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_698_),
    .B(_701_),
    .C(_643_),
    .Y(_705_)
);

AOI21X1 _1140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_218_),
    .B(_240_),
    .C(_229_),
    .Y(_290_)
);

FILL FILL_1__922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1197_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_756_),
    .B(_754_),
    .Y(_760_)
);

FILL FILL_0__944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1020_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf1),
    .B(XinHL[0]),
    .Y(_125_)
);

FILL FILL_1__1778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1916_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf1),
    .B(_190_),
    .C(_101_),
    .Y(_53_)
);

OAI21X1 _1425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_453_),
    .B(_570_),
    .C(_463_),
    .Y(_571_)
);

INVX1 _1005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[14]),
    .Y(_161_)
);

FILL FILL_1__1587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1305_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_796_),
    .Y(_797_)
);

NOR2X1 _1234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_375_),
    .B(_381_),
    .Y(_382_)
);

FILL FILL_0__982_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_y[6]),
    .Y(_149_)
);

FILL FILL_1__1396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1114_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1883_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_33_),
    .CLK(clk_bF$buf6),
    .Q(_y[13])
);

NAND3X1 _1463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_494_),
    .B(_496_),
    .C(_601_),
    .Y(_609_)
);

NOR2X1 _1043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_192_),
    .B(_194_),
    .Y(_195_)
);

FILL FILL_4__1603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1274_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_570_),
    .B(_663_),
    .C(_565_),
    .Y(_664_)
);

FILL FILL_3__1763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1343_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_774_),
    .Y(_835_)
);

XOR2X1 _1272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_374_),
    .B(_376_),
    .Y(_420_)
);

FILL FILL_4__1832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1819_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_875_),
    .B(_851_),
    .C(_878_),
    .Y(_889_)
);

NAND3X1 _1328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[1]),
    .B(Cin[2]),
    .C(_474_),
    .Y(_475_)
);

FILL FILL_3__1572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1152_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_218_),
    .Y(_232_)
);

FILL FILL_4__1641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL101250x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_698_),
    .B(_701_),
    .C(_697_),
    .Y(_702_)
);

OAI21X1 _1137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_280_),
    .B(_281_),
    .C(_278_),
    .Y(_287_)
);

FILL FILL_3__1381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1017_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_61_),
    .B(_916_),
    .Y(_62_)
);

AND2X2 _1366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_466_),
    .B(_469_),
    .Y(_513_)
);

FILL FILL_3__1190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1246_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_726_),
    .B(_728_),
    .C(_725_),
    .Y(_739_)
);

NAND2X1 _1175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[0]),
    .B(Cin[1]),
    .Y(_324_)
);

FILL FILL_1__957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1635_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__931_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_827_),
    .B(_794_),
    .Y(_832_)
);

AOI21X1 _1269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_407_),
    .B(_401_),
    .C(_390_),
    .Y(_417_)
);

FILL FILL_3__1093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1062_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1901_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_51_),
    .CLK(clk_bF$buf2),
    .Q(Yin0[3])
);

FILL FILL_3__953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1149_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_614_),
    .B(_616_),
    .C(_642_),
    .Y(_643_)
);

INVX1 _1078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_228_),
    .Y(_229_)
);

FILL FILL_2__1712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1291_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_756_),
    .B(_817_),
    .C(_825_),
    .Y(_852_)
);

FILL FILL_1__1452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1385_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[3]),
    .B(_77_),
    .C(_104_),
    .Y(_78_)
);

FILL FILL_1__1546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100050x70350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1194_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_754_),
    .B(_756_),
    .Y(_757_)
);

FILL FILL_0__941_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf4),
    .B(y[3]),
    .C(_110_),
    .D(y[7]),
    .Y(_123_)
);

FILL FILL_1__1775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1913_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf3),
    .B(Xin[0]),
    .Y(_100_)
);

NAND3X1 _1422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_565_),
    .B(_564_),
    .C(_567_),
    .Y(_568_)
);

INVX1 _1002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_y[13]),
    .Y(_159_)
);

FILL FILL_4__928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1302_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_792_),
    .B(_761_),
    .C(_793_),
    .Y(_794_)
);

AOI21X1 _1231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_340_),
    .B(_342_),
    .C(_378_),
    .Y(_379_)
);

NAND2X1 _982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf4),
    .B(_y[5]),
    .Y(_147_)
);

FILL FILL_1__1393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1288_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_846_),
    .B(_848_),
    .Y(_849_)
);

FILL FILL_3__1531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1029_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1880_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_30_),
    .CLK(clk_bF$buf5),
    .Q(_y[10])
);

AOI21X1 _1460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_492_),
    .B(_496_),
    .C(_485_),
    .Y(_606_)
);

AOI21X1 _1040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[2]),
    .B(Cin_0_bF$buf1),
    .C(Yin0[2]),
    .Y(_192_)
);

FILL FILL_4__1600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1097_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_658_),
    .B(_660_),
    .C(_659_),
    .Y(_661_)
);

FILL FILL_3__988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100950x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1816_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148__bF$buf0),
    .B(_886_),
    .C(_844_),
    .Y(_32_)
);

AOI21X1 _1325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_409_),
    .B(_411_),
    .C(_471_),
    .Y(_472_)
);

FILL FILL_1__1487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1205_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_683_),
    .B(_684_),
    .C(_670_),
    .Y(_699_)
);

AOI21X1 _1134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_283_),
    .B(_279_),
    .C(_251_),
    .Y(_284_)
);

FILL FILL_1__1296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1014_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_58_),
    .B(_57_),
    .Y(_59_)
);

AOI21X1 _1363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_500_),
    .B(_497_),
    .C(_484_),
    .Y(_510_)
);

FILL FILL_0__1823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1174_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf2),
    .B(_82_),
    .C(_98_),
    .Y(_50_)
);

NAND3X1 _1419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_556_),
    .B(_551_),
    .C(_554_),
    .Y(_565_)
);

FILL FILL_3__1663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1243_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_671_),
    .B(_735_),
    .C(_677_),
    .Y(_736_)
);

NAND2X1 _1172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_320_),
    .B(_316_),
    .Y(_321_)
);

FILL FILL_1__954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1719_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_790_),
    .Y(_791_)
);

OAI21X1 _1228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_307_),
    .B(_375_),
    .C(_320_),
    .Y(_376_)
);

FILL FILL_0__976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1052_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf4),
    .B(_y[4]),
    .Y(_145_)
);

FILL FILL_0__1441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1108_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1877_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_27_),
    .CLK(clk_bF$buf1),
    .Q(_y[7])
);

INVX1 _1457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_597_),
    .Y(_603_)
);

INVX1 _1037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_188_),
    .Y(_189_)
);

FILL FILL_3__1281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1268_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1337_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_791_),
    .B(_828_),
    .C(_826_),
    .Y(_829_)
);

AOI21X1 _1266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_328_),
    .B(_331_),
    .C(_322_),
    .Y(_414_)
);

FILL FILL_3__1090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1146_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_572_),
    .B(_574_),
    .Y(_640_)
);

INVX1 _1075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_223_),
    .Y(_226_)
);

FILL FILL_4__1635_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100050x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1314_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_651_),
    .B(_732_),
    .Y(_733_)
);

NAND2X1 _1169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_312_),
    .B(_314_),
    .Y(_318_)
);

FILL FILL_2__1803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1382_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148__bF$buf1),
    .B(_163_),
    .C(_75_),
    .D(_73_),
    .Y(_35_)
);

FILL FILL100650x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1049_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_446_),
    .B(_543_),
    .C(_525_),
    .Y(_544_)
);

FILL FILL_2__1612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100350x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1191_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_753_),
    .B(_752_),
    .C(_750_),
    .Y(_754_)
);

INVX1 _941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[11]),
    .Y(_120_)
);

FILL FILL_1__1772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1285_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_716_),
    .B(_845_),
    .C(_542_),
    .Y(_846_)
);

FILL FILL_1__1446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1094_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_650_),
    .B(_653_),
    .C(_652_),
    .Y(_658_)
);

FILL FILL_3__985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1813_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882_),
    .B(_883_),
    .Y(_884_)
);

NAND3X1 _1322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_373_),
    .B(_467_),
    .C(_468_),
    .Y(_469_)
);

FILL FILL_1__1484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100050x23550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1202_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_604_),
    .B(_598_),
    .C(_607_),
    .Y(_696_)
);

AOI21X1 _1131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_258_),
    .B(_261_),
    .C(_253_),
    .Y(_281_)
);

FILL FILL_1__1293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1188_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[3]),
    .B(Cin[4]),
    .Y(_751_)
);

FILL FILL_0__935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1011_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[2]),
    .B(y[14]),
    .C(_117_),
    .Y(_118_)
);

FILL FILL_1__1769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1349_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin3[1]),
    .B(_896_),
    .Y(_56_)
);

AOI21X1 _1360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_397_),
    .B(_400_),
    .C(_391_),
    .Y(_507_)
);

FILL FILL_0__1820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1171_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf3),
    .B(Yin0[1]),
    .Y(_97_)
);

OAI21X1 _1416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_473_),
    .B(_561_),
    .C(_481_),
    .Y(_562_)
);

FILL FILL_3__1660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1716_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_763_),
    .B(_767_),
    .C(_769_),
    .Y(_788_)
);

INVX1 _1225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_372_),
    .Y(_373_)
);

FILL FILL_0__973_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf3),
    .B(_y[3]),
    .Y(_143_)
);

FILL FILL_1__1387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1105_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1874_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_24_),
    .CLK(clk_bF$buf1),
    .Q(_y[4])
);

INVX1 _1454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_590_),
    .Y(_600_)
);

INVX1 _1034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_181_),
    .Y(_186_)
);

FILL FILL_1__1196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100950x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1334_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_821_),
    .B(_825_),
    .C(_794_),
    .Y(_826_)
);

OAI21X1 _1263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_402_),
    .B(_406_),
    .C(_392_),
    .Y(_411_)
);

FILL FILL_4__1823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1074_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_850_),
    .B(_876_),
    .C(_880_),
    .Y(_881_)
);

NAND3X1 _1319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_372_),
    .B(_465_),
    .C(_461_),
    .Y(_466_)
);

FILL FILL_3__1563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1143_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_542_),
    .B(_633_),
    .C(_636_),
    .Y(_637_)
);

AOI21X1 _1072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[3]),
    .B(Cin_0_bF$buf2),
    .C(Yin0[3]),
    .Y(_223_)
);

FILL FILL_4__1632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1619_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_670_),
    .B(_685_),
    .Y(_693_)
);

AND2X2 _1128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_277_),
    .B(_273_),
    .Y(_278_)
);

FILL FILL_3__1792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100350x39150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1008_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_890_),
    .B(_895_),
    .Y(_917_)
);

OAI21X1 _1357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_498_),
    .B(_499_),
    .C(_486_),
    .Y(_504_)
);

FILL FILL_3__1181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1657_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1237_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_725_),
    .Y(_730_)
);

OAI21X1 _1166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_271_),
    .B(_275_),
    .C(_314_),
    .Y(_315_)
);

FILL FILL_1__948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1046_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert6 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert7 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert8 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert9 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf2)
);

AND2X2 _1395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_533_),
    .B(_435_),
    .Y(_541_)
);

FILL FILL100650x78150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1214_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_542_),
    .B(_634_),
    .Y(_635_)
);

NAND2X1 _1069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[2]),
    .B(Cin[1]),
    .Y(_220_)
);

FILL FILL_2__1703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100950x31350 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf0),
    .B(_786_),
    .C(_843_),
    .Y(_31_)
);

FILL FILL_1__1443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1369_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_431_),
    .B(_433_),
    .C(_444_),
    .Y(_445_)
);

FILL FILL_2__1512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1919_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_579_),
    .B(_581_),
    .Y(_655_)
);

FILL FILL_3__982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100350x27450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1185_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin2[1]),
    .Y(_748_)
);

FILL FILL_0__932_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_105_),
    .B(_114_),
    .C(_115_),
    .Y(_921_[1])
);

FILL FILL_1__1766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1415_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_84_),
    .B(_91_),
    .C(_95_),
    .Y(_47_)
);

OAI21X1 _1413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237_),
    .B(_304_),
    .C(_552_),
    .Y(_559_)
);

FILL FILL_1__1575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL100650x66450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL101250x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1713_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_785_),
    .B(_784_),
    .C(_714_),
    .Y(_30_)
);

AOI22X1 _1222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[0]),
    .B(Cin[6]),
    .C(XinHL[1]),
    .D(Cin[5]),
    .Y(_370_)
);

FILL FILL_0__970_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf3),
    .B(_y[2]),
    .Y(_141_)
);

FILL FILL_1__1384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1102_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1871_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_21_),
    .CLK(clk_bF$buf4),
    .Q(_y[1])
);

OAI21X1 _1451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_590_),
    .B(_592_),
    .C(_596_),
    .Y(_597_)
);

NAND2X1 _1031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_y[1]),
    .B(_148__bF$buf1),
    .Y(_184_)
);

FILL FILL_1__1193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1088_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_553_),
    .B(_651_),
    .Y(_652_)
);

FILL FILL_3__979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1249_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_795_),
    .B(_806_),
    .C(_810_),
    .Y(_823_)
);

NAND3X1 _1260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_390_),
    .B(_401_),
    .C(_407_),
    .Y(_408_)
);

FILL FILL_4__1820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1807_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_873_),
    .Y(_878_)
);

NAND3X1 _1316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_454_),
    .B(_450_),
    .C(_452_),
    .Y(_463_)
);

FILL FILL_3__1560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1616_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_689_),
    .B(_686_),
    .C(_668_),
    .Y(_690_)
);

INVX2 _1125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[3]),
    .Y(_275_)
);

FILL FILL_1__1287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1005_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_889_),
    .B(_904_),
    .C(_913_),
    .Y(_914_)
);

NAND3X1 _1354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_484_),
    .B(_497_),
    .C(_500_),
    .Y(_501_)
);

FILL FILL100350x15750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1234_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[1]),
    .B(Cin[5]),
    .Y(_727_)
);

AND2X2 _1163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[2]),
    .B(Cin[3]),
    .Y(_312_)
);

FILL FILL_1__945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1394_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_777_),
    .B(_782_),
    .Y(_783_)
);

NAND2X1 _1219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_305_),
    .B(_308_),
    .Y(_367_)
);

FILL FILL_0__967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1043_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148__bF$buf4),
    .B(_151_),
    .C(_538_),
    .D(_535_),
    .Y(_27_)
);

FILL FILL_0__1432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1519_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1868_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_18_),
    .CLK(clk_bF$buf4),
    .Q(y[14])
);

NAND3X1 _1448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_494_),
    .B(_496_),
    .C(_593_),
    .Y(_594_)
);

OR2X2 _1028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_180_),
    .B(_165_),
    .Y(_181_)
);

FILL FILL_3__1692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1761_ (
    .gnd(gnd),
    .vdd(vdd)
);

endmodule

magic
tech scmos
magscale 1 2
timestamp 1711577914
<< metal1 >>
rect -63 6258 -3 6518
rect 6750 6502 6843 6518
rect 5907 6457 5933 6463
rect 4767 6437 4873 6443
rect 5407 6437 5493 6443
rect 5547 6437 5633 6443
rect 6187 6437 6293 6443
rect 1487 6417 1533 6423
rect 2627 6417 2653 6423
rect 3267 6417 3293 6423
rect 3587 6417 3633 6423
rect 1767 6357 1893 6363
rect 1987 6357 2113 6363
rect 2167 6357 2253 6363
rect 3187 6357 3313 6363
rect 3847 6357 3953 6363
rect 5027 6357 5073 6363
rect 5647 6357 5693 6363
rect 5747 6357 5773 6363
rect 5847 6357 5913 6363
rect 6247 6357 6353 6363
rect 2627 6337 2673 6343
rect -63 6242 30 6258
rect -63 5738 -3 6242
rect 1627 6173 1633 6187
rect 3767 6177 3793 6183
rect 1587 6157 1653 6163
rect 3173 6143 3187 6153
rect 3087 6140 3187 6143
rect 3087 6137 3183 6140
rect 4807 6137 4893 6143
rect 5767 6137 5833 6143
rect 6047 6137 6153 6143
rect 6247 6137 6373 6143
rect 6567 6137 6613 6143
rect 6657 6137 6713 6143
rect 3760 6123 3773 6127
rect 3757 6113 3773 6123
rect 6657 6123 6663 6137
rect 6607 6117 6663 6123
rect 3757 6083 3763 6113
rect 3707 6077 3763 6083
rect 827 6057 933 6063
rect 6783 5998 6843 6502
rect 6750 5982 6843 5998
rect 1447 5937 1473 5943
rect 3207 5937 3253 5943
rect 3933 5943 3947 5953
rect 3887 5940 3947 5943
rect 3887 5937 3943 5940
rect 1567 5917 1713 5923
rect 3167 5917 3313 5923
rect 6407 5917 6493 5923
rect 1427 5897 1473 5903
rect 1607 5837 1773 5843
rect 1947 5837 2013 5843
rect 2967 5837 3013 5843
rect 3407 5837 3473 5843
rect 3607 5837 3633 5843
rect 4027 5837 4153 5843
rect 5347 5837 5393 5843
rect 6047 5797 6093 5803
rect -63 5722 30 5738
rect -63 5218 -3 5722
rect 4647 5617 4693 5623
rect 5807 5617 5973 5623
rect 6287 5617 6353 5623
rect 6547 5617 6573 5623
rect 5900 5603 5913 5607
rect 5897 5593 5913 5603
rect 6027 5603 6040 5607
rect 6027 5593 6043 5603
rect 6187 5597 6233 5603
rect 6607 5603 6620 5607
rect 6607 5593 6623 5603
rect 3927 5557 3953 5563
rect 5897 5563 5903 5593
rect 6037 5567 6043 5593
rect 6407 5577 6483 5583
rect 5867 5557 5903 5563
rect 6027 5557 6043 5567
rect 6477 5567 6483 5577
rect 6477 5557 6493 5567
rect 6027 5553 6040 5557
rect 6480 5553 6493 5557
rect 5167 5537 5273 5543
rect 6617 5543 6623 5593
rect 6547 5537 6623 5543
rect 5127 5517 5213 5523
rect 6783 5478 6843 5982
rect 6750 5462 6843 5478
rect 2167 5437 2213 5443
rect 2307 5397 2353 5403
rect 6487 5397 6553 5403
rect 2400 5383 2413 5387
rect 2397 5373 2413 5383
rect 3520 5383 3533 5387
rect 3517 5373 3533 5383
rect 5820 5383 5833 5387
rect 5817 5373 5833 5383
rect 6277 5377 6313 5383
rect 2397 5343 2403 5373
rect 2347 5337 2403 5343
rect 3517 5347 3523 5373
rect 5817 5347 5823 5373
rect 6277 5347 6283 5377
rect 6373 5383 6387 5393
rect 6600 5383 6613 5387
rect 6373 5380 6403 5383
rect 6377 5377 6403 5380
rect 6397 5347 6403 5377
rect 3517 5337 3533 5347
rect 3520 5333 3533 5337
rect 3647 5337 3673 5343
rect 5817 5337 5833 5347
rect 5820 5333 5833 5337
rect 6267 5337 6283 5347
rect 6267 5333 6280 5337
rect 6387 5337 6403 5347
rect 6597 5373 6613 5383
rect 6387 5333 6400 5337
rect 507 5317 633 5323
rect 2207 5317 2233 5323
rect 4687 5317 4753 5323
rect 4827 5317 4893 5323
rect 6597 5323 6603 5373
rect 6547 5317 6603 5323
rect 6727 5277 6753 5283
rect -63 5202 30 5218
rect -63 4698 -3 5202
rect 3407 5137 3493 5143
rect 67 5097 113 5103
rect 2267 5097 2293 5103
rect 4687 5097 4793 5103
rect 4907 5097 4933 5103
rect 5067 5097 5133 5103
rect 5647 5097 5713 5103
rect 5947 5097 6013 5103
rect 6147 5097 6193 5103
rect 1993 5083 2007 5093
rect 4600 5083 4613 5087
rect 1993 5080 2023 5083
rect 1997 5077 2023 5080
rect 2017 5043 2023 5077
rect 4597 5073 4613 5083
rect 6187 5083 6200 5087
rect 6187 5073 6203 5083
rect 2017 5037 2053 5043
rect 4597 5043 4603 5073
rect 6197 5047 6203 5073
rect 4547 5037 4603 5043
rect 5347 5037 5373 5043
rect 6187 5037 6203 5047
rect 6187 5033 6200 5037
rect 2287 5017 2353 5023
rect 3927 5017 3953 5023
rect 187 4997 273 5003
rect 2727 4997 2753 5003
rect 6783 4958 6843 5462
rect 6750 4942 6843 4958
rect 2527 4897 2573 4903
rect 5227 4897 5253 4903
rect 167 4877 233 4883
rect 707 4877 733 4883
rect 2547 4877 2593 4883
rect 4707 4877 4773 4883
rect 5027 4877 5053 4883
rect 6187 4877 6213 4883
rect 747 4797 793 4803
rect 1737 4766 1743 4873
rect 6347 4877 6413 4883
rect 2380 4863 2393 4867
rect 2377 4853 2393 4863
rect 3627 4863 3640 4867
rect 5540 4863 5553 4867
rect 3627 4853 3643 4863
rect 2377 4827 2383 4853
rect 2377 4817 2393 4827
rect 2380 4813 2393 4817
rect 3637 4823 3643 4853
rect 5537 4853 5553 4863
rect 5847 4863 5860 4867
rect 5847 4853 5863 4863
rect 6527 4863 6540 4867
rect 6560 4863 6573 4867
rect 6527 4853 6543 4863
rect 3637 4817 3673 4823
rect 5537 4823 5543 4853
rect 5507 4817 5543 4823
rect 5667 4817 5713 4823
rect 5857 4823 5863 4853
rect 6537 4827 6543 4853
rect 5857 4817 5893 4823
rect 6527 4817 6543 4827
rect 6557 4853 6573 4863
rect 6667 4863 6680 4867
rect 6667 4853 6683 4863
rect 6557 4827 6563 4853
rect 6557 4817 6573 4827
rect 6527 4813 6540 4817
rect 6560 4813 6573 4817
rect 6677 4823 6683 4853
rect 6657 4817 6683 4823
rect 6657 4807 6663 4817
rect 3787 4797 3873 4803
rect 4287 4797 4353 4803
rect 4747 4797 4853 4803
rect 6640 4805 6663 4807
rect 6647 4797 6663 4805
rect 6647 4793 6660 4797
rect 4267 4777 4313 4783
rect 4407 4777 4453 4783
rect -63 4682 30 4698
rect -63 4178 -3 4682
rect 6227 4657 6253 4663
rect 4647 4637 4693 4643
rect 6387 4597 6433 4603
rect 3447 4577 3473 4583
rect 3627 4577 3713 4583
rect 4407 4577 4433 4583
rect 5147 4577 5213 4583
rect 5307 4577 5413 4583
rect 5520 4583 5533 4587
rect 5517 4573 5533 4583
rect 6047 4577 6073 4583
rect 6227 4577 6313 4583
rect 2367 4563 2380 4567
rect 2367 4553 2383 4563
rect 4827 4563 4840 4567
rect 5517 4563 5523 4573
rect 5780 4563 5793 4567
rect 4827 4553 4843 4563
rect 2377 4543 2383 4553
rect 2377 4537 2403 4543
rect 2397 4527 2403 4537
rect 4837 4527 4843 4553
rect 5497 4557 5523 4563
rect 5497 4527 5503 4557
rect 5777 4553 5793 4563
rect 2397 4517 2413 4527
rect 2400 4513 2413 4517
rect 4427 4517 4453 4523
rect 4827 4517 4843 4527
rect 4827 4513 4840 4517
rect 5127 4517 5153 4523
rect 5497 4517 5513 4527
rect 5500 4513 5513 4517
rect 5777 4523 5783 4553
rect 5747 4517 5783 4523
rect 6187 4517 6213 4523
rect 2507 4497 2573 4503
rect 5467 4497 5493 4503
rect 6237 4503 6243 4533
rect 6393 4523 6407 4533
rect 6367 4520 6407 4523
rect 6367 4517 6403 4520
rect 6507 4517 6533 4523
rect 6237 4497 6313 4503
rect 6487 4497 6593 4503
rect 6667 4497 6693 4503
rect 6507 4477 6533 4483
rect 6783 4438 6843 4942
rect 6750 4422 6843 4438
rect 5947 4397 5973 4403
rect 6467 4397 6503 4403
rect 5117 4377 5153 4383
rect 2207 4357 2293 4363
rect 3707 4357 3753 4363
rect 867 4343 880 4347
rect 5117 4343 5123 4377
rect 5147 4357 5173 4363
rect 6177 4357 6233 4363
rect 867 4333 883 4343
rect 5117 4337 5153 4343
rect 5797 4337 5833 4343
rect 877 4323 883 4333
rect 877 4317 903 4323
rect 897 4307 903 4317
rect 5797 4307 5803 4337
rect 5947 4343 5960 4347
rect 6177 4343 6183 4357
rect 5947 4333 5963 4343
rect 897 4297 913 4307
rect 900 4293 913 4297
rect 5327 4303 5340 4307
rect 5327 4293 5343 4303
rect 5787 4297 5803 4307
rect 5813 4307 5827 4313
rect 5957 4307 5963 4333
rect 5813 4300 5833 4307
rect 5817 4297 5833 4300
rect 5787 4293 5800 4297
rect 5820 4293 5833 4297
rect 5947 4297 5963 4307
rect 6157 4337 6183 4343
rect 6157 4307 6163 4337
rect 6307 4337 6353 4343
rect 6157 4297 6173 4307
rect 5947 4293 5960 4297
rect 6160 4293 6173 4297
rect 6497 4303 6503 4397
rect 6660 4343 6673 4347
rect 6657 4333 6673 4343
rect 6497 4297 6523 4303
rect 847 4277 893 4283
rect 3167 4277 3273 4283
rect 4307 4277 4393 4283
rect 4927 4277 4993 4283
rect 5337 4283 5343 4293
rect 6517 4287 6523 4297
rect 6657 4287 6663 4333
rect 5227 4277 5393 4283
rect 6067 4277 6113 4283
rect 6127 4277 6233 4283
rect 6277 4277 6373 4283
rect 5307 4257 5393 4263
rect 6277 4243 6283 4277
rect 6517 4285 6540 4287
rect 6517 4277 6533 4285
rect 6520 4273 6533 4277
rect 6307 4257 6353 4263
rect 6277 4237 6333 4243
rect -63 4162 30 4178
rect -63 3658 -3 4162
rect 3847 4097 3913 4103
rect 3687 4077 3793 4083
rect 3687 4057 3713 4063
rect 4220 4063 4233 4067
rect 4217 4053 4233 4063
rect 4987 4057 5033 4063
rect 5227 4057 5253 4063
rect 5847 4057 5903 4063
rect 3900 4043 3913 4047
rect 3897 4033 3913 4043
rect 4007 4043 4020 4047
rect 4217 4043 4223 4053
rect 4500 4043 4513 4047
rect 4007 4033 4023 4043
rect 3897 3986 3903 4033
rect 4017 4007 4023 4033
rect 4007 3997 4023 4007
rect 4197 4037 4223 4043
rect 4197 4007 4203 4037
rect 4497 4033 4513 4043
rect 4197 3997 4213 4007
rect 4007 3993 4020 3997
rect 4200 3993 4213 3997
rect 4187 3977 4233 3983
rect 4497 3983 4503 4033
rect 5897 4007 5903 4057
rect 6247 4057 6313 4063
rect 6547 4043 6560 4047
rect 6547 4033 6563 4043
rect 5897 3997 5913 4007
rect 5900 3993 5913 3997
rect 6387 3997 6433 4003
rect 6557 4003 6563 4033
rect 6557 3997 6593 4003
rect 4497 3977 4533 3983
rect 4767 3977 4813 3983
rect 3547 3957 3573 3963
rect 6783 3918 6843 4422
rect 6750 3902 6843 3918
rect 2267 3857 2313 3863
rect 3880 3823 3893 3827
rect 3877 3813 3893 3823
rect 4547 3823 4560 3827
rect 4740 3823 4753 3827
rect 4547 3813 4563 3823
rect 3877 3783 3883 3813
rect 3827 3777 3883 3783
rect 4557 3783 4563 3813
rect 4737 3813 4753 3823
rect 4993 3823 5007 3832
rect 4993 3820 5043 3823
rect 4997 3817 5043 3820
rect 4737 3787 4743 3813
rect 5037 3787 5043 3817
rect 5827 3823 5840 3827
rect 6320 3823 6333 3827
rect 5827 3813 5843 3823
rect 4557 3777 4593 3783
rect 4737 3777 4753 3787
rect 4740 3773 4753 3777
rect 5037 3777 5053 3787
rect 5040 3773 5053 3777
rect 5837 3783 5843 3813
rect 6317 3813 6333 3823
rect 6607 3823 6620 3827
rect 6640 3823 6653 3827
rect 6607 3813 6623 3823
rect 6317 3803 6323 3813
rect 6277 3797 6323 3803
rect 6277 3787 6283 3797
rect 5837 3777 5893 3783
rect 6267 3777 6283 3787
rect 6267 3773 6280 3777
rect 6307 3777 6333 3783
rect 6617 3767 6623 3813
rect 6637 3813 6653 3823
rect 1227 3757 1253 3763
rect 3527 3757 3633 3763
rect 3687 3757 3753 3763
rect 4547 3757 4653 3763
rect 4707 3757 4773 3763
rect 6147 3757 6213 3763
rect 6637 3763 6643 3813
rect 6637 3757 6673 3763
rect 3567 3737 3633 3743
rect -63 3642 30 3658
rect -63 3138 -3 3642
rect 3307 3577 3333 3583
rect 567 3537 593 3543
rect 1607 3537 1633 3543
rect 4627 3537 4693 3543
rect 4767 3537 4813 3543
rect 5227 3537 5293 3543
rect 1060 3523 1073 3527
rect 1057 3513 1073 3523
rect 2780 3523 2793 3527
rect 2777 3513 2793 3523
rect 4620 3523 4633 3527
rect 4617 3513 4633 3523
rect 5527 3523 5540 3527
rect 5880 3523 5893 3527
rect 5527 3513 5543 3523
rect 433 3487 447 3493
rect 1057 3487 1063 3513
rect 427 3480 447 3487
rect 427 3477 443 3480
rect 427 3473 440 3477
rect 1047 3477 1063 3487
rect 2777 3487 2783 3513
rect 4617 3487 4623 3513
rect 5537 3487 5543 3513
rect 2777 3477 2793 3487
rect 1047 3473 1060 3477
rect 2780 3473 2793 3477
rect 4617 3477 4633 3487
rect 4620 3473 4633 3477
rect 5067 3477 5093 3483
rect 5527 3477 5543 3487
rect 5877 3513 5893 3523
rect 5527 3473 5540 3477
rect 1067 3457 1093 3463
rect 3327 3457 3373 3463
rect 4187 3457 4313 3463
rect 5877 3463 5883 3513
rect 6037 3483 6043 3533
rect 6220 3523 6233 3527
rect 6217 3513 6233 3523
rect 6007 3477 6043 3483
rect 6217 3483 6223 3513
rect 6167 3477 6223 3483
rect 6327 3477 6353 3483
rect 5847 3457 5883 3463
rect 5867 3437 5893 3443
rect 6783 3398 6843 3902
rect 6750 3382 6843 3398
rect 6667 3357 6733 3363
rect 5833 3323 5847 3333
rect 5833 3320 5863 3323
rect 5837 3317 5863 3320
rect 1067 3303 1080 3307
rect 4180 3303 4193 3307
rect 1067 3300 1083 3303
rect 1067 3293 1087 3300
rect 1073 3286 1087 3293
rect 4177 3293 4193 3303
rect 4177 3267 4183 3293
rect 4177 3257 4193 3267
rect 4180 3253 4193 3257
rect 4607 3237 4633 3243
rect 5327 3237 5453 3243
rect 5857 3246 5863 3317
rect 6040 3303 6053 3307
rect 6037 3293 6053 3303
rect 6167 3303 6180 3307
rect 6360 3303 6373 3307
rect 6167 3293 6183 3303
rect 6037 3267 6043 3293
rect 6020 3266 6043 3267
rect 6027 3257 6043 3266
rect 6027 3253 6040 3257
rect 6177 3246 6183 3293
rect 6357 3293 6373 3303
rect 6540 3303 6553 3307
rect 6537 3293 6553 3303
rect 6357 3263 6363 3293
rect 6327 3257 6363 3263
rect 6537 3267 6543 3293
rect 6537 3257 6553 3267
rect 6540 3253 6553 3257
rect 5687 3237 5733 3243
rect 6507 3237 6573 3243
rect 4907 3197 4993 3203
rect -63 3122 30 3138
rect -63 2618 -3 3122
rect 1087 3100 1143 3103
rect 1087 3097 1147 3100
rect 1133 3087 1147 3097
rect 4567 3037 4713 3043
rect 6227 3037 6273 3043
rect 2827 3017 2953 3023
rect 3227 3017 3273 3023
rect 3327 3017 3413 3023
rect 3987 3017 4013 3023
rect 4027 3017 4053 3023
rect 4107 3017 4253 3023
rect 4657 3017 4693 3023
rect 4307 3003 4320 3007
rect 4657 3003 4663 3017
rect 4927 3017 4993 3023
rect 6247 3017 6313 3023
rect 4307 2993 4323 3003
rect 787 2957 813 2963
rect 4127 2957 4173 2963
rect 4317 2963 4323 2993
rect 4637 2997 4663 3003
rect 4917 3003 4923 3013
rect 6397 3017 6473 3023
rect 4917 2997 4943 3003
rect 4317 2957 4353 2963
rect 4637 2947 4643 2997
rect 4937 2967 4943 2997
rect 6187 3003 6200 3007
rect 6187 2993 6203 3003
rect 4927 2957 4943 2967
rect 6197 2963 6203 2993
rect 6397 2967 6403 3017
rect 6197 2957 6253 2963
rect 4927 2953 4940 2957
rect 6397 2957 6413 2967
rect 6400 2953 6413 2957
rect 3007 2937 3113 2943
rect 4487 2937 4513 2943
rect 4620 2946 4643 2947
rect 4627 2937 4643 2946
rect 4627 2933 4640 2937
rect 5867 2937 5933 2943
rect 6783 2878 6843 3382
rect 6750 2862 6843 2878
rect 2967 2797 3013 2803
rect 4067 2797 4113 2803
rect 6627 2797 6693 2803
rect 3687 2783 3700 2787
rect 3687 2773 3703 2783
rect 4347 2777 4373 2783
rect 6087 2783 6100 2787
rect 6120 2783 6133 2787
rect 6087 2773 6103 2783
rect 3697 2747 3703 2773
rect 3687 2737 3703 2747
rect 3717 2747 3723 2773
rect 6097 2747 6103 2773
rect 3717 2737 3733 2747
rect 3687 2733 3700 2737
rect 3720 2733 3733 2737
rect 6087 2737 6103 2747
rect 6117 2773 6133 2783
rect 6280 2783 6293 2787
rect 6277 2773 6293 2783
rect 6417 2777 6453 2783
rect 6117 2747 6123 2773
rect 6277 2747 6283 2773
rect 6117 2737 6133 2747
rect 6087 2733 6100 2737
rect 6120 2733 6133 2737
rect 6277 2737 6293 2747
rect 6280 2733 6293 2737
rect 6417 2743 6423 2777
rect 6397 2737 6423 2743
rect 6397 2727 6403 2737
rect 1047 2717 1113 2723
rect 1767 2717 1833 2723
rect 1947 2717 1973 2723
rect 1987 2723 2000 2727
rect 1987 2717 2003 2723
rect 1987 2713 2000 2717
rect 3547 2717 3593 2723
rect 4527 2717 4573 2723
rect 5687 2717 5813 2723
rect 6227 2717 6253 2723
rect 6387 2717 6403 2727
rect 6387 2713 6400 2717
rect 1887 2697 1953 2703
rect 6387 2697 6433 2703
rect -63 2602 30 2618
rect -63 2098 -3 2602
rect 5607 2517 5633 2523
rect 807 2497 933 2503
rect 2357 2497 2413 2503
rect 887 2477 913 2483
rect 2357 2447 2363 2497
rect 2927 2497 3013 2503
rect 4497 2497 4533 2503
rect 2380 2483 2393 2487
rect 2347 2437 2363 2447
rect 2377 2473 2393 2483
rect 4497 2483 4503 2497
rect 5813 2503 5827 2513
rect 5747 2500 5827 2503
rect 5747 2497 5823 2500
rect 6007 2497 6133 2503
rect 6527 2497 6573 2503
rect 5920 2483 5933 2487
rect 4477 2477 4503 2483
rect 2377 2447 2383 2473
rect 4477 2447 4483 2477
rect 5917 2473 5933 2483
rect 6080 2483 6093 2487
rect 6077 2473 6093 2483
rect 6580 2483 6593 2487
rect 6577 2473 6593 2483
rect 2377 2437 2393 2447
rect 2347 2433 2360 2437
rect 2380 2433 2393 2437
rect 4477 2437 4493 2447
rect 4480 2433 4493 2437
rect 5267 2437 5293 2443
rect 5917 2443 5923 2473
rect 5887 2437 5923 2443
rect 6077 2447 6083 2473
rect 6577 2447 6583 2473
rect 6077 2437 6093 2447
rect 6080 2433 6093 2437
rect 6577 2437 6593 2447
rect 6580 2433 6593 2437
rect 827 2417 873 2423
rect 4727 2417 4793 2423
rect 6227 2397 6253 2403
rect 6783 2358 6843 2862
rect 6750 2342 6843 2358
rect 5833 2303 5847 2313
rect 5807 2300 5847 2303
rect 5807 2297 5843 2300
rect 4247 2277 4313 2283
rect 6467 2277 6533 2283
rect 4493 2263 4507 2273
rect 4493 2260 4523 2263
rect 4497 2257 4523 2260
rect 4517 2227 4523 2257
rect 5087 2257 5143 2263
rect 4507 2217 4523 2227
rect 5137 2227 5143 2257
rect 5607 2257 5633 2263
rect 5980 2263 5993 2267
rect 5977 2253 5993 2263
rect 6087 2257 6123 2263
rect 5137 2217 5153 2227
rect 4507 2213 4520 2217
rect 5140 2213 5153 2217
rect 5977 2223 5983 2253
rect 5947 2217 5983 2223
rect 6117 2227 6123 2257
rect 6117 2217 6133 2227
rect 6120 2213 6133 2217
rect 407 2197 513 2203
rect 4247 2197 4333 2203
rect 4807 2197 4893 2203
rect 5587 2197 5673 2203
rect 6227 2197 6273 2203
rect 2687 2157 2733 2163
rect -63 2082 30 2098
rect -63 1578 -3 2082
rect 6547 2057 6573 2063
rect 1347 1997 1453 2003
rect 4867 1997 4913 2003
rect 6567 1997 6653 2003
rect 827 1977 913 1983
rect 927 1977 993 1983
rect 1367 1977 1413 1983
rect 4077 1977 4113 1983
rect 2227 1957 2253 1963
rect 3160 1963 3173 1967
rect 3157 1953 3173 1963
rect 4077 1963 4083 1977
rect 4187 1977 4213 1983
rect 4347 1977 4393 1983
rect 4687 1977 4763 1983
rect 4057 1957 4083 1963
rect 407 1917 473 1923
rect 3157 1923 3163 1953
rect 3127 1917 3163 1923
rect 3647 1897 3733 1903
rect 4057 1903 4063 1957
rect 4577 1907 4583 1973
rect 4707 1963 4720 1967
rect 4707 1953 4723 1963
rect 4717 1927 4723 1953
rect 4707 1917 4723 1927
rect 4757 1927 4763 1977
rect 4987 1977 5043 1983
rect 4887 1957 4913 1963
rect 5007 1963 5020 1967
rect 5007 1953 5023 1963
rect 5017 1927 5023 1953
rect 4757 1917 4773 1927
rect 4707 1913 4720 1917
rect 4760 1913 4773 1917
rect 5007 1917 5023 1927
rect 5007 1913 5020 1917
rect 4057 1897 4113 1903
rect 4560 1906 4583 1907
rect 4567 1897 4583 1906
rect 4567 1893 4580 1897
rect 5037 1903 5043 1977
rect 6707 1963 6720 1967
rect 6707 1953 6723 1963
rect 6717 1927 6723 1953
rect 6707 1917 6723 1927
rect 6707 1913 6720 1917
rect 4987 1897 5043 1903
rect 5607 1897 5673 1903
rect 5727 1897 5773 1903
rect 6267 1897 6373 1903
rect 6783 1838 6843 2342
rect 6750 1822 6843 1838
rect 4067 1757 4103 1763
rect 2800 1743 2813 1747
rect 2797 1733 2813 1743
rect 3627 1737 3663 1743
rect 2797 1707 2803 1733
rect 3657 1707 3663 1737
rect 4097 1743 4103 1757
rect 6507 1757 6613 1763
rect 3947 1737 3983 1743
rect 4097 1737 4123 1743
rect 2797 1697 2813 1707
rect 2800 1693 2813 1697
rect 3657 1697 3673 1707
rect 3660 1693 3673 1697
rect 847 1677 893 1683
rect 3347 1677 3393 1683
rect 3927 1677 3953 1683
rect 3977 1667 3983 1737
rect 4117 1707 4123 1737
rect 6327 1737 6393 1743
rect 6667 1737 6733 1743
rect 4107 1697 4123 1707
rect 4107 1693 4120 1697
rect 4047 1677 4073 1683
rect 4087 1677 4193 1683
rect 5667 1677 5793 1683
rect 3960 1666 3983 1667
rect 3967 1657 3983 1666
rect 3967 1653 3980 1657
rect 4733 1663 4747 1673
rect 4687 1660 4747 1663
rect 4687 1657 4743 1660
rect 3807 1597 3833 1603
rect -63 1562 30 1578
rect -63 1058 -3 1562
rect 3987 1497 4073 1503
rect 4653 1503 4667 1513
rect 4653 1500 4713 1503
rect 4657 1497 4713 1500
rect 3267 1457 3313 1463
rect 3527 1457 3613 1463
rect 3667 1457 3813 1463
rect 4647 1457 4713 1463
rect 5367 1457 5513 1463
rect 6347 1457 6412 1463
rect 3507 1437 3533 1443
rect 6437 1407 6443 1453
rect 6747 1443 6760 1447
rect 6747 1433 6763 1443
rect 6757 1407 6763 1433
rect 4507 1397 4553 1403
rect 6437 1397 6453 1407
rect 6440 1393 6453 1397
rect 6567 1397 6613 1403
rect 6747 1397 6763 1407
rect 6747 1393 6760 1397
rect 3487 1377 3533 1383
rect 5607 1377 5653 1383
rect 5427 1337 5453 1343
rect 5727 1337 5753 1343
rect 6783 1318 6843 1822
rect 6750 1302 6843 1318
rect 347 1217 373 1223
rect 1087 1217 1113 1223
rect 1387 1217 1413 1223
rect 3977 1217 4033 1223
rect 2167 1177 2193 1183
rect 3977 1183 3983 1217
rect 4147 1223 4160 1227
rect 4147 1213 4163 1223
rect 5747 1223 5760 1227
rect 5747 1213 5763 1223
rect 4157 1187 4163 1213
rect 4360 1203 4373 1207
rect 4357 1193 4373 1203
rect 4357 1187 4363 1193
rect 5757 1187 5763 1213
rect 3957 1177 3983 1183
rect 527 1157 593 1163
rect 2007 1157 2073 1163
rect 2307 1157 2353 1163
rect 2627 1157 2673 1163
rect 3487 1157 3553 1163
rect 3957 1163 3963 1177
rect 4147 1177 4163 1187
rect 4147 1173 4160 1177
rect 4347 1177 4363 1187
rect 4347 1173 4360 1177
rect 5747 1177 5763 1187
rect 5917 1217 5953 1223
rect 5917 1183 5923 1217
rect 6207 1217 6253 1223
rect 5897 1177 5923 1183
rect 5747 1173 5760 1177
rect 3907 1157 3963 1163
rect 4307 1157 4373 1163
rect 4767 1157 4873 1163
rect 5897 1163 5903 1177
rect 5867 1157 5903 1163
rect 3967 1117 4013 1123
rect -63 1042 30 1058
rect -63 538 -3 1042
rect 1687 957 1813 963
rect 1027 937 1073 943
rect 1247 937 1293 943
rect 1447 937 1473 943
rect 4147 937 4273 943
rect 4967 937 4993 943
rect 5927 937 6073 943
rect 2527 857 2573 863
rect 2627 857 2673 863
rect 2867 857 2953 863
rect 6167 857 6233 863
rect 6783 798 6843 1302
rect 6750 782 6843 798
rect 1387 717 1413 723
rect 2127 717 2253 723
rect 2467 717 2513 723
rect 3817 707 3823 733
rect 3847 717 3873 723
rect 4307 717 4373 723
rect 5127 717 5193 723
rect 2147 697 2173 703
rect 4107 697 4143 703
rect 4137 667 4143 697
rect 4137 657 4153 667
rect 4140 653 4153 657
rect 627 637 753 643
rect 1967 637 2013 643
rect 3787 637 3853 643
rect 3947 637 4053 643
rect 4267 637 4373 643
rect 4587 637 4713 643
rect 5087 637 5193 643
rect 5387 637 5513 643
rect 6067 637 6153 643
rect 6647 637 6673 643
rect 587 617 693 623
rect 5407 617 5493 623
rect 4313 603 4327 613
rect 4267 600 4327 603
rect 4267 597 4323 600
rect -63 522 30 538
rect -63 18 -3 522
rect 4347 437 4393 443
rect 327 417 413 423
rect 4287 417 4413 423
rect 4487 417 4573 423
rect 5387 417 5443 423
rect 2837 397 2873 403
rect 2837 367 2843 397
rect 4987 397 5033 403
rect 5437 367 5443 417
rect 6487 417 6523 423
rect 6517 403 6523 417
rect 6517 397 6543 403
rect 2827 357 2843 367
rect 2827 353 2840 357
rect 5427 357 5443 367
rect 6537 363 6543 397
rect 6537 357 6573 363
rect 5427 353 5440 357
rect 3627 337 3713 343
rect 4267 337 4313 343
rect 4327 337 4353 343
rect 5647 337 5713 343
rect 6783 278 6843 782
rect 6750 262 6843 278
rect 647 240 683 243
rect 647 237 687 240
rect 673 227 687 237
rect 4587 237 4633 243
rect 4453 183 4467 193
rect 4437 180 4467 183
rect 4437 177 4463 180
rect 1407 163 1420 167
rect 1407 153 1423 163
rect 1417 147 1423 153
rect 1417 137 1433 147
rect 1420 133 1433 137
rect 1727 137 1753 143
rect 3287 137 3313 143
rect 4437 143 4443 177
rect 4407 137 4443 143
rect 6307 137 6333 143
rect 407 117 553 123
rect 1407 117 1493 123
rect 4267 117 4293 123
rect 4447 117 4513 123
rect 6007 117 6053 123
rect 627 97 713 103
rect -63 2 30 18
rect 6783 2 6843 262
<< m2contact >>
rect 5893 6453 5907 6467
rect 5933 6453 5947 6467
rect 4753 6433 4767 6447
rect 4873 6433 4887 6447
rect 5393 6433 5407 6447
rect 5493 6434 5507 6448
rect 5533 6434 5547 6448
rect 5633 6433 5647 6447
rect 6173 6433 6187 6447
rect 6293 6433 6307 6447
rect 1473 6413 1487 6427
rect 1533 6413 1547 6427
rect 2613 6413 2627 6427
rect 2653 6413 2667 6427
rect 3253 6413 3267 6427
rect 3293 6413 3307 6427
rect 3573 6413 3587 6427
rect 3633 6413 3647 6427
rect 1753 6353 1767 6367
rect 1893 6353 1907 6367
rect 1973 6353 1987 6367
rect 2113 6351 2127 6365
rect 2153 6351 2167 6365
rect 2253 6351 2267 6365
rect 3173 6353 3187 6367
rect 3313 6353 3327 6367
rect 3833 6353 3847 6367
rect 3953 6353 3967 6367
rect 5013 6353 5027 6367
rect 5073 6353 5087 6367
rect 5633 6353 5647 6367
rect 5693 6351 5707 6365
rect 5733 6353 5747 6367
rect 5773 6353 5787 6367
rect 5833 6353 5847 6367
rect 5913 6352 5927 6366
rect 6233 6353 6247 6367
rect 6353 6353 6367 6367
rect 2613 6333 2627 6347
rect 2673 6333 2687 6347
rect 1613 6173 1627 6187
rect 1633 6173 1647 6187
rect 3753 6173 3767 6187
rect 3793 6173 3807 6187
rect 1573 6153 1587 6167
rect 1653 6152 1667 6166
rect 3173 6153 3187 6167
rect 3073 6133 3087 6147
rect 4793 6133 4807 6147
rect 4893 6133 4907 6147
rect 5753 6133 5767 6147
rect 5833 6133 5847 6147
rect 6033 6133 6047 6147
rect 6153 6134 6167 6148
rect 6233 6133 6247 6147
rect 6373 6133 6387 6147
rect 6553 6133 6567 6147
rect 6613 6133 6627 6147
rect 3773 6113 3787 6127
rect 6593 6113 6607 6127
rect 6713 6133 6727 6147
rect 3693 6073 3707 6087
rect 813 6053 827 6067
rect 933 6053 947 6067
rect 3933 5953 3947 5967
rect 1433 5933 1447 5947
rect 1473 5933 1487 5947
rect 3193 5933 3207 5947
rect 3253 5933 3267 5947
rect 3873 5933 3887 5947
rect 1553 5913 1567 5927
rect 1713 5913 1727 5927
rect 3153 5913 3167 5927
rect 3313 5913 3327 5927
rect 6393 5913 6407 5927
rect 6493 5913 6507 5927
rect 1413 5893 1427 5907
rect 1473 5892 1487 5906
rect 1593 5833 1607 5847
rect 1773 5833 1787 5847
rect 1933 5833 1947 5847
rect 2013 5833 2027 5847
rect 2953 5833 2967 5847
rect 3013 5833 3027 5847
rect 3393 5833 3407 5847
rect 3473 5833 3487 5847
rect 3593 5833 3607 5847
rect 3633 5833 3647 5847
rect 4013 5833 4027 5847
rect 4153 5833 4167 5847
rect 5333 5833 5347 5847
rect 5393 5833 5407 5847
rect 6033 5793 6047 5807
rect 6093 5793 6107 5807
rect 4633 5614 4647 5628
rect 4693 5613 4707 5627
rect 5793 5613 5807 5627
rect 5973 5613 5987 5627
rect 6273 5613 6287 5627
rect 6353 5613 6367 5627
rect 6533 5614 6547 5628
rect 6573 5613 6587 5627
rect 5913 5593 5927 5607
rect 6013 5593 6027 5607
rect 6173 5593 6187 5607
rect 6233 5593 6247 5607
rect 6593 5593 6607 5607
rect 3913 5553 3927 5567
rect 3953 5553 3967 5567
rect 5853 5553 5867 5567
rect 6393 5573 6407 5587
rect 6013 5553 6027 5567
rect 6493 5553 6507 5567
rect 5153 5533 5167 5547
rect 5273 5533 5287 5547
rect 6533 5533 6547 5547
rect 5113 5513 5127 5527
rect 5213 5513 5227 5527
rect 2153 5433 2167 5447
rect 2213 5433 2227 5447
rect 2293 5393 2307 5407
rect 2353 5393 2367 5407
rect 6373 5393 6387 5407
rect 6473 5393 6487 5407
rect 6553 5393 6567 5407
rect 2413 5373 2427 5387
rect 3533 5373 3547 5387
rect 5833 5373 5847 5387
rect 2333 5333 2347 5347
rect 6313 5373 6327 5387
rect 3533 5333 3547 5347
rect 3633 5333 3647 5347
rect 3673 5333 3687 5347
rect 5833 5333 5847 5347
rect 6253 5333 6267 5347
rect 6373 5333 6387 5347
rect 6613 5373 6627 5387
rect 493 5313 507 5327
rect 633 5313 647 5327
rect 2193 5312 2207 5326
rect 2233 5313 2247 5327
rect 4673 5313 4687 5327
rect 4753 5313 4767 5327
rect 4813 5313 4827 5327
rect 4893 5313 4907 5327
rect 6533 5313 6547 5327
rect 6713 5273 6727 5287
rect 6753 5273 6767 5287
rect 3393 5133 3407 5147
rect 3493 5133 3507 5147
rect 53 5093 67 5107
rect 113 5093 127 5107
rect 1993 5093 2007 5107
rect 2253 5094 2267 5108
rect 2293 5093 2307 5107
rect 4673 5093 4687 5107
rect 4793 5093 4807 5107
rect 4893 5093 4907 5107
rect 4933 5093 4947 5107
rect 5053 5093 5067 5107
rect 5133 5093 5147 5107
rect 5633 5093 5647 5107
rect 5713 5093 5727 5107
rect 5933 5093 5947 5107
rect 6013 5093 6027 5107
rect 6133 5094 6147 5108
rect 6193 5093 6207 5107
rect 4613 5073 4627 5087
rect 6173 5073 6187 5087
rect 2053 5033 2067 5047
rect 4533 5033 4547 5047
rect 5333 5033 5347 5047
rect 5373 5033 5387 5047
rect 6173 5033 6187 5047
rect 2273 5013 2287 5027
rect 2353 5013 2367 5027
rect 3913 5013 3927 5027
rect 3953 5013 3967 5027
rect 173 4993 187 5007
rect 273 4993 287 5007
rect 2713 4993 2727 5007
rect 2753 4993 2767 5007
rect 2513 4893 2527 4907
rect 2573 4893 2587 4907
rect 5213 4893 5227 4907
rect 5253 4893 5267 4907
rect 153 4873 167 4887
rect 233 4873 247 4887
rect 693 4873 707 4887
rect 733 4873 747 4887
rect 1733 4873 1747 4887
rect 2533 4873 2547 4887
rect 2593 4873 2607 4887
rect 4693 4873 4707 4887
rect 4773 4873 4787 4887
rect 5013 4873 5027 4887
rect 5053 4873 5067 4887
rect 6173 4873 6187 4887
rect 733 4793 747 4807
rect 793 4793 807 4807
rect 6213 4872 6227 4886
rect 6333 4873 6347 4887
rect 6413 4873 6427 4887
rect 2393 4853 2407 4867
rect 3613 4853 3627 4867
rect 2393 4813 2407 4827
rect 5553 4853 5567 4867
rect 5833 4853 5847 4867
rect 6513 4853 6527 4867
rect 3673 4813 3687 4827
rect 5493 4813 5507 4827
rect 5653 4813 5667 4827
rect 5713 4813 5727 4827
rect 5893 4813 5907 4827
rect 6513 4813 6527 4827
rect 6573 4853 6587 4867
rect 6653 4853 6667 4867
rect 6573 4813 6587 4827
rect 3773 4793 3787 4807
rect 3873 4793 3887 4807
rect 4273 4793 4287 4807
rect 4353 4793 4367 4807
rect 4733 4793 4747 4807
rect 4853 4793 4867 4807
rect 6633 4791 6647 4805
rect 4253 4773 4267 4787
rect 4313 4773 4327 4787
rect 4393 4773 4407 4787
rect 4453 4773 4467 4787
rect 1733 4752 1747 4766
rect 6213 4653 6227 4667
rect 6253 4652 6267 4666
rect 4633 4633 4647 4647
rect 4693 4633 4707 4647
rect 6373 4592 6387 4606
rect 6433 4593 6447 4607
rect 3433 4573 3447 4587
rect 3473 4572 3487 4586
rect 3613 4573 3627 4587
rect 3713 4573 3727 4587
rect 4393 4573 4407 4587
rect 4433 4573 4447 4587
rect 5133 4573 5147 4587
rect 5213 4574 5227 4588
rect 5293 4573 5307 4587
rect 5413 4573 5427 4587
rect 5533 4573 5547 4587
rect 6033 4573 6047 4587
rect 6073 4573 6087 4587
rect 6213 4573 6227 4587
rect 6313 4573 6327 4587
rect 2353 4553 2367 4567
rect 4813 4553 4827 4567
rect 5793 4553 5807 4567
rect 2413 4513 2427 4527
rect 4413 4513 4427 4527
rect 4453 4513 4467 4527
rect 4813 4513 4827 4527
rect 5113 4513 5127 4527
rect 5153 4513 5167 4527
rect 5513 4513 5527 4527
rect 5733 4513 5747 4527
rect 6233 4533 6247 4547
rect 6393 4533 6407 4547
rect 6173 4513 6187 4527
rect 6213 4513 6227 4527
rect 2493 4493 2507 4507
rect 2573 4493 2587 4507
rect 5453 4493 5467 4507
rect 5493 4493 5507 4507
rect 6353 4513 6367 4527
rect 6493 4513 6507 4527
rect 6533 4513 6547 4527
rect 6313 4493 6327 4507
rect 6473 4493 6487 4507
rect 6593 4493 6607 4507
rect 6653 4493 6667 4507
rect 6693 4493 6707 4507
rect 6493 4473 6507 4487
rect 6533 4473 6547 4487
rect 5933 4393 5947 4407
rect 5973 4393 5987 4407
rect 6453 4393 6467 4407
rect 2193 4353 2207 4367
rect 2293 4353 2307 4367
rect 3693 4353 3707 4367
rect 3753 4353 3767 4367
rect 853 4333 867 4347
rect 5153 4373 5167 4387
rect 5133 4353 5147 4367
rect 5173 4353 5187 4367
rect 5153 4333 5167 4347
rect 5833 4333 5847 4347
rect 5933 4333 5947 4347
rect 6233 4353 6247 4367
rect 913 4293 927 4307
rect 5313 4293 5327 4307
rect 5773 4293 5787 4307
rect 5813 4313 5827 4327
rect 5833 4293 5847 4307
rect 5933 4293 5947 4307
rect 6293 4333 6307 4347
rect 6353 4333 6367 4347
rect 6173 4293 6187 4307
rect 6673 4333 6687 4347
rect 833 4273 847 4287
rect 893 4273 907 4287
rect 3153 4273 3167 4287
rect 3273 4271 3287 4285
rect 4293 4273 4307 4287
rect 4393 4273 4407 4287
rect 4913 4273 4927 4287
rect 4993 4273 5007 4287
rect 5213 4273 5227 4287
rect 5393 4273 5407 4287
rect 6053 4273 6067 4287
rect 6113 4273 6127 4287
rect 6233 4273 6247 4287
rect 5293 4253 5307 4267
rect 5393 4252 5407 4266
rect 6373 4273 6387 4287
rect 6533 4271 6547 4285
rect 6653 4273 6667 4287
rect 6293 4253 6307 4267
rect 6353 4253 6367 4267
rect 6333 4232 6347 4246
rect 3833 4093 3847 4107
rect 3913 4093 3927 4107
rect 3673 4073 3687 4087
rect 3793 4073 3807 4087
rect 3673 4052 3687 4066
rect 3713 4052 3727 4066
rect 4233 4053 4247 4067
rect 4973 4053 4987 4067
rect 5033 4053 5047 4067
rect 5213 4053 5227 4067
rect 5253 4053 5267 4067
rect 5833 4054 5847 4068
rect 3913 4033 3927 4047
rect 3993 4033 4007 4047
rect 3993 3993 4007 4007
rect 4513 4033 4527 4047
rect 4213 3993 4227 4007
rect 3893 3972 3907 3986
rect 4173 3973 4187 3987
rect 4233 3973 4247 3987
rect 6233 4053 6247 4067
rect 6313 4054 6327 4068
rect 6533 4033 6547 4047
rect 5913 3993 5927 4007
rect 6373 3993 6387 4007
rect 6433 3993 6447 4007
rect 6593 3993 6607 4007
rect 4533 3973 4547 3987
rect 4753 3973 4767 3987
rect 4813 3973 4827 3987
rect 3533 3953 3547 3967
rect 3573 3953 3587 3967
rect 2253 3853 2267 3867
rect 2313 3853 2327 3867
rect 4993 3832 5007 3846
rect 3893 3813 3907 3827
rect 4533 3813 4547 3827
rect 3813 3773 3827 3787
rect 4753 3813 4767 3827
rect 5813 3813 5827 3827
rect 4593 3773 4607 3787
rect 4753 3773 4767 3787
rect 5053 3773 5067 3787
rect 6333 3813 6347 3827
rect 6593 3813 6607 3827
rect 5893 3773 5907 3787
rect 6253 3773 6267 3787
rect 6293 3773 6307 3787
rect 6333 3773 6347 3787
rect 6653 3813 6667 3827
rect 1213 3753 1227 3767
rect 1253 3753 1267 3767
rect 3513 3753 3527 3767
rect 3633 3753 3647 3767
rect 3673 3753 3687 3767
rect 3753 3753 3767 3767
rect 4533 3753 4547 3767
rect 4653 3753 4667 3767
rect 4693 3753 4707 3767
rect 4773 3753 4787 3767
rect 6133 3753 6147 3767
rect 6213 3753 6227 3767
rect 6613 3753 6627 3767
rect 6673 3753 6687 3767
rect 3553 3733 3567 3747
rect 3633 3732 3647 3746
rect 3293 3573 3307 3587
rect 3333 3573 3347 3587
rect 553 3533 567 3547
rect 593 3533 607 3547
rect 1593 3533 1607 3547
rect 1633 3533 1647 3547
rect 4613 3533 4627 3547
rect 4693 3533 4707 3547
rect 4753 3533 4767 3547
rect 4813 3533 4827 3547
rect 5213 3533 5227 3547
rect 5293 3533 5307 3547
rect 6033 3533 6047 3547
rect 1073 3513 1087 3527
rect 2793 3513 2807 3527
rect 4633 3513 4647 3527
rect 5513 3513 5527 3527
rect 433 3493 447 3507
rect 413 3473 427 3487
rect 1033 3473 1047 3487
rect 2793 3473 2807 3487
rect 4633 3473 4647 3487
rect 5053 3473 5067 3487
rect 5093 3473 5107 3487
rect 5513 3473 5527 3487
rect 5893 3513 5907 3527
rect 1053 3453 1067 3467
rect 1093 3453 1107 3467
rect 3313 3453 3327 3467
rect 3373 3453 3387 3467
rect 4173 3453 4187 3467
rect 4313 3453 4327 3467
rect 5833 3452 5847 3466
rect 5993 3473 6007 3487
rect 6233 3513 6247 3527
rect 6153 3473 6167 3487
rect 6313 3473 6327 3487
rect 6353 3473 6367 3487
rect 5853 3433 5867 3447
rect 5893 3433 5907 3447
rect 6653 3353 6667 3367
rect 6733 3352 6747 3366
rect 5833 3333 5847 3347
rect 1053 3293 1067 3307
rect 1073 3272 1087 3286
rect 4193 3293 4207 3307
rect 4193 3253 4207 3267
rect 4593 3233 4607 3247
rect 4633 3233 4647 3247
rect 5313 3233 5327 3247
rect 5453 3233 5467 3247
rect 5673 3233 5687 3247
rect 6053 3293 6067 3307
rect 6153 3293 6167 3307
rect 6013 3252 6027 3266
rect 6373 3293 6387 3307
rect 6553 3293 6567 3307
rect 6313 3253 6327 3267
rect 6553 3253 6567 3267
rect 5733 3232 5747 3246
rect 5853 3232 5867 3246
rect 6173 3232 6187 3246
rect 6493 3233 6507 3247
rect 6573 3231 6587 3245
rect 4893 3193 4907 3207
rect 4993 3193 5007 3207
rect 1073 3093 1087 3107
rect 1133 3073 1147 3087
rect 4553 3033 4567 3047
rect 4713 3033 4727 3047
rect 6213 3033 6227 3047
rect 6273 3033 6287 3047
rect 2813 3013 2827 3027
rect 2953 3013 2967 3027
rect 3213 3013 3227 3027
rect 3273 3013 3287 3027
rect 3313 3013 3327 3027
rect 3413 3013 3427 3027
rect 3973 3012 3987 3026
rect 4013 3013 4027 3027
rect 4053 3013 4067 3027
rect 4093 3013 4107 3027
rect 4253 3013 4267 3027
rect 4293 2993 4307 3007
rect 4693 3013 4707 3027
rect 4913 3013 4927 3027
rect 4993 3013 5007 3027
rect 6233 3013 6247 3027
rect 773 2953 787 2967
rect 813 2953 827 2967
rect 4113 2953 4127 2967
rect 4173 2953 4187 2967
rect 6313 3012 6327 3026
rect 4353 2953 4367 2967
rect 6173 2993 6187 3007
rect 4913 2953 4927 2967
rect 6473 3014 6487 3028
rect 6253 2953 6267 2967
rect 6413 2953 6427 2967
rect 2993 2933 3007 2947
rect 3113 2933 3127 2947
rect 4473 2933 4487 2947
rect 4513 2933 4527 2947
rect 4613 2932 4627 2946
rect 5853 2933 5867 2947
rect 5933 2933 5947 2947
rect 2953 2793 2967 2807
rect 3013 2793 3027 2807
rect 4053 2793 4067 2807
rect 4113 2793 4127 2807
rect 6613 2793 6627 2807
rect 6693 2793 6707 2807
rect 3673 2773 3687 2787
rect 3713 2773 3727 2787
rect 4333 2773 4347 2787
rect 4373 2773 4387 2787
rect 6073 2773 6087 2787
rect 3673 2733 3687 2747
rect 3733 2733 3747 2747
rect 6073 2733 6087 2747
rect 6133 2773 6147 2787
rect 6293 2773 6307 2787
rect 6133 2733 6147 2747
rect 6293 2733 6307 2747
rect 6453 2773 6467 2787
rect 1033 2713 1047 2727
rect 1113 2713 1127 2727
rect 1753 2713 1767 2727
rect 1833 2711 1847 2725
rect 1933 2713 1947 2727
rect 1973 2713 1987 2727
rect 3533 2713 3547 2727
rect 3593 2713 3607 2727
rect 4513 2713 4527 2727
rect 4573 2713 4587 2727
rect 5673 2713 5687 2727
rect 5813 2713 5827 2727
rect 6213 2713 6227 2727
rect 6253 2713 6267 2727
rect 6373 2713 6387 2727
rect 1873 2693 1887 2707
rect 1953 2692 1967 2706
rect 6373 2692 6387 2706
rect 6433 2693 6447 2707
rect 5593 2513 5607 2527
rect 5633 2513 5647 2527
rect 5813 2513 5827 2527
rect 793 2493 807 2507
rect 933 2493 947 2507
rect 873 2473 887 2487
rect 913 2473 927 2487
rect 2413 2493 2427 2507
rect 2913 2493 2927 2507
rect 3013 2493 3027 2507
rect 2333 2433 2347 2447
rect 2393 2473 2407 2487
rect 4533 2493 4547 2507
rect 5733 2493 5747 2507
rect 5993 2493 6007 2507
rect 6133 2493 6147 2507
rect 6513 2493 6527 2507
rect 6573 2493 6587 2507
rect 5933 2473 5947 2487
rect 6093 2473 6107 2487
rect 6593 2473 6607 2487
rect 2393 2433 2407 2447
rect 4493 2433 4507 2447
rect 5253 2433 5267 2447
rect 5293 2433 5307 2447
rect 5873 2433 5887 2447
rect 6093 2433 6107 2447
rect 6593 2433 6607 2447
rect 813 2413 827 2427
rect 873 2413 887 2427
rect 4713 2411 4727 2425
rect 4793 2413 4807 2427
rect 6213 2392 6227 2406
rect 6253 2393 6267 2407
rect 5833 2313 5847 2327
rect 5793 2293 5807 2307
rect 4233 2273 4247 2287
rect 4313 2273 4327 2287
rect 4493 2273 4507 2287
rect 6453 2274 6467 2288
rect 6533 2273 6547 2287
rect 5073 2253 5087 2267
rect 4493 2213 4507 2227
rect 5593 2253 5607 2267
rect 5633 2253 5647 2267
rect 5993 2253 6007 2267
rect 6073 2253 6087 2267
rect 5153 2213 5167 2227
rect 5933 2213 5947 2227
rect 6133 2213 6147 2227
rect 393 2193 407 2207
rect 513 2193 527 2207
rect 4233 2193 4247 2207
rect 4333 2193 4347 2207
rect 4793 2191 4807 2205
rect 4893 2193 4907 2207
rect 5573 2193 5587 2207
rect 5673 2193 5687 2207
rect 6213 2192 6227 2206
rect 6273 2193 6287 2207
rect 2673 2153 2687 2167
rect 2733 2152 2747 2166
rect 6533 2053 6547 2067
rect 6573 2053 6587 2067
rect 1333 1993 1347 2007
rect 1453 1993 1467 2007
rect 4853 1993 4867 2007
rect 4913 1993 4927 2007
rect 6553 1993 6567 2007
rect 6653 1993 6667 2007
rect 813 1973 827 1987
rect 913 1973 927 1987
rect 993 1973 1007 1987
rect 1353 1973 1367 1987
rect 1413 1973 1427 1987
rect 2213 1953 2227 1967
rect 2253 1953 2267 1967
rect 3173 1953 3187 1967
rect 4113 1973 4127 1987
rect 4173 1973 4187 1987
rect 4213 1973 4227 1987
rect 4333 1973 4347 1987
rect 4393 1973 4407 1987
rect 4573 1973 4587 1987
rect 4673 1973 4687 1987
rect 393 1913 407 1927
rect 473 1913 487 1927
rect 3113 1913 3127 1927
rect 3633 1893 3647 1907
rect 3733 1891 3747 1905
rect 4693 1953 4707 1967
rect 4693 1913 4707 1927
rect 4973 1973 4987 1987
rect 4873 1953 4887 1967
rect 4913 1952 4927 1966
rect 4993 1953 5007 1967
rect 4773 1913 4787 1927
rect 4993 1913 5007 1927
rect 4113 1893 4127 1907
rect 4553 1892 4567 1906
rect 4973 1893 4987 1907
rect 6693 1953 6707 1967
rect 6693 1913 6707 1927
rect 5593 1893 5607 1907
rect 5673 1893 5687 1907
rect 5713 1891 5727 1905
rect 5773 1893 5787 1907
rect 6253 1893 6267 1907
rect 6373 1893 6387 1907
rect 4053 1754 4067 1768
rect 2813 1733 2827 1747
rect 3613 1733 3627 1747
rect 3933 1733 3947 1747
rect 6493 1753 6507 1767
rect 6613 1753 6627 1767
rect 2813 1693 2827 1707
rect 3673 1693 3687 1707
rect 833 1673 847 1687
rect 893 1673 907 1687
rect 3333 1673 3347 1687
rect 3393 1673 3407 1687
rect 3913 1671 3927 1685
rect 3953 1673 3967 1687
rect 6313 1733 6327 1747
rect 6393 1733 6407 1747
rect 6653 1733 6667 1747
rect 6733 1733 6747 1747
rect 4093 1693 4107 1707
rect 4033 1671 4047 1685
rect 4073 1673 4087 1687
rect 4193 1673 4207 1687
rect 4733 1673 4747 1687
rect 5653 1673 5667 1687
rect 5793 1673 5807 1687
rect 3953 1652 3967 1666
rect 4673 1653 4687 1667
rect 3793 1593 3807 1607
rect 3833 1593 3847 1607
rect 4653 1513 4667 1527
rect 3973 1493 3987 1507
rect 4073 1493 4087 1507
rect 4713 1493 4727 1507
rect 3253 1453 3267 1467
rect 3313 1452 3327 1466
rect 3513 1453 3527 1467
rect 3613 1454 3627 1468
rect 3653 1453 3667 1467
rect 3813 1453 3827 1467
rect 4633 1453 4647 1467
rect 4713 1453 4727 1467
rect 5353 1453 5367 1467
rect 5513 1453 5527 1467
rect 6333 1452 6347 1466
rect 6412 1453 6426 1467
rect 6433 1453 6447 1467
rect 3493 1433 3507 1447
rect 3533 1433 3547 1447
rect 6733 1433 6747 1447
rect 4493 1393 4507 1407
rect 4553 1393 4567 1407
rect 6453 1393 6467 1407
rect 6553 1393 6567 1407
rect 6613 1393 6627 1407
rect 6733 1393 6747 1407
rect 3473 1373 3487 1387
rect 3533 1373 3547 1387
rect 5593 1373 5607 1387
rect 5653 1373 5667 1387
rect 5413 1333 5427 1347
rect 5453 1332 5467 1346
rect 5713 1333 5727 1347
rect 5753 1333 5767 1347
rect 333 1213 347 1227
rect 373 1213 387 1227
rect 1073 1213 1087 1227
rect 1113 1213 1127 1227
rect 1373 1213 1387 1227
rect 1413 1213 1427 1227
rect 2153 1173 2167 1187
rect 2193 1173 2207 1187
rect 4033 1213 4047 1227
rect 4133 1213 4147 1227
rect 5733 1213 5747 1227
rect 4373 1193 4387 1207
rect 513 1153 527 1167
rect 593 1153 607 1167
rect 1993 1153 2007 1167
rect 2073 1151 2087 1165
rect 2293 1153 2307 1167
rect 2353 1153 2367 1167
rect 2613 1153 2627 1167
rect 2673 1153 2687 1167
rect 3473 1153 3487 1167
rect 3553 1153 3567 1167
rect 3893 1153 3907 1167
rect 4133 1173 4147 1187
rect 4333 1173 4347 1187
rect 5733 1173 5747 1187
rect 5953 1213 5967 1227
rect 6193 1213 6207 1227
rect 6253 1212 6267 1226
rect 4293 1153 4307 1167
rect 4373 1153 4387 1167
rect 4753 1153 4767 1167
rect 4873 1153 4887 1167
rect 5853 1153 5867 1167
rect 3953 1113 3967 1127
rect 4013 1113 4027 1127
rect 1673 953 1687 967
rect 1813 953 1827 967
rect 1013 933 1027 947
rect 1073 933 1087 947
rect 1233 933 1247 947
rect 1293 933 1307 947
rect 1433 933 1447 947
rect 1473 934 1487 948
rect 4133 933 4147 947
rect 4273 933 4287 947
rect 4953 933 4967 947
rect 4993 933 5007 947
rect 5913 933 5927 947
rect 6073 933 6087 947
rect 2513 853 2527 867
rect 2573 853 2587 867
rect 2613 853 2627 867
rect 2673 853 2687 867
rect 2853 853 2867 867
rect 2953 853 2967 867
rect 6153 853 6167 867
rect 6233 853 6247 867
rect 3813 733 3827 747
rect 1373 713 1387 727
rect 1413 713 1427 727
rect 2113 713 2127 727
rect 2253 713 2267 727
rect 2453 713 2467 727
rect 2513 713 2527 727
rect 3833 713 3847 727
rect 3873 713 3887 727
rect 4293 713 4307 727
rect 4373 713 4387 727
rect 5113 713 5127 727
rect 5193 713 5207 727
rect 2133 693 2147 707
rect 2173 693 2187 707
rect 3813 693 3827 707
rect 4093 693 4107 707
rect 4153 653 4167 667
rect 613 633 627 647
rect 753 633 767 647
rect 1953 633 1967 647
rect 2013 631 2027 645
rect 3773 633 3787 647
rect 3853 633 3867 647
rect 3933 633 3947 647
rect 4053 633 4067 647
rect 4253 633 4267 647
rect 4373 633 4387 647
rect 4573 633 4587 647
rect 4713 631 4727 645
rect 5073 633 5087 647
rect 5193 633 5207 647
rect 5373 633 5387 647
rect 5513 633 5527 647
rect 6053 633 6067 647
rect 6153 633 6167 647
rect 6633 633 6647 647
rect 6673 633 6687 647
rect 573 613 587 627
rect 693 613 707 627
rect 4313 613 4327 627
rect 5393 613 5407 627
rect 4253 592 4267 606
rect 5493 612 5507 626
rect 4333 433 4347 447
rect 4393 433 4407 447
rect 313 413 327 427
rect 413 413 427 427
rect 4273 413 4287 427
rect 4413 412 4427 426
rect 4473 413 4487 427
rect 4573 413 4587 427
rect 5373 413 5387 427
rect 2873 393 2887 407
rect 4973 393 4987 407
rect 5033 393 5047 407
rect 6473 413 6487 427
rect 2813 353 2827 367
rect 5413 353 5427 367
rect 6573 353 6587 367
rect 3613 331 3627 345
rect 3713 333 3727 347
rect 4253 333 4267 347
rect 4313 333 4327 347
rect 4353 333 4367 347
rect 5633 333 5647 347
rect 5713 333 5727 347
rect 633 233 647 247
rect 4573 233 4587 247
rect 4633 233 4647 247
rect 673 213 687 227
rect 4453 193 4467 207
rect 1393 153 1407 167
rect 1433 133 1447 147
rect 1713 133 1727 147
rect 1753 133 1767 147
rect 3273 133 3287 147
rect 3313 133 3327 147
rect 4393 133 4407 147
rect 6293 133 6307 147
rect 6333 133 6347 147
rect 393 113 407 127
rect 553 113 567 127
rect 1393 113 1407 127
rect 1493 113 1507 127
rect 4253 113 4267 127
rect 4293 113 4307 127
rect 4433 113 4447 127
rect 4513 113 4527 127
rect 5993 112 6007 126
rect 6053 113 6067 127
rect 613 93 627 107
rect 713 93 727 107
<< metal2 >>
rect 76 6376 103 6383
rect 76 6367 83 6376
rect 76 6027 83 6353
rect 156 6327 163 6383
rect 176 6116 183 6453
rect 216 6128 223 6414
rect 536 6427 543 6493
rect 576 6416 583 6453
rect 816 6416 863 6423
rect 376 6386 383 6413
rect 256 6127 263 6383
rect 296 6380 303 6383
rect 293 6367 307 6380
rect 456 6327 463 6372
rect 596 6227 603 6383
rect 116 6027 123 6083
rect 116 5827 123 5863
rect 216 5843 223 6114
rect 296 6116 303 6153
rect 453 6120 467 6133
rect 456 6116 463 6120
rect 496 6116 543 6123
rect 536 6107 543 6116
rect 356 6080 363 6083
rect 353 6067 367 6080
rect 236 5863 243 5894
rect 236 5856 283 5863
rect 216 5836 243 5843
rect 236 5627 243 5836
rect 216 5596 243 5603
rect 56 5347 63 5552
rect 216 5387 223 5533
rect 236 5507 243 5596
rect 256 5483 263 5856
rect 316 5707 323 5852
rect 356 5727 363 6013
rect 536 5987 543 6093
rect 556 6087 563 6213
rect 596 6116 603 6173
rect 436 5896 443 5933
rect 376 5866 383 5893
rect 516 5866 523 5933
rect 576 5896 583 5973
rect 656 5967 663 6133
rect 736 6116 743 6153
rect 796 6143 803 6413
rect 816 6187 823 6416
rect 1276 6416 1283 6493
rect 1396 6416 1403 6453
rect 1476 6427 1483 6453
rect 916 6380 923 6383
rect 913 6367 927 6380
rect 776 6136 803 6143
rect 776 6128 783 6136
rect 856 6086 863 6153
rect 936 6116 943 6173
rect 956 6167 963 6413
rect 1016 6380 1023 6383
rect 1013 6367 1027 6380
rect 1056 6207 1063 6373
rect 1136 6347 1143 6383
rect 1176 6380 1183 6383
rect 1173 6367 1187 6380
rect 1336 6367 1343 6413
rect 1516 6386 1523 6453
rect 1736 6416 1743 6453
rect 1536 6367 1543 6413
rect 1596 6287 1603 6383
rect 1676 6347 1683 6414
rect 1056 6116 1063 6193
rect 1196 6116 1203 6173
rect 1236 6116 1243 6193
rect 796 6067 803 6083
rect 956 6076 983 6083
rect 796 6056 813 6067
rect 800 6053 813 6056
rect 947 6053 953 6067
rect 456 5827 463 5863
rect 596 5827 603 5863
rect 276 5567 283 5693
rect 456 5667 463 5813
rect 356 5596 403 5603
rect 396 5507 403 5596
rect 416 5566 423 5653
rect 453 5600 467 5613
rect 456 5596 463 5600
rect 616 5596 623 5653
rect 656 5627 663 5953
rect 716 5896 723 5933
rect 796 5867 803 5913
rect 836 5896 843 5953
rect 873 5900 887 5913
rect 876 5896 883 5900
rect 896 5860 903 5863
rect 893 5847 907 5860
rect 656 5596 663 5613
rect 776 5608 783 5813
rect 516 5547 523 5563
rect 236 5476 263 5483
rect 76 5336 93 5343
rect 56 4707 63 5093
rect 76 5087 83 5336
rect 116 5107 123 5133
rect 113 5080 127 5093
rect 116 5076 123 5080
rect 116 4856 123 5013
rect 153 4867 167 4873
rect 96 4567 103 4823
rect 136 4707 143 4823
rect 176 4647 183 4993
rect 196 4767 203 5074
rect 216 5047 223 5332
rect 236 5267 243 5476
rect 516 5383 523 5533
rect 556 5483 563 5594
rect 636 5487 643 5563
rect 547 5476 563 5483
rect 496 5376 523 5383
rect 236 5027 243 5193
rect 296 5076 303 5253
rect 336 5247 343 5343
rect 476 5327 483 5343
rect 476 5316 493 5327
rect 480 5313 493 5316
rect 536 5303 543 5473
rect 676 5407 683 5563
rect 613 5380 627 5393
rect 616 5376 623 5380
rect 656 5376 703 5383
rect 636 5340 643 5343
rect 633 5327 647 5340
rect 696 5307 703 5376
rect 736 5346 743 5593
rect 836 5563 843 5833
rect 956 5596 963 5833
rect 976 5603 983 6076
rect 1016 6067 1023 6114
rect 1076 6047 1083 6083
rect 1216 6080 1223 6083
rect 1213 6067 1227 6080
rect 1056 5896 1063 5933
rect 1236 5896 1243 5933
rect 1256 5903 1263 6083
rect 1296 6047 1303 6193
rect 1376 6116 1383 6153
rect 1356 6007 1363 6083
rect 1456 5947 1463 6114
rect 1476 6087 1483 6233
rect 1696 6227 1703 6372
rect 1756 6367 1763 6383
rect 1576 6167 1583 6193
rect 1607 6173 1613 6187
rect 1647 6173 1653 6187
rect 1676 6167 1683 6193
rect 1736 6167 1743 6273
rect 1756 6247 1763 6353
rect 1836 6307 1843 6414
rect 1896 6380 1903 6383
rect 1893 6367 1907 6380
rect 1973 6367 1987 6372
rect 2016 6347 2023 6393
rect 1660 6166 1683 6167
rect 1536 6116 1543 6153
rect 1667 6156 1683 6166
rect 1667 6153 1680 6156
rect 1516 6007 1523 6083
rect 1427 5933 1433 5947
rect 1473 5927 1487 5933
rect 1256 5896 1283 5903
rect 1096 5867 1103 5894
rect 1076 5807 1083 5863
rect 1156 5807 1163 5894
rect 1276 5703 1283 5896
rect 1400 5903 1413 5907
rect 1396 5896 1413 5903
rect 1400 5893 1413 5896
rect 1296 5847 1303 5893
rect 1336 5807 1343 5863
rect 1476 5807 1483 5892
rect 1516 5867 1523 5993
rect 1616 5987 1623 6152
rect 1736 6087 1743 6153
rect 1696 5967 1703 6083
rect 1756 6067 1763 6113
rect 1776 6087 1783 6293
rect 1876 6116 1923 6123
rect 1856 6080 1863 6083
rect 1853 6067 1867 6080
rect 1916 6007 1923 6116
rect 1936 6087 1943 6333
rect 2036 6327 2043 6413
rect 2076 6167 2083 6383
rect 2127 6355 2153 6362
rect 2176 6287 2183 6372
rect 2216 6327 2223 6372
rect 2313 6362 2327 6373
rect 2336 6367 2343 6493
rect 2267 6360 2327 6362
rect 2267 6355 2323 6360
rect 2356 6287 2363 6414
rect 2656 6427 2663 6563
rect 2836 6527 2843 6563
rect 2996 6527 3003 6563
rect 2696 6428 2703 6473
rect 2456 6327 2463 6413
rect 2516 6347 2523 6383
rect 2616 6347 2623 6413
rect 2636 6347 2643 6414
rect 2736 6416 2743 6453
rect 2116 6227 2123 6273
rect 2036 6116 2083 6123
rect 2136 6116 2143 6193
rect 2016 6007 2023 6083
rect 1547 5913 1553 5927
rect 1727 5913 1733 5927
rect 1640 5903 1653 5907
rect 1636 5896 1653 5903
rect 1640 5893 1653 5896
rect 1793 5900 1807 5913
rect 1796 5896 1803 5900
rect 1916 5896 1923 5972
rect 2076 5967 2083 6116
rect 1596 5860 1603 5863
rect 1593 5847 1607 5860
rect 1776 5847 1783 5863
rect 1787 5836 1803 5843
rect 1336 5743 1343 5793
rect 1336 5736 1363 5743
rect 1256 5696 1283 5703
rect 976 5596 1003 5603
rect 796 5556 843 5563
rect 896 5560 903 5563
rect 893 5547 907 5560
rect 876 5536 893 5543
rect 796 5407 803 5453
rect 793 5380 807 5393
rect 796 5376 803 5380
rect 876 5346 883 5536
rect 936 5407 943 5563
rect 996 5527 1003 5596
rect 1136 5596 1143 5673
rect 1096 5467 1103 5563
rect 1116 5443 1123 5553
rect 1236 5547 1243 5673
rect 1256 5667 1263 5696
rect 1096 5436 1123 5443
rect 896 5346 903 5393
rect 1096 5376 1103 5436
rect 1136 5376 1143 5413
rect 976 5307 983 5343
rect 516 5296 543 5303
rect 276 5007 283 5043
rect 240 4943 253 4947
rect 236 4933 253 4943
rect 236 4887 243 4933
rect 233 4860 247 4873
rect 236 4856 243 4860
rect 256 4783 263 4823
rect 256 4776 283 4783
rect 36 4067 43 4353
rect 96 4336 103 4553
rect 116 4367 123 4633
rect 216 4556 223 4653
rect 256 4507 263 4753
rect 96 4007 103 4273
rect 116 4247 123 4303
rect 156 4287 163 4493
rect 276 4487 283 4776
rect 296 4667 303 5013
rect 316 4627 323 5033
rect 336 5027 343 5233
rect 356 5047 363 5074
rect 416 4927 423 5043
rect 516 5007 523 5296
rect 1016 5287 1023 5373
rect 647 5076 663 5083
rect 656 5007 663 5076
rect 736 5076 763 5083
rect 416 4863 423 4913
rect 676 4907 683 5073
rect 696 4947 703 4973
rect 416 4856 443 4863
rect 436 4823 443 4856
rect 456 4826 463 4853
rect 576 4826 583 4893
rect 680 4883 693 4887
rect 676 4873 693 4883
rect 676 4856 683 4873
rect 716 4867 723 4933
rect 736 4927 743 5076
rect 776 5023 783 5032
rect 756 5016 783 5023
rect 356 4767 363 4823
rect 396 4816 443 4823
rect 616 4807 623 4853
rect 656 4820 663 4823
rect 653 4807 667 4820
rect 736 4807 743 4873
rect 756 4807 763 5016
rect 856 4856 863 4933
rect 956 4887 963 5043
rect 996 4947 1003 5043
rect 996 4856 1003 4912
rect 1036 4868 1043 5353
rect 1076 5207 1083 5343
rect 1116 5143 1123 5332
rect 1196 5247 1203 5533
rect 1316 5376 1323 5473
rect 1356 5467 1363 5736
rect 1416 5427 1423 5633
rect 1476 5596 1483 5633
rect 1536 5547 1543 5713
rect 1636 5596 1643 5673
rect 1556 5567 1563 5594
rect 1716 5566 1723 5733
rect 1776 5596 1783 5773
rect 1796 5747 1803 5836
rect 1816 5827 1823 5863
rect 1876 5787 1883 5894
rect 1936 5860 1943 5863
rect 1933 5847 1947 5860
rect 1976 5827 1983 5852
rect 2016 5847 2023 5913
rect 2096 5896 2103 6093
rect 2216 6087 2223 6173
rect 2156 6047 2163 6083
rect 2133 5900 2147 5913
rect 2136 5896 2143 5900
rect 2316 5896 2323 5993
rect 2356 5987 2363 6273
rect 2416 6116 2423 6253
rect 2456 6116 2463 6313
rect 2516 6083 2523 6193
rect 2476 6076 2523 6083
rect 1896 5627 1903 5673
rect 1916 5596 1923 5673
rect 1976 5567 1983 5813
rect 2156 5787 2163 5863
rect 2176 5807 2183 5852
rect 2016 5727 2023 5753
rect 2056 5727 2063 5753
rect 2036 5596 2043 5673
rect 2056 5627 2063 5673
rect 2176 5596 2183 5793
rect 2236 5747 2243 5894
rect 2376 5867 2383 5913
rect 1616 5560 1623 5563
rect 1613 5547 1627 5560
rect 1456 5346 1463 5373
rect 1256 5167 1263 5343
rect 1356 5247 1363 5343
rect 1576 5167 1583 5374
rect 1656 5376 1663 5513
rect 1876 5416 1883 5453
rect 1916 5376 1943 5383
rect 1107 5136 1123 5143
rect 1096 5076 1103 5133
rect 1176 5047 1183 5153
rect 1616 5127 1623 5373
rect 1676 5287 1683 5343
rect 1716 5227 1723 5343
rect 1273 5080 1287 5093
rect 1276 5076 1283 5080
rect 1196 4987 1203 5074
rect 1376 5043 1383 5093
rect 1496 5076 1523 5083
rect 1516 5067 1523 5076
rect 1256 4947 1263 5043
rect 1376 5036 1403 5043
rect 1516 4947 1523 5053
rect 796 4820 803 4823
rect 793 4807 807 4820
rect 836 4807 843 4823
rect 756 4767 763 4793
rect 296 4616 313 4623
rect 296 4526 303 4616
rect 353 4560 367 4573
rect 356 4556 363 4560
rect 436 4527 443 4554
rect 336 4487 343 4523
rect 456 4487 463 4693
rect 836 4687 843 4793
rect 936 4787 943 4853
rect 1016 4787 1023 4823
rect 516 4556 523 4613
rect 336 4447 343 4473
rect 196 4306 203 4353
rect 276 4127 283 4292
rect 116 3967 123 4034
rect 136 3816 143 3993
rect 116 3727 123 3783
rect 196 3727 203 3772
rect 256 3767 263 4034
rect 296 4007 303 4213
rect 316 4087 323 4333
rect 336 4307 343 4393
rect 396 4348 403 4473
rect 476 4407 483 4554
rect 576 4306 583 4333
rect 376 4227 383 4303
rect 416 4300 423 4303
rect 413 4287 427 4300
rect 476 4227 483 4303
rect 596 4227 603 4653
rect 1056 4568 1063 4873
rect 1076 4826 1083 4853
rect 1116 4787 1123 4812
rect 1176 4787 1183 4823
rect 976 4560 1003 4563
rect 976 4556 1007 4560
rect 993 4547 1007 4556
rect 1236 4556 1243 4893
rect 1316 4856 1323 4893
rect 1476 4856 1483 4913
rect 1636 4887 1643 5043
rect 1656 4856 1663 5033
rect 1676 4863 1683 5073
rect 1696 5046 1703 5113
rect 1756 5076 1763 5332
rect 1936 5187 1943 5376
rect 1996 5183 2003 5573
rect 2156 5487 2163 5552
rect 2146 5473 2147 5480
rect 2133 5463 2147 5473
rect 2133 5460 2163 5463
rect 2136 5456 2167 5460
rect 2153 5447 2167 5456
rect 2176 5388 2183 5513
rect 2216 5447 2223 5513
rect 2236 5427 2243 5733
rect 2256 5727 2263 5773
rect 2396 5747 2403 5953
rect 2296 5608 2303 5713
rect 2256 5447 2263 5593
rect 2376 5527 2383 5673
rect 2436 5596 2443 5633
rect 2476 5596 2483 5733
rect 2496 5727 2503 5933
rect 2396 5563 2403 5594
rect 2396 5556 2423 5563
rect 2336 5467 2343 5513
rect 2016 5336 2043 5343
rect 2016 5287 2023 5336
rect 1996 5176 2023 5183
rect 1736 4927 1743 5043
rect 1776 5007 1783 5043
rect 1816 4987 1823 5093
rect 1993 5088 2007 5093
rect 1856 5007 1863 5074
rect 1936 4987 1943 5043
rect 1733 4887 1747 4892
rect 1676 4856 1703 4863
rect 1396 4826 1403 4853
rect 1696 4826 1703 4856
rect 776 4516 803 4523
rect 796 4487 803 4516
rect 856 4516 883 4523
rect 736 4480 743 4483
rect 733 4467 747 4480
rect 656 4336 663 4413
rect 356 4048 363 4113
rect 396 4036 403 4073
rect 336 3783 343 3992
rect 376 3967 383 4003
rect 296 3780 303 3783
rect 293 3767 307 3780
rect 316 3776 343 3783
rect 156 3467 163 3713
rect 167 3456 183 3463
rect 136 3296 143 3373
rect 113 3000 127 3013
rect 116 2996 123 3000
rect 176 2863 183 3456
rect 196 3307 203 3673
rect 256 3516 263 3553
rect 236 3480 243 3483
rect 233 3467 247 3480
rect 296 3447 303 3473
rect 276 3263 283 3293
rect 256 3256 283 3263
rect 256 3127 263 3256
rect 156 2856 183 2863
rect 36 2687 43 2743
rect 16 2183 23 2633
rect 36 2347 43 2673
rect 56 2527 63 2573
rect 136 2476 143 2853
rect 156 2487 163 2856
rect 216 2788 223 2893
rect 316 2867 323 3776
rect 356 3528 363 3833
rect 396 3567 403 3933
rect 436 3847 443 4133
rect 476 4067 483 4213
rect 556 4036 563 4093
rect 593 4040 607 4053
rect 596 4036 603 4040
rect 496 3947 503 4003
rect 416 3687 423 3783
rect 476 3780 483 3783
rect 473 3767 487 3780
rect 536 3776 563 3783
rect 433 3507 447 3514
rect 336 3427 343 3473
rect 413 3467 427 3473
rect 436 3447 443 3472
rect 456 3447 463 3553
rect 556 3547 563 3776
rect 576 3687 583 3853
rect 596 3727 603 3973
rect 696 3827 703 4433
rect 836 4348 843 4413
rect 856 4347 863 4516
rect 1076 4467 1083 4523
rect 1216 4427 1223 4523
rect 716 3987 723 4334
rect 836 4247 843 4273
rect 876 4247 883 4334
rect 896 4287 903 4353
rect 933 4340 947 4353
rect 936 4336 943 4340
rect 976 4336 983 4373
rect 1036 4306 1043 4333
rect 1296 4306 1303 4373
rect 816 4236 833 4243
rect 716 3816 723 3913
rect 816 3823 823 4236
rect 836 4006 843 4033
rect 876 4007 883 4093
rect 916 4048 923 4293
rect 956 4287 963 4303
rect 1116 4300 1123 4303
rect 1113 4287 1127 4300
rect 956 4048 963 4273
rect 1196 4227 1203 4303
rect 1276 4048 1283 4253
rect 1316 4147 1323 4633
rect 1356 4556 1363 4773
rect 1396 4556 1403 4812
rect 1436 4787 1443 4823
rect 1596 4787 1603 4812
rect 1736 4787 1743 4852
rect 1376 4467 1383 4523
rect 1416 4443 1423 4523
rect 1456 4507 1463 4673
rect 1416 4436 1443 4443
rect 1416 4227 1423 4413
rect 1436 4143 1443 4436
rect 1456 4347 1463 4453
rect 1436 4136 1463 4143
rect 996 3967 1003 4034
rect 1196 4036 1223 4043
rect 796 3816 823 3823
rect 696 3647 703 3773
rect 576 3528 583 3553
rect 776 3543 783 3813
rect 756 3536 783 3543
rect 596 3487 603 3533
rect 376 3260 383 3263
rect 373 3247 387 3260
rect 216 2643 223 2713
rect 276 2687 283 2743
rect 336 2740 343 2743
rect 333 2727 347 2740
rect 196 2636 223 2643
rect 36 2227 43 2293
rect 16 2176 43 2183
rect 16 1447 23 1833
rect 36 1507 43 2176
rect 56 2007 63 2473
rect 196 2447 203 2636
rect 256 2476 263 2533
rect 116 2307 123 2443
rect 216 2436 243 2443
rect 96 2220 103 2223
rect 93 2207 107 2220
rect 76 1967 83 2053
rect 96 1956 103 1993
rect 136 1956 143 2212
rect 176 2107 183 2333
rect 216 2223 223 2436
rect 276 2256 283 2293
rect 216 2216 233 2223
rect 176 1956 183 2093
rect 296 1968 303 2273
rect 336 2187 343 2533
rect 356 2307 363 2733
rect 376 2687 383 3233
rect 396 2788 403 3413
rect 436 3260 443 3263
rect 433 3247 447 3260
rect 436 3207 443 3233
rect 536 3147 543 3413
rect 556 3407 563 3472
rect 616 3427 623 3514
rect 656 3447 663 3483
rect 556 3266 563 3393
rect 756 3303 763 3536
rect 776 3487 783 3514
rect 756 3296 783 3303
rect 556 3087 563 3252
rect 676 3207 683 3263
rect 747 3256 763 3263
rect 756 3227 763 3256
rect 556 3047 563 3073
rect 416 2996 423 3033
rect 456 2907 463 2963
rect 516 2947 523 3013
rect 556 2996 563 3033
rect 576 2960 583 2963
rect 573 2947 587 2960
rect 376 2527 383 2673
rect 396 2647 403 2774
rect 496 2707 503 2773
rect 516 2667 523 2813
rect 576 2776 583 2853
rect 636 2827 643 2994
rect 656 2967 663 3093
rect 693 3000 707 3013
rect 696 2996 703 3000
rect 736 2996 743 3053
rect 776 3007 783 3296
rect 760 2963 773 2967
rect 756 2956 773 2963
rect 760 2953 773 2956
rect 796 2966 803 3816
rect 936 3783 943 3893
rect 896 3776 943 3783
rect 836 3516 843 3633
rect 896 3407 903 3483
rect 856 3296 863 3333
rect 896 3308 903 3393
rect 816 2967 823 3073
rect 836 3027 843 3133
rect 936 3067 943 3653
rect 956 3487 963 3953
rect 1036 3907 1043 4033
rect 976 3786 983 3873
rect 1016 3528 1023 3753
rect 1036 3727 1043 3783
rect 1096 3687 1103 3913
rect 1196 3867 1203 4036
rect 1356 4043 1363 4113
rect 1456 4087 1463 4136
rect 1336 4036 1363 4043
rect 1476 4043 1483 4693
rect 1516 4647 1523 4713
rect 1536 4556 1543 4653
rect 1716 4556 1723 4653
rect 1736 4627 1743 4752
rect 1796 4556 1823 4563
rect 1876 4556 1883 4933
rect 1896 4827 1903 4913
rect 1976 4907 1983 5043
rect 2016 4987 2023 5176
rect 2036 5046 2043 5173
rect 2056 5083 2063 5253
rect 2156 5207 2163 5353
rect 2196 5347 2203 5413
rect 2296 5407 2303 5433
rect 2253 5380 2267 5393
rect 2256 5376 2263 5380
rect 2296 5376 2303 5393
rect 2236 5340 2243 5343
rect 2233 5327 2247 5340
rect 2176 5127 2183 5253
rect 2196 5247 2203 5312
rect 2316 5287 2323 5343
rect 2056 5076 2083 5083
rect 2053 5027 2067 5033
rect 1976 4856 1983 4893
rect 1996 4887 2003 4933
rect 2096 4868 2103 5032
rect 2156 4883 2163 5073
rect 2136 4876 2163 4883
rect 2136 4856 2143 4876
rect 2096 4587 2103 4854
rect 2196 4827 2203 5233
rect 2216 5088 2223 5253
rect 2336 5247 2343 5333
rect 2356 5267 2363 5393
rect 2376 5227 2383 5373
rect 2396 5307 2403 5393
rect 2416 5387 2423 5556
rect 2496 5447 2503 5563
rect 2253 5108 2267 5113
rect 2293 5088 2307 5093
rect 2336 5047 2343 5173
rect 2396 5076 2403 5272
rect 2436 5207 2443 5343
rect 2487 5336 2503 5343
rect 2433 5080 2447 5093
rect 2436 5076 2443 5080
rect 2216 4987 2223 5033
rect 2236 5007 2243 5043
rect 2276 5040 2283 5043
rect 2273 5027 2287 5040
rect 2356 5043 2363 5074
rect 2356 5036 2383 5043
rect 2353 5007 2367 5013
rect 2180 4823 2193 4827
rect 2116 4787 2123 4823
rect 2176 4816 2193 4823
rect 2180 4813 2193 4816
rect 2216 4787 2223 4973
rect 2316 4907 2323 4933
rect 2296 4856 2303 4893
rect 2116 4667 2123 4773
rect 2276 4767 2283 4823
rect 2356 4767 2363 4993
rect 2376 4807 2383 5036
rect 2476 5007 2483 5293
rect 2496 5046 2503 5336
rect 2516 5267 2523 5453
rect 2536 5307 2543 6033
rect 2556 6027 2563 6073
rect 2596 5987 2603 6083
rect 2636 6080 2643 6083
rect 2633 6067 2647 6080
rect 2576 5827 2583 5863
rect 2616 5807 2623 5863
rect 2676 5807 2683 6333
rect 2716 6207 2723 6383
rect 2756 6116 2763 6173
rect 2736 6080 2743 6083
rect 2733 6067 2747 6080
rect 2736 5896 2743 5993
rect 2796 5907 2803 6513
rect 2856 6416 2863 6473
rect 2896 6416 2903 6473
rect 2876 6347 2883 6383
rect 3016 6207 3023 6383
rect 3056 6327 3063 6383
rect 3056 6187 3063 6313
rect 2876 6116 2883 6153
rect 2816 6047 2823 6114
rect 2916 6086 2923 6153
rect 2996 6143 3003 6173
rect 2996 6136 3023 6143
rect 3016 6128 3023 6136
rect 2936 6116 2983 6123
rect 2856 6047 2863 6083
rect 2936 6007 2943 6116
rect 2933 5900 2947 5913
rect 2936 5896 2943 5900
rect 2716 5707 2723 5863
rect 2756 5767 2763 5863
rect 2556 5567 2563 5633
rect 2596 5527 2603 5563
rect 2636 5527 2643 5563
rect 2627 5476 2653 5483
rect 2656 5343 2663 5413
rect 2696 5388 2703 5653
rect 2756 5596 2763 5732
rect 2796 5687 2803 5852
rect 2836 5847 2843 5894
rect 2996 5866 3003 6051
rect 3036 5947 3043 6083
rect 3056 5967 3063 6033
rect 3076 6007 3083 6133
rect 3056 5908 3063 5953
rect 3096 5928 3103 6513
rect 3196 6428 3203 6473
rect 3116 6416 3163 6423
rect 3116 6307 3123 6416
rect 3216 6380 3223 6383
rect 3173 6367 3187 6372
rect 3213 6367 3227 6380
rect 3116 6267 3123 6293
rect 3156 6116 3163 6153
rect 3173 6147 3187 6153
rect 3116 6086 3123 6113
rect 3216 5987 3223 6083
rect 3256 6027 3263 6413
rect 3276 6347 3283 6453
rect 3296 6427 3303 6563
rect 3316 6380 3323 6383
rect 3356 6380 3363 6383
rect 3313 6367 3327 6380
rect 3353 6367 3367 6380
rect 3276 6087 3283 6253
rect 3316 6116 3323 6173
rect 3356 6116 3363 6233
rect 3416 6086 3423 6153
rect 3216 5976 3233 5987
rect 3220 5973 3233 5976
rect 2956 5860 2963 5863
rect 2953 5847 2967 5860
rect 2827 5596 2843 5603
rect 2716 5447 2723 5573
rect 2776 5527 2783 5563
rect 2676 5376 2693 5383
rect 2676 5346 2683 5376
rect 2736 5376 2743 5413
rect 2636 5336 2663 5343
rect 2636 5207 2643 5336
rect 2756 5307 2763 5343
rect 2636 5046 2643 5193
rect 2656 5107 2663 5233
rect 2676 5167 2683 5213
rect 2407 4863 2420 4867
rect 2407 4856 2423 4863
rect 2456 4856 2463 4913
rect 2407 4853 2420 4856
rect 2356 4647 2363 4713
rect 2376 4707 2383 4793
rect 1516 4467 1523 4523
rect 1536 4376 1543 4493
rect 1636 4407 1643 4554
rect 1796 4527 1803 4556
rect 1973 4560 1987 4573
rect 1976 4556 1983 4560
rect 2316 4556 2323 4613
rect 2353 4567 2367 4573
rect 2376 4568 2383 4653
rect 2396 4623 2403 4813
rect 2436 4667 2443 4823
rect 2396 4616 2423 4623
rect 1616 4303 1623 4333
rect 1676 4306 1683 4393
rect 1776 4336 1783 4433
rect 1596 4296 1623 4303
rect 1756 4187 1763 4303
rect 1476 4036 1503 4043
rect 1136 3587 1143 3813
rect 1176 3687 1183 3783
rect 1216 3780 1223 3783
rect 1213 3767 1227 3780
rect 1256 3767 1263 3833
rect 1336 3816 1343 3873
rect 1376 3847 1383 3953
rect 1376 3816 1383 3833
rect 1276 3786 1283 3813
rect 1416 3786 1423 3913
rect 1256 3607 1263 3753
rect 1087 3513 1093 3527
rect 996 3447 1003 3483
rect 996 3347 1003 3433
rect 1036 3347 1043 3473
rect 1056 3467 1063 3513
rect 1047 3336 1063 3343
rect 1056 3307 1063 3336
rect 1076 3303 1083 3492
rect 1156 3463 1163 3483
rect 1107 3456 1163 3463
rect 1076 3296 1093 3303
rect 1016 3260 1023 3263
rect 1013 3247 1027 3260
rect 1076 3247 1083 3272
rect 1096 3263 1103 3294
rect 1096 3256 1123 3263
rect 1067 3093 1073 3107
rect 1096 3087 1103 3113
rect 776 2746 783 2853
rect 636 2647 643 2743
rect 396 2476 403 2573
rect 436 2476 443 2613
rect 476 2476 483 2513
rect 373 2260 387 2273
rect 376 2256 383 2260
rect 416 2256 423 2293
rect 476 2226 483 2253
rect 396 2220 403 2223
rect 436 2220 443 2223
rect 393 2207 407 2220
rect 433 2207 447 2220
rect 447 2196 463 2203
rect 396 1927 403 2172
rect 116 1767 123 1923
rect 356 1867 363 1923
rect 136 1736 163 1743
rect 156 1627 163 1736
rect 216 1687 223 1753
rect 276 1736 283 1813
rect 416 1807 423 1913
rect 416 1767 423 1793
rect 313 1740 327 1753
rect 436 1747 443 2093
rect 456 1926 463 2196
rect 496 2187 503 2353
rect 576 2307 583 2553
rect 596 2447 603 2613
rect 676 2527 683 2743
rect 736 2740 743 2743
rect 733 2727 747 2740
rect 656 2440 663 2443
rect 596 2283 603 2433
rect 653 2427 667 2440
rect 696 2407 703 2474
rect 736 2367 743 2653
rect 796 2567 803 2952
rect 836 2867 843 3013
rect 896 2996 923 3003
rect 856 2927 863 2963
rect 916 2827 923 2996
rect 1013 3000 1027 3013
rect 1016 2996 1023 3000
rect 936 2803 943 2993
rect 996 2847 1003 2913
rect 1036 2887 1043 2963
rect 916 2796 943 2803
rect 896 2746 903 2774
rect 793 2480 807 2493
rect 796 2476 803 2480
rect 776 2407 783 2443
rect 816 2440 823 2443
rect 813 2427 827 2440
rect 876 2427 883 2473
rect 596 2276 623 2283
rect 616 2256 623 2276
rect 516 1956 523 2193
rect 596 2187 603 2223
rect 576 2147 583 2173
rect 316 1736 323 1740
rect 256 1700 263 1703
rect 253 1687 267 1700
rect 136 1436 163 1443
rect 16 1406 23 1433
rect 156 1367 163 1436
rect 136 1047 143 1183
rect 176 1047 183 1493
rect 196 1087 203 1213
rect 216 1186 223 1453
rect 296 1447 303 1703
rect 416 1700 423 1703
rect 413 1687 427 1700
rect 456 1687 463 1813
rect 376 1436 383 1493
rect 256 1400 263 1403
rect 253 1387 267 1400
rect 296 1147 303 1183
rect 136 916 143 973
rect 176 916 183 1033
rect 336 1007 343 1213
rect 316 927 323 973
rect 116 708 123 883
rect 156 880 163 883
rect 153 867 167 880
rect 236 847 243 913
rect 336 886 343 953
rect 356 927 363 1373
rect 396 1367 403 1403
rect 396 1247 403 1353
rect 387 1223 400 1227
rect 387 1216 403 1223
rect 436 1216 443 1403
rect 476 1307 483 1913
rect 536 1867 543 1923
rect 496 1387 503 1434
rect 387 1213 400 1216
rect 496 1186 503 1313
rect 416 967 423 1172
rect 516 1167 523 1553
rect 536 1467 543 1493
rect 556 1448 563 1693
rect 576 1687 583 2133
rect 656 2107 663 2223
rect 596 1436 603 2033
rect 636 1923 643 1993
rect 696 1956 723 1963
rect 716 1926 723 1956
rect 756 1927 763 2273
rect 776 2027 783 2313
rect 813 1960 827 1973
rect 816 1956 823 1960
rect 636 1916 663 1923
rect 616 1567 623 1853
rect 636 1847 643 1916
rect 796 1807 803 1923
rect 836 1887 843 1912
rect 656 1736 663 1793
rect 813 1763 827 1773
rect 796 1760 827 1763
rect 836 1763 843 1873
rect 796 1756 823 1760
rect 836 1756 863 1763
rect 796 1743 803 1756
rect 776 1736 803 1743
rect 656 1447 663 1673
rect 676 1587 683 1703
rect 756 1627 763 1734
rect 776 1706 783 1736
rect 856 1736 863 1756
rect 896 1747 903 2732
rect 916 2707 923 2796
rect 916 2487 923 2693
rect 936 2647 943 2773
rect 1036 2740 1043 2743
rect 1033 2727 1047 2740
rect 947 2503 960 2507
rect 947 2493 963 2503
rect 956 2476 963 2493
rect 1016 2446 1023 2473
rect 976 2407 983 2443
rect 916 1987 923 2393
rect 1016 2227 1023 2254
rect 976 2187 983 2223
rect 976 2127 983 2173
rect 1036 2007 1043 2533
rect 1076 2488 1083 2733
rect 1096 2567 1103 3073
rect 1116 2867 1123 3256
rect 1156 3227 1163 3252
rect 1196 3123 1203 3473
rect 1216 3266 1223 3333
rect 1276 3296 1283 3353
rect 1296 3327 1303 3473
rect 1316 3367 1323 3573
rect 1436 3483 1443 3833
rect 1476 3816 1483 3893
rect 1496 3847 1503 4036
rect 1736 4036 1743 4113
rect 1636 4006 1643 4033
rect 1636 3927 1643 3992
rect 1656 3967 1663 4034
rect 1396 3476 1443 3483
rect 1336 3347 1343 3453
rect 1393 3300 1407 3313
rect 1456 3303 1463 3533
rect 1396 3296 1403 3300
rect 1436 3296 1463 3303
rect 1376 3243 1383 3263
rect 1376 3236 1403 3243
rect 1196 3116 1213 3123
rect 1133 3087 1147 3093
rect 1156 3027 1163 3053
rect 1153 3000 1167 3013
rect 1156 2996 1163 3000
rect 1216 2996 1223 3113
rect 1396 3027 1403 3236
rect 1416 3007 1423 3263
rect 1476 3207 1483 3353
rect 1456 3127 1463 3173
rect 1496 3147 1503 3593
rect 1536 3547 1543 3853
rect 1656 3843 1663 3932
rect 1816 3867 1823 4353
rect 1836 4307 1843 4393
rect 1893 4340 1907 4353
rect 1896 4336 1903 4340
rect 1936 4336 1943 4553
rect 2036 4447 2043 4523
rect 2156 4520 2163 4523
rect 2153 4507 2167 4520
rect 2256 4467 2263 4513
rect 2196 4327 2203 4353
rect 2216 4306 2223 4334
rect 2156 4267 2163 4303
rect 1836 4006 1843 4213
rect 1936 4036 1943 4073
rect 1636 3836 1663 3843
rect 1636 3816 1643 3836
rect 1556 3516 1563 3673
rect 1593 3520 1607 3533
rect 1616 3528 1623 3772
rect 1696 3767 1703 3814
rect 1716 3786 1723 3813
rect 1856 3786 1863 3853
rect 1776 3780 1783 3783
rect 1773 3767 1787 3780
rect 1736 3587 1743 3633
rect 1876 3543 1883 3813
rect 1896 3767 1903 4003
rect 1976 3927 1983 4003
rect 2036 3907 2043 4253
rect 2156 4036 2163 4253
rect 2056 3947 2063 4033
rect 2216 3927 2223 4292
rect 1996 3827 2003 3893
rect 1936 3767 1943 3783
rect 1936 3647 1943 3753
rect 1976 3747 1983 3783
rect 2136 3747 2143 3913
rect 2236 3707 2243 4433
rect 2296 4367 2303 4523
rect 2336 4487 2343 4523
rect 2376 4487 2383 4554
rect 2396 4526 2403 4593
rect 2416 4563 2423 4616
rect 2516 4607 2523 4893
rect 2536 4887 2543 5032
rect 2556 4967 2563 5013
rect 2576 4907 2583 5043
rect 2616 5036 2633 5043
rect 2616 4927 2623 5036
rect 2593 4860 2607 4873
rect 2596 4856 2603 4860
rect 2636 4856 2643 4953
rect 2656 4867 2663 5093
rect 2756 5007 2763 5193
rect 2816 5107 2823 5373
rect 2836 5167 2843 5596
rect 2856 5247 2863 5793
rect 2876 5608 2883 5831
rect 2953 5827 2967 5833
rect 2956 5596 2963 5673
rect 2876 5407 2883 5594
rect 2936 5487 2943 5552
rect 2996 5507 3003 5852
rect 3016 5727 3023 5833
rect 3076 5827 3083 5863
rect 3156 5827 3163 5913
rect 2976 5347 2983 5433
rect 2896 5307 2903 5343
rect 2416 4556 2443 4563
rect 2473 4560 2487 4573
rect 2476 4556 2483 4560
rect 2316 4336 2323 4453
rect 2416 4427 2423 4513
rect 2496 4520 2503 4523
rect 2493 4507 2507 4520
rect 2556 4507 2563 4853
rect 2676 4847 2683 4993
rect 2576 4507 2583 4553
rect 2576 4447 2583 4493
rect 2636 4427 2643 4523
rect 2476 4306 2483 4413
rect 2556 4336 2563 4413
rect 2676 4367 2683 4812
rect 2716 4647 2723 4993
rect 2776 4927 2783 5093
rect 2796 5076 2823 5083
rect 2796 4967 2803 5076
rect 2896 5007 2903 5173
rect 2916 4987 2923 5074
rect 2956 5046 2963 5343
rect 3016 5147 3023 5713
rect 3076 5596 3083 5813
rect 3176 5807 3183 5913
rect 3196 5907 3203 5933
rect 3216 5866 3223 5953
rect 3253 5947 3267 5953
rect 3313 5900 3327 5913
rect 3316 5896 3323 5900
rect 3356 5860 3363 5863
rect 3353 5847 3367 5860
rect 3136 5608 3143 5773
rect 3156 5563 3163 5673
rect 3193 5608 3207 5613
rect 3236 5596 3243 5653
rect 3276 5566 3283 5593
rect 3316 5566 3323 5613
rect 3336 5596 3343 5653
rect 3376 5627 3383 5713
rect 3396 5707 3403 5833
rect 3396 5596 3403 5693
rect 3156 5556 3183 5563
rect 3076 5376 3083 5493
rect 3056 5247 3063 5343
rect 3096 5207 3103 5343
rect 3156 5223 3163 5374
rect 3176 5287 3183 5556
rect 3216 5507 3223 5563
rect 3236 5376 3243 5413
rect 3336 5388 3343 5413
rect 3136 5216 3163 5223
rect 2967 5036 2983 5043
rect 2836 4826 2843 4913
rect 3016 4903 3023 5003
rect 2996 4896 3023 4903
rect 2876 4856 2883 4893
rect 2756 4820 2763 4823
rect 2753 4807 2767 4820
rect 2976 4727 2983 4854
rect 2996 4667 3003 4896
rect 2756 4556 2763 4653
rect 2896 4556 2923 4563
rect 2976 4556 3003 4563
rect 2736 4487 2743 4523
rect 2696 4347 2703 4453
rect 2336 4207 2343 4303
rect 2376 4267 2383 4303
rect 2616 4267 2623 4303
rect 2293 4040 2307 4053
rect 2296 4036 2303 4040
rect 2276 3867 2283 3992
rect 2327 3853 2333 3867
rect 2256 3786 2263 3853
rect 2236 3667 2243 3693
rect 1876 3536 1903 3543
rect 1596 3516 1603 3520
rect 1636 3487 1643 3533
rect 1736 3516 1783 3523
rect 1536 3447 1543 3483
rect 1576 3403 1583 3483
rect 1776 3447 1783 3516
rect 1896 3516 1903 3536
rect 1936 3486 1943 3633
rect 2256 3516 2263 3673
rect 1556 3396 1583 3403
rect 1536 3296 1543 3353
rect 1556 3327 1563 3396
rect 1576 3296 1583 3373
rect 1736 3263 1743 3433
rect 1816 3347 1823 3373
rect 1816 3296 1823 3333
rect 1876 3327 1883 3483
rect 2016 3407 2023 3483
rect 2056 3296 2063 3393
rect 1636 3187 1643 3263
rect 1696 3256 1743 3263
rect 1176 2907 1183 2963
rect 1116 2727 1123 2853
rect 1196 2847 1203 2953
rect 1296 2907 1303 2933
rect 1176 2776 1183 2833
rect 1296 2746 1303 2893
rect 1316 2887 1323 2994
rect 1456 2996 1463 3113
rect 1513 3000 1527 3013
rect 1516 2996 1523 3000
rect 1396 2956 1423 2963
rect 1373 2943 1387 2953
rect 1373 2940 1403 2943
rect 1376 2936 1403 2940
rect 1396 2887 1403 2936
rect 1356 2776 1363 2873
rect 1336 2587 1343 2743
rect 1376 2667 1383 2732
rect 1416 2647 1423 2956
rect 1556 2883 1563 2973
rect 1576 2907 1583 3013
rect 1636 2960 1643 2963
rect 1633 2947 1647 2960
rect 1676 2887 1683 3053
rect 1696 2887 1703 3093
rect 1716 2966 1723 3133
rect 1756 3127 1763 3252
rect 1876 3187 1883 3263
rect 1796 2907 1803 2963
rect 1856 2947 1863 2993
rect 1876 2927 1883 3173
rect 1956 2996 1963 3133
rect 1996 2966 2003 3193
rect 2096 3087 2103 3514
rect 2176 3447 2183 3514
rect 2116 3023 2123 3293
rect 2136 3266 2143 3393
rect 2176 3296 2183 3433
rect 2256 3307 2263 3413
rect 2276 3347 2283 3813
rect 2396 3627 2403 4173
rect 2496 4123 2503 4253
rect 2496 4116 2523 4123
rect 2516 4036 2523 4116
rect 2556 4007 2563 4034
rect 2436 3816 2443 3873
rect 2476 3816 2483 3853
rect 2516 3827 2523 3913
rect 2616 3827 2623 4253
rect 2673 4040 2687 4053
rect 2676 4036 2683 4040
rect 2716 4036 2723 4413
rect 2736 4207 2743 4473
rect 2776 4467 2783 4523
rect 2636 3786 2643 3893
rect 2656 3767 2663 4003
rect 2756 3828 2763 4033
rect 2776 3887 2783 4093
rect 2836 4036 2843 4433
rect 2856 4247 2863 4373
rect 2876 4367 2883 4554
rect 2896 4347 2903 4556
rect 2996 4487 3003 4556
rect 2936 4336 2943 4413
rect 2976 4336 2983 4393
rect 2876 4267 2883 4313
rect 2916 4147 2923 4303
rect 3016 4227 3023 4873
rect 3076 4856 3083 4973
rect 3096 4887 3103 5133
rect 3136 5047 3143 5216
rect 3096 4727 3103 4823
rect 3156 4807 3163 5093
rect 3176 4747 3183 5273
rect 3216 5187 3223 5343
rect 3196 5076 3203 5173
rect 3256 5127 3263 5153
rect 3256 5076 3263 5113
rect 3296 5107 3303 5332
rect 3236 4856 3243 4893
rect 3196 4807 3203 4823
rect 3036 4526 3043 4633
rect 3093 4560 3107 4573
rect 3096 4556 3103 4560
rect 3116 4487 3123 4523
rect 3093 4340 3107 4353
rect 3096 4336 3103 4340
rect 3076 4267 3083 4303
rect 3116 4263 3123 4303
rect 3156 4287 3163 4493
rect 3176 4407 3183 4573
rect 3116 4256 3143 4263
rect 2916 4107 2923 4133
rect 3036 4067 3043 4193
rect 3076 4187 3083 4253
rect 2873 4040 2887 4053
rect 2876 4036 2883 4040
rect 2916 4007 2923 4053
rect 3033 4040 3047 4053
rect 3036 4036 3043 4040
rect 2816 3967 2823 4003
rect 2436 3516 2443 3593
rect 2416 3427 2423 3483
rect 2356 3307 2363 3373
rect 2276 3187 2283 3263
rect 2396 3247 2403 3333
rect 2456 3296 2463 3333
rect 2096 3016 2123 3023
rect 2096 2996 2103 3016
rect 2136 2996 2143 3033
rect 2233 3008 2247 3013
rect 2276 2996 2283 3113
rect 1556 2876 1583 2883
rect 1436 2746 1443 2853
rect 1496 2776 1503 2833
rect 1536 2776 1543 2813
rect 1476 2647 1483 2743
rect 1576 2743 1583 2876
rect 1596 2746 1603 2873
rect 1556 2736 1583 2743
rect 1096 2476 1103 2553
rect 1276 2488 1283 2513
rect 1176 2367 1183 2473
rect 1093 2260 1107 2273
rect 1096 2256 1103 2260
rect 1176 2226 1183 2353
rect 1256 2256 1263 2293
rect 1336 2226 1343 2293
rect 1396 2256 1403 2474
rect 1436 2256 1443 2353
rect 1456 2343 1463 2443
rect 1456 2336 1483 2343
rect 1076 2207 1083 2223
rect 993 1960 1007 1973
rect 996 1956 1003 1960
rect 976 1887 983 1923
rect 833 1687 847 1692
rect 756 1436 763 1553
rect 576 1327 583 1403
rect 616 1307 623 1403
rect 573 1220 587 1233
rect 576 1216 583 1220
rect 556 1147 563 1183
rect 596 1180 603 1183
rect 593 1167 607 1180
rect 456 916 463 1033
rect 176 527 183 693
rect 136 396 143 513
rect 196 403 203 713
rect 253 708 267 713
rect 296 696 303 813
rect 236 607 243 652
rect 276 627 283 663
rect 336 427 343 872
rect 356 666 363 833
rect 396 723 403 883
rect 436 880 443 883
rect 433 867 447 880
rect 496 747 503 1073
rect 576 916 583 993
rect 636 967 643 1173
rect 656 1147 663 1433
rect 736 1400 743 1403
rect 733 1387 747 1400
rect 776 1327 783 1403
rect 556 827 563 883
rect 596 787 603 883
rect 396 716 423 723
rect 416 708 423 716
rect 356 627 363 652
rect 436 607 443 663
rect 300 423 313 427
rect 296 413 313 423
rect 176 396 223 403
rect 296 396 303 413
rect 216 366 223 396
rect 336 387 343 413
rect 356 366 363 513
rect 413 400 427 413
rect 453 400 467 413
rect 416 396 423 400
rect 456 396 463 400
rect 116 176 123 313
rect 156 267 163 363
rect 496 327 503 733
rect 536 707 543 753
rect 596 696 603 752
rect 576 627 583 663
rect 616 660 623 663
rect 613 647 627 660
rect 576 467 583 613
rect 516 367 523 453
rect 636 427 643 653
rect 656 507 663 773
rect 676 647 683 1273
rect 776 1228 783 1313
rect 756 1216 773 1223
rect 736 1127 743 1183
rect 716 827 723 883
rect 796 867 803 1253
rect 736 696 743 753
rect 816 723 823 1673
rect 836 1387 843 1453
rect 896 1436 903 1673
rect 916 1467 923 1873
rect 1016 1787 1023 1923
rect 1056 1867 1063 2013
rect 996 1736 1003 1773
rect 1016 1700 1023 1703
rect 936 1607 943 1692
rect 1013 1687 1027 1700
rect 936 1436 943 1593
rect 1056 1587 1063 1813
rect 1076 1706 1083 2193
rect 1236 2087 1243 2223
rect 1416 2167 1423 2223
rect 1476 2207 1483 2336
rect 1516 2223 1523 2474
rect 1556 2447 1563 2736
rect 1616 2707 1623 2774
rect 1716 2707 1723 2743
rect 1756 2727 1763 2773
rect 1776 2746 1783 2853
rect 1816 2776 1823 2813
rect 1833 2703 1847 2711
rect 1916 2707 1923 2773
rect 1936 2727 1943 2913
rect 2116 2887 2123 2963
rect 1996 2776 2003 2853
rect 2036 2776 2043 2813
rect 1956 2746 1963 2773
rect 1987 2713 1993 2727
rect 1833 2700 1873 2703
rect 1836 2696 1873 2700
rect 1960 2706 1980 2707
rect 1967 2693 1973 2706
rect 2016 2667 2023 2743
rect 2076 2727 2083 2743
rect 2136 2736 2163 2743
rect 1776 2476 1783 2553
rect 1716 2256 1723 2474
rect 1516 2216 1543 2223
rect 1176 1956 1183 2013
rect 1236 1968 1243 2073
rect 1320 2003 1333 2007
rect 1316 1993 1333 2003
rect 1316 1956 1323 1993
rect 1076 1527 1083 1692
rect 1096 1448 1103 1953
rect 1356 1923 1363 1973
rect 1413 1960 1427 1973
rect 1416 1956 1423 1960
rect 1456 1956 1463 1993
rect 1156 1887 1163 1923
rect 1156 1736 1163 1852
rect 1296 1807 1303 1923
rect 1336 1916 1363 1923
rect 1276 1748 1283 1773
rect 1336 1747 1343 1916
rect 1476 1920 1483 1923
rect 1473 1907 1487 1920
rect 1116 1700 1123 1703
rect 1113 1687 1127 1700
rect 876 1287 883 1403
rect 916 1267 923 1403
rect 876 1167 883 1183
rect 876 1007 883 1153
rect 876 916 883 993
rect 916 907 923 953
rect 956 928 963 1313
rect 976 1186 983 1433
rect 996 1227 1003 1253
rect 1076 1227 1083 1253
rect 1016 1127 1023 1183
rect 976 916 983 953
rect 1013 928 1027 933
rect 996 827 1003 883
rect 1076 867 1083 933
rect 1096 928 1103 1393
rect 1116 1267 1123 1673
rect 1176 1448 1183 1633
rect 1216 1448 1223 1493
rect 1336 1436 1343 1733
rect 1356 1463 1363 1793
rect 1396 1736 1403 1793
rect 1436 1736 1443 1853
rect 1496 1707 1503 1912
rect 1516 1767 1523 2216
rect 1636 2187 1643 2253
rect 1687 2216 1703 2223
rect 1556 1956 1603 1963
rect 1536 1867 1543 1954
rect 1556 1907 1563 1956
rect 1676 1927 1683 2212
rect 1736 2187 1743 2223
rect 1796 2027 1803 2653
rect 2076 2527 2083 2713
rect 2156 2707 2163 2736
rect 2176 2667 2183 2994
rect 2196 2827 2203 2973
rect 2256 2907 2263 2963
rect 2296 2807 2303 2963
rect 2376 2947 2383 3093
rect 2496 3087 2503 3613
rect 2456 2996 2463 3033
rect 2493 3000 2507 3013
rect 2516 3003 2523 3693
rect 2756 3647 2763 3753
rect 2536 3027 2543 3353
rect 2576 3327 2583 3483
rect 2636 3447 2643 3493
rect 2596 3296 2603 3353
rect 2636 3296 2643 3433
rect 2656 3427 2663 3513
rect 2716 3476 2743 3483
rect 2716 3263 2723 3453
rect 2736 3367 2743 3476
rect 2756 3467 2763 3633
rect 2776 3567 2783 3873
rect 2776 3487 2783 3553
rect 2796 3527 2803 3813
rect 2816 3667 2823 3953
rect 2856 3907 2863 4003
rect 2856 3567 2863 3783
rect 2896 3727 2903 3783
rect 2896 3567 2903 3593
rect 2916 3547 2923 3773
rect 2996 3727 3003 3814
rect 3016 3786 3023 3893
rect 3116 3847 3123 4213
rect 3136 4207 3143 4256
rect 3196 4187 3203 4793
rect 3256 4787 3263 4823
rect 3276 4607 3283 5073
rect 3296 4787 3303 4973
rect 3316 4826 3323 5133
rect 3336 5107 3343 5374
rect 3376 5343 3383 5513
rect 3416 5388 3423 6013
rect 3436 5787 3443 6473
rect 3516 6416 3523 6473
rect 3696 6428 3703 6493
rect 3576 6386 3583 6413
rect 3536 6347 3543 6383
rect 3616 6267 3623 6414
rect 3647 6423 3660 6427
rect 3647 6416 3663 6423
rect 3647 6413 3660 6416
rect 3756 6386 3763 6433
rect 3776 6383 3783 6414
rect 3916 6386 3923 6433
rect 3976 6416 3983 6493
rect 4907 6476 4933 6483
rect 4156 6416 4163 6473
rect 4876 6460 4913 6463
rect 4873 6456 4913 6460
rect 4436 6416 4443 6453
rect 4873 6447 4887 6456
rect 4473 6420 4487 6433
rect 4740 6443 4753 6447
rect 4476 6416 4483 6420
rect 4613 6420 4627 6433
rect 4736 6433 4753 6443
rect 4616 6416 4623 6420
rect 4736 6416 4743 6433
rect 3776 6380 3803 6383
rect 3773 6376 3803 6380
rect 3773 6367 3787 6376
rect 3496 6116 3503 6153
rect 3556 6087 3563 6193
rect 3576 6083 3583 6213
rect 3636 6116 3643 6153
rect 3676 6116 3683 6153
rect 3576 6076 3623 6083
rect 3516 6063 3523 6072
rect 3496 6056 3523 6063
rect 3496 5896 3503 6056
rect 3596 5987 3603 6013
rect 3656 6007 3663 6083
rect 3696 6047 3703 6073
rect 3476 5860 3483 5863
rect 3473 5847 3487 5860
rect 3516 5856 3543 5863
rect 3436 5567 3443 5713
rect 3496 5608 3503 5633
rect 3536 5608 3543 5856
rect 3556 5827 3563 5953
rect 3596 5847 3603 5973
rect 3656 5896 3663 5953
rect 3696 5896 3703 6033
rect 3636 5860 3643 5863
rect 3633 5847 3647 5860
rect 3456 5507 3463 5594
rect 3576 5467 3583 5653
rect 3376 5336 3403 5343
rect 3356 5088 3363 5293
rect 3476 5247 3483 5373
rect 3496 5267 3503 5413
rect 3396 5076 3403 5133
rect 3336 5007 3343 5032
rect 3376 4856 3383 5043
rect 3436 4947 3443 5173
rect 3493 5147 3507 5153
rect 3516 5147 3523 5393
rect 3536 5387 3543 5453
rect 3556 5376 3563 5413
rect 3596 5376 3603 5594
rect 3616 5407 3623 5773
rect 3736 5667 3743 6273
rect 3756 6227 3763 6253
rect 3796 6187 3803 6376
rect 3956 6380 3963 6383
rect 3816 6367 3823 6372
rect 3953 6367 3967 6380
rect 3816 6356 3833 6367
rect 3820 6353 3833 6356
rect 4056 6287 4063 6413
rect 4516 6386 4523 6413
rect 4796 6386 4803 6433
rect 4893 6420 4907 6433
rect 4896 6416 4903 6420
rect 5093 6420 5107 6433
rect 5096 6416 5103 6420
rect 5216 6416 5223 6473
rect 5247 6436 5273 6443
rect 4836 6387 4843 6414
rect 5393 6420 5407 6433
rect 5396 6416 5403 6420
rect 4176 6307 4183 6383
rect 3756 6107 3763 6173
rect 3787 6123 3800 6127
rect 3787 6116 3803 6123
rect 3787 6113 3800 6116
rect 3876 6087 3883 6114
rect 3976 6047 3983 6083
rect 3816 5896 3823 5953
rect 3873 5947 3887 5953
rect 3896 5866 3903 5933
rect 3676 5596 3683 5633
rect 3696 5467 3703 5563
rect 3756 5483 3763 5852
rect 3796 5667 3803 5793
rect 3776 5507 3783 5594
rect 3796 5567 3803 5632
rect 3876 5596 3883 5693
rect 3916 5647 3923 5993
rect 3933 5947 3947 5953
rect 3996 5896 4003 6053
rect 4036 5987 4043 6114
rect 4056 6007 4063 6233
rect 4076 6086 4083 6133
rect 4096 6116 4103 6153
rect 4156 6116 4173 6123
rect 4176 6067 4183 6114
rect 4196 6047 4203 6353
rect 4276 6247 4283 6383
rect 4316 6207 4323 6372
rect 4596 6267 4603 6383
rect 5296 6386 5303 6413
rect 5076 6380 5083 6383
rect 4276 6128 4283 6153
rect 4496 6116 4503 6193
rect 4596 6187 4603 6253
rect 4656 6127 4663 6333
rect 4016 5860 4023 5863
rect 4013 5847 4027 5860
rect 4056 5827 4063 5894
rect 4076 5866 4083 6013
rect 4156 5860 4163 5863
rect 4153 5847 4167 5860
rect 4236 5827 4243 5933
rect 4276 5896 4283 6053
rect 4336 6007 4343 6083
rect 4376 6027 4383 6114
rect 4676 6086 4683 6173
rect 4793 6120 4807 6133
rect 4796 6116 4803 6120
rect 4436 6047 4443 6083
rect 4476 6047 4483 6083
rect 3936 5567 3943 5793
rect 4036 5596 4043 5713
rect 4156 5627 4163 5713
rect 4196 5667 4203 5693
rect 4153 5600 4167 5613
rect 4156 5596 4163 5600
rect 4196 5596 4203 5653
rect 3956 5567 3963 5594
rect 3900 5563 3913 5567
rect 3756 5476 3783 5483
rect 3676 5456 3693 5463
rect 3656 5347 3663 5413
rect 3676 5347 3683 5456
rect 3696 5387 3703 5413
rect 3620 5343 3633 5347
rect 3536 5167 3543 5333
rect 3576 5287 3583 5343
rect 3616 5336 3633 5343
rect 3620 5333 3633 5336
rect 3776 5267 3783 5476
rect 3856 5467 3863 5563
rect 3896 5556 3913 5563
rect 3900 5553 3913 5556
rect 3876 5376 3883 5493
rect 4013 5380 4027 5393
rect 4016 5376 4023 5380
rect 3816 5346 3823 5373
rect 4056 5343 4063 5393
rect 4047 5336 4063 5343
rect 3516 5103 3523 5133
rect 3496 5096 3523 5103
rect 3496 5076 3503 5096
rect 3536 5076 3543 5153
rect 3436 4803 3443 4823
rect 3416 4796 3443 4803
rect 3236 4556 3243 4593
rect 3256 4487 3263 4523
rect 3296 4520 3303 4523
rect 3293 4507 3307 4520
rect 3336 4467 3343 4533
rect 3356 4526 3363 4633
rect 3416 4568 3423 4796
rect 3436 4587 3443 4713
rect 3456 4707 3463 4813
rect 3476 4607 3483 4873
rect 3516 4863 3523 5043
rect 3576 5027 3583 5113
rect 3676 5076 3683 5113
rect 3596 4987 3603 5074
rect 3716 5047 3723 5074
rect 3736 5047 3743 5253
rect 3816 5227 3823 5332
rect 3993 5327 4007 5332
rect 4036 5287 4043 5332
rect 3776 5088 3783 5173
rect 3496 4856 3523 4863
rect 3533 4860 3547 4873
rect 3536 4856 3543 4860
rect 3496 4647 3503 4856
rect 3616 4867 3623 4893
rect 3516 4747 3523 4812
rect 3476 4527 3483 4572
rect 3436 4507 3443 4523
rect 3496 4507 3503 4553
rect 3296 4336 3303 4433
rect 3436 4427 3443 4493
rect 3416 4416 3433 4423
rect 3236 4187 3243 4303
rect 3156 4036 3163 4173
rect 3196 4036 3203 4133
rect 3176 3927 3183 4003
rect 3256 3827 3263 3913
rect 3116 3687 3123 3772
rect 2873 3520 2887 3533
rect 3096 3528 3103 3673
rect 2876 3516 2883 3520
rect 2776 3296 2783 3333
rect 2796 3323 2803 3473
rect 2816 3387 2823 3472
rect 2836 3427 2843 3453
rect 2796 3316 2823 3323
rect 2616 3260 2623 3263
rect 2613 3247 2627 3260
rect 2716 3256 2743 3263
rect 2496 2996 2503 3000
rect 2516 2996 2543 3003
rect 2436 2927 2443 2963
rect 2476 2943 2483 2963
rect 2476 2936 2503 2943
rect 2496 2847 2503 2936
rect 2536 2867 2543 2996
rect 2556 2966 2563 3193
rect 2796 3043 2803 3293
rect 2816 3266 2823 3316
rect 2876 3296 2883 3433
rect 2916 3367 2923 3483
rect 2976 3266 2983 3313
rect 2996 3263 3003 3433
rect 3136 3347 3143 3513
rect 3053 3300 3067 3313
rect 3096 3308 3103 3333
rect 3056 3296 3063 3300
rect 3107 3296 3123 3303
rect 2996 3256 3043 3263
rect 3076 3167 3083 3263
rect 3116 3123 3123 3296
rect 3156 3263 3163 3653
rect 3276 3647 3283 4271
rect 3336 4167 3343 4334
rect 3356 4303 3363 4373
rect 3416 4336 3423 4416
rect 3356 4296 3373 4303
rect 3376 4247 3383 4292
rect 3313 4040 3327 4053
rect 3316 4036 3323 4040
rect 3356 3847 3363 3992
rect 3376 3867 3383 4133
rect 3476 4127 3483 4303
rect 3516 4243 3523 4733
rect 3556 4727 3563 4823
rect 3596 4820 3603 4823
rect 3593 4807 3607 4820
rect 3636 4807 3643 5013
rect 3836 4987 3843 5043
rect 3876 5027 3883 5093
rect 3536 4567 3543 4593
rect 3576 4556 3583 4613
rect 3613 4560 3627 4573
rect 3616 4556 3623 4560
rect 3547 4523 3560 4527
rect 3547 4516 3563 4523
rect 3596 4520 3603 4523
rect 3547 4513 3560 4516
rect 3593 4507 3607 4520
rect 3496 4236 3523 4243
rect 3496 4067 3503 4236
rect 3516 4087 3523 4193
rect 3296 3587 3303 3833
rect 3376 3823 3383 3853
rect 3356 3816 3383 3823
rect 3356 3627 3363 3753
rect 3396 3587 3403 4053
rect 3516 4036 3523 4073
rect 3536 4006 3543 4333
rect 3556 4306 3563 4453
rect 3616 4336 3623 4413
rect 3567 4296 3583 4303
rect 3556 4167 3563 4253
rect 3236 3516 3243 3553
rect 3216 3463 3223 3472
rect 3216 3456 3243 3463
rect 3216 3296 3223 3433
rect 3156 3256 3183 3263
rect 3096 3116 3123 3123
rect 2776 3036 2803 3043
rect 2613 3000 2627 3013
rect 2616 2996 2623 3000
rect 2776 2996 2783 3036
rect 2813 3000 2827 3013
rect 2816 2996 2823 3000
rect 2636 2960 2643 2963
rect 2633 2947 2647 2960
rect 2493 2780 2507 2793
rect 2496 2776 2503 2780
rect 1907 2476 1923 2483
rect 1916 2307 1923 2476
rect 1796 1983 1803 2013
rect 1776 1976 1803 1983
rect 1776 1956 1783 1976
rect 1836 1956 1843 2173
rect 1856 2127 1863 2223
rect 1896 2087 1903 2223
rect 1956 2167 1963 2254
rect 1976 2187 1983 2293
rect 2096 2226 2103 2253
rect 2016 2220 2023 2223
rect 2013 2207 2027 2220
rect 1896 2047 1903 2073
rect 1696 1887 1703 1954
rect 1673 1740 1687 1753
rect 1676 1736 1683 1740
rect 1456 1687 1463 1703
rect 1616 1687 1623 1734
rect 1756 1706 1763 1853
rect 1796 1827 1803 1923
rect 1936 1867 1943 2093
rect 1956 1987 1963 2153
rect 1356 1456 1383 1463
rect 1376 1436 1383 1456
rect 1456 1407 1463 1673
rect 1536 1436 1543 1513
rect 1576 1447 1583 1533
rect 1696 1467 1703 1703
rect 1633 1440 1647 1453
rect 1636 1436 1643 1440
rect 1356 1287 1363 1403
rect 1127 1214 1133 1227
rect 1156 1216 1163 1273
rect 1127 1213 1140 1214
rect 1156 916 1163 993
rect 1236 947 1243 1193
rect 1256 928 1263 1273
rect 1360 1223 1373 1227
rect 1356 1216 1373 1223
rect 1360 1213 1373 1216
rect 1516 1216 1523 1313
rect 1576 1287 1583 1433
rect 1596 1247 1603 1392
rect 1696 1367 1703 1403
rect 1736 1367 1743 1553
rect 1707 1356 1723 1363
rect 1696 1287 1703 1313
rect 1336 1180 1343 1183
rect 1333 1167 1347 1180
rect 1396 1167 1403 1213
rect 1416 1107 1423 1213
rect 1456 1127 1463 1183
rect 1296 947 1303 973
rect 1487 934 1493 947
rect 1480 933 1493 934
rect 1293 920 1307 933
rect 1296 916 1303 920
rect 1096 886 1103 914
rect 1436 887 1443 933
rect 1516 916 1523 973
rect 1596 887 1603 1233
rect 1676 1223 1683 1273
rect 1656 1216 1683 1223
rect 1656 916 1663 1093
rect 1673 947 1687 953
rect 1696 916 1703 953
rect 1716 923 1723 1356
rect 1756 1347 1763 1633
rect 1796 1567 1803 1703
rect 1876 1627 1883 1833
rect 1956 1807 1963 1973
rect 2016 1847 2023 1923
rect 1896 1683 1903 1734
rect 1916 1703 1923 1793
rect 2056 1767 2063 2173
rect 2136 2167 2143 2353
rect 2196 2347 2203 2774
rect 2316 2740 2323 2743
rect 2313 2727 2327 2740
rect 2376 2723 2383 2743
rect 2376 2716 2403 2723
rect 2276 2647 2283 2673
rect 2396 2487 2403 2716
rect 2236 2387 2243 2473
rect 2296 2440 2303 2443
rect 2293 2427 2307 2440
rect 2333 2427 2347 2433
rect 2176 2256 2183 2293
rect 2356 2267 2363 2474
rect 2376 2447 2383 2474
rect 2413 2480 2427 2493
rect 2416 2476 2423 2480
rect 2456 2476 2463 2573
rect 2436 2440 2443 2443
rect 2393 2427 2407 2433
rect 2433 2427 2447 2440
rect 2236 2167 2243 2223
rect 2276 2187 2283 2223
rect 2200 1963 2213 1967
rect 2196 1956 2213 1963
rect 2096 1923 2103 1954
rect 2200 1953 2213 1956
rect 2236 1947 2243 2053
rect 2296 1956 2303 2053
rect 2316 1987 2323 2093
rect 2356 1963 2363 2213
rect 2376 1987 2383 2333
rect 2476 2303 2483 2432
rect 2476 2296 2503 2303
rect 2396 2067 2403 2293
rect 2496 2167 2503 2296
rect 2516 2287 2523 2533
rect 2536 2307 2543 2713
rect 2576 2488 2583 2893
rect 2633 2780 2647 2793
rect 2636 2776 2643 2780
rect 2616 2587 2623 2743
rect 2596 2440 2603 2443
rect 2593 2427 2607 2440
rect 2656 2427 2663 2474
rect 2596 2256 2603 2353
rect 2616 2287 2623 2313
rect 2616 2220 2623 2223
rect 2576 2187 2583 2212
rect 2613 2207 2627 2220
rect 2456 2087 2463 2133
rect 2496 2127 2503 2153
rect 2347 1956 2363 1963
rect 2096 1916 2123 1923
rect 2116 1807 2123 1916
rect 2176 1887 2183 1923
rect 2236 1867 2243 1933
rect 2256 1927 2263 1953
rect 2436 1887 2443 1954
rect 1916 1696 1943 1703
rect 1896 1676 1923 1683
rect 1876 1587 1883 1613
rect 1776 1216 1783 1473
rect 1833 1440 1847 1453
rect 1836 1436 1843 1440
rect 1916 1407 1923 1676
rect 1936 1507 1943 1696
rect 2016 1667 2023 1703
rect 2056 1700 2063 1703
rect 2053 1687 2067 1700
rect 1756 1107 1763 1183
rect 1716 916 1743 923
rect 1136 880 1143 883
rect 1133 867 1147 880
rect 1496 880 1503 883
rect 1536 880 1543 883
rect 1313 867 1327 872
rect 1493 867 1507 880
rect 1533 867 1547 880
rect 1676 880 1683 883
rect 816 716 843 723
rect 696 656 723 663
rect 216 176 223 233
rect 316 146 323 313
rect 536 207 543 353
rect 656 247 663 433
rect 676 366 683 633
rect 696 627 703 656
rect 753 647 767 652
rect 816 627 823 693
rect 836 666 843 716
rect 856 687 863 813
rect 896 696 903 733
rect 936 696 943 753
rect 1367 713 1373 727
rect 1427 713 1433 727
rect 1233 700 1247 713
rect 1236 696 1243 700
rect 1436 696 1483 703
rect 916 660 923 663
rect 816 467 823 613
rect 836 447 843 652
rect 913 647 927 660
rect 716 396 723 433
rect 873 400 887 413
rect 876 396 883 400
rect 916 396 923 453
rect 736 327 743 363
rect 776 287 783 363
rect 633 227 647 233
rect 413 180 427 193
rect 416 176 423 180
rect 536 176 543 193
rect 576 176 583 213
rect 96 87 103 143
rect 236 107 243 143
rect 396 127 403 143
rect 496 127 503 173
rect 556 140 563 143
rect 553 127 567 140
rect 393 107 407 113
rect 596 87 603 143
rect 613 107 627 113
rect 636 87 643 174
rect 656 146 663 233
rect 673 227 687 233
rect 816 146 823 393
rect 976 363 983 473
rect 1036 427 1043 694
rect 1136 627 1143 694
rect 1216 627 1223 652
rect 1056 396 1063 473
rect 1116 363 1123 453
rect 1156 366 1163 413
rect 1196 396 1203 473
rect 1236 396 1243 493
rect 1296 367 1303 593
rect 1336 507 1343 694
rect 1376 467 1383 652
rect 1416 627 1423 663
rect 896 327 903 363
rect 936 356 983 363
rect 1076 356 1123 363
rect 1316 366 1323 413
rect 1356 396 1363 453
rect 1396 396 1403 493
rect 1476 487 1483 696
rect 1496 666 1503 713
rect 1556 696 1563 773
rect 1536 627 1543 663
rect 1536 613 1553 627
rect 1536 607 1543 613
rect 1636 587 1643 872
rect 1673 867 1687 880
rect 1736 747 1743 916
rect 1796 927 1803 1183
rect 1836 1107 1843 1293
rect 1856 1247 1863 1403
rect 1936 1387 1943 1493
rect 1976 1436 1983 1473
rect 2016 1436 2023 1553
rect 2056 1443 2063 1673
rect 2156 1667 2163 1833
rect 2176 1687 2183 1753
rect 2276 1607 2283 1793
rect 2296 1647 2303 1813
rect 2316 1706 2323 1853
rect 2396 1736 2403 1833
rect 2456 1807 2463 2073
rect 2556 1968 2563 2173
rect 2676 2167 2683 2933
rect 2696 2787 2703 2994
rect 2796 2746 2803 2813
rect 2756 2567 2763 2743
rect 2696 2387 2703 2433
rect 2696 2207 2703 2373
rect 2736 2367 2743 2443
rect 2756 2256 2763 2413
rect 2776 2387 2783 2443
rect 2796 2323 2803 2433
rect 2816 2343 2823 2913
rect 2836 2443 2843 2952
rect 2876 2827 2883 2994
rect 2876 2607 2883 2743
rect 2896 2667 2903 3033
rect 2967 3023 2980 3027
rect 2967 3013 2983 3023
rect 2976 2996 2983 3013
rect 3016 2996 3023 3033
rect 2956 2907 2963 2963
rect 2996 2960 3003 2963
rect 2993 2947 3007 2960
rect 2976 2847 2983 2873
rect 3096 2827 3103 3116
rect 3136 2996 3143 3093
rect 3216 2967 3223 3013
rect 3236 3008 3243 3456
rect 3256 3407 3263 3483
rect 3316 3467 3323 3514
rect 3336 3447 3343 3573
rect 3416 3516 3423 3853
rect 3436 3643 3443 3813
rect 3536 3787 3543 3953
rect 3496 3767 3503 3783
rect 3496 3756 3513 3767
rect 3500 3753 3513 3756
rect 3556 3747 3563 4153
rect 3576 3967 3583 4213
rect 3636 4036 3643 4303
rect 3656 4227 3663 4933
rect 3716 4856 3723 4973
rect 3676 4647 3683 4813
rect 3676 4427 3683 4573
rect 3696 4427 3703 4753
rect 3736 4687 3743 4823
rect 3776 4807 3783 4853
rect 3796 4826 3803 4973
rect 3836 4947 3843 4973
rect 3896 4856 3903 5193
rect 3916 5027 3923 5113
rect 3956 5040 3963 5043
rect 3953 5027 3967 5040
rect 3876 4820 3883 4823
rect 3873 4807 3887 4820
rect 3916 4727 3923 4753
rect 3713 4587 3727 4593
rect 3713 4567 3727 4573
rect 3756 4556 3763 4693
rect 3796 4568 3803 4613
rect 3716 4387 3723 4513
rect 3736 4467 3743 4523
rect 3696 4267 3703 4353
rect 3753 4340 3767 4353
rect 3756 4336 3763 4340
rect 3796 4336 3803 4473
rect 3736 4207 3743 4303
rect 3776 4247 3783 4303
rect 3667 4073 3673 4087
rect 3673 4040 3687 4052
rect 3696 4047 3703 4193
rect 3716 4087 3723 4133
rect 3676 4036 3683 4040
rect 3656 3927 3663 4003
rect 3696 3963 3703 3993
rect 3716 3987 3723 4052
rect 3696 3956 3723 3963
rect 3616 3867 3623 3893
rect 3656 3816 3663 3873
rect 3576 3776 3603 3783
rect 3436 3636 3463 3643
rect 3436 3583 3443 3613
rect 3456 3607 3463 3636
rect 3436 3576 3463 3583
rect 3396 3467 3403 3483
rect 3387 3456 3403 3467
rect 3387 3453 3400 3456
rect 3316 3436 3333 3443
rect 3316 3227 3323 3436
rect 3273 3000 3287 3013
rect 3313 3000 3327 3013
rect 3276 2996 3283 3000
rect 3316 2996 3323 3000
rect 2913 2480 2927 2493
rect 2956 2487 2963 2793
rect 3013 2780 3027 2793
rect 3016 2776 3023 2780
rect 3076 2667 3083 2743
rect 2916 2476 2923 2480
rect 2836 2436 2863 2443
rect 2816 2336 2843 2343
rect 2796 2316 2823 2323
rect 2736 2187 2743 2223
rect 2776 2167 2783 2212
rect 2816 2167 2823 2316
rect 2476 1847 2483 1913
rect 2073 1443 2087 1453
rect 2056 1440 2087 1443
rect 2056 1436 2083 1440
rect 2036 1400 2043 1403
rect 2033 1387 2047 1400
rect 2076 1323 2083 1373
rect 2076 1316 2103 1323
rect 1876 1186 1883 1253
rect 1956 1147 1963 1183
rect 1996 1167 2003 1213
rect 2016 1186 2023 1293
rect 2056 1228 2063 1253
rect 2076 1247 2083 1293
rect 2096 1216 2103 1316
rect 2156 1187 2163 1393
rect 2116 1163 2123 1183
rect 2087 1156 2123 1163
rect 2176 1147 2183 1573
rect 2196 1407 2203 1593
rect 2316 1527 2323 1692
rect 2336 1687 2343 1734
rect 2556 1736 2563 1873
rect 2616 1807 2623 1853
rect 2496 1706 2503 1733
rect 2616 1706 2623 1753
rect 2376 1700 2383 1703
rect 2373 1687 2387 1700
rect 2636 1667 2643 1813
rect 2716 1767 2723 2153
rect 2736 1843 2743 2152
rect 2796 1920 2803 1923
rect 2793 1907 2807 1920
rect 2836 1907 2843 2336
rect 2736 1836 2763 1843
rect 2756 1703 2763 1836
rect 2816 1747 2823 1853
rect 2856 1827 2863 2436
rect 2896 2367 2903 2443
rect 2936 2223 2943 2443
rect 2976 2226 2983 2653
rect 3116 2647 3123 2933
rect 3236 2927 3243 2994
rect 3336 2943 3343 2963
rect 3296 2936 3343 2943
rect 3296 2927 3303 2936
rect 3136 2587 3143 2813
rect 3156 2707 3163 2774
rect 2996 2268 3003 2573
rect 3027 2503 3040 2507
rect 3027 2493 3043 2503
rect 3036 2476 3043 2493
rect 3156 2407 3163 2533
rect 3036 2256 3043 2393
rect 3156 2323 3163 2353
rect 3176 2347 3183 2633
rect 3216 2587 3223 2673
rect 3256 2667 3263 2853
rect 3296 2747 3303 2913
rect 3316 2776 3323 2813
rect 3376 2788 3383 3213
rect 3396 3147 3403 3433
rect 3416 3308 3423 3353
rect 3416 3267 3423 3294
rect 3396 2727 3403 3133
rect 3416 3087 3423 3193
rect 3436 3067 3443 3473
rect 3456 3127 3463 3576
rect 3476 3447 3483 3573
rect 3496 3527 3503 3733
rect 3556 3667 3563 3693
rect 3576 3627 3583 3776
rect 3633 3767 3647 3772
rect 3673 3767 3687 3773
rect 3596 3727 3603 3753
rect 3516 3516 3523 3553
rect 3536 3476 3583 3483
rect 3636 3447 3643 3732
rect 3696 3707 3703 3814
rect 3716 3723 3723 3956
rect 3736 3947 3743 4093
rect 3756 4003 3763 4133
rect 3836 4107 3843 4554
rect 3856 4447 3863 4613
rect 3916 4568 3923 4713
rect 3936 4687 3943 5013
rect 3996 4967 4003 5043
rect 3976 4956 3993 4963
rect 3956 4627 3963 4893
rect 3976 4826 3983 4956
rect 4036 4907 4043 5273
rect 4076 5227 4083 5273
rect 4096 5103 4103 5533
rect 4176 5416 4183 5513
rect 4136 5187 4143 5213
rect 4156 5127 4163 5153
rect 4076 5096 4103 5103
rect 4056 4947 4063 5033
rect 4076 4907 4083 5096
rect 4156 5076 4163 5113
rect 4116 4967 4123 5043
rect 4196 5027 4203 5253
rect 4136 4927 4143 4993
rect 3856 4167 3863 4412
rect 3876 4207 3883 4513
rect 3896 4387 3903 4523
rect 3976 4516 4003 4523
rect 3916 4227 3923 4303
rect 3936 4187 3943 4253
rect 3796 4048 3803 4073
rect 3836 4036 3843 4072
rect 3756 3996 3783 4003
rect 3816 4000 3823 4003
rect 3776 3816 3783 3996
rect 3813 3987 3827 4000
rect 3876 3983 3883 4053
rect 3896 4007 3903 4113
rect 3913 4087 3927 4093
rect 3956 4087 3963 4292
rect 3976 4083 3983 4433
rect 3996 4427 4003 4516
rect 3996 4348 4003 4413
rect 3996 4107 4003 4334
rect 3976 4076 4003 4083
rect 3916 4047 3923 4073
rect 3933 4040 3947 4053
rect 3936 4036 3943 4040
rect 3996 4047 4003 4076
rect 3856 3976 3883 3983
rect 3756 3780 3763 3783
rect 3753 3767 3767 3780
rect 3716 3716 3733 3723
rect 3736 3627 3743 3713
rect 3756 3607 3763 3673
rect 3796 3607 3803 3633
rect 3796 3523 3803 3553
rect 3756 3516 3803 3523
rect 3496 3227 3503 3263
rect 3427 3023 3440 3027
rect 3427 3013 3443 3023
rect 3436 2996 3443 3013
rect 3476 3007 3483 3053
rect 3416 2627 3423 2953
rect 3456 2907 3463 2952
rect 3213 2480 3227 2493
rect 3276 2488 3283 2593
rect 3427 2583 3440 2587
rect 3427 2580 3443 2583
rect 3427 2573 3447 2580
rect 3433 2567 3447 2573
rect 3416 2503 3423 2533
rect 3396 2496 3423 2503
rect 3216 2476 3223 2480
rect 3396 2476 3403 2496
rect 3216 2323 3223 2413
rect 3416 2347 3423 2433
rect 3156 2316 3223 2323
rect 3076 2256 3083 2293
rect 3096 2267 3103 2313
rect 3173 2260 3187 2273
rect 3176 2256 3183 2260
rect 2927 2216 2943 2223
rect 2936 2007 2943 2216
rect 2996 2107 3003 2133
rect 3016 2047 3023 2223
rect 3056 2003 3063 2212
rect 3116 2087 3123 2113
rect 3036 1996 3063 2003
rect 2876 1887 2883 1954
rect 2976 1887 2983 1923
rect 3016 1887 3023 1993
rect 2856 1736 2863 1773
rect 2896 1748 2903 1853
rect 2296 1406 2303 1513
rect 2256 1347 2263 1403
rect 2307 1396 2323 1403
rect 2267 1336 2283 1343
rect 2236 1216 2243 1273
rect 2276 1227 2283 1336
rect 1827 963 1840 967
rect 1827 953 1843 963
rect 1836 943 1843 953
rect 1836 936 1863 943
rect 1756 867 1763 914
rect 1856 916 1863 936
rect 1976 916 1983 953
rect 1756 696 1763 853
rect 1836 708 1843 883
rect 1996 787 2003 872
rect 1916 696 1923 773
rect 1656 627 1663 694
rect 1776 587 1783 663
rect 1896 660 1903 663
rect 1893 647 1907 660
rect 1956 647 1963 733
rect 2056 696 2063 914
rect 1976 667 1983 694
rect 2116 667 2123 713
rect 2176 707 2183 1133
rect 2196 887 2203 1173
rect 2256 1027 2263 1172
rect 2296 1167 2303 1273
rect 2316 928 2323 1396
rect 2336 1247 2343 1573
rect 2416 1436 2423 1473
rect 2416 1216 2423 1253
rect 2456 1186 2463 1253
rect 2356 1180 2363 1183
rect 2276 807 2283 883
rect 2276 747 2283 793
rect 2253 700 2267 713
rect 2256 696 2263 700
rect 2076 660 2083 663
rect 2073 647 2087 660
rect 2020 645 2040 647
rect 2027 633 2033 645
rect 1513 400 1527 413
rect 1516 396 1523 400
rect 1556 396 1563 493
rect 1576 287 1583 363
rect 1636 287 1643 394
rect 1656 327 1663 433
rect 1736 396 1743 473
rect 1796 367 1803 473
rect 2036 396 2043 433
rect 916 176 923 233
rect 976 146 983 253
rect 1176 176 1183 253
rect 1256 146 1263 273
rect 1316 176 1323 213
rect 1396 167 1403 273
rect 1716 227 1723 352
rect 1476 176 1483 213
rect 1513 180 1527 193
rect 1516 176 1523 180
rect 1676 176 1683 213
rect 1416 146 1423 173
rect 856 140 863 143
rect 853 127 867 140
rect 896 107 903 143
rect 1016 107 1023 143
rect 1196 140 1203 143
rect 1193 127 1207 140
rect 1336 140 1343 143
rect 1333 127 1347 140
rect 1447 143 1460 147
rect 1447 136 1463 143
rect 1496 140 1503 143
rect 1447 133 1460 136
rect 1493 127 1507 140
rect 1700 143 1713 147
rect 1696 136 1713 143
rect 1700 133 1713 136
rect 1736 146 1743 193
rect 1756 147 1763 313
rect 1796 176 1803 273
rect 1816 207 1823 394
rect 1836 176 1843 253
rect 1896 247 1903 363
rect 1976 327 1983 373
rect 2096 307 2103 363
rect 1896 146 1903 233
rect 2016 176 2023 233
rect 1387 113 1393 127
rect 727 93 733 107
rect 1656 87 1663 132
rect 1916 107 1923 173
rect 1996 107 2003 132
rect 2016 83 2023 113
rect 1987 76 2023 83
rect 2056 27 2063 213
rect 2076 187 2083 253
rect 2136 227 2143 693
rect 2316 663 2323 733
rect 2236 660 2243 663
rect 2233 647 2247 660
rect 2296 656 2323 663
rect 2256 396 2263 433
rect 2156 176 2163 394
rect 2216 143 2223 233
rect 2336 227 2343 1173
rect 2353 1167 2367 1180
rect 2436 916 2443 953
rect 2476 943 2483 1433
rect 2516 1407 2523 1653
rect 2676 1607 2683 1703
rect 2716 1647 2723 1703
rect 2736 1696 2763 1703
rect 2613 1440 2627 1453
rect 2616 1436 2623 1440
rect 2496 1187 2503 1373
rect 2696 1216 2703 1393
rect 2716 1243 2723 1513
rect 2736 1327 2743 1696
rect 2776 1607 2783 1713
rect 2796 1706 2803 1733
rect 2816 1667 2823 1693
rect 2796 1527 2803 1653
rect 2796 1400 2803 1403
rect 2793 1387 2807 1400
rect 2716 1236 2743 1243
rect 2736 1228 2743 1236
rect 2616 1167 2623 1213
rect 2676 1180 2683 1183
rect 2673 1167 2687 1180
rect 2556 1027 2563 1073
rect 2476 936 2503 943
rect 2416 787 2423 883
rect 2476 747 2483 913
rect 2416 696 2423 733
rect 2453 700 2467 713
rect 2456 696 2463 700
rect 2356 367 2363 433
rect 2376 408 2383 473
rect 2396 396 2403 533
rect 2436 467 2443 663
rect 2476 403 2483 473
rect 2496 427 2503 936
rect 2516 867 2523 953
rect 2556 916 2563 1013
rect 2633 920 2647 933
rect 2636 916 2643 920
rect 2576 880 2583 883
rect 2616 880 2623 883
rect 2573 867 2587 880
rect 2613 867 2627 880
rect 2587 860 2603 863
rect 2587 856 2607 860
rect 2593 847 2607 856
rect 2536 747 2543 793
rect 2516 547 2523 713
rect 2556 696 2563 773
rect 2596 696 2603 793
rect 2576 547 2583 663
rect 2476 396 2503 403
rect 2313 180 2327 193
rect 2316 176 2323 180
rect 2396 146 2403 313
rect 2416 307 2423 363
rect 2456 307 2463 363
rect 2456 176 2463 213
rect 2496 207 2503 396
rect 2516 366 2523 533
rect 2136 140 2143 143
rect 2133 127 2147 140
rect 2176 136 2223 143
rect 2336 107 2343 143
rect 2436 107 2443 173
rect 1936 -24 1943 13
rect 2436 -24 2443 13
rect 2496 -17 2503 143
rect 2536 27 2543 413
rect 2616 396 2623 493
rect 2636 487 2643 833
rect 2656 663 2663 873
rect 2676 867 2683 1033
rect 2696 887 2703 1153
rect 2716 787 2723 1183
rect 2776 1167 2783 1313
rect 2836 1267 2843 1593
rect 2856 1327 2863 1653
rect 2876 1647 2883 1703
rect 2876 1387 2883 1434
rect 2896 1407 2903 1673
rect 2936 1667 2943 1773
rect 2956 1687 2963 1793
rect 3036 1767 3043 1996
rect 3096 1920 3103 1923
rect 3093 1907 3107 1920
rect 3136 1926 3143 2093
rect 3116 1827 3123 1913
rect 3156 1747 3163 2033
rect 3187 1963 3200 1967
rect 3187 1956 3203 1963
rect 3236 1956 3243 2013
rect 3187 1953 3200 1956
rect 3296 1927 3303 2333
rect 3356 2256 3363 2333
rect 3256 1807 3263 1912
rect 2996 1647 3003 1703
rect 2976 1436 2983 1613
rect 3036 1607 3043 1703
rect 3136 1700 3143 1703
rect 3133 1687 3147 1700
rect 3146 1680 3147 1687
rect 3156 1627 3163 1673
rect 3176 1647 3183 1753
rect 3196 1687 3203 1793
rect 3316 1706 3323 2173
rect 3336 1967 3343 2212
rect 3356 1956 3363 2013
rect 3376 1987 3383 2223
rect 3436 2187 3443 2473
rect 3456 2407 3463 2713
rect 3496 2583 3503 2743
rect 3516 2607 3523 2833
rect 3496 2576 3523 2583
rect 3516 2507 3523 2576
rect 3536 2487 3543 2713
rect 3516 2367 3523 2443
rect 3556 2427 3563 3433
rect 3576 2927 3583 3413
rect 3656 3407 3663 3513
rect 3796 3483 3803 3516
rect 3776 3476 3803 3483
rect 3776 3407 3783 3476
rect 3816 3447 3823 3773
rect 3836 3667 3843 3933
rect 3856 3767 3863 3976
rect 3993 3983 4007 3993
rect 3976 3980 4007 3983
rect 3976 3976 4003 3980
rect 3876 3747 3883 3953
rect 3896 3827 3903 3972
rect 3936 3828 3943 3913
rect 3976 3827 3983 3976
rect 4016 3967 4023 4554
rect 4036 4527 4043 4713
rect 4056 4567 4063 4823
rect 4076 4556 4083 4613
rect 4116 4588 4123 4893
rect 4216 4856 4223 5133
rect 4236 4887 4243 5313
rect 4256 5267 4263 5833
rect 4296 5827 4303 5863
rect 4376 5807 4383 6013
rect 4696 6007 4703 6114
rect 4776 6047 4783 6083
rect 4856 6047 4863 6233
rect 4876 6147 4883 6372
rect 4896 6147 4903 6213
rect 4916 6167 4923 6372
rect 5073 6367 5087 6380
rect 4956 6116 4963 6293
rect 4936 6047 4943 6083
rect 4436 5947 4443 5973
rect 4436 5896 4443 5933
rect 4756 5896 4763 5933
rect 4396 5707 4403 5893
rect 4276 5567 4283 5653
rect 4316 5527 4323 5563
rect 4276 5346 4283 5513
rect 4376 5467 4383 5493
rect 4376 5376 4383 5453
rect 4336 5127 4343 5213
rect 4356 5207 4363 5332
rect 4416 5267 4423 5374
rect 4396 5107 4403 5193
rect 4276 5040 4283 5043
rect 4273 5027 4287 5040
rect 4416 5043 4423 5253
rect 4436 5187 4443 5513
rect 4456 5467 4463 5563
rect 4496 5376 4503 5553
rect 4516 5527 4523 5594
rect 4536 5527 4543 5833
rect 4556 5767 4563 5863
rect 4556 5647 4563 5753
rect 4616 5727 4623 5863
rect 4636 5767 4643 5894
rect 4576 5603 4583 5713
rect 4636 5628 4643 5653
rect 4676 5647 4683 5894
rect 4736 5860 4743 5863
rect 4733 5847 4747 5860
rect 4736 5807 4743 5833
rect 4556 5596 4583 5603
rect 4516 5267 4523 5343
rect 4556 5247 4563 5596
rect 4596 5447 4603 5533
rect 4616 5527 4623 5563
rect 4676 5487 4683 5633
rect 4696 5547 4703 5613
rect 4736 5596 4743 5693
rect 4776 5687 4783 5863
rect 4576 5346 4583 5413
rect 4636 5376 4643 5473
rect 4656 5267 4663 5343
rect 4676 5287 4683 5313
rect 4696 5267 4703 5493
rect 4716 5307 4723 5473
rect 4756 5447 4763 5563
rect 4816 5487 4823 5693
rect 4836 5427 4843 5753
rect 4856 5608 4863 5953
rect 4916 5860 4923 5863
rect 4913 5847 4927 5860
rect 4956 5687 4963 6053
rect 4996 6047 5003 6173
rect 5016 6027 5023 6353
rect 5196 6347 5203 6383
rect 5076 6080 5083 6083
rect 5073 6067 5087 6080
rect 5116 5927 5123 6113
rect 5136 6086 5143 6333
rect 5376 6307 5383 6383
rect 5416 6380 5423 6383
rect 5413 6367 5427 6380
rect 5456 6367 5463 6453
rect 5507 6438 5533 6445
rect 5176 6247 5183 6273
rect 5176 6116 5183 6233
rect 5196 6187 5203 6253
rect 5216 6167 5223 6193
rect 5216 6116 5223 6153
rect 5376 6116 5383 6193
rect 5476 6167 5483 6413
rect 5576 6207 5583 6493
rect 5647 6436 5693 6443
rect 5716 6416 5723 6473
rect 5893 6467 5907 6473
rect 5947 6453 5953 6467
rect 5807 6436 5863 6443
rect 5856 6428 5863 6436
rect 5916 6387 5923 6453
rect 5656 6380 5663 6383
rect 5633 6367 5647 6373
rect 5653 6367 5667 6380
rect 5836 6380 5843 6383
rect 5707 6356 5733 6363
rect 5756 6287 5763 6372
rect 5833 6367 5847 6380
rect 5787 6353 5793 6367
rect 5836 6307 5843 6353
rect 5053 5900 5067 5913
rect 5056 5896 5063 5900
rect 5096 5896 5143 5903
rect 5076 5807 5083 5863
rect 5136 5787 5143 5896
rect 5156 5707 5163 5993
rect 5396 5967 5403 6083
rect 5213 5900 5227 5913
rect 5216 5896 5223 5900
rect 5196 5807 5203 5863
rect 4776 5376 4783 5413
rect 4756 5340 4763 5343
rect 4476 5076 4483 5113
rect 4416 5036 4463 5043
rect 4136 4743 4143 4854
rect 4136 4736 4163 4743
rect 4096 4520 4103 4523
rect 4093 4507 4107 4520
rect 4156 4427 4163 4736
rect 4176 4507 4183 4773
rect 4196 4767 4203 4823
rect 4276 4807 4283 4913
rect 4256 4727 4263 4773
rect 4296 4747 4303 4812
rect 4316 4787 4323 5032
rect 4533 5023 4547 5033
rect 4516 5020 4547 5023
rect 4513 5016 4543 5020
rect 4513 5007 4527 5016
rect 4376 4868 4383 4933
rect 4356 4807 4363 4823
rect 4356 4683 4363 4793
rect 4336 4676 4363 4683
rect 4196 4523 4203 4673
rect 4336 4563 4343 4676
rect 4316 4556 4343 4563
rect 4376 4556 4383 4593
rect 4396 4587 4403 4773
rect 4436 4763 4443 4854
rect 4456 4787 4463 4993
rect 4476 4767 4483 4873
rect 4536 4868 4543 4973
rect 4556 4947 4563 5093
rect 4416 4756 4443 4763
rect 4416 4647 4423 4756
rect 4416 4607 4423 4633
rect 4196 4520 4223 4523
rect 4196 4516 4227 4520
rect 4213 4507 4227 4516
rect 4236 4487 4243 4523
rect 4036 4303 4043 4333
rect 4036 4296 4053 4303
rect 4176 4247 4183 4393
rect 4196 4348 4203 4413
rect 4036 3907 4043 4233
rect 4076 4107 4083 4213
rect 4093 4040 4107 4053
rect 4096 4036 4103 4040
rect 4136 4036 4143 4113
rect 4116 3903 4123 4003
rect 4176 3987 4183 4193
rect 4216 4067 4223 4373
rect 4276 4336 4283 4393
rect 4296 4367 4303 4553
rect 4316 4447 4323 4556
rect 4400 4523 4413 4527
rect 4356 4427 4363 4523
rect 4396 4516 4413 4523
rect 4400 4513 4413 4516
rect 4356 4387 4363 4413
rect 4256 4123 4263 4303
rect 4296 4300 4303 4303
rect 4293 4287 4307 4300
rect 4236 4116 4263 4123
rect 4236 4067 4243 4116
rect 4276 4048 4283 4273
rect 4376 4267 4383 4493
rect 4436 4447 4443 4573
rect 4456 4527 4463 4693
rect 4456 4336 4463 4393
rect 4476 4367 4483 4753
rect 4556 4747 4563 4823
rect 4576 4807 4583 5213
rect 4596 5023 4603 5173
rect 4616 5087 4623 5253
rect 4667 5094 4673 5107
rect 4660 5093 4673 5094
rect 4636 5040 4643 5043
rect 4633 5027 4647 5040
rect 4596 5016 4623 5023
rect 4596 4747 4603 4853
rect 4616 4667 4623 5016
rect 4696 4887 4703 5074
rect 4673 4860 4687 4873
rect 4716 4867 4723 5272
rect 4736 5227 4743 5333
rect 4753 5327 4767 5340
rect 4796 5327 4803 5343
rect 4796 5316 4813 5327
rect 4800 5313 4813 5316
rect 4756 5127 4763 5313
rect 4776 5147 4783 5293
rect 4836 5247 4843 5343
rect 4793 5088 4807 5093
rect 4776 4987 4783 5043
rect 4876 5027 4883 5563
rect 4916 5560 4923 5563
rect 4913 5547 4927 5560
rect 4956 5507 4963 5673
rect 5076 5596 5083 5633
rect 5016 5507 5023 5552
rect 5116 5527 5123 5633
rect 5156 5547 5163 5593
rect 5176 5567 5183 5653
rect 5316 5647 5323 5893
rect 5216 5527 5223 5563
rect 5276 5560 5283 5563
rect 5273 5547 5287 5560
rect 4896 5327 4903 5493
rect 4956 5388 4963 5433
rect 4996 5383 5003 5413
rect 4996 5376 5023 5383
rect 4936 5247 4943 5343
rect 4976 5263 4983 5343
rect 4956 5256 4983 5263
rect 4956 5207 4963 5256
rect 4893 5087 4907 5093
rect 4836 4947 4843 4973
rect 4896 4967 4903 5033
rect 4736 4887 4743 4933
rect 4676 4856 4683 4860
rect 4656 4747 4663 4823
rect 4696 4816 4713 4823
rect 4396 4287 4403 4333
rect 4496 4303 4503 4653
rect 4636 4607 4643 4633
rect 4636 4543 4643 4593
rect 4656 4568 4663 4653
rect 4636 4536 4663 4543
rect 4196 4036 4243 4043
rect 4096 3896 4123 3903
rect 4076 3827 4083 3893
rect 4096 3867 4103 3896
rect 3916 3707 3923 3783
rect 3916 3527 3923 3633
rect 3836 3423 3843 3514
rect 3936 3487 3943 3733
rect 3956 3727 3963 3783
rect 3816 3416 3843 3423
rect 3736 3347 3743 3393
rect 3636 3087 3643 3333
rect 3676 3167 3683 3263
rect 3613 3000 3627 3013
rect 3616 2996 3623 3000
rect 3676 2996 3683 3073
rect 3796 2967 3803 3373
rect 3816 3227 3823 3416
rect 3936 3303 3943 3473
rect 3956 3427 3963 3692
rect 3976 3647 3983 3773
rect 3976 3527 3983 3593
rect 3996 3567 4003 3783
rect 4096 3727 4103 3832
rect 4116 3747 4123 3873
rect 4196 3823 4203 4036
rect 4213 3987 4227 3993
rect 4176 3816 4223 3823
rect 4216 3607 4223 3816
rect 3993 3520 4007 3532
rect 3996 3516 4003 3520
rect 4036 3516 4043 3593
rect 4016 3363 4023 3483
rect 4076 3387 4083 3533
rect 4096 3487 4103 3553
rect 4216 3487 4223 3514
rect 3996 3356 4023 3363
rect 3936 3296 3963 3303
rect 3916 3087 3923 3263
rect 3916 2996 3923 3073
rect 3613 2780 3627 2793
rect 3616 2776 3623 2780
rect 3676 2787 3683 2913
rect 3696 2788 3703 2953
rect 3736 2927 3743 2963
rect 3736 2887 3743 2913
rect 3816 2827 3823 2993
rect 3713 2787 3727 2793
rect 3696 2747 3703 2774
rect 3596 2740 3603 2743
rect 3593 2727 3607 2740
rect 3493 2260 3507 2273
rect 3496 2256 3503 2260
rect 3536 2227 3543 2273
rect 3396 2007 3403 2113
rect 3476 2087 3483 2223
rect 3396 1867 3403 1893
rect 3336 1748 3343 1773
rect 2996 1487 3003 1593
rect 3016 1327 3023 1403
rect 3076 1327 3083 1553
rect 2796 1167 2803 1213
rect 2816 967 2823 1213
rect 3076 1183 3083 1273
rect 2856 1180 2863 1183
rect 2853 1167 2867 1180
rect 2896 1027 2903 1183
rect 2996 1147 3003 1183
rect 3036 1176 3083 1183
rect 3096 1147 3103 1593
rect 3196 1527 3203 1633
rect 3253 1467 3267 1473
rect 3236 1456 3253 1463
rect 3116 1307 3123 1393
rect 3236 1367 3243 1456
rect 3276 1448 3283 1693
rect 3336 1687 3343 1734
rect 3356 1667 3363 1813
rect 3476 1807 3483 2032
rect 3516 1983 3523 2093
rect 3536 2047 3543 2213
rect 3576 2107 3583 2713
rect 3636 2687 3643 2743
rect 3673 2727 3687 2733
rect 3716 2707 3723 2752
rect 3733 2727 3747 2733
rect 3756 2687 3763 2743
rect 3596 2367 3603 2613
rect 3616 2467 3623 2653
rect 3676 2476 3683 2513
rect 3616 2327 3623 2453
rect 3636 2287 3643 2443
rect 3593 2268 3607 2273
rect 3516 1976 3543 1983
rect 3496 1827 3503 1973
rect 3536 1956 3543 1976
rect 3596 1956 3603 2173
rect 3636 1907 3643 2053
rect 3416 1736 3423 1793
rect 3516 1767 3523 1833
rect 3596 1807 3603 1833
rect 3616 1787 3623 1853
rect 3396 1700 3403 1703
rect 3393 1687 3407 1700
rect 3296 1467 3303 1493
rect 3316 1487 3323 1573
rect 3313 1440 3327 1452
rect 3316 1436 3323 1440
rect 3356 1436 3363 1533
rect 3376 1443 3383 1593
rect 3396 1583 3403 1652
rect 3416 1607 3423 1633
rect 3396 1576 3423 1583
rect 3376 1436 3403 1443
rect 3176 1216 3183 1293
rect 3216 1216 3223 1273
rect 3116 1186 3123 1213
rect 3007 1136 3023 1143
rect 2776 867 2783 883
rect 2776 747 2783 853
rect 2816 747 2823 883
rect 2856 867 2863 914
rect 2693 700 2707 713
rect 2696 696 2703 700
rect 2656 656 2683 663
rect 2636 203 2643 363
rect 2636 196 2663 203
rect 2476 -24 2503 -17
rect 2556 -24 2563 193
rect 2656 146 2663 196
rect 2676 187 2683 656
rect 2696 366 2703 493
rect 2716 408 2723 663
rect 2776 587 2783 673
rect 2876 663 2883 872
rect 2956 696 2963 853
rect 2976 847 2983 883
rect 2856 656 2883 663
rect 2756 396 2763 453
rect 2776 360 2783 363
rect 2773 347 2787 360
rect 2816 183 2823 353
rect 2836 307 2843 413
rect 2856 363 2863 656
rect 2976 627 2983 663
rect 2876 407 2883 533
rect 2916 396 2923 453
rect 2856 356 2883 363
rect 2876 327 2883 356
rect 2796 176 2823 183
rect 2916 176 2923 313
rect 2996 287 3003 394
rect 3016 183 3023 1136
rect 3036 547 3043 1053
rect 3136 916 3143 953
rect 3236 916 3243 1053
rect 3276 967 3283 1434
rect 3336 1387 3343 1403
rect 3336 1243 3343 1373
rect 3316 1236 3343 1243
rect 3316 1228 3323 1236
rect 3336 1007 3343 1183
rect 3376 1027 3383 1393
rect 3396 1067 3403 1436
rect 3416 1407 3423 1576
rect 3436 1487 3443 1533
rect 3496 1447 3503 1733
rect 3516 1707 3523 1753
rect 3573 1740 3587 1753
rect 3616 1747 3623 1773
rect 3576 1736 3583 1740
rect 3516 1667 3523 1693
rect 3556 1547 3563 1613
rect 3616 1587 3623 1673
rect 3616 1468 3623 1513
rect 3636 1507 3643 1733
rect 3656 1567 3663 2413
rect 3676 2123 3683 2413
rect 3696 2387 3703 2493
rect 3716 2488 3723 2593
rect 3696 2147 3703 2333
rect 3676 2116 3703 2123
rect 3676 1947 3683 2093
rect 3696 1867 3703 2116
rect 3716 2067 3723 2474
rect 3756 2256 3763 2453
rect 3796 2440 3803 2443
rect 3793 2427 3807 2440
rect 3876 2427 3883 2873
rect 3896 2407 3903 2853
rect 3916 2787 3923 2913
rect 3956 2867 3963 3296
rect 3996 3266 4003 3356
rect 3976 3047 3983 3113
rect 3976 2907 3983 3012
rect 3996 2807 4003 3073
rect 4016 3027 4023 3333
rect 4116 3296 4123 3373
rect 4036 3127 4043 3193
rect 4076 3027 4083 3213
rect 4096 3167 4103 3263
rect 4116 3127 4123 3173
rect 4053 3000 4067 3013
rect 4093 3000 4107 3013
rect 4056 2996 4063 3000
rect 4096 2996 4103 3000
rect 4036 2847 4043 2963
rect 4113 2947 4127 2953
rect 4036 2746 4043 2793
rect 4056 2687 4063 2793
rect 3916 2476 3923 2673
rect 4056 2607 4063 2673
rect 3976 2447 3983 2553
rect 3956 2440 3963 2443
rect 3953 2427 3967 2440
rect 3756 2107 3763 2153
rect 3756 1956 3763 2093
rect 3776 2087 3783 2223
rect 3856 2187 3863 2223
rect 3856 2027 3863 2173
rect 3956 2167 3963 2392
rect 3976 2287 3983 2433
rect 4016 2387 4023 2493
rect 4056 2476 4063 2572
rect 4076 2527 4083 2913
rect 4096 2827 4103 2853
rect 4116 2807 4123 2873
rect 4136 2847 4143 3253
rect 4156 2927 4163 3413
rect 4176 3107 4183 3453
rect 4196 3307 4203 3473
rect 4236 3363 4243 3973
rect 4256 3427 4263 3953
rect 4316 3927 4323 4253
rect 4416 4227 4423 4303
rect 4476 4296 4503 4303
rect 4416 4036 4423 4073
rect 4276 3827 4283 3913
rect 4336 3867 4343 4034
rect 4396 3967 4403 3992
rect 4376 3787 4383 3853
rect 4336 3763 4343 3783
rect 4316 3756 4343 3763
rect 4316 3687 4323 3756
rect 4316 3480 4323 3483
rect 4216 3360 4243 3363
rect 4213 3356 4243 3360
rect 4213 3347 4227 3356
rect 4176 2967 4183 3093
rect 4196 3027 4203 3253
rect 4216 3187 4223 3263
rect 4216 3087 4223 3133
rect 4216 2996 4223 3073
rect 4256 3027 4263 3253
rect 4276 3127 4283 3473
rect 4313 3467 4327 3480
rect 4296 3387 4303 3453
rect 4356 3407 4363 3483
rect 4376 3347 4383 3473
rect 4396 3463 4403 3913
rect 4416 3487 4423 3933
rect 4476 3927 4483 4296
rect 4496 4007 4503 4093
rect 4516 4047 4523 4433
rect 4556 4347 4563 4483
rect 4573 4340 4587 4353
rect 4576 4336 4583 4340
rect 4616 4336 4623 4453
rect 4536 4227 4543 4253
rect 4596 4227 4603 4303
rect 4576 4048 4583 4073
rect 4476 3828 4483 3873
rect 4536 3827 4543 3973
rect 4396 3456 4423 3463
rect 4296 3267 4303 3333
rect 4416 3227 4423 3456
rect 4436 3447 4443 3773
rect 4456 3747 4463 3783
rect 4496 3707 4503 3783
rect 4533 3747 4547 3753
rect 4556 3587 4563 3913
rect 4576 3667 4583 3973
rect 4596 3927 4603 4003
rect 4636 3987 4643 4034
rect 4636 3816 4643 3873
rect 4656 3867 4663 4536
rect 4676 4427 4683 4793
rect 4696 4647 4703 4733
rect 4696 4587 4703 4612
rect 4716 4563 4723 4813
rect 4736 4807 4743 4873
rect 4756 4767 4763 4853
rect 4776 4827 4783 4873
rect 4836 4856 4843 4893
rect 4876 4856 4883 4913
rect 4856 4820 4863 4823
rect 4853 4807 4867 4820
rect 4736 4583 4743 4753
rect 4736 4576 4763 4583
rect 4696 4556 4723 4563
rect 4756 4556 4763 4576
rect 4676 4287 4683 4413
rect 4676 4167 4683 4273
rect 4676 3987 4683 4153
rect 4696 4127 4703 4556
rect 4816 4567 4823 4753
rect 4736 4467 4743 4523
rect 4736 4300 4743 4303
rect 4733 4287 4747 4300
rect 4776 4267 4783 4303
rect 4716 4036 4723 4173
rect 4756 4036 4763 4113
rect 4816 4063 4823 4513
rect 4836 4487 4843 4653
rect 4856 4343 4863 4733
rect 4916 4667 4923 5113
rect 4933 5080 4947 5093
rect 4936 5076 4943 5080
rect 4996 5076 5003 5113
rect 4936 4747 4943 5013
rect 4976 4987 4983 5043
rect 4996 4856 5003 4993
rect 5016 4887 5023 5376
rect 5036 5167 5043 5353
rect 5196 5347 5203 5374
rect 5216 5367 5223 5492
rect 5256 5376 5263 5433
rect 5336 5347 5343 5833
rect 5356 5787 5363 5863
rect 5396 5860 5403 5863
rect 5393 5847 5407 5860
rect 5436 5667 5443 5853
rect 5456 5727 5463 6114
rect 5476 6087 5483 6153
rect 5496 6116 5543 6123
rect 5496 5907 5503 6116
rect 5676 6116 5683 6153
rect 5616 6083 5623 6114
rect 5596 6076 5623 6083
rect 5696 6080 5703 6083
rect 5596 6047 5603 6076
rect 5693 6067 5707 6080
rect 5756 6067 5763 6133
rect 5596 5896 5603 6033
rect 5376 5566 5383 5633
rect 5396 5427 5403 5593
rect 5436 5376 5443 5552
rect 5536 5527 5543 5863
rect 5576 5843 5583 5863
rect 5656 5847 5663 6053
rect 5776 6043 5783 6173
rect 5796 6127 5803 6153
rect 5833 6120 5847 6133
rect 5873 6120 5887 6133
rect 5836 6116 5843 6120
rect 5876 6116 5883 6120
rect 5916 6087 5923 6352
rect 6016 6347 6023 6383
rect 5936 6247 5943 6333
rect 6076 6287 6083 6433
rect 6136 6416 6143 6493
rect 6173 6420 6187 6433
rect 6293 6428 6307 6433
rect 6176 6416 6183 6420
rect 6496 6416 6503 6453
rect 6236 6386 6243 6413
rect 6416 6386 6423 6413
rect 6156 6380 6163 6383
rect 6153 6367 6167 6380
rect 6316 6380 6323 6383
rect 6356 6380 6363 6383
rect 6233 6367 6247 6372
rect 6313 6367 6327 6380
rect 6353 6367 6367 6380
rect 5936 6087 5943 6233
rect 5996 6116 6003 6173
rect 6033 6120 6047 6133
rect 6036 6116 6043 6120
rect 5776 6036 5803 6043
rect 5716 5896 5723 5933
rect 5756 5908 5763 5993
rect 5796 5867 5803 6036
rect 5816 6007 5823 6083
rect 5696 5860 5703 5863
rect 5736 5860 5743 5863
rect 5693 5847 5707 5860
rect 5556 5836 5583 5843
rect 5556 5567 5563 5836
rect 5733 5847 5747 5860
rect 5786 5853 5787 5860
rect 5707 5836 5723 5843
rect 5616 5596 5623 5773
rect 5656 5596 5663 5653
rect 5696 5607 5703 5693
rect 5056 5247 5063 5293
rect 5076 5287 5083 5343
rect 5036 4867 5043 5153
rect 5056 4927 5063 5093
rect 5096 5088 5103 5313
rect 5156 5247 5163 5343
rect 5476 5346 5483 5413
rect 5276 5127 5283 5332
rect 5266 5113 5267 5120
rect 5253 5103 5267 5113
rect 5253 5100 5283 5103
rect 5256 5096 5283 5100
rect 5133 5080 5147 5093
rect 5136 5076 5143 5080
rect 5216 5047 5223 5093
rect 5276 5076 5283 5096
rect 5116 4967 5123 5043
rect 5333 5027 5347 5033
rect 5356 5007 5363 5074
rect 5376 5047 5383 5332
rect 5496 5307 5503 5513
rect 5556 5376 5563 5532
rect 5576 5507 5583 5594
rect 5596 5376 5603 5553
rect 5636 5507 5643 5563
rect 5676 5560 5683 5563
rect 5673 5547 5687 5560
rect 5636 5346 5643 5453
rect 5536 5323 5543 5343
rect 5536 5316 5563 5323
rect 5396 5046 5403 5233
rect 5436 5076 5443 5113
rect 5016 4767 5023 4823
rect 5056 4723 5063 4873
rect 5156 4856 5163 4913
rect 5267 4893 5273 4907
rect 5216 4867 5223 4893
rect 5096 4787 5103 4853
rect 5136 4787 5143 4823
rect 5036 4716 5063 4723
rect 4876 4367 4883 4653
rect 4916 4556 4923 4613
rect 4936 4407 4943 4523
rect 4976 4487 4983 4523
rect 4847 4336 4863 4343
rect 4896 4336 4903 4393
rect 4796 4056 4823 4063
rect 4616 3780 4623 3783
rect 4656 3780 4663 3783
rect 4556 3523 4563 3573
rect 4576 3528 4583 3593
rect 4536 3516 4563 3523
rect 4467 3476 4483 3483
rect 4436 3308 4443 3333
rect 4456 3307 4463 3473
rect 4576 3483 4583 3514
rect 4556 3476 4583 3483
rect 4487 3313 4513 3327
rect 4316 3047 4323 3133
rect 4256 2996 4263 3013
rect 4293 3007 4307 3013
rect 4316 2967 4323 2994
rect 4196 2827 4203 2933
rect 4236 2887 4243 2952
rect 4276 2907 4283 2963
rect 4276 2776 4283 2853
rect 4336 2787 4343 3173
rect 4376 3008 4383 3193
rect 4416 2996 4423 3073
rect 4436 3007 4443 3294
rect 4496 3296 4503 3313
rect 4536 3308 4543 3333
rect 4456 2967 4463 3253
rect 4476 3147 4483 3263
rect 4356 2807 4363 2953
rect 4476 2947 4483 3133
rect 4516 3087 4523 3263
rect 4536 3163 4543 3213
rect 4556 3187 4563 3476
rect 4576 3207 4583 3433
rect 4596 3247 4603 3773
rect 4613 3767 4627 3780
rect 4653 3767 4667 3780
rect 4616 3707 4623 3753
rect 4616 3367 4623 3533
rect 4636 3527 4643 3713
rect 4696 3587 4703 3753
rect 4716 3727 4723 3973
rect 4736 3867 4743 4003
rect 4736 3767 4743 3853
rect 4756 3827 4763 3973
rect 4796 3907 4803 4056
rect 4836 4043 4843 4333
rect 4876 4300 4883 4303
rect 4916 4300 4923 4303
rect 4873 4287 4887 4300
rect 4913 4287 4927 4300
rect 4956 4267 4963 4353
rect 4976 4287 4983 4393
rect 4996 4287 5003 4513
rect 5016 4347 5023 4653
rect 5036 4427 5043 4716
rect 5136 4667 5143 4773
rect 5136 4526 5143 4573
rect 5156 4527 5163 4713
rect 5176 4547 5183 4812
rect 5216 4647 5223 4853
rect 5236 4787 5243 4854
rect 5356 4827 5363 4854
rect 5296 4767 5303 4823
rect 5376 4727 5383 4973
rect 5436 4856 5443 4893
rect 5216 4588 5223 4612
rect 5253 4560 5267 4573
rect 5293 4567 5307 4573
rect 5256 4556 5263 4560
rect 5053 4340 5067 4353
rect 5056 4336 5063 4340
rect 5096 4336 5103 4433
rect 5116 4347 5123 4513
rect 5156 4387 5163 4413
rect 5176 4367 5183 4533
rect 5236 4520 5243 4523
rect 5196 4447 5203 4513
rect 5233 4507 5247 4520
rect 5276 4467 5283 4523
rect 4896 4187 4903 4213
rect 4956 4048 4963 4253
rect 5036 4107 5043 4303
rect 5076 4187 5083 4292
rect 4836 4036 4863 4043
rect 4816 3987 4823 4034
rect 4876 4000 4883 4003
rect 4873 3987 4887 4000
rect 4856 3976 4873 3983
rect 4796 3816 4803 3872
rect 4836 3827 4843 3893
rect 4776 3780 4783 3783
rect 4756 3607 4763 3773
rect 4773 3767 4787 3780
rect 4816 3763 4823 3783
rect 4796 3756 4823 3763
rect 4653 3520 4667 3533
rect 4693 3520 4707 3533
rect 4656 3516 4663 3520
rect 4696 3516 4703 3520
rect 4636 3347 4643 3473
rect 4673 3467 4687 3472
rect 4716 3427 4723 3483
rect 4756 3467 4763 3533
rect 4707 3396 4733 3403
rect 4616 3263 4623 3313
rect 4616 3256 4643 3263
rect 4536 3156 4563 3163
rect 4556 3047 4563 3156
rect 4496 2907 4503 2953
rect 4216 2746 4223 2773
rect 4116 2740 4123 2743
rect 4113 2727 4127 2740
rect 4156 2707 4163 2743
rect 4056 2367 4063 2413
rect 4033 2260 4047 2273
rect 4036 2256 4043 2260
rect 3736 1847 3743 1891
rect 3716 1787 3723 1813
rect 3776 1787 3783 1853
rect 3856 1847 3863 1933
rect 3846 1833 3847 1840
rect 3833 1823 3847 1833
rect 3833 1820 3863 1823
rect 3836 1816 3863 1820
rect 3716 1736 3723 1773
rect 3687 1703 3700 1707
rect 3687 1693 3703 1703
rect 3696 1587 3703 1693
rect 3796 1667 3803 1713
rect 3816 1707 3823 1753
rect 3856 1736 3863 1816
rect 3876 1767 3883 2073
rect 3976 1956 3983 2013
rect 3996 2007 4003 2033
rect 4016 1867 4023 2113
rect 3896 1736 3903 1773
rect 3936 1747 3943 1773
rect 4036 1767 4043 2153
rect 4056 2067 4063 2212
rect 4053 2027 4067 2032
rect 4053 2020 4073 2027
rect 4056 2016 4073 2020
rect 4060 2013 4073 2016
rect 4056 1768 4063 1993
rect 4096 1956 4103 2373
rect 4116 2227 4123 2653
rect 4136 2446 4143 2513
rect 4156 2507 4163 2693
rect 4296 2667 4303 2743
rect 4356 2707 4363 2772
rect 4176 2547 4183 2613
rect 4376 2607 4383 2773
rect 4456 2740 4463 2743
rect 4453 2727 4467 2740
rect 4176 2476 4183 2533
rect 4216 2476 4223 2573
rect 4136 2127 4143 2313
rect 4236 2287 4243 2443
rect 4316 2327 4323 2593
rect 4356 2476 4363 2533
rect 4356 2367 4363 2393
rect 4376 2307 4383 2443
rect 4173 2260 4187 2273
rect 4176 2256 4183 2260
rect 4313 2260 4327 2273
rect 4316 2256 4323 2260
rect 4196 2187 4203 2212
rect 4116 1987 4123 2093
rect 4156 2007 4163 2153
rect 4236 2067 4243 2193
rect 4173 1960 4187 1973
rect 4196 1967 4203 2053
rect 4213 1987 4227 1993
rect 4176 1956 4183 1960
rect 4236 1963 4243 2053
rect 4256 1967 4263 2253
rect 4336 2220 4343 2223
rect 4333 2207 4347 2220
rect 4216 1956 4243 1963
rect 4116 1920 4123 1923
rect 4113 1907 4127 1920
rect 4156 1887 4163 1923
rect 3956 1687 3963 1733
rect 3816 1607 3823 1672
rect 3787 1593 3793 1607
rect 3833 1587 3847 1593
rect 3476 1400 3483 1403
rect 3473 1387 3487 1400
rect 3516 1347 3523 1453
rect 3653 1448 3667 1453
rect 3536 1387 3543 1433
rect 3696 1427 3703 1493
rect 3716 1487 3723 1533
rect 3796 1507 3803 1572
rect 3776 1436 3783 1473
rect 3813 1440 3827 1453
rect 3816 1436 3823 1440
rect 3456 1216 3463 1333
rect 3536 1186 3543 1373
rect 3596 1267 3603 1403
rect 3476 1180 3483 1183
rect 3473 1167 3487 1180
rect 3316 916 3323 953
rect 3176 887 3183 914
rect 3076 847 3083 883
rect 3116 880 3123 883
rect 3113 867 3127 880
rect 3136 736 3143 773
rect 3196 747 3203 914
rect 3416 847 3423 1013
rect 3436 867 3443 914
rect 3496 847 3503 883
rect 3536 867 3543 1172
rect 3556 1167 3563 1253
rect 3596 1216 3603 1253
rect 3636 1223 3643 1403
rect 3656 1307 3663 1353
rect 3636 1216 3663 1223
rect 3616 1107 3623 1183
rect 3616 928 3623 1033
rect 3636 943 3643 1073
rect 3656 967 3663 1216
rect 3676 1067 3683 1313
rect 3736 1267 3743 1433
rect 3876 1427 3883 1613
rect 3896 1507 3903 1613
rect 3916 1467 3923 1671
rect 3936 1436 3943 1533
rect 3956 1487 3963 1652
rect 3976 1563 3983 1753
rect 4096 1747 4103 1853
rect 4116 1707 4123 1833
rect 4076 1700 4083 1703
rect 4073 1687 4087 1700
rect 4036 1627 4043 1671
rect 4056 1607 4063 1653
rect 3976 1556 4003 1563
rect 3976 1507 3983 1533
rect 3996 1507 4003 1556
rect 4076 1507 4083 1613
rect 4007 1496 4023 1503
rect 3973 1440 3987 1453
rect 3976 1436 3983 1440
rect 3796 1307 3803 1353
rect 3836 1307 3843 1403
rect 3753 1220 3767 1233
rect 3756 1216 3763 1220
rect 3916 1216 3923 1253
rect 3956 1223 3963 1403
rect 3956 1216 3983 1223
rect 3736 1067 3743 1183
rect 3636 936 3663 943
rect 3656 916 3663 936
rect 3636 807 3643 883
rect 3736 787 3743 953
rect 3756 923 3763 993
rect 3776 987 3783 1183
rect 3816 1027 3823 1093
rect 3756 916 3783 923
rect 3816 916 3823 1013
rect 3836 967 3843 1213
rect 3976 1186 3983 1216
rect 3896 1180 3903 1183
rect 3893 1167 3907 1180
rect 3976 1127 3983 1172
rect 3947 1113 3953 1127
rect 3996 1087 4003 1313
rect 4016 1167 4023 1496
rect 4096 1463 4103 1693
rect 4136 1683 4143 1713
rect 4087 1456 4103 1463
rect 4116 1676 4143 1683
rect 4073 1440 4087 1453
rect 4116 1448 4123 1676
rect 4136 1487 4143 1533
rect 4076 1436 4083 1440
rect 4036 1327 4043 1434
rect 4096 1400 4103 1403
rect 4033 1227 4047 1233
rect 4056 1216 4063 1393
rect 4093 1387 4107 1400
rect 4136 1227 4143 1293
rect 4076 1180 4083 1183
rect 4073 1167 4087 1180
rect 4013 1107 4027 1113
rect 4116 1027 4123 1183
rect 3793 867 3807 872
rect 3076 703 3083 733
rect 3076 696 3103 703
rect 3213 663 3227 673
rect 3196 660 3227 663
rect 3196 656 3223 660
rect 3256 627 3263 694
rect 3356 647 3363 673
rect 3376 667 3383 694
rect 3436 660 3443 663
rect 3433 647 3447 660
rect 3116 527 3123 573
rect 3036 407 3043 493
rect 3076 427 3083 453
rect 3073 400 3087 413
rect 3076 396 3083 400
rect 3116 396 3123 513
rect 3056 327 3063 363
rect 3093 347 3107 352
rect 3156 347 3163 613
rect 3256 487 3263 613
rect 3496 487 3503 694
rect 3516 666 3523 733
rect 3716 727 3723 753
rect 3716 696 3723 713
rect 3756 707 3763 813
rect 3616 627 3623 663
rect 3676 627 3683 693
rect 3776 647 3783 773
rect 3816 747 3823 773
rect 3836 727 3843 883
rect 3876 787 3883 953
rect 3936 916 3943 1013
rect 3976 916 3983 993
rect 4136 947 4143 1173
rect 4156 1147 4163 1793
rect 4216 1736 4223 1956
rect 4296 1956 4303 2173
rect 4376 2167 4383 2213
rect 4396 2147 4403 2393
rect 4416 2367 4423 2443
rect 4456 2268 4463 2692
rect 4476 2587 4483 2733
rect 4496 2707 4503 2893
rect 4516 2727 4523 2933
rect 4576 2776 4583 2833
rect 4596 2807 4603 3073
rect 4616 3047 4623 3113
rect 4616 2967 4623 2994
rect 4616 2788 4623 2932
rect 4636 2867 4643 3233
rect 4696 3207 4703 3263
rect 4716 3183 4723 3313
rect 4776 3308 4783 3653
rect 4796 3527 4803 3756
rect 4836 3607 4843 3773
rect 4856 3727 4863 3976
rect 4916 3947 4923 4003
rect 4876 3627 4883 3893
rect 4936 3863 4943 3973
rect 4956 3907 4963 4034
rect 4976 3927 4983 4053
rect 5033 4040 5047 4053
rect 5036 4036 5043 4040
rect 5076 4036 5083 4093
rect 5136 4007 5143 4353
rect 5233 4348 5247 4353
rect 5156 4247 5163 4333
rect 5216 4300 5223 4303
rect 5213 4287 5227 4300
rect 5216 4067 5223 4233
rect 5256 4107 5263 4292
rect 5296 4267 5303 4334
rect 5316 4307 5323 4633
rect 5413 4560 5427 4573
rect 5416 4556 5423 4560
rect 5336 4507 5343 4554
rect 5396 4520 5403 4523
rect 5393 4507 5407 4520
rect 5436 4427 5443 4523
rect 5476 4507 5483 4573
rect 5496 4507 5503 4813
rect 5516 4587 5523 4873
rect 5536 4587 5543 5293
rect 5556 4867 5563 5316
rect 5656 5207 5663 5393
rect 5676 5147 5683 5413
rect 5716 5407 5723 5836
rect 5773 5843 5787 5853
rect 5756 5840 5787 5843
rect 5756 5836 5783 5840
rect 5736 5507 5743 5613
rect 5756 5607 5763 5836
rect 5816 5647 5823 5894
rect 5936 5787 5943 5933
rect 5956 5767 5963 5973
rect 6016 5896 6023 6072
rect 6076 5908 6083 6133
rect 6096 6027 6103 6173
rect 6116 5903 6123 6273
rect 6220 6145 6233 6147
rect 6167 6138 6233 6145
rect 6216 6133 6233 6138
rect 6216 6116 6223 6133
rect 6196 6047 6203 6083
rect 6096 5896 6123 5903
rect 6156 5896 6163 6033
rect 5793 5600 5807 5613
rect 5796 5596 5803 5600
rect 5816 5543 5823 5552
rect 5796 5536 5823 5543
rect 5736 5376 5743 5413
rect 5796 5388 5803 5536
rect 5696 5336 5723 5343
rect 5696 5307 5703 5336
rect 5796 5307 5803 5374
rect 5696 5267 5703 5293
rect 5593 5080 5607 5093
rect 5727 5093 5733 5107
rect 5633 5088 5647 5093
rect 5596 5076 5603 5080
rect 5696 5046 5703 5093
rect 5716 5076 5743 5083
rect 5793 5080 5807 5093
rect 5796 5076 5803 5080
rect 5616 4888 5623 5043
rect 5716 4927 5723 5076
rect 5816 5023 5823 5493
rect 5836 5387 5843 5533
rect 5856 5427 5863 5553
rect 5876 5547 5883 5753
rect 5996 5647 6003 5863
rect 6036 5843 6043 5852
rect 6016 5836 6043 5843
rect 5916 5607 5923 5633
rect 5896 5467 5903 5594
rect 5973 5600 5987 5613
rect 6016 5607 6023 5836
rect 5976 5596 5983 5600
rect 5956 5347 5963 5453
rect 5796 5016 5823 5023
rect 5640 4823 5653 4827
rect 5596 4820 5603 4823
rect 5593 4807 5607 4820
rect 5636 4816 5653 4823
rect 5640 4813 5653 4816
rect 5676 4826 5683 4913
rect 5716 4827 5723 4913
rect 5753 4860 5767 4873
rect 5756 4856 5763 4860
rect 5796 4856 5803 5016
rect 5836 4867 5843 5333
rect 5776 4803 5783 4823
rect 5756 4796 5783 4803
rect 5556 4556 5563 4793
rect 5416 4336 5423 4373
rect 5396 4300 5403 4303
rect 5393 4287 5407 4300
rect 5213 4040 5227 4053
rect 5216 4036 5223 4040
rect 4996 3996 5023 4003
rect 4996 3967 5003 3996
rect 4996 3867 5003 3953
rect 4936 3856 4963 3863
rect 4956 3816 4963 3856
rect 4993 3827 5007 3832
rect 5016 3786 5023 3873
rect 4936 3647 4943 3783
rect 5036 3647 5043 3814
rect 4813 3520 4827 3533
rect 4853 3520 4867 3533
rect 4816 3516 4823 3520
rect 4856 3516 4863 3520
rect 4696 3176 4723 3183
rect 4656 3027 4663 3093
rect 4676 2996 4683 3113
rect 4696 3027 4703 3176
rect 4713 3047 4727 3053
rect 4756 3007 4763 3273
rect 4696 2887 4703 2963
rect 4696 2747 4703 2852
rect 4516 2476 4523 2533
rect 4536 2507 4543 2733
rect 4556 2707 4563 2743
rect 4576 2527 4583 2713
rect 4596 2567 4603 2743
rect 4636 2723 4643 2743
rect 4716 2727 4723 2933
rect 4776 2847 4783 3294
rect 4796 3263 4803 3473
rect 4836 3367 4843 3483
rect 4876 3480 4883 3483
rect 4873 3467 4887 3480
rect 4796 3256 4823 3263
rect 4876 3260 4883 3263
rect 4816 3103 4823 3256
rect 4873 3247 4887 3260
rect 4887 3193 4893 3207
rect 4816 3096 4843 3103
rect 4796 2963 4803 3053
rect 4816 3007 4823 3073
rect 4836 2996 4843 3096
rect 4856 3027 4863 3073
rect 4916 3027 4923 3613
rect 4936 3486 4943 3533
rect 4996 3516 5003 3633
rect 5036 3447 5043 3593
rect 5056 3587 5063 3773
rect 5076 3727 5083 3783
rect 5056 3487 5063 3573
rect 5096 3567 5103 3753
rect 5176 3667 5183 3973
rect 5196 3786 5203 4003
rect 5256 3987 5263 4053
rect 5296 4003 5303 4232
rect 5296 3996 5323 4003
rect 5276 3816 5283 3873
rect 5216 3783 5223 3813
rect 5316 3783 5323 3996
rect 5336 3967 5343 4003
rect 5396 3987 5403 4252
rect 5416 4006 5423 4033
rect 5436 4003 5443 4293
rect 5456 4247 5463 4493
rect 5516 4483 5523 4513
rect 5573 4503 5587 4512
rect 5556 4500 5587 4503
rect 5556 4496 5583 4500
rect 5556 4483 5563 4496
rect 5496 4476 5523 4483
rect 5536 4476 5563 4483
rect 5476 4306 5483 4413
rect 5496 4347 5503 4476
rect 5536 4467 5543 4476
rect 5527 4456 5543 4467
rect 5527 4453 5540 4456
rect 5536 4336 5543 4433
rect 5576 4336 5583 4473
rect 5596 4387 5603 4633
rect 5636 4563 5643 4793
rect 5756 4767 5763 4796
rect 5856 4787 5863 5293
rect 5896 5087 5903 5332
rect 5976 5307 5983 5493
rect 6016 5467 6023 5553
rect 6036 5507 6043 5793
rect 6076 5607 6083 5894
rect 6096 5807 6103 5896
rect 6236 5907 6243 6073
rect 6136 5827 6143 5863
rect 6136 5707 6143 5813
rect 6116 5608 6123 5633
rect 6176 5607 6183 5863
rect 6256 5827 6263 6113
rect 6296 5987 6303 6213
rect 6436 6187 6443 6413
rect 6516 6363 6523 6383
rect 6516 6356 6543 6363
rect 6313 6123 6327 6133
rect 6313 6120 6343 6123
rect 6373 6120 6387 6133
rect 6316 6116 6343 6120
rect 6376 6116 6383 6120
rect 6396 5927 6403 6083
rect 6456 6067 6463 6153
rect 6536 6147 6543 6356
rect 6576 6167 6583 6413
rect 6616 6287 6623 6473
rect 6696 6416 6703 6473
rect 6636 6227 6643 6372
rect 6716 6307 6723 6383
rect 6553 6120 6567 6133
rect 6556 6116 6563 6120
rect 6353 5900 6367 5913
rect 6393 5907 6407 5913
rect 6356 5896 6363 5900
rect 6276 5627 6283 5893
rect 6296 5607 6303 5852
rect 6076 5388 6083 5553
rect 6096 5447 6103 5563
rect 6136 5487 6143 5563
rect 6196 5507 6203 5594
rect 6316 5596 6323 5633
rect 6347 5613 6353 5627
rect 6376 5596 6383 5653
rect 6416 5643 6423 6053
rect 6496 6047 6503 6083
rect 6456 5907 6463 6032
rect 6493 5908 6507 5913
rect 6536 5896 6543 6033
rect 6396 5636 6423 5643
rect 6236 5547 6243 5593
rect 6396 5587 6403 5636
rect 6276 5560 6283 5563
rect 6273 5547 6287 5560
rect 6236 5447 6243 5533
rect 6236 5376 6243 5433
rect 6116 5346 6123 5373
rect 6016 5323 6023 5343
rect 6016 5316 6043 5323
rect 5933 5080 5947 5093
rect 5936 5076 5943 5080
rect 5956 5023 5963 5043
rect 5936 5016 5963 5023
rect 5936 4868 5943 5016
rect 5996 4923 6003 5033
rect 6016 4987 6023 5093
rect 6036 5047 6043 5316
rect 6056 5207 6063 5343
rect 6096 5076 6103 5133
rect 6136 5108 6143 5373
rect 6176 5287 6183 5343
rect 6176 5087 6183 5273
rect 5996 4916 6013 4923
rect 5773 4723 5787 4733
rect 5756 4720 5787 4723
rect 5756 4716 5783 4720
rect 5616 4556 5663 4563
rect 5616 4348 5623 4556
rect 5756 4527 5763 4716
rect 5796 4567 5803 4713
rect 5876 4647 5883 4854
rect 6016 4826 6023 4913
rect 5720 4523 5733 4527
rect 5676 4427 5683 4523
rect 5716 4516 5733 4523
rect 5720 4513 5733 4516
rect 5776 4443 5783 4554
rect 5836 4556 5843 4593
rect 5896 4567 5903 4813
rect 5816 4467 5823 4512
rect 5776 4436 5793 4443
rect 5656 4416 5673 4423
rect 5616 4306 5623 4334
rect 5636 4247 5643 4393
rect 5656 4306 5663 4416
rect 5476 4036 5483 4093
rect 5516 4036 5523 4133
rect 5616 4043 5623 4093
rect 5596 4036 5623 4043
rect 5636 4036 5643 4133
rect 5596 4006 5603 4036
rect 5436 3996 5463 4003
rect 5456 3816 5463 3996
rect 5536 4000 5543 4003
rect 5533 3987 5547 4000
rect 5216 3776 5243 3783
rect 5296 3776 5323 3783
rect 5236 3707 5243 3776
rect 5476 3707 5483 3783
rect 5496 3747 5503 3772
rect 5207 3533 5213 3547
rect 5133 3528 5147 3533
rect 5176 3516 5223 3523
rect 5076 3467 5083 3514
rect 5107 3483 5120 3487
rect 5107 3476 5123 3483
rect 5107 3473 5120 3476
rect 4936 2967 4943 3353
rect 4956 3227 4963 3433
rect 5216 3407 5223 3516
rect 5236 3487 5243 3613
rect 5256 3527 5263 3573
rect 5336 3567 5343 3593
rect 5293 3520 5307 3533
rect 5296 3516 5303 3520
rect 5196 3347 5203 3373
rect 5036 3227 5043 3263
rect 5076 3247 5083 3273
rect 5096 3223 5103 3294
rect 5196 3263 5203 3333
rect 5296 3296 5303 3453
rect 5316 3447 5323 3483
rect 5376 3447 5383 3553
rect 5436 3516 5443 3693
rect 5516 3527 5523 3814
rect 5536 3727 5543 3973
rect 5573 3820 5587 3833
rect 5576 3816 5583 3820
rect 5636 3747 5643 3783
rect 5396 3407 5403 3514
rect 5456 3427 5463 3472
rect 5496 3427 5503 3483
rect 5356 3263 5363 3294
rect 5376 3266 5383 3333
rect 5476 3296 5483 3333
rect 5156 3256 5203 3263
rect 5076 3216 5103 3223
rect 5007 3196 5053 3203
rect 5076 3127 5083 3216
rect 5276 3207 5283 3263
rect 5316 3260 5323 3263
rect 5313 3247 5327 3260
rect 5336 3256 5363 3263
rect 4993 3000 5007 3013
rect 4996 2996 5003 3000
rect 5036 2996 5043 3053
rect 4796 2956 4823 2963
rect 4816 2743 4823 2956
rect 4896 2943 4903 2963
rect 4956 2963 4963 2994
rect 5076 2967 5083 3113
rect 5136 2996 5143 3033
rect 4956 2956 4983 2963
rect 4616 2716 4643 2723
rect 4616 2627 4623 2716
rect 4553 2480 4567 2493
rect 4556 2476 4563 2480
rect 4476 2427 4483 2473
rect 4496 2287 4503 2433
rect 4493 2268 4507 2273
rect 4316 2027 4323 2073
rect 4416 1983 4423 2253
rect 4416 1976 4443 1983
rect 4333 1960 4347 1973
rect 4336 1956 4343 1960
rect 4196 1700 4203 1703
rect 4193 1687 4207 1700
rect 4236 1567 4243 1703
rect 4276 1667 4283 1923
rect 4396 1923 4403 1973
rect 4176 1403 4183 1453
rect 4196 1447 4203 1533
rect 4236 1436 4243 1493
rect 4276 1436 4283 1493
rect 4296 1467 4303 1893
rect 4176 1396 4203 1403
rect 4176 947 4183 1273
rect 4056 916 4103 923
rect 4136 916 4143 933
rect 3873 727 3887 733
rect 3796 666 3803 713
rect 3873 700 3887 713
rect 3876 696 3883 700
rect 2996 176 3023 183
rect 3056 176 3063 213
rect 2596 -17 2603 143
rect 2756 -17 2763 143
rect 2896 87 2903 143
rect 2996 -17 3003 176
rect 3196 176 3203 473
rect 3276 396 3283 453
rect 3396 396 3403 453
rect 3316 367 3323 394
rect 3516 387 3523 513
rect 3596 396 3603 473
rect 3816 408 3823 693
rect 3856 660 3863 663
rect 3853 647 3867 660
rect 3956 643 3963 833
rect 3996 827 4003 883
rect 4036 867 4043 913
rect 3976 787 3983 813
rect 4036 708 4043 733
rect 4056 727 4063 916
rect 4116 767 4123 883
rect 4156 827 4163 883
rect 4196 867 4203 1396
rect 4216 1223 4223 1403
rect 4316 1367 4323 1813
rect 4356 1807 4363 1923
rect 4376 1916 4403 1923
rect 4376 1736 4383 1916
rect 4396 1807 4403 1853
rect 4416 1747 4423 1953
rect 4356 1667 4363 1703
rect 4396 1607 4403 1703
rect 4416 1647 4423 1693
rect 4436 1687 4443 1976
rect 4456 1967 4463 2193
rect 4476 2187 4483 2223
rect 4493 2207 4507 2213
rect 4476 2087 4483 2173
rect 4473 1960 4487 1973
rect 4476 1956 4483 1960
rect 4516 1956 4523 2373
rect 4536 2307 4543 2443
rect 4536 2087 4543 2272
rect 4556 2187 4563 2413
rect 4576 2287 4583 2443
rect 4596 2327 4603 2353
rect 4616 2307 4623 2513
rect 4636 2443 4643 2693
rect 4696 2476 4703 2513
rect 4636 2436 4663 2443
rect 4636 2287 4643 2353
rect 4556 1963 4563 2152
rect 4576 2127 4583 2223
rect 4636 2220 4643 2223
rect 4633 2207 4647 2220
rect 4656 2167 4663 2436
rect 4676 2347 4683 2443
rect 4576 1987 4583 2113
rect 4556 1956 4583 1963
rect 4540 1924 4553 1927
rect 4536 1917 4553 1924
rect 4540 1913 4553 1917
rect 4540 1906 4560 1907
rect 4540 1903 4553 1906
rect 4536 1893 4553 1903
rect 4456 1667 4463 1733
rect 4476 1627 4483 1873
rect 4536 1827 4543 1893
rect 4576 1887 4583 1956
rect 4596 1927 4603 1993
rect 4616 1967 4623 2033
rect 4656 2007 4663 2132
rect 4676 1987 4683 2273
rect 4696 2207 4703 2373
rect 4716 2247 4723 2411
rect 4756 2387 4763 2713
rect 4776 2687 4783 2743
rect 4796 2736 4823 2743
rect 4876 2936 4903 2943
rect 4776 2446 4783 2673
rect 4796 2427 4803 2736
rect 4876 2727 4883 2936
rect 4916 2867 4923 2953
rect 4976 2927 4983 2956
rect 4896 2667 4903 2743
rect 4856 2476 4863 2593
rect 4896 2476 4903 2653
rect 4816 2407 4823 2433
rect 4776 2256 4783 2353
rect 4756 2220 4763 2223
rect 4653 1960 4667 1972
rect 4696 1967 4703 1993
rect 4656 1956 4663 1960
rect 4636 1887 4643 1923
rect 4536 1736 4543 1813
rect 4576 1706 4583 1833
rect 4336 1387 4343 1513
rect 4356 1347 4363 1593
rect 4456 1436 4463 1513
rect 4496 1407 4503 1593
rect 4216 1216 4233 1223
rect 4276 1216 4283 1253
rect 4336 1247 4343 1273
rect 4256 1180 4263 1183
rect 4296 1180 4303 1183
rect 4253 1167 4267 1180
rect 4293 1167 4307 1180
rect 4296 1067 4303 1153
rect 4336 1107 4343 1173
rect 4356 1067 4363 1253
rect 4376 1228 4383 1353
rect 4396 1327 4403 1403
rect 4493 1387 4507 1393
rect 4373 1207 4387 1214
rect 4396 1183 4403 1273
rect 4456 1247 4463 1353
rect 4516 1267 4523 1671
rect 4576 1567 4583 1692
rect 4496 1256 4513 1263
rect 4456 1216 4463 1233
rect 4496 1207 4503 1256
rect 4536 1228 4543 1513
rect 4596 1448 4603 1813
rect 4676 1803 4683 1912
rect 4696 1827 4703 1913
rect 4676 1796 4703 1803
rect 4636 1547 4643 1703
rect 4676 1667 4683 1693
rect 4656 1607 4663 1653
rect 4696 1587 4703 1796
rect 4716 1687 4723 2212
rect 4753 2207 4767 2220
rect 4793 2187 4807 2191
rect 4836 2187 4843 2443
rect 4876 2387 4883 2443
rect 4856 2127 4863 2293
rect 4916 2256 4923 2313
rect 4936 2287 4943 2713
rect 4956 2663 4963 2732
rect 4976 2687 4983 2913
rect 5096 2847 5103 2994
rect 5216 2947 5223 3033
rect 5256 2967 5263 3013
rect 5316 2996 5323 3153
rect 5336 3087 5343 3256
rect 5456 3260 5463 3263
rect 5453 3247 5467 3260
rect 5516 3167 5523 3473
rect 5536 3087 5543 3633
rect 5556 3407 5563 3593
rect 5596 3516 5603 3693
rect 5636 3647 5643 3733
rect 5676 3527 5683 3973
rect 5696 3847 5703 4003
rect 5736 3967 5743 4153
rect 5756 3907 5763 4273
rect 5776 4047 5783 4293
rect 5796 4287 5803 4433
rect 5836 4347 5843 4493
rect 5856 4387 5863 4523
rect 5916 4503 5923 4773
rect 5936 4523 5943 4793
rect 6036 4647 6043 4853
rect 6056 4747 6063 5053
rect 6136 4856 6143 4993
rect 6156 4987 6163 5043
rect 6196 5046 6203 5093
rect 6176 5007 6183 5033
rect 6176 4887 6183 4933
rect 6216 4907 6223 5153
rect 6116 4727 6123 4823
rect 5996 4607 6003 4633
rect 5996 4556 6003 4593
rect 6156 4587 6163 4823
rect 6216 4667 6223 4872
rect 6236 4867 6243 5313
rect 6256 5127 6263 5333
rect 6276 5327 6283 5493
rect 6296 5347 6303 5413
rect 6316 5387 6323 5533
rect 6336 5507 6343 5563
rect 6376 5407 6383 5513
rect 6373 5388 6387 5393
rect 6376 5287 6383 5333
rect 6256 5083 6263 5113
rect 6376 5088 6383 5273
rect 6256 5076 6283 5083
rect 6376 5043 6383 5074
rect 6293 5027 6307 5032
rect 6336 5007 6343 5043
rect 6356 5036 6383 5043
rect 6356 4983 6363 5036
rect 6336 4976 6363 4983
rect 6336 4947 6343 4976
rect 6256 4856 6263 4913
rect 6333 4887 6347 4893
rect 6236 4607 6243 4813
rect 6256 4687 6263 4793
rect 6276 4767 6283 4823
rect 6276 4707 6283 4753
rect 6316 4747 6323 4823
rect 6356 4787 6363 4953
rect 6376 4707 6383 4913
rect 6396 4907 6403 5552
rect 6416 5527 6423 5613
rect 6436 5503 6443 5793
rect 6416 5496 6443 5503
rect 6416 5307 6423 5496
rect 6456 5427 6463 5853
rect 6476 5787 6483 5863
rect 6516 5807 6523 5863
rect 6556 5767 6563 5853
rect 6576 5767 6583 6013
rect 6596 5863 6603 6113
rect 6616 6027 6623 6133
rect 6713 6120 6727 6133
rect 6716 6116 6723 6120
rect 6636 6067 6643 6114
rect 6696 6063 6703 6083
rect 6736 6076 6763 6083
rect 6696 6056 6723 6063
rect 6696 5896 6703 6013
rect 6716 5907 6723 6056
rect 6736 5863 6743 6053
rect 6756 5883 6763 6076
rect 6776 5907 6783 6293
rect 6756 5876 6783 5883
rect 6596 5856 6623 5863
rect 6476 5527 6483 5752
rect 6496 5607 6503 5653
rect 6527 5614 6533 5627
rect 6520 5613 6540 5614
rect 6573 5600 6587 5613
rect 6596 5607 6603 5713
rect 6576 5596 6583 5600
rect 6616 5567 6623 5856
rect 6636 5807 6643 5863
rect 6676 5787 6683 5863
rect 6736 5856 6763 5863
rect 6496 5463 6503 5553
rect 6516 5547 6523 5563
rect 6516 5536 6533 5547
rect 6520 5533 6533 5536
rect 6556 5487 6563 5563
rect 6496 5456 6523 5463
rect 6460 5403 6473 5407
rect 6456 5393 6473 5403
rect 6456 5376 6463 5393
rect 6496 5376 6503 5433
rect 6516 5407 6523 5456
rect 6416 4927 6423 5173
rect 6456 5076 6463 5113
rect 6476 5103 6483 5332
rect 6496 5187 6503 5313
rect 6536 5143 6543 5313
rect 6556 5167 6563 5393
rect 6536 5136 6563 5143
rect 6476 5096 6503 5103
rect 6496 5076 6503 5096
rect 6476 5040 6483 5043
rect 6473 5027 6487 5040
rect 6516 5007 6523 5043
rect 6436 4887 6443 4993
rect 6556 4967 6563 5136
rect 6413 4860 6427 4873
rect 6416 4856 6423 4860
rect 6496 4856 6503 4953
rect 6516 4867 6523 4913
rect 6476 4803 6483 4823
rect 6476 4796 6503 4803
rect 6256 4583 6263 4652
rect 6376 4627 6383 4693
rect 6436 4607 6443 4713
rect 6456 4627 6463 4773
rect 6236 4576 6263 4583
rect 6033 4560 6047 4573
rect 6036 4556 6043 4560
rect 6076 4523 6083 4573
rect 5936 4516 5963 4523
rect 5916 4496 5943 4503
rect 5936 4407 5943 4496
rect 5936 4347 5943 4372
rect 5813 4327 5827 4333
rect 5816 4127 5823 4292
rect 5796 4036 5803 4073
rect 5836 4068 5843 4293
rect 5856 4227 5863 4303
rect 5896 4287 5903 4303
rect 5733 3820 5747 3833
rect 5736 3816 5743 3820
rect 5816 3827 5823 3953
rect 5656 3387 5663 3483
rect 5640 3263 5653 3267
rect 5596 3207 5603 3263
rect 5636 3256 5653 3263
rect 5640 3253 5653 3256
rect 5676 3247 5683 3473
rect 5596 3107 5603 3193
rect 5496 2996 5503 3033
rect 5096 2776 5103 2833
rect 4956 2656 4983 2663
rect 4956 2427 4963 2513
rect 4976 2487 4983 2656
rect 5056 2627 5063 2743
rect 5056 2476 5103 2483
rect 4996 2423 5003 2443
rect 4996 2416 5023 2423
rect 4896 2220 4903 2223
rect 4893 2207 4907 2220
rect 4876 2196 4893 2203
rect 4836 2067 4843 2093
rect 4856 2007 4863 2113
rect 4736 1887 4743 1954
rect 4736 1747 4743 1873
rect 4756 1867 4763 1973
rect 4853 1960 4867 1972
rect 4876 1967 4883 2196
rect 4856 1956 4863 1960
rect 4776 1887 4783 1913
rect 4896 1923 4903 2172
rect 4916 2067 4923 2153
rect 4976 2103 4983 2273
rect 4956 2096 4983 2103
rect 4956 2003 4963 2096
rect 4913 1987 4927 1993
rect 4936 1996 4963 2003
rect 4936 1967 4943 1996
rect 4976 1987 4983 2053
rect 4976 1956 4983 1973
rect 4996 1967 5003 2393
rect 5016 2267 5023 2416
rect 5036 2407 5043 2443
rect 5036 2256 5043 2313
rect 5076 2267 5083 2433
rect 5016 2107 5023 2213
rect 5056 2147 5063 2223
rect 5016 1967 5023 2093
rect 5096 2087 5103 2476
rect 5116 2387 5123 2432
rect 5136 2383 5143 2853
rect 5176 2627 5183 2933
rect 5236 2776 5243 2833
rect 5176 2476 5183 2513
rect 5216 2476 5223 2732
rect 5256 2667 5263 2743
rect 5296 2667 5303 2963
rect 5396 2927 5403 2973
rect 5556 2966 5563 3033
rect 5616 2996 5623 3153
rect 5636 3147 5643 3233
rect 5696 3047 5703 3793
rect 5796 3707 5803 3783
rect 5836 3567 5843 3813
rect 5796 3516 5803 3553
rect 5716 3247 5723 3514
rect 5820 3484 5833 3487
rect 5776 3427 5783 3483
rect 5816 3477 5833 3484
rect 5820 3473 5833 3477
rect 5796 3387 5803 3433
rect 5816 3347 5823 3393
rect 5836 3347 5843 3452
rect 5856 3447 5863 3893
rect 5876 3487 5883 4073
rect 5896 4047 5903 4273
rect 5936 4227 5943 4293
rect 5956 4287 5963 4516
rect 5976 4467 5983 4523
rect 5936 4068 5943 4213
rect 5976 4167 5983 4393
rect 6016 4387 6023 4523
rect 6056 4516 6083 4523
rect 6036 4336 6043 4393
rect 6056 4367 6063 4516
rect 6096 4503 6103 4553
rect 6096 4496 6143 4503
rect 6076 4336 6083 4373
rect 6116 4347 6123 4473
rect 6136 4463 6143 4496
rect 6156 4487 6163 4512
rect 6176 4463 6183 4513
rect 6136 4456 6183 4463
rect 6196 4447 6203 4554
rect 6216 4527 6223 4573
rect 6236 4547 6243 4576
rect 6313 4560 6327 4573
rect 6316 4556 6323 4560
rect 6340 4523 6353 4527
rect 6233 4503 6247 4512
rect 6216 4500 6247 4503
rect 6216 4496 6243 4500
rect 5996 4207 6003 4333
rect 6056 4300 6063 4303
rect 6053 4287 6067 4300
rect 6136 4283 6143 4433
rect 6216 4423 6223 4496
rect 6196 4416 6223 4423
rect 6127 4276 6143 4283
rect 5973 4040 5987 4053
rect 5976 4036 5983 4040
rect 5896 4007 5903 4033
rect 5956 4000 5963 4003
rect 5913 3987 5927 3993
rect 5953 3987 5967 4000
rect 5996 3996 6023 4003
rect 5936 3816 5943 3853
rect 5996 3787 6003 3973
rect 6016 3927 6023 3996
rect 6036 3987 6043 4013
rect 6056 3887 6063 4252
rect 6076 3947 6083 4213
rect 6096 3983 6103 4113
rect 6116 4036 6123 4273
rect 6156 4107 6163 4393
rect 6196 4367 6203 4416
rect 6216 4336 6223 4373
rect 6236 4367 6243 4393
rect 6296 4387 6303 4523
rect 6336 4516 6353 4523
rect 6340 4513 6353 4516
rect 6176 4267 6183 4293
rect 6236 4300 6243 4303
rect 6233 4287 6247 4300
rect 6176 4036 6183 4073
rect 6136 4000 6143 4003
rect 6133 3987 6147 4000
rect 6096 3976 6123 3983
rect 5896 3527 5903 3773
rect 5916 3547 5923 3772
rect 5936 3516 5943 3593
rect 5956 3547 5963 3783
rect 6016 3783 6023 3873
rect 6016 3776 6043 3783
rect 6036 3547 6043 3776
rect 6056 3707 6063 3783
rect 6096 3747 6103 3773
rect 6056 3607 6063 3693
rect 6116 3687 6123 3976
rect 6196 3967 6203 4093
rect 6136 3767 6143 3933
rect 6156 3827 6163 3913
rect 6196 3816 6203 3953
rect 6216 3867 6223 4173
rect 6256 4107 6263 4273
rect 6276 4187 6283 4293
rect 6296 4283 6303 4333
rect 6316 4307 6323 4493
rect 6296 4276 6323 4283
rect 6293 4247 6307 4253
rect 6316 4068 6323 4276
rect 6336 4267 6343 4433
rect 6356 4347 6363 4453
rect 6376 4407 6383 4592
rect 6396 4547 6403 4593
rect 6456 4556 6463 4613
rect 6496 4527 6503 4796
rect 6396 4447 6403 4512
rect 6396 4336 6403 4433
rect 6436 4427 6443 4523
rect 6476 4427 6483 4493
rect 6440 4404 6453 4407
rect 6436 4393 6453 4404
rect 6436 4367 6443 4393
rect 6433 4340 6447 4353
rect 6456 4347 6463 4372
rect 6436 4336 6443 4340
rect 6376 4300 6383 4303
rect 6356 4267 6363 4293
rect 6373 4287 6387 4300
rect 6416 4283 6423 4303
rect 6416 4276 6443 4283
rect 6396 4243 6403 4273
rect 6333 4227 6347 4232
rect 6376 4236 6403 4243
rect 6236 3867 6243 4053
rect 6376 4007 6383 4236
rect 6256 3927 6263 3993
rect 6296 3983 6303 4003
rect 6276 3980 6303 3983
rect 6273 3976 6303 3980
rect 6273 3967 6287 3976
rect 6286 3960 6287 3967
rect 6216 3767 6223 3783
rect 6216 3727 6223 3753
rect 6256 3743 6263 3773
rect 6236 3736 6263 3743
rect 6096 3516 6103 3593
rect 5953 3467 5967 3472
rect 5736 3267 5743 3333
rect 5796 3316 5843 3323
rect 5796 3296 5803 3316
rect 5747 3256 5763 3263
rect 5436 2907 5443 2963
rect 5416 2776 5423 2893
rect 5476 2867 5483 2963
rect 5696 2887 5703 2994
rect 5736 2887 5743 3232
rect 5447 2783 5460 2787
rect 5447 2773 5463 2783
rect 5396 2687 5403 2743
rect 5256 2447 5263 2613
rect 5276 2447 5283 2513
rect 5316 2476 5323 2573
rect 5136 2376 5163 2383
rect 5116 2167 5123 2253
rect 5136 2226 5143 2353
rect 5156 2267 5163 2376
rect 5196 2367 5203 2443
rect 5216 2343 5223 2373
rect 5196 2336 5223 2343
rect 5196 2256 5203 2336
rect 5236 2268 5243 2313
rect 4653 1507 4667 1513
rect 4716 1507 4723 1673
rect 4733 1667 4747 1673
rect 4666 1500 4667 1507
rect 4633 1440 4647 1453
rect 4636 1436 4643 1440
rect 4567 1403 4580 1407
rect 4567 1396 4583 1403
rect 4567 1393 4580 1396
rect 4676 1367 4683 1493
rect 4727 1453 4733 1467
rect 4756 1436 4763 1573
rect 4816 1507 4823 1873
rect 4836 1807 4843 1923
rect 4876 1916 4903 1923
rect 4876 1903 4883 1916
rect 4856 1896 4883 1903
rect 4396 1176 4423 1183
rect 4373 1167 4387 1172
rect 4376 1047 4383 1132
rect 4273 920 4287 933
rect 4276 916 4283 920
rect 4336 927 4343 973
rect 4216 883 4223 914
rect 4416 916 4423 1073
rect 4476 1027 4483 1183
rect 4596 1107 4603 1183
rect 4636 1027 4643 1313
rect 4696 1307 4703 1433
rect 4776 1400 4783 1403
rect 4773 1387 4787 1400
rect 4836 1367 4843 1734
rect 4856 1567 4863 1896
rect 4896 1736 4903 1873
rect 4916 1767 4923 1952
rect 4876 1687 4883 1703
rect 4876 1523 4883 1673
rect 4956 1627 4963 1912
rect 4976 1706 4983 1893
rect 4976 1567 4983 1692
rect 4856 1516 4883 1523
rect 4856 1443 4863 1516
rect 4856 1436 4883 1443
rect 4656 1186 4663 1293
rect 4696 1216 4703 1253
rect 4896 1247 4903 1403
rect 4956 1287 4963 1453
rect 4756 1180 4763 1183
rect 4753 1167 4767 1180
rect 4476 967 4483 1013
rect 4636 916 4643 953
rect 4216 876 4243 883
rect 4156 707 4163 773
rect 4080 703 4093 707
rect 4076 696 4093 703
rect 4080 693 4093 696
rect 4196 696 4203 832
rect 4236 787 4243 876
rect 4256 827 4263 883
rect 3947 636 3963 643
rect 3856 607 3863 633
rect 3936 607 3943 633
rect 3976 607 3983 693
rect 4056 660 4063 663
rect 4053 647 4067 660
rect 3636 396 3683 403
rect 3256 360 3263 363
rect 3253 347 3267 360
rect 3236 227 3243 313
rect 3616 307 3623 331
rect 3676 327 3683 396
rect 3716 396 3743 403
rect 3796 396 3813 403
rect 3716 347 3723 396
rect 3836 366 3843 533
rect 3676 287 3683 313
rect 3236 176 3243 213
rect 3076 140 3083 143
rect 3073 127 3087 140
rect 3136 47 3143 174
rect 3260 143 3273 147
rect 3216 87 3223 143
rect 3256 136 3273 143
rect 3260 133 3273 136
rect 3296 127 3303 173
rect 3316 147 3323 273
rect 3576 207 3583 253
rect 3596 176 3603 253
rect 3376 87 3383 143
rect 3536 87 3543 143
rect 3573 127 3587 132
rect 3636 127 3643 173
rect 3656 146 3663 193
rect 3753 180 3767 193
rect 3756 176 3763 180
rect 3836 146 3843 273
rect 3856 267 3863 433
rect 3876 287 3883 473
rect 3956 396 3963 533
rect 3873 180 3887 193
rect 3876 176 3883 180
rect 3916 176 3923 333
rect 3936 247 3943 363
rect 3996 207 4003 373
rect 4016 366 4023 553
rect 4156 527 4163 653
rect 4253 627 4267 633
rect 4240 606 4260 607
rect 4247 593 4253 606
rect 4056 396 4063 433
rect 4096 396 4103 493
rect 4276 427 4283 753
rect 4296 727 4303 883
rect 4456 847 4463 883
rect 4696 847 4703 933
rect 4756 916 4763 1132
rect 4816 1067 4823 1214
rect 4856 1107 4863 1183
rect 4716 887 4723 914
rect 4856 886 4863 913
rect 4376 727 4383 753
rect 4373 700 4387 713
rect 4376 696 4383 700
rect 4276 396 4283 413
rect 4296 403 4303 692
rect 4336 660 4363 663
rect 4336 656 4367 660
rect 4313 607 4327 613
rect 4336 527 4343 656
rect 4353 647 4367 656
rect 4373 627 4387 633
rect 4367 596 4393 603
rect 4296 396 4323 403
rect 4116 327 4123 363
rect 4256 360 4263 363
rect 4253 347 4267 360
rect 4316 347 4323 396
rect 4336 347 4343 433
rect 4376 408 4383 573
rect 4456 487 4463 693
rect 4407 433 4413 447
rect 4476 427 4483 693
rect 4496 666 4503 733
rect 4576 696 4583 753
rect 4596 660 4603 663
rect 4593 647 4607 660
rect 4656 643 4663 833
rect 4736 696 4743 833
rect 4756 660 4763 663
rect 4636 636 4663 643
rect 4573 627 4587 633
rect 4413 400 4427 412
rect 4416 396 4423 400
rect 4353 347 4367 352
rect 4096 276 4133 283
rect 4096 227 4103 276
rect 4073 180 4087 193
rect 4116 187 4123 253
rect 4076 176 4083 180
rect 4136 167 4143 193
rect 4236 176 4243 233
rect 3936 107 3943 143
rect 4056 107 4063 143
rect 4156 47 4163 173
rect 4256 140 4263 143
rect 4253 127 4267 140
rect 4296 127 4303 333
rect 4396 227 4403 273
rect 4316 87 4323 193
rect 4353 180 4367 193
rect 4356 176 4363 180
rect 4416 146 4423 273
rect 4436 267 4443 363
rect 4476 287 4483 413
rect 4573 400 4587 413
rect 4576 396 4583 400
rect 4496 267 4503 394
rect 4393 127 4407 133
rect 4436 127 4443 213
rect 4453 187 4467 193
rect 4496 176 4503 253
rect 4556 227 4563 363
rect 4516 140 4523 143
rect 4513 127 4527 140
rect 4576 27 4583 233
rect 4596 227 4603 363
rect 4636 247 4643 636
rect 4676 607 4683 652
rect 4753 647 4767 660
rect 4716 607 4723 631
rect 4796 587 4803 694
rect 4816 647 4823 883
rect 4876 807 4883 1153
rect 4896 886 4903 1113
rect 4956 947 4963 1213
rect 4976 1107 4983 1353
rect 4996 1227 5003 1913
rect 5016 1887 5023 1932
rect 5036 1763 5043 2073
rect 5076 1956 5083 2033
rect 5096 1916 5123 1923
rect 5116 1867 5123 1916
rect 5036 1756 5063 1763
rect 5056 1736 5063 1756
rect 5076 1627 5083 1653
rect 5096 1463 5103 1753
rect 5087 1456 5103 1463
rect 5076 1436 5083 1453
rect 5016 1216 5023 1333
rect 5036 1267 5043 1403
rect 5056 1216 5063 1353
rect 5096 1216 5103 1433
rect 5116 1347 5123 1853
rect 5136 1847 5143 1873
rect 5156 1867 5163 2213
rect 5216 2187 5223 2223
rect 5276 2147 5283 2273
rect 5276 2107 5283 2133
rect 5253 1960 5267 1973
rect 5256 1956 5263 1960
rect 5156 1736 5163 1853
rect 5176 1787 5183 1953
rect 5256 1706 5263 1773
rect 5136 1367 5143 1633
rect 5296 1627 5303 2433
rect 5376 2367 5383 2443
rect 5416 2307 5423 2553
rect 5456 2488 5463 2773
rect 5476 2587 5483 2774
rect 5576 2746 5583 2833
rect 5536 2707 5543 2743
rect 5596 2607 5603 2873
rect 5656 2776 5663 2873
rect 5616 2707 5623 2774
rect 5673 2727 5687 2732
rect 5436 2476 5453 2483
rect 5436 2446 5443 2476
rect 5476 2476 5483 2513
rect 5516 2476 5523 2573
rect 5536 2440 5543 2443
rect 5533 2427 5547 2440
rect 5576 2327 5583 2553
rect 5596 2527 5603 2593
rect 5636 2476 5643 2513
rect 5733 2487 5747 2493
rect 5616 2387 5623 2433
rect 5656 2367 5663 2443
rect 5756 2407 5763 3113
rect 5776 2996 5783 3233
rect 5816 3167 5823 3263
rect 5836 3207 5843 3316
rect 5856 3267 5863 3333
rect 5776 2746 5783 2853
rect 5796 2847 5803 2963
rect 5856 2947 5863 3232
rect 5876 2967 5883 3413
rect 5896 3387 5903 3433
rect 5936 3296 5943 3393
rect 5996 3363 6003 3473
rect 6016 3427 6023 3514
rect 5996 3356 6023 3363
rect 6016 3287 6023 3356
rect 5896 2867 5903 3233
rect 5916 3207 5923 3252
rect 5956 3187 5963 3263
rect 5956 3127 5963 3173
rect 5916 3007 5923 3073
rect 5936 2996 5943 3033
rect 5976 3008 5983 3133
rect 6016 3087 6023 3252
rect 6036 2966 6043 3333
rect 6056 3307 6063 3413
rect 6076 3347 6083 3483
rect 6176 3486 6183 3713
rect 6116 3296 6123 3373
rect 6156 3307 6163 3473
rect 6176 3407 6183 3472
rect 6176 3367 6183 3393
rect 6176 3267 6183 3313
rect 6096 3260 6103 3263
rect 6056 3147 6063 3253
rect 6093 3247 6107 3260
rect 6136 3147 6143 3252
rect 5956 2960 5963 2963
rect 5836 2776 5843 2853
rect 5916 2743 5923 2953
rect 5953 2947 5967 2960
rect 5816 2740 5823 2743
rect 5813 2727 5827 2740
rect 5856 2707 5863 2743
rect 5896 2736 5923 2743
rect 5776 2507 5783 2533
rect 5796 2476 5803 2593
rect 5813 2507 5827 2513
rect 5836 2476 5843 2553
rect 5776 2383 5783 2413
rect 5756 2376 5783 2383
rect 5353 2260 5367 2273
rect 5356 2256 5363 2260
rect 5580 2263 5593 2267
rect 5576 2256 5593 2263
rect 5580 2253 5593 2256
rect 5336 2067 5343 2223
rect 5376 1956 5383 1993
rect 5356 1887 5363 1923
rect 5396 1920 5403 1923
rect 5393 1907 5407 1920
rect 5456 1907 5463 2053
rect 5476 2047 5483 2253
rect 5516 2147 5523 2173
rect 5556 2147 5563 2223
rect 5516 1956 5523 2133
rect 5576 2107 5583 2193
rect 5596 2007 5603 2213
rect 5616 2067 5623 2254
rect 5736 2256 5743 2313
rect 5756 2283 5763 2376
rect 5816 2367 5823 2443
rect 5787 2293 5793 2307
rect 5816 2287 5823 2332
rect 5856 2323 5863 2443
rect 5876 2387 5883 2433
rect 5896 2347 5903 2736
rect 5916 2427 5923 2713
rect 5936 2647 5943 2933
rect 5956 2727 5963 2873
rect 5996 2807 6003 2963
rect 6056 2827 6063 3073
rect 6136 2996 6143 3033
rect 6176 3007 6183 3232
rect 6196 2927 6203 3613
rect 6236 3527 6243 3736
rect 6276 3627 6283 3853
rect 6296 3787 6303 3953
rect 6336 3907 6343 4003
rect 6396 4006 6403 4193
rect 6356 3883 6363 3993
rect 6416 3907 6423 4213
rect 6436 4207 6443 4276
rect 6456 4167 6463 4253
rect 6476 4227 6483 4413
rect 6496 4207 6503 4473
rect 6516 4467 6523 4813
rect 6536 4727 6543 4893
rect 6556 4826 6563 4893
rect 6576 4867 6583 5513
rect 6596 5147 6603 5413
rect 6616 5387 6623 5513
rect 6636 5427 6643 5673
rect 6656 5447 6663 5753
rect 6696 5596 6703 5673
rect 6736 5607 6743 5833
rect 6716 5527 6723 5563
rect 6736 5503 6743 5553
rect 6716 5496 6743 5503
rect 6656 5403 6663 5433
rect 6656 5396 6683 5403
rect 6676 5376 6683 5396
rect 6716 5387 6723 5496
rect 6616 5127 6623 5333
rect 6656 5287 6663 5343
rect 6696 5340 6703 5343
rect 6693 5327 6707 5340
rect 6716 5287 6723 5333
rect 6736 5327 6743 5473
rect 6756 5303 6763 5856
rect 6736 5296 6763 5303
rect 6656 5076 6663 5113
rect 6636 4907 6643 5043
rect 6676 5007 6683 5043
rect 6653 4867 6667 4873
rect 6596 4820 6603 4823
rect 6576 4687 6583 4813
rect 6593 4807 6607 4820
rect 6596 4747 6603 4793
rect 6636 4767 6643 4791
rect 6536 4567 6543 4673
rect 6596 4556 6603 4613
rect 6536 4487 6543 4513
rect 6656 4523 6663 4813
rect 6616 4516 6663 4523
rect 6516 4347 6523 4393
rect 6556 4336 6563 4373
rect 6576 4367 6583 4491
rect 6596 4447 6603 4493
rect 6616 4407 6623 4493
rect 6636 4303 6643 4473
rect 6536 4147 6543 4271
rect 6476 4036 6483 4133
rect 6536 4047 6543 4093
rect 6436 3967 6443 3993
rect 6336 3876 6363 3883
rect 6336 3827 6343 3876
rect 6393 3820 6407 3833
rect 6396 3816 6403 3820
rect 6316 3767 6323 3813
rect 6216 3307 6223 3514
rect 6276 3516 6283 3553
rect 6296 3527 6303 3573
rect 6316 3487 6323 3673
rect 6256 3463 6263 3483
rect 6256 3456 6283 3463
rect 6256 3296 6263 3353
rect 6276 3327 6283 3456
rect 6296 3347 6303 3473
rect 6336 3427 6343 3773
rect 6356 3527 6363 3673
rect 6376 3667 6383 3783
rect 6413 3767 6427 3772
rect 6456 3747 6463 3933
rect 6396 3516 6403 3553
rect 6436 3516 6443 3553
rect 6456 3527 6463 3712
rect 6367 3483 6380 3487
rect 6367 3476 6383 3483
rect 6367 3473 6380 3476
rect 6287 3316 6303 3323
rect 6296 3296 6303 3316
rect 6336 3267 6343 3373
rect 6236 3187 6243 3263
rect 6276 3207 6283 3252
rect 6316 3047 6323 3253
rect 6356 3087 6363 3313
rect 6376 3307 6383 3453
rect 6416 3347 6423 3483
rect 6476 3467 6483 3973
rect 6496 3847 6503 4003
rect 6556 3987 6563 4273
rect 6576 4207 6583 4303
rect 6616 4296 6643 4303
rect 6656 4303 6663 4493
rect 6676 4347 6683 4953
rect 6696 4827 6703 5033
rect 6696 4507 6703 4693
rect 6716 4367 6723 5133
rect 6736 4487 6743 5296
rect 6756 4607 6763 5273
rect 6736 4336 6743 4433
rect 6776 4347 6783 5876
rect 6656 4296 6683 4303
rect 6616 4187 6623 4296
rect 6576 3947 6583 4172
rect 6636 4163 6643 4253
rect 6656 4223 6663 4273
rect 6676 4247 6683 4296
rect 6716 4283 6723 4292
rect 6696 4276 6723 4283
rect 6656 4216 6683 4223
rect 6636 4156 6653 4163
rect 6616 4048 6623 4073
rect 6656 4036 6663 4153
rect 6676 4063 6683 4216
rect 6696 4087 6703 4276
rect 6676 4060 6703 4063
rect 6676 4056 6707 4060
rect 6693 4047 6707 4056
rect 6593 3983 6607 3993
rect 6593 3980 6623 3983
rect 6596 3976 6623 3980
rect 6516 3816 6523 3873
rect 6553 3820 6567 3833
rect 6596 3827 6603 3913
rect 6556 3816 6563 3820
rect 6616 3783 6623 3976
rect 6636 3907 6643 4003
rect 6656 3883 6663 3973
rect 6576 3763 6583 3783
rect 6556 3756 6583 3763
rect 6596 3776 6623 3783
rect 6636 3876 6663 3883
rect 6393 3300 6407 3313
rect 6396 3296 6403 3300
rect 6436 3296 6443 3333
rect 6216 2967 6223 3033
rect 6216 2927 6223 2953
rect 6236 2947 6243 3013
rect 6256 3007 6263 3033
rect 6276 2996 6283 3033
rect 6313 3008 6327 3012
rect 6376 2967 6383 3253
rect 6416 3167 6423 3263
rect 6456 3147 6463 3252
rect 6496 3247 6503 3733
rect 6556 3667 6563 3756
rect 6596 3687 6603 3776
rect 6616 3707 6623 3753
rect 6153 2907 6167 2913
rect 6147 2900 6167 2907
rect 6147 2896 6163 2900
rect 6147 2893 6160 2896
rect 5996 2776 6003 2793
rect 6076 2787 6083 2893
rect 5976 2507 5983 2733
rect 6016 2687 6023 2743
rect 6056 2740 6063 2743
rect 6053 2727 6067 2740
rect 6096 2746 6103 2813
rect 6136 2787 6143 2853
rect 6256 2847 6263 2953
rect 6153 2780 6167 2793
rect 6193 2780 6207 2793
rect 6156 2776 6163 2780
rect 6196 2776 6203 2780
rect 5993 2488 6007 2493
rect 5947 2483 5960 2487
rect 5947 2476 5963 2483
rect 5947 2473 5960 2476
rect 6036 2483 6043 2633
rect 6076 2603 6083 2733
rect 6096 2687 6103 2732
rect 6116 2607 6123 2773
rect 6136 2707 6143 2733
rect 6216 2740 6223 2743
rect 6213 2727 6227 2740
rect 6256 2727 6263 2753
rect 6276 2727 6283 2933
rect 6296 2907 6303 2963
rect 6396 2907 6403 3053
rect 6436 2996 6443 3053
rect 6476 3028 6483 3113
rect 6516 3087 6523 3533
rect 6556 3516 6563 3653
rect 6576 3547 6583 3633
rect 6576 3463 6583 3472
rect 6556 3456 6583 3463
rect 6556 3307 6563 3456
rect 6616 3347 6623 3553
rect 6636 3487 6643 3876
rect 6676 3843 6683 4003
rect 6696 3927 6703 3993
rect 6656 3840 6683 3843
rect 6653 3836 6683 3840
rect 6653 3827 6667 3836
rect 6696 3816 6703 3873
rect 6716 3843 6723 4233
rect 6736 4223 6743 4273
rect 6756 4267 6763 4303
rect 6736 4216 6763 4223
rect 6736 3867 6743 4193
rect 6716 3836 6743 3843
rect 6736 3816 6743 3836
rect 6756 3827 6763 4216
rect 6676 3780 6683 3783
rect 6656 3527 6663 3772
rect 6673 3767 6687 3780
rect 6696 3516 6703 3553
rect 6736 3528 6743 3693
rect 6756 3527 6763 3773
rect 6776 3647 6783 4293
rect 6656 3367 6663 3453
rect 6676 3387 6683 3483
rect 6776 3483 6783 3553
rect 6756 3476 6783 3483
rect 6696 3403 6703 3453
rect 6696 3396 6723 3403
rect 6593 3300 6607 3313
rect 6596 3296 6603 3300
rect 6536 3067 6543 3273
rect 6516 3008 6523 3033
rect 6307 2783 6320 2787
rect 6307 2776 6323 2783
rect 6356 2776 6363 2893
rect 6307 2773 6320 2776
rect 6076 2596 6103 2603
rect 6056 2527 6063 2553
rect 6036 2476 6063 2483
rect 5856 2316 5883 2323
rect 5833 2307 5847 2313
rect 5756 2276 5783 2283
rect 5636 2207 5643 2253
rect 5676 2220 5683 2223
rect 5673 2207 5687 2220
rect 5716 2203 5723 2223
rect 5707 2196 5723 2203
rect 5587 1956 5603 1963
rect 5596 1907 5603 1956
rect 5336 1736 5343 1853
rect 5456 1736 5463 1773
rect 5636 1748 5643 2073
rect 5696 1956 5703 2193
rect 5676 1907 5683 1923
rect 5776 1907 5783 2276
rect 5816 2226 5823 2273
rect 5876 2256 5883 2316
rect 5976 2283 5983 2443
rect 6056 2387 6063 2476
rect 6076 2407 6083 2573
rect 6096 2487 6103 2596
rect 6133 2480 6147 2493
rect 6136 2476 6143 2480
rect 6176 2476 6183 2513
rect 5956 2276 5983 2283
rect 5896 2220 5903 2223
rect 5893 2207 5907 2220
rect 5836 1968 5843 2033
rect 5876 1956 5883 1993
rect 5687 1896 5703 1903
rect 5396 1627 5403 1733
rect 5476 1700 5483 1703
rect 5473 1687 5487 1700
rect 5536 1667 5543 1713
rect 5316 1436 5323 1493
rect 5356 1467 5363 1593
rect 5356 1436 5363 1453
rect 5036 1107 5043 1183
rect 5056 1007 5063 1153
rect 5096 1027 5103 1053
rect 4916 696 4923 793
rect 4956 666 4963 813
rect 4856 660 4863 663
rect 4656 363 4663 553
rect 4816 547 4823 633
rect 4836 467 4843 653
rect 4853 647 4867 660
rect 4976 627 4983 713
rect 4716 408 4723 433
rect 4836 403 4843 453
rect 4996 408 5003 933
rect 5056 928 5063 993
rect 5096 916 5103 1013
rect 5136 947 5143 1253
rect 5156 1227 5163 1373
rect 5216 1327 5223 1403
rect 5276 1127 5283 1313
rect 5336 1223 5343 1403
rect 5376 1400 5383 1403
rect 5373 1387 5387 1400
rect 5416 1347 5423 1473
rect 5316 1216 5343 1223
rect 5376 1216 5383 1333
rect 5196 916 5223 923
rect 5276 916 5283 1053
rect 5016 886 5023 913
rect 5033 700 5047 713
rect 5076 703 5083 883
rect 5113 727 5127 733
rect 5036 696 5043 700
rect 5076 696 5103 703
rect 5056 647 5063 663
rect 5056 636 5073 647
rect 5060 633 5073 636
rect 5096 587 5103 696
rect 5116 666 5123 713
rect 5176 696 5183 753
rect 5196 727 5203 916
rect 5296 707 5303 1214
rect 5316 1067 5323 1216
rect 5316 696 5323 1013
rect 5336 787 5343 1093
rect 5356 1087 5363 1172
rect 5396 1127 5403 1183
rect 5393 920 5407 933
rect 5396 916 5403 920
rect 5436 916 5443 1553
rect 5556 1527 5563 1733
rect 5616 1700 5623 1703
rect 5613 1687 5627 1700
rect 5656 1687 5663 1703
rect 5653 1667 5667 1673
rect 5456 1367 5463 1513
rect 5513 1440 5527 1453
rect 5516 1436 5523 1440
rect 5496 1367 5503 1403
rect 5456 927 5463 1332
rect 5536 1247 5543 1403
rect 5596 1387 5603 1493
rect 5516 1236 5533 1243
rect 5516 1216 5523 1236
rect 5556 1216 5563 1253
rect 5496 1147 5503 1183
rect 5536 1180 5543 1183
rect 5533 1167 5547 1180
rect 5596 1127 5603 1293
rect 5616 1186 5623 1533
rect 5696 1487 5703 1896
rect 5716 1703 5723 1891
rect 5856 1847 5863 1923
rect 5936 1887 5943 2213
rect 5956 2207 5963 2276
rect 5996 2267 6003 2373
rect 6096 2323 6103 2433
rect 6156 2407 6163 2443
rect 6076 2316 6103 2323
rect 6016 2256 6023 2293
rect 6076 2267 6083 2316
rect 5976 2147 5983 2253
rect 6036 2187 6043 2223
rect 6047 1996 6063 2003
rect 5976 1956 5983 1993
rect 6036 1956 6043 1993
rect 5956 1926 5963 1953
rect 5867 1836 5883 1843
rect 5716 1696 5743 1703
rect 5756 1700 5763 1703
rect 5796 1700 5803 1703
rect 5656 1400 5663 1403
rect 5653 1387 5667 1400
rect 5716 1347 5723 1553
rect 5676 1247 5683 1333
rect 5673 1220 5687 1233
rect 5676 1216 5683 1220
rect 5736 1227 5743 1696
rect 5753 1687 5767 1700
rect 5793 1687 5807 1700
rect 5836 1436 5843 1693
rect 5856 1567 5863 1773
rect 5776 1367 5783 1403
rect 5656 1147 5663 1183
rect 5736 1107 5743 1173
rect 5756 1147 5763 1333
rect 5876 1307 5883 1836
rect 5976 1787 5983 1813
rect 5976 1736 5983 1773
rect 5916 1687 5923 1703
rect 5896 1427 5903 1613
rect 5916 1507 5923 1673
rect 5956 1627 5963 1703
rect 6016 1607 6023 1873
rect 6056 1743 6063 1996
rect 6096 1807 6103 2293
rect 6116 2047 6123 2333
rect 6153 2260 6167 2273
rect 6196 2267 6203 2433
rect 6216 2427 6223 2533
rect 6156 2256 6163 2260
rect 6216 2227 6223 2392
rect 6136 2027 6143 2213
rect 6216 2147 6223 2192
rect 6236 2167 6243 2713
rect 6256 2407 6263 2713
rect 6296 2527 6303 2733
rect 6376 2740 6383 2743
rect 6373 2727 6387 2740
rect 6367 2706 6380 2707
rect 6367 2693 6373 2706
rect 6336 2476 6343 2573
rect 6316 2440 6323 2443
rect 6313 2427 6327 2440
rect 6296 2256 6303 2333
rect 6316 2307 6323 2353
rect 6356 2327 6363 2443
rect 6396 2367 6403 2733
rect 6416 2667 6423 2953
rect 6436 2747 6443 2933
rect 6456 2907 6463 2963
rect 6496 2927 6503 2963
rect 6536 2927 6543 3013
rect 6556 2947 6563 3253
rect 6456 2787 6463 2893
rect 6476 2807 6483 2853
rect 6496 2788 6503 2813
rect 6433 2687 6447 2693
rect 6416 2427 6423 2593
rect 6476 2488 6483 2513
rect 6536 2503 6543 2892
rect 6576 2867 6583 3231
rect 6616 3167 6623 3263
rect 6676 3167 6683 3333
rect 6656 2996 6663 3033
rect 6696 3007 6703 3353
rect 6716 2963 6723 3396
rect 6736 3387 6743 3453
rect 6527 2496 6543 2503
rect 6556 2856 6573 2863
rect 6513 2480 6527 2493
rect 6516 2476 6523 2480
rect 6336 2316 6353 2323
rect 6336 2267 6343 2316
rect 6376 2283 6383 2333
rect 6436 2307 6443 2433
rect 6456 2288 6463 2443
rect 6496 2440 6503 2443
rect 6493 2427 6507 2440
rect 6533 2423 6547 2433
rect 6516 2420 6547 2423
rect 6516 2416 6543 2420
rect 6356 2276 6383 2283
rect 6356 2226 6363 2276
rect 6496 2267 6503 2413
rect 6276 2220 6283 2223
rect 6116 1923 6123 1954
rect 6116 1916 6143 1923
rect 6036 1736 6063 1743
rect 6036 1547 6043 1736
rect 6136 1736 6143 1916
rect 6156 1847 6163 1923
rect 6256 1907 6263 2213
rect 6273 2207 6287 2220
rect 6276 1927 6283 2153
rect 6076 1627 6083 1703
rect 6116 1700 6123 1703
rect 6113 1687 6127 1700
rect 5976 1436 5983 1493
rect 6056 1406 6063 1473
rect 5516 916 5563 923
rect 5496 887 5503 914
rect 5516 827 5523 916
rect 5616 886 5623 973
rect 5736 916 5743 1013
rect 5536 696 5543 773
rect 5196 660 5203 663
rect 5193 647 5207 660
rect 5236 607 5243 652
rect 5256 627 5263 693
rect 5376 647 5383 663
rect 5416 647 5423 694
rect 5596 666 5603 833
rect 5676 827 5683 883
rect 5696 696 5703 773
rect 5476 660 5483 663
rect 5516 660 5523 663
rect 5473 647 5487 660
rect 5513 647 5527 660
rect 5376 567 5383 633
rect 5393 607 5407 613
rect 5416 527 5423 633
rect 5500 626 5520 627
rect 5507 613 5513 626
rect 4836 396 4863 403
rect 4656 356 4703 363
rect 4676 176 4683 333
rect 4716 176 4723 233
rect 4736 187 4743 363
rect 4616 107 4623 173
rect 4776 107 4783 233
rect 4836 227 4843 373
rect 4976 363 4983 393
rect 4996 366 5003 394
rect 5047 403 5060 407
rect 5047 396 5063 403
rect 5176 396 5183 453
rect 5047 393 5060 396
rect 4956 356 4983 363
rect 4836 176 4843 213
rect 4896 146 4903 213
rect 4916 188 4923 323
rect 4996 176 5003 213
rect 5136 176 5143 313
rect 5196 267 5203 363
rect 5276 287 5283 513
rect 5373 400 5387 413
rect 5376 396 5383 400
rect 5296 327 5303 394
rect 5356 360 5363 363
rect 5353 347 5367 360
rect 5416 323 5423 353
rect 5436 347 5443 553
rect 5633 408 5647 413
rect 5416 316 5443 323
rect 4976 140 4983 143
rect 4973 127 4987 140
rect 5216 47 5223 213
rect 5316 203 5323 293
rect 5296 196 5323 203
rect 5296 176 5303 196
rect 5336 176 5343 273
rect 5376 146 5383 213
rect 5396 146 5403 253
rect 5436 176 5443 316
rect 5496 267 5503 363
rect 5656 360 5663 363
rect 5653 347 5667 360
rect 5636 307 5643 333
rect 5696 327 5703 353
rect 5713 347 5727 353
rect 5736 307 5743 853
rect 5776 703 5783 1253
rect 5836 1216 5843 1293
rect 5873 1220 5887 1233
rect 5876 1216 5883 1220
rect 5796 967 5803 1172
rect 5796 887 5803 953
rect 5816 867 5823 1183
rect 5856 1180 5863 1183
rect 5853 1167 5867 1180
rect 5916 1007 5923 1353
rect 5913 920 5927 933
rect 5936 928 5943 1293
rect 5956 1227 5963 1403
rect 6076 1347 6083 1553
rect 6176 1487 6183 1733
rect 6196 1507 6203 1793
rect 6296 1767 6303 2173
rect 6376 2007 6383 2253
rect 6516 2227 6523 2416
rect 6476 2087 6483 2223
rect 6536 2067 6543 2273
rect 6447 2043 6460 2047
rect 6447 2033 6463 2043
rect 6336 1956 6343 1993
rect 6416 1987 6423 2013
rect 6316 1847 6323 1912
rect 6300 1743 6313 1747
rect 6296 1736 6313 1743
rect 6300 1733 6313 1736
rect 6236 1527 6243 1703
rect 6096 1387 6103 1473
rect 6196 1448 6203 1493
rect 6136 1287 6143 1403
rect 6176 1400 6183 1403
rect 6173 1387 6187 1400
rect 5976 1260 6013 1263
rect 5973 1256 6013 1260
rect 5973 1247 5987 1256
rect 5986 1240 5987 1247
rect 5993 1220 6007 1233
rect 5996 1216 6003 1220
rect 6016 1180 6023 1183
rect 6013 1167 6027 1180
rect 5916 916 5923 920
rect 5856 787 5863 883
rect 5956 883 5963 1093
rect 5976 886 5983 993
rect 6036 987 6043 1173
rect 6056 1087 6063 1213
rect 6076 1186 6083 1273
rect 6156 1216 6163 1333
rect 6196 1227 6203 1253
rect 6176 1163 6183 1183
rect 6236 1167 6243 1473
rect 6256 1287 6263 1434
rect 6276 1403 6283 1593
rect 6336 1487 6343 1753
rect 6356 1567 6363 1923
rect 6396 1907 6403 1923
rect 6387 1896 6403 1907
rect 6387 1893 6400 1896
rect 6436 1847 6443 1993
rect 6456 1867 6463 2033
rect 6556 2007 6563 2856
rect 6596 2827 6603 2953
rect 6636 2883 6643 2963
rect 6616 2876 6643 2883
rect 6656 2883 6663 2933
rect 6676 2907 6683 2963
rect 6696 2956 6723 2963
rect 6656 2876 6683 2883
rect 6616 2847 6623 2876
rect 6600 2803 6613 2807
rect 6596 2793 6613 2803
rect 6596 2776 6603 2793
rect 6636 2776 6643 2853
rect 6676 2783 6683 2876
rect 6696 2807 6703 2956
rect 6676 2776 6703 2783
rect 6656 2723 6663 2743
rect 6636 2716 6663 2723
rect 6636 2687 6643 2716
rect 6636 2507 6643 2673
rect 6656 2567 6663 2693
rect 6576 2347 6583 2493
rect 6607 2483 6620 2487
rect 6607 2476 6623 2483
rect 6656 2476 6663 2532
rect 6676 2487 6683 2733
rect 6607 2473 6620 2476
rect 6636 2440 6643 2443
rect 6596 2323 6603 2433
rect 6633 2427 6647 2440
rect 6596 2316 6613 2323
rect 6616 2256 6623 2313
rect 6576 2147 6583 2223
rect 6556 1907 6563 1972
rect 6376 1706 6383 1833
rect 6393 1747 6407 1753
rect 6436 1736 6443 1793
rect 6493 1743 6507 1753
rect 6487 1740 6507 1743
rect 6487 1736 6503 1740
rect 6333 1440 6347 1452
rect 6376 1448 6383 1593
rect 6416 1467 6423 1703
rect 6516 1587 6523 1853
rect 6536 1607 6543 1753
rect 6556 1747 6563 1872
rect 6576 1767 6583 2053
rect 6616 1956 6623 2013
rect 6636 1987 6643 2212
rect 6656 2087 6663 2293
rect 6676 2027 6683 2433
rect 6696 2427 6703 2776
rect 6716 2707 6723 2933
rect 6656 1956 6663 1993
rect 6696 1967 6703 2392
rect 6596 1736 6603 1793
rect 6613 1767 6627 1773
rect 6636 1736 6643 1833
rect 6656 1747 6663 1893
rect 6676 1887 6683 1923
rect 6436 1467 6443 1553
rect 6336 1436 6343 1440
rect 6276 1396 6303 1403
rect 6276 1307 6283 1333
rect 6256 1247 6263 1273
rect 6296 1267 6303 1396
rect 6416 1403 6423 1453
rect 6496 1448 6503 1513
rect 6536 1507 6543 1593
rect 6556 1443 6563 1693
rect 6576 1607 6583 1703
rect 6676 1627 6683 1793
rect 6536 1436 6583 1443
rect 6356 1347 6363 1403
rect 6396 1396 6423 1403
rect 6260 1226 6280 1227
rect 6267 1223 6280 1226
rect 6267 1216 6283 1223
rect 6267 1213 6280 1216
rect 6156 1156 6183 1163
rect 5936 876 5963 883
rect 5756 696 5783 703
rect 5796 696 5803 773
rect 5936 747 5943 876
rect 5836 696 5843 733
rect 5756 666 5763 696
rect 5956 696 5963 753
rect 5996 708 6003 973
rect 6076 947 6083 1053
rect 6076 916 6083 933
rect 6096 703 6103 872
rect 6136 847 6143 914
rect 6156 867 6163 1156
rect 6296 1087 6303 1183
rect 6196 916 6203 973
rect 6316 928 6323 1153
rect 6376 1027 6383 1253
rect 6396 1127 6403 1396
rect 6436 1327 6443 1432
rect 6467 1403 6480 1407
rect 6467 1393 6483 1403
rect 6436 1216 6443 1292
rect 6476 1228 6483 1393
rect 6496 1180 6523 1183
rect 6496 1176 6527 1180
rect 6496 1087 6503 1176
rect 6513 1167 6527 1176
rect 6336 883 6343 953
rect 6076 696 6103 703
rect 6136 696 6143 833
rect 5856 627 5863 663
rect 5916 467 5923 693
rect 5976 627 5983 663
rect 6056 647 6063 693
rect 6076 666 6083 696
rect 6156 660 6163 663
rect 6153 647 6167 660
rect 5853 400 5867 413
rect 5856 396 5863 400
rect 6013 400 6027 413
rect 6016 396 6023 400
rect 6176 396 6183 453
rect 5756 363 5763 394
rect 5756 356 5783 363
rect 5516 227 5523 273
rect 5556 146 5563 213
rect 5596 176 5603 273
rect 5696 143 5703 253
rect 5756 176 5763 333
rect 5776 247 5783 356
rect 5796 307 5803 363
rect 5836 327 5843 363
rect 5916 327 5923 394
rect 6216 366 6223 753
rect 6236 627 6243 853
rect 6256 843 6263 883
rect 6336 876 6353 883
rect 6256 836 6283 843
rect 6276 696 6283 836
rect 6316 696 6323 833
rect 6376 666 6383 693
rect 6296 607 6303 663
rect 6276 596 6293 603
rect 6276 408 6283 596
rect 6316 396 6323 453
rect 5996 360 6003 363
rect 5993 347 6007 360
rect 5816 147 5823 233
rect 5956 176 5963 273
rect 5996 147 6003 233
rect 6076 176 6083 313
rect 6116 303 6123 363
rect 6096 296 6123 303
rect 6096 247 6103 296
rect 6116 176 6123 273
rect 6236 247 6243 273
rect 6216 176 6223 213
rect 6336 147 6343 363
rect 6376 307 6383 652
rect 6396 607 6403 843
rect 6476 707 6483 1013
rect 6536 847 6543 1313
rect 6556 1167 6563 1393
rect 6576 1387 6583 1436
rect 6576 1347 6583 1373
rect 6596 1283 6603 1613
rect 6616 1407 6623 1593
rect 6696 1567 6703 1913
rect 6716 1747 6723 2653
rect 6736 1847 6743 3352
rect 6656 1467 6663 1493
rect 6676 1436 6683 1513
rect 6713 1440 6727 1453
rect 6736 1447 6743 1733
rect 6716 1436 6723 1440
rect 6756 1407 6763 3476
rect 6776 3127 6783 3453
rect 6776 1767 6783 3073
rect 6696 1400 6703 1403
rect 6693 1387 6707 1400
rect 6576 1276 6603 1283
rect 6576 1227 6583 1276
rect 6596 1216 6603 1253
rect 6616 1180 6623 1183
rect 6613 1167 6627 1180
rect 6556 823 6563 1113
rect 6556 816 6583 823
rect 6460 666 6480 667
rect 6460 663 6473 666
rect 6456 656 6473 663
rect 6460 653 6473 656
rect 6473 400 6487 413
rect 6536 408 6543 733
rect 6576 696 6583 816
rect 6616 767 6623 843
rect 6593 723 6607 733
rect 6593 720 6623 723
rect 6596 716 6623 720
rect 6616 696 6623 716
rect 6636 660 6643 663
rect 6633 647 6647 660
rect 6676 647 6683 753
rect 6616 636 6633 643
rect 6476 396 6483 400
rect 6396 347 6403 394
rect 6556 367 6563 613
rect 6616 396 6623 636
rect 6396 176 6403 333
rect 6496 267 6503 363
rect 6576 176 6583 353
rect 6596 247 6603 363
rect 6636 307 6643 363
rect 6736 188 6743 1393
rect 6776 767 6783 1573
rect 5656 136 5703 143
rect 5896 47 5903 143
rect 5993 107 6007 112
rect 6036 107 6043 133
rect 6053 127 6067 132
rect 6096 107 6103 143
rect 6280 143 6293 147
rect 6276 136 6293 143
rect 6280 133 6293 136
rect 6456 47 6463 143
rect 6596 47 6603 143
rect 2596 -24 2623 -17
rect 2756 -24 2783 -17
rect 2996 -24 3023 -17
rect 4456 -24 4463 13
<< m3contact >>
rect 533 6493 547 6507
rect 1273 6493 1287 6507
rect 2333 6493 2347 6507
rect 173 6453 187 6467
rect 113 6414 127 6428
rect 73 6353 87 6367
rect 153 6313 167 6327
rect 133 6114 147 6128
rect 213 6414 227 6428
rect 273 6414 287 6428
rect 373 6413 387 6427
rect 433 6414 447 6428
rect 573 6453 587 6467
rect 533 6413 547 6427
rect 613 6414 627 6428
rect 733 6414 747 6428
rect 793 6413 807 6427
rect 213 6114 227 6128
rect 373 6372 387 6386
rect 413 6372 427 6386
rect 453 6372 467 6386
rect 553 6372 567 6386
rect 293 6353 307 6367
rect 453 6313 467 6327
rect 753 6372 767 6386
rect 553 6213 567 6227
rect 593 6213 607 6227
rect 293 6153 307 6167
rect 153 6072 167 6086
rect 73 6013 87 6027
rect 113 6013 127 6027
rect 153 5894 167 5908
rect 173 5852 187 5866
rect 253 6113 267 6127
rect 453 6133 467 6147
rect 333 6114 347 6128
rect 533 6093 547 6107
rect 313 6072 327 6086
rect 473 6072 487 6086
rect 353 6053 367 6067
rect 353 6013 367 6027
rect 233 5894 247 5908
rect 293 5894 307 5908
rect 113 5813 127 5827
rect 233 5613 247 5627
rect 53 5552 67 5566
rect 113 5552 127 5566
rect 213 5533 227 5547
rect 153 5513 167 5527
rect 113 5374 127 5388
rect 153 5374 167 5388
rect 233 5493 247 5507
rect 313 5852 327 5866
rect 593 6173 607 6187
rect 733 6153 747 6167
rect 653 6133 667 6147
rect 553 6073 567 6087
rect 613 6072 627 6086
rect 533 5973 547 5987
rect 573 5973 587 5987
rect 433 5933 447 5947
rect 513 5933 527 5947
rect 373 5893 387 5907
rect 893 6414 907 6428
rect 953 6413 967 6427
rect 1033 6414 1047 6428
rect 1153 6414 1167 6428
rect 1393 6453 1407 6467
rect 1473 6453 1487 6467
rect 1513 6453 1527 6467
rect 1733 6453 1747 6467
rect 1333 6413 1347 6427
rect 1433 6414 1447 6428
rect 873 6372 887 6386
rect 913 6353 927 6367
rect 813 6173 827 6187
rect 933 6173 947 6187
rect 853 6153 867 6167
rect 773 6114 787 6128
rect 893 6114 907 6128
rect 1053 6373 1067 6387
rect 1013 6353 1027 6367
rect 1293 6372 1307 6386
rect 1573 6414 1587 6428
rect 1613 6414 1627 6428
rect 1673 6414 1687 6428
rect 1773 6414 1787 6428
rect 1833 6414 1847 6428
rect 1913 6414 1927 6428
rect 1953 6414 1967 6428
rect 1413 6372 1427 6386
rect 1453 6372 1467 6386
rect 1513 6372 1527 6386
rect 1173 6353 1187 6367
rect 1333 6353 1347 6367
rect 1533 6353 1547 6367
rect 1133 6333 1147 6347
rect 1633 6372 1647 6386
rect 1693 6372 1707 6386
rect 1673 6333 1687 6347
rect 1593 6273 1607 6287
rect 1473 6233 1487 6247
rect 1053 6193 1067 6207
rect 1233 6193 1247 6207
rect 1293 6193 1307 6207
rect 953 6153 967 6167
rect 1013 6114 1027 6128
rect 1193 6173 1207 6187
rect 1093 6114 1107 6128
rect 753 6072 767 6086
rect 853 6072 867 6086
rect 913 6072 927 6086
rect 953 6053 967 6067
rect 653 5953 667 5967
rect 833 5953 847 5967
rect 613 5894 627 5908
rect 373 5852 387 5866
rect 413 5852 427 5866
rect 513 5852 527 5866
rect 553 5852 567 5866
rect 453 5813 467 5827
rect 593 5813 607 5827
rect 353 5713 367 5727
rect 273 5693 287 5707
rect 313 5693 327 5707
rect 413 5653 427 5667
rect 453 5653 467 5667
rect 613 5653 627 5667
rect 313 5594 327 5608
rect 273 5553 287 5567
rect 333 5552 347 5566
rect 453 5613 467 5627
rect 493 5594 507 5608
rect 553 5594 567 5608
rect 713 5933 727 5947
rect 793 5913 807 5927
rect 873 5913 887 5927
rect 733 5852 747 5866
rect 793 5853 807 5867
rect 853 5852 867 5866
rect 833 5833 847 5847
rect 893 5833 907 5847
rect 953 5833 967 5847
rect 773 5813 787 5827
rect 653 5613 667 5627
rect 413 5552 427 5566
rect 473 5552 487 5566
rect 513 5533 527 5547
rect 393 5493 407 5507
rect 213 5373 227 5387
rect 53 5333 67 5347
rect 93 5332 107 5346
rect 213 5332 227 5346
rect 113 5133 127 5147
rect 73 5073 87 5087
rect 153 5074 167 5088
rect 193 5074 207 5088
rect 93 5032 107 5046
rect 133 5032 147 5046
rect 113 5013 127 5027
rect 153 4853 167 4867
rect 53 4693 67 4707
rect 133 4693 147 4707
rect 533 5473 547 5487
rect 733 5593 747 5607
rect 773 5594 787 5608
rect 633 5473 647 5487
rect 273 5332 287 5346
rect 233 5253 247 5267
rect 293 5253 307 5267
rect 233 5193 247 5207
rect 213 5033 227 5047
rect 613 5393 627 5407
rect 673 5393 687 5407
rect 593 5332 607 5346
rect 913 5594 927 5608
rect 1013 6053 1027 6067
rect 1213 6053 1227 6067
rect 1073 6033 1087 6047
rect 1053 5933 1067 5947
rect 1233 5933 1247 5947
rect 1093 5894 1107 5908
rect 1153 5894 1167 5908
rect 1193 5894 1207 5908
rect 1373 6153 1387 6167
rect 1413 6114 1427 6128
rect 1453 6114 1467 6128
rect 1293 6033 1307 6047
rect 1393 6072 1407 6086
rect 1353 5993 1367 6007
rect 1793 6372 1807 6386
rect 1733 6273 1747 6287
rect 1693 6213 1707 6227
rect 1573 6193 1587 6207
rect 1673 6193 1687 6207
rect 1593 6173 1607 6187
rect 1653 6173 1667 6187
rect 2033 6413 2047 6427
rect 2093 6414 2107 6428
rect 2133 6414 2147 6428
rect 2233 6414 2247 6428
rect 2273 6414 2287 6428
rect 2013 6393 2027 6407
rect 1933 6372 1947 6386
rect 1973 6372 1987 6386
rect 1933 6333 1947 6347
rect 2013 6333 2027 6347
rect 1773 6293 1787 6307
rect 1833 6293 1847 6307
rect 1753 6233 1767 6247
rect 1533 6153 1547 6167
rect 1613 6152 1627 6166
rect 1733 6153 1747 6167
rect 1573 6114 1587 6128
rect 1473 6073 1487 6087
rect 1553 6072 1567 6086
rect 1513 5993 1527 6007
rect 1413 5933 1427 5947
rect 1453 5933 1467 5947
rect 1473 5913 1487 5927
rect 1013 5852 1027 5866
rect 1093 5853 1107 5867
rect 1213 5852 1227 5866
rect 1073 5793 1087 5807
rect 1153 5793 1167 5807
rect 1293 5893 1307 5907
rect 1353 5894 1367 5908
rect 1473 5892 1487 5906
rect 1293 5833 1307 5847
rect 1373 5852 1387 5866
rect 1673 6114 1687 6128
rect 1753 6113 1767 6127
rect 1613 5973 1627 5987
rect 1733 6073 1747 6087
rect 1833 6114 1847 6128
rect 1773 6073 1787 6087
rect 1813 6072 1827 6086
rect 1753 6053 1767 6067
rect 1853 6053 1867 6067
rect 2033 6313 2047 6327
rect 2113 6372 2127 6386
rect 2173 6372 2187 6386
rect 2213 6372 2227 6386
rect 2253 6372 2267 6386
rect 2292 6372 2306 6386
rect 2313 6373 2327 6387
rect 2353 6414 2367 6428
rect 2393 6414 2407 6428
rect 2333 6353 2347 6367
rect 2213 6313 2227 6327
rect 2453 6413 2467 6427
rect 2533 6414 2547 6428
rect 2633 6414 2647 6428
rect 2793 6513 2807 6527
rect 2833 6513 2847 6527
rect 2993 6513 3007 6527
rect 3093 6513 3107 6527
rect 2693 6473 2707 6487
rect 2733 6453 2747 6467
rect 2413 6372 2427 6386
rect 2553 6372 2567 6386
rect 2693 6414 2707 6428
rect 2673 6372 2687 6386
rect 2513 6333 2527 6347
rect 2633 6333 2647 6347
rect 2453 6313 2467 6327
rect 2113 6273 2127 6287
rect 2173 6273 2187 6287
rect 2353 6273 2367 6287
rect 2113 6213 2127 6227
rect 2133 6193 2147 6207
rect 2073 6153 2087 6167
rect 1993 6114 2007 6128
rect 2213 6173 2227 6187
rect 1933 6073 1947 6087
rect 1973 6072 1987 6086
rect 1913 5993 1927 6007
rect 2013 5993 2027 6007
rect 1913 5972 1927 5986
rect 1693 5953 1707 5967
rect 1533 5913 1547 5927
rect 1733 5913 1747 5927
rect 1793 5913 1807 5927
rect 1573 5894 1587 5908
rect 1653 5893 1667 5907
rect 1753 5894 1767 5908
rect 1873 5894 1887 5908
rect 2173 6114 2187 6128
rect 2093 6093 2107 6107
rect 2073 5953 2087 5967
rect 2013 5913 2027 5927
rect 1953 5894 1967 5908
rect 1513 5853 1527 5867
rect 1533 5852 1547 5866
rect 1333 5793 1347 5807
rect 1473 5793 1487 5807
rect 1773 5773 1787 5787
rect 1133 5673 1147 5687
rect 1233 5673 1247 5687
rect 793 5453 807 5467
rect 793 5393 807 5407
rect 833 5374 847 5388
rect 893 5533 907 5547
rect 1073 5594 1087 5608
rect 1193 5594 1207 5608
rect 993 5513 1007 5527
rect 1113 5553 1127 5567
rect 1093 5453 1107 5467
rect 1253 5653 1267 5667
rect 1313 5552 1327 5566
rect 1193 5533 1207 5547
rect 1233 5533 1247 5547
rect 893 5393 907 5407
rect 933 5393 947 5407
rect 953 5374 967 5388
rect 1013 5373 1027 5387
rect 1133 5413 1147 5427
rect 733 5332 747 5346
rect 773 5332 787 5346
rect 813 5332 827 5346
rect 872 5332 886 5346
rect 893 5332 907 5346
rect 933 5332 947 5346
rect 333 5233 347 5247
rect 233 5013 247 5027
rect 313 5033 327 5047
rect 293 5013 307 5027
rect 253 4933 267 4947
rect 193 4753 207 4767
rect 253 4753 267 4767
rect 213 4653 227 4667
rect 113 4633 127 4647
rect 173 4633 187 4647
rect 93 4553 107 4567
rect 33 4512 47 4526
rect 33 4353 47 4367
rect 153 4554 167 4568
rect 153 4493 167 4507
rect 253 4493 267 4507
rect 113 4353 127 4367
rect 93 4273 107 4287
rect 33 4053 47 4067
rect 293 4653 307 4667
rect 353 5074 367 5088
rect 393 5074 407 5088
rect 433 5074 447 5088
rect 353 5033 367 5047
rect 333 5013 347 5027
rect 693 5293 707 5307
rect 973 5293 987 5307
rect 1033 5353 1047 5367
rect 1013 5273 1027 5287
rect 633 5074 647 5088
rect 533 5032 547 5046
rect 673 5073 687 5087
rect 513 4993 527 5007
rect 573 4993 587 5007
rect 653 4993 667 5007
rect 413 4913 427 4927
rect 373 4854 387 4868
rect 693 4973 707 4987
rect 692 4933 706 4947
rect 713 4933 727 4947
rect 573 4893 587 4907
rect 673 4893 687 4907
rect 453 4853 467 4867
rect 513 4854 527 4868
rect 613 4853 627 4867
rect 813 5074 827 5088
rect 933 5074 947 5088
rect 973 5074 987 5088
rect 773 5032 787 5046
rect 733 4913 747 4927
rect 713 4853 727 4867
rect 453 4812 467 4826
rect 493 4812 507 4826
rect 533 4812 547 4826
rect 573 4812 587 4826
rect 693 4812 707 4826
rect 853 4933 867 4947
rect 813 4854 827 4868
rect 993 4933 1007 4947
rect 993 4912 1007 4926
rect 953 4873 967 4887
rect 933 4853 947 4867
rect 1113 5332 1127 5346
rect 1073 5193 1087 5207
rect 1093 5133 1107 5147
rect 1313 5473 1327 5487
rect 1273 5374 1287 5388
rect 1713 5733 1727 5747
rect 1533 5713 1547 5727
rect 1413 5633 1427 5647
rect 1473 5633 1487 5647
rect 1353 5453 1367 5467
rect 1453 5552 1467 5566
rect 1633 5673 1647 5687
rect 1553 5594 1567 5608
rect 1593 5594 1607 5608
rect 1553 5553 1567 5567
rect 1813 5813 1827 5827
rect 1973 5852 1987 5866
rect 2293 6114 2307 6128
rect 2213 6073 2227 6087
rect 2313 6072 2327 6086
rect 2153 6033 2167 6047
rect 2313 5993 2327 6007
rect 2133 5913 2147 5927
rect 2233 5894 2247 5908
rect 2273 5894 2287 5908
rect 2413 6253 2427 6267
rect 2513 6193 2527 6207
rect 2433 6072 2447 6086
rect 2573 6114 2587 6128
rect 2613 6114 2627 6128
rect 2553 6073 2567 6087
rect 2533 6033 2547 6047
rect 2353 5973 2367 5987
rect 2393 5953 2407 5967
rect 2373 5913 2387 5927
rect 2113 5852 2127 5866
rect 1973 5813 1987 5827
rect 1873 5773 1887 5787
rect 1793 5733 1807 5747
rect 1892 5673 1906 5687
rect 1913 5673 1927 5687
rect 1893 5613 1907 5627
rect 1873 5594 1887 5608
rect 2173 5852 2187 5866
rect 2173 5793 2187 5807
rect 2153 5773 2167 5787
rect 2013 5753 2027 5767
rect 2053 5753 2067 5767
rect 2013 5713 2027 5727
rect 2053 5713 2067 5727
rect 2032 5673 2046 5687
rect 2053 5673 2067 5687
rect 2053 5613 2067 5627
rect 2293 5852 2307 5866
rect 2333 5852 2347 5866
rect 2373 5853 2387 5867
rect 2253 5773 2267 5787
rect 2233 5733 2247 5747
rect 1993 5573 2007 5587
rect 1713 5552 1727 5566
rect 1753 5552 1767 5566
rect 1893 5552 1907 5566
rect 1973 5553 1987 5567
rect 1533 5533 1547 5547
rect 1613 5533 1627 5547
rect 1653 5513 1667 5527
rect 1413 5413 1427 5427
rect 1453 5373 1467 5387
rect 1533 5374 1547 5388
rect 1573 5374 1587 5388
rect 1193 5233 1207 5247
rect 1293 5332 1307 5346
rect 1413 5332 1427 5346
rect 1453 5332 1467 5346
rect 1353 5233 1367 5247
rect 1613 5373 1627 5387
rect 1873 5453 1887 5467
rect 1693 5374 1707 5388
rect 1173 5153 1187 5167
rect 1253 5153 1267 5167
rect 1573 5153 1587 5167
rect 1133 5074 1147 5088
rect 1673 5273 1687 5287
rect 1753 5332 1767 5346
rect 1813 5332 1827 5346
rect 1713 5213 1727 5227
rect 1613 5113 1627 5127
rect 1693 5113 1707 5127
rect 1273 5093 1287 5107
rect 1373 5093 1387 5107
rect 1193 5074 1207 5088
rect 1233 5074 1247 5088
rect 1113 5032 1127 5046
rect 1173 5033 1187 5047
rect 1613 5074 1627 5088
rect 1673 5073 1687 5087
rect 1513 5053 1527 5067
rect 1193 4973 1207 4987
rect 1433 4993 1447 5007
rect 1593 5032 1607 5046
rect 1253 4933 1267 4947
rect 1513 4933 1527 4947
rect 1473 4913 1487 4927
rect 1233 4893 1247 4907
rect 1313 4893 1327 4907
rect 1053 4873 1067 4887
rect 1033 4854 1047 4868
rect 613 4793 627 4807
rect 653 4793 667 4807
rect 753 4793 767 4807
rect 833 4793 847 4807
rect 353 4753 367 4767
rect 753 4753 767 4767
rect 453 4693 467 4707
rect 313 4613 327 4627
rect 353 4573 367 4587
rect 393 4554 407 4568
rect 433 4554 447 4568
rect 293 4512 307 4526
rect 373 4512 387 4526
rect 433 4513 447 4527
rect 973 4812 987 4826
rect 933 4773 947 4787
rect 1013 4773 1027 4787
rect 833 4673 847 4687
rect 593 4653 607 4667
rect 513 4613 527 4627
rect 473 4554 487 4568
rect 553 4554 567 4568
rect 273 4473 287 4487
rect 333 4473 347 4487
rect 393 4473 407 4487
rect 453 4473 467 4487
rect 333 4433 347 4447
rect 333 4393 347 4407
rect 193 4353 207 4367
rect 253 4334 267 4348
rect 313 4333 327 4347
rect 193 4292 207 4306
rect 233 4292 247 4306
rect 273 4292 287 4306
rect 153 4273 167 4287
rect 113 4233 127 4247
rect 293 4213 307 4227
rect 273 4113 287 4127
rect 113 4034 127 4048
rect 153 4034 167 4048
rect 213 4034 227 4048
rect 253 4034 267 4048
rect 33 3992 47 4006
rect 93 3993 107 4007
rect 133 3993 147 4007
rect 113 3953 127 3967
rect 153 3772 167 3786
rect 193 3772 207 3786
rect 533 4512 547 4526
rect 473 4393 487 4407
rect 393 4334 407 4348
rect 433 4334 447 4348
rect 573 4333 587 4347
rect 333 4293 347 4307
rect 413 4273 427 4287
rect 533 4292 547 4306
rect 573 4292 587 4306
rect 1073 4853 1087 4867
rect 1133 4854 1147 4868
rect 1073 4812 1087 4826
rect 1113 4812 1127 4826
rect 1113 4773 1127 4787
rect 1173 4773 1187 4787
rect 673 4554 687 4568
rect 1053 4554 1067 4568
rect 1093 4554 1107 4568
rect 1193 4554 1207 4568
rect 1273 4854 1287 4868
rect 1393 4853 1407 4867
rect 1653 5033 1667 5047
rect 1633 4873 1647 4887
rect 1613 4854 1627 4868
rect 1933 5173 1947 5187
rect 2053 5552 2067 5566
rect 2153 5552 2167 5566
rect 2193 5552 2207 5566
rect 2173 5513 2187 5527
rect 2213 5513 2227 5527
rect 2132 5473 2146 5487
rect 2153 5473 2167 5487
rect 2093 5413 2107 5427
rect 2493 5933 2507 5947
rect 2453 5894 2467 5908
rect 2433 5852 2447 5866
rect 2393 5733 2407 5747
rect 2473 5733 2487 5747
rect 2253 5713 2267 5727
rect 2293 5713 2307 5727
rect 2373 5673 2387 5687
rect 2253 5593 2267 5607
rect 2293 5594 2307 5608
rect 2333 5594 2347 5608
rect 2313 5552 2327 5566
rect 2433 5633 2447 5647
rect 2393 5594 2407 5608
rect 2493 5713 2507 5727
rect 2333 5513 2347 5527
rect 2373 5513 2387 5527
rect 2333 5453 2347 5467
rect 2253 5433 2267 5447
rect 2293 5433 2307 5447
rect 2193 5413 2207 5427
rect 2233 5413 2247 5427
rect 2133 5374 2147 5388
rect 2173 5374 2187 5388
rect 2153 5353 2167 5367
rect 2013 5273 2027 5287
rect 2053 5253 2067 5267
rect 1813 5093 1827 5107
rect 1693 5032 1707 5046
rect 1773 4993 1787 5007
rect 1853 5074 1867 5088
rect 1913 5074 1927 5088
rect 1953 5074 1967 5088
rect 1993 5074 2007 5088
rect 1893 5032 1907 5046
rect 1853 4993 1867 5007
rect 1813 4973 1827 4987
rect 1933 4973 1947 4987
rect 1873 4933 1887 4947
rect 1733 4913 1747 4927
rect 1733 4892 1747 4906
rect 1813 4893 1827 4907
rect 1733 4852 1747 4866
rect 1853 4854 1867 4868
rect 1293 4812 1307 4826
rect 1333 4812 1347 4826
rect 1393 4812 1407 4826
rect 1353 4773 1367 4787
rect 1313 4633 1327 4647
rect 993 4533 1007 4547
rect 793 4473 807 4487
rect 733 4453 747 4467
rect 693 4433 707 4447
rect 653 4413 667 4427
rect 373 4213 387 4227
rect 473 4213 487 4227
rect 593 4213 607 4227
rect 433 4133 447 4147
rect 353 4113 367 4127
rect 313 4073 327 4087
rect 393 4073 407 4087
rect 353 4034 367 4048
rect 293 3993 307 4007
rect 333 3992 347 4006
rect 373 3953 387 3967
rect 393 3933 407 3947
rect 353 3833 367 3847
rect 253 3753 267 3767
rect 293 3753 307 3767
rect 113 3713 127 3727
rect 153 3713 167 3727
rect 193 3713 207 3727
rect 93 3514 107 3528
rect 133 3472 147 3486
rect 193 3673 207 3687
rect 153 3453 167 3467
rect 133 3373 147 3387
rect 93 3252 107 3266
rect 113 3013 127 3027
rect 153 2952 167 2966
rect 133 2853 147 2867
rect 253 3553 267 3567
rect 293 3473 307 3487
rect 233 3453 247 3467
rect 293 3433 307 3447
rect 193 3293 207 3307
rect 273 3293 287 3307
rect 253 3113 267 3127
rect 253 2994 267 3008
rect 293 2952 307 2966
rect 213 2893 227 2907
rect 93 2732 107 2746
rect 33 2673 47 2687
rect 13 2633 27 2647
rect 53 2573 67 2587
rect 53 2513 67 2527
rect 53 2473 67 2487
rect 553 4093 567 4107
rect 473 4053 487 4067
rect 513 4034 527 4048
rect 593 4053 607 4067
rect 653 4034 667 4048
rect 533 3992 547 4006
rect 593 3973 607 3987
rect 493 3933 507 3947
rect 573 3853 587 3867
rect 433 3833 447 3847
rect 473 3753 487 3767
rect 413 3673 427 3687
rect 393 3553 407 3567
rect 453 3553 467 3567
rect 353 3514 367 3528
rect 393 3514 407 3528
rect 433 3514 447 3528
rect 333 3473 347 3487
rect 373 3472 387 3486
rect 433 3472 447 3486
rect 413 3453 427 3467
rect 653 3814 667 3828
rect 833 4413 847 4427
rect 713 4334 727 4348
rect 793 4334 807 4348
rect 833 4334 847 4348
rect 913 4473 927 4487
rect 1073 4453 1087 4467
rect 1213 4413 1227 4427
rect 973 4373 987 4387
rect 1293 4373 1307 4387
rect 893 4353 907 4367
rect 933 4353 947 4367
rect 873 4334 887 4348
rect 813 4292 827 4306
rect 1033 4333 1047 4347
rect 1133 4334 1147 4348
rect 773 3992 787 4006
rect 713 3973 727 3987
rect 713 3913 727 3927
rect 693 3813 707 3827
rect 773 3813 787 3827
rect 833 4233 847 4247
rect 873 4233 887 4247
rect 873 4093 887 4107
rect 833 4033 847 4047
rect 993 4292 1007 4306
rect 1033 4292 1047 4306
rect 1153 4292 1167 4306
rect 953 4273 967 4287
rect 1113 4273 1127 4287
rect 1253 4292 1267 4306
rect 1293 4292 1307 4306
rect 1273 4253 1287 4267
rect 1193 4213 1207 4227
rect 1493 4812 1507 4826
rect 1593 4812 1607 4826
rect 1633 4812 1647 4826
rect 1693 4812 1707 4826
rect 1753 4812 1767 4826
rect 1433 4773 1447 4787
rect 1593 4773 1607 4787
rect 1733 4773 1747 4787
rect 1513 4713 1527 4727
rect 1473 4693 1487 4707
rect 1453 4673 1467 4687
rect 1373 4453 1387 4467
rect 1453 4493 1467 4507
rect 1453 4453 1467 4467
rect 1413 4413 1427 4427
rect 1373 4334 1387 4348
rect 1413 4213 1427 4227
rect 1313 4133 1327 4147
rect 1453 4333 1467 4347
rect 1353 4113 1367 4127
rect 913 4034 927 4048
rect 953 4034 967 4048
rect 993 4034 1007 4048
rect 833 3992 847 4006
rect 873 3993 887 4007
rect 933 3992 947 4006
rect 1033 4033 1047 4047
rect 1093 4034 1107 4048
rect 953 3953 967 3967
rect 993 3953 1007 3967
rect 933 3893 947 3907
rect 693 3773 707 3787
rect 593 3713 607 3727
rect 573 3673 587 3687
rect 693 3633 707 3647
rect 573 3553 587 3567
rect 493 3514 507 3528
rect 533 3514 547 3528
rect 573 3514 587 3528
rect 613 3514 627 3528
rect 673 3514 687 3528
rect 713 3514 727 3528
rect 513 3472 527 3486
rect 553 3472 567 3486
rect 593 3473 607 3487
rect 432 3433 446 3447
rect 453 3433 467 3447
rect 333 3413 347 3427
rect 393 3413 407 3427
rect 533 3413 547 3427
rect 373 3233 387 3247
rect 313 2853 327 2867
rect 213 2774 227 2788
rect 213 2713 227 2727
rect 353 2733 367 2747
rect 333 2713 347 2727
rect 273 2673 287 2687
rect 153 2473 167 2487
rect 33 2333 47 2347
rect 33 2293 47 2307
rect 33 2213 47 2227
rect 13 1833 27 1847
rect 253 2533 267 2547
rect 333 2533 347 2547
rect 293 2474 307 2488
rect 193 2433 207 2447
rect 173 2333 187 2347
rect 113 2293 127 2307
rect 113 2254 127 2268
rect 133 2212 147 2226
rect 93 2193 107 2207
rect 73 2053 87 2067
rect 53 1993 67 2007
rect 93 1993 107 2007
rect 73 1953 87 1967
rect 273 2432 287 2446
rect 273 2293 287 2307
rect 293 2273 307 2287
rect 233 2212 247 2226
rect 173 2093 187 2107
rect 493 3252 507 3266
rect 433 3233 447 3247
rect 433 3193 447 3207
rect 693 3472 707 3486
rect 653 3433 667 3447
rect 613 3413 627 3427
rect 553 3393 567 3407
rect 613 3294 627 3308
rect 773 3514 787 3528
rect 773 3473 787 3487
rect 553 3252 567 3266
rect 533 3133 547 3147
rect 733 3252 747 3266
rect 753 3213 767 3227
rect 673 3193 687 3207
rect 653 3093 667 3107
rect 553 3073 567 3087
rect 413 3033 427 3047
rect 553 3033 567 3047
rect 513 3013 527 3027
rect 593 2994 607 3008
rect 633 2994 647 3008
rect 513 2933 527 2947
rect 573 2933 587 2947
rect 453 2893 467 2907
rect 573 2853 587 2867
rect 513 2813 527 2827
rect 393 2774 407 2788
rect 453 2774 467 2788
rect 373 2673 387 2687
rect 493 2773 507 2787
rect 493 2693 507 2707
rect 733 3053 747 3067
rect 693 3013 707 3027
rect 773 2993 787 3007
rect 653 2953 667 2967
rect 713 2952 727 2966
rect 833 3772 847 3786
rect 933 3653 947 3667
rect 833 3633 847 3647
rect 873 3514 887 3528
rect 853 3472 867 3486
rect 893 3393 907 3407
rect 853 3333 867 3347
rect 893 3294 907 3308
rect 833 3133 847 3147
rect 813 3073 827 3087
rect 1093 3913 1107 3927
rect 1033 3893 1047 3907
rect 973 3873 987 3887
rect 1013 3814 1027 3828
rect 1053 3814 1067 3828
rect 973 3772 987 3786
rect 1013 3753 1027 3767
rect 1033 3713 1047 3727
rect 1273 4034 1287 4048
rect 1453 4073 1467 4087
rect 1533 4653 1547 4667
rect 1713 4653 1727 4667
rect 1513 4633 1527 4647
rect 1573 4554 1587 4568
rect 1633 4554 1647 4568
rect 1673 4554 1687 4568
rect 1733 4613 1747 4627
rect 1893 4913 1907 4927
rect 2033 5173 2047 5187
rect 2253 5393 2267 5407
rect 2393 5393 2407 5407
rect 2193 5333 2207 5347
rect 2273 5332 2287 5346
rect 2173 5253 2187 5267
rect 2153 5193 2167 5207
rect 2313 5273 2327 5287
rect 2213 5253 2227 5267
rect 2193 5233 2207 5247
rect 2173 5113 2187 5127
rect 2113 5074 2127 5088
rect 2153 5073 2167 5087
rect 2032 5032 2046 5046
rect 2093 5032 2107 5046
rect 2053 5013 2067 5027
rect 2013 4973 2027 4987
rect 1993 4933 2007 4947
rect 1973 4893 1987 4907
rect 1993 4873 2007 4887
rect 2013 4854 2027 4868
rect 2093 4854 2107 4868
rect 1893 4813 1907 4827
rect 1993 4812 2007 4826
rect 2373 5373 2387 5387
rect 2353 5253 2367 5267
rect 2333 5233 2347 5247
rect 2453 5552 2467 5566
rect 2513 5453 2527 5467
rect 2493 5433 2507 5447
rect 2453 5374 2467 5388
rect 2393 5293 2407 5307
rect 2393 5272 2407 5286
rect 2373 5213 2387 5227
rect 2333 5173 2347 5187
rect 2253 5113 2267 5127
rect 2213 5074 2227 5088
rect 2253 5073 2267 5087
rect 2293 5074 2307 5088
rect 2353 5074 2367 5088
rect 2473 5332 2487 5346
rect 2473 5293 2487 5307
rect 2433 5193 2447 5207
rect 2433 5093 2447 5107
rect 2213 5033 2227 5047
rect 2333 5033 2347 5047
rect 2233 4993 2247 5007
rect 2353 4993 2367 5007
rect 2213 4973 2227 4987
rect 2193 4813 2207 4827
rect 2313 4933 2327 4947
rect 2292 4893 2306 4907
rect 2313 4893 2327 4907
rect 2113 4773 2127 4787
rect 2213 4773 2227 4787
rect 2313 4812 2327 4826
rect 2413 5032 2427 5046
rect 2553 6013 2567 6027
rect 2633 6053 2647 6067
rect 2593 5973 2607 5987
rect 2593 5894 2607 5908
rect 2573 5813 2587 5827
rect 2713 6193 2727 6207
rect 2753 6173 2767 6187
rect 2733 6053 2747 6067
rect 2733 5993 2747 6007
rect 2853 6473 2867 6487
rect 2893 6473 2907 6487
rect 3033 6414 3047 6428
rect 2833 6372 2847 6386
rect 2873 6333 2887 6347
rect 3053 6313 3067 6327
rect 3013 6193 3027 6207
rect 2993 6173 3007 6187
rect 3053 6173 3067 6187
rect 2873 6153 2887 6167
rect 2913 6153 2927 6167
rect 2813 6114 2827 6128
rect 2913 6072 2927 6086
rect 2813 6033 2827 6047
rect 2853 6033 2867 6047
rect 3013 6114 3027 6128
rect 2993 6072 3007 6086
rect 2993 6051 3007 6065
rect 2933 5993 2947 6007
rect 2933 5913 2947 5927
rect 2793 5893 2807 5907
rect 2833 5894 2847 5908
rect 2893 5894 2907 5908
rect 2613 5793 2627 5807
rect 2673 5793 2687 5807
rect 2793 5852 2807 5866
rect 2753 5753 2767 5767
rect 2753 5732 2767 5746
rect 2713 5693 2727 5707
rect 2693 5653 2707 5667
rect 2553 5633 2567 5647
rect 2613 5594 2627 5608
rect 2653 5594 2667 5608
rect 2553 5553 2567 5567
rect 2593 5513 2607 5527
rect 2633 5513 2647 5527
rect 2613 5473 2627 5487
rect 2653 5473 2667 5487
rect 2653 5413 2667 5427
rect 2613 5374 2627 5388
rect 2593 5332 2607 5346
rect 3053 6033 3067 6047
rect 3073 5993 3087 6007
rect 3053 5953 3067 5967
rect 3033 5933 3047 5947
rect 3193 6473 3207 6487
rect 3273 6453 3287 6467
rect 3193 6414 3207 6428
rect 3173 6372 3187 6386
rect 3213 6353 3227 6367
rect 3113 6293 3127 6307
rect 3113 6253 3127 6267
rect 3153 6153 3167 6167
rect 3113 6113 3127 6127
rect 3173 6133 3187 6147
rect 3193 6114 3207 6128
rect 3113 6072 3127 6086
rect 3173 6072 3187 6086
rect 3693 6493 3707 6507
rect 3973 6493 3987 6507
rect 5573 6493 5587 6507
rect 6133 6493 6147 6507
rect 3433 6473 3447 6487
rect 3513 6473 3527 6487
rect 3333 6414 3347 6428
rect 3373 6414 3387 6428
rect 3353 6353 3367 6367
rect 3273 6333 3287 6347
rect 3273 6253 3287 6267
rect 3353 6233 3367 6247
rect 3313 6173 3327 6187
rect 3413 6153 3427 6167
rect 3273 6073 3287 6087
rect 3333 6072 3347 6086
rect 3373 6072 3387 6086
rect 3413 6072 3427 6086
rect 3253 6013 3267 6027
rect 3413 6013 3427 6027
rect 3233 5973 3247 5987
rect 3213 5953 3227 5967
rect 3253 5953 3267 5967
rect 3093 5914 3107 5928
rect 3173 5913 3187 5927
rect 3053 5894 3067 5908
rect 3093 5893 3107 5907
rect 2873 5852 2887 5866
rect 2913 5852 2927 5866
rect 2993 5852 3007 5866
rect 2833 5833 2847 5847
rect 2873 5831 2887 5845
rect 2853 5793 2867 5807
rect 2793 5673 2807 5687
rect 2813 5594 2827 5608
rect 2713 5573 2727 5587
rect 2773 5513 2787 5527
rect 2713 5433 2727 5447
rect 2733 5413 2747 5427
rect 2693 5374 2707 5388
rect 2773 5374 2787 5388
rect 2813 5373 2827 5387
rect 2533 5293 2547 5307
rect 2513 5253 2527 5267
rect 2673 5332 2687 5346
rect 2713 5332 2727 5346
rect 2753 5293 2767 5307
rect 2653 5233 2667 5247
rect 2633 5193 2647 5207
rect 2553 5074 2567 5088
rect 2593 5074 2607 5088
rect 2673 5213 2687 5227
rect 2753 5193 2767 5207
rect 2673 5153 2687 5167
rect 2653 5093 2667 5107
rect 2493 5032 2507 5046
rect 2533 5032 2547 5046
rect 2473 4993 2487 5007
rect 2453 4913 2467 4927
rect 2373 4793 2387 4807
rect 2273 4753 2287 4767
rect 2353 4753 2367 4767
rect 2353 4713 2367 4727
rect 2113 4653 2127 4667
rect 2373 4693 2387 4707
rect 2373 4653 2387 4667
rect 2353 4633 2367 4647
rect 2313 4613 2327 4627
rect 1973 4573 1987 4587
rect 2093 4573 2107 4587
rect 1553 4512 1567 4526
rect 1533 4493 1547 4507
rect 1513 4453 1527 4467
rect 1933 4553 1947 4567
rect 2013 4554 2027 4568
rect 2133 4554 2147 4568
rect 2273 4554 2287 4568
rect 2353 4573 2367 4587
rect 2473 4812 2487 4826
rect 2433 4653 2447 4667
rect 2393 4593 2407 4607
rect 2373 4554 2387 4568
rect 1693 4512 1707 4526
rect 1793 4513 1807 4527
rect 1853 4512 1867 4526
rect 1773 4433 1787 4447
rect 1633 4393 1647 4407
rect 1673 4393 1687 4407
rect 1493 4334 1507 4348
rect 1613 4333 1627 4347
rect 1733 4334 1747 4348
rect 1833 4393 1847 4407
rect 1813 4353 1827 4367
rect 1673 4292 1687 4306
rect 1713 4292 1727 4306
rect 1753 4173 1767 4187
rect 1733 4113 1747 4127
rect 1453 3992 1467 4006
rect 1373 3953 1387 3967
rect 1333 3873 1347 3887
rect 1193 3853 1207 3867
rect 1253 3833 1267 3847
rect 1133 3813 1147 3827
rect 1193 3814 1207 3828
rect 1093 3673 1107 3687
rect 1273 3813 1287 3827
rect 1413 3913 1427 3927
rect 1373 3833 1387 3847
rect 1473 3893 1487 3907
rect 1433 3833 1447 3847
rect 1273 3772 1287 3786
rect 1313 3772 1327 3786
rect 1353 3772 1367 3786
rect 1413 3772 1427 3786
rect 1173 3673 1187 3687
rect 1253 3593 1267 3607
rect 1133 3573 1147 3587
rect 1313 3573 1327 3587
rect 1013 3514 1027 3528
rect 1053 3513 1067 3527
rect 1093 3513 1107 3527
rect 1133 3514 1147 3528
rect 1173 3514 1187 3528
rect 1213 3514 1227 3528
rect 1273 3514 1287 3528
rect 953 3473 967 3487
rect 993 3433 1007 3447
rect 1073 3492 1087 3506
rect 993 3333 1007 3347
rect 1033 3333 1047 3347
rect 993 3294 1007 3308
rect 1033 3294 1047 3308
rect 1113 3472 1127 3486
rect 1193 3473 1207 3487
rect 1293 3473 1307 3487
rect 1093 3294 1107 3308
rect 1133 3294 1147 3308
rect 1013 3233 1027 3247
rect 1073 3233 1087 3247
rect 1093 3113 1107 3127
rect 1053 3093 1067 3107
rect 1093 3073 1107 3087
rect 933 3053 947 3067
rect 833 3013 847 3027
rect 1013 3013 1027 3027
rect 793 2952 807 2966
rect 773 2853 787 2867
rect 633 2813 647 2827
rect 613 2774 627 2788
rect 593 2732 607 2746
rect 513 2653 527 2667
rect 393 2633 407 2647
rect 633 2633 647 2647
rect 433 2613 447 2627
rect 593 2613 607 2627
rect 393 2573 407 2587
rect 373 2513 387 2527
rect 573 2553 587 2567
rect 473 2513 487 2527
rect 533 2474 547 2488
rect 413 2432 427 2446
rect 493 2353 507 2367
rect 353 2293 367 2307
rect 413 2293 427 2307
rect 373 2273 387 2287
rect 473 2253 487 2267
rect 473 2212 487 2226
rect 433 2193 447 2207
rect 333 2173 347 2187
rect 393 2172 407 2186
rect 233 1954 247 1968
rect 293 1954 307 1968
rect 433 2093 447 2107
rect 413 1913 427 1927
rect 353 1853 367 1867
rect 273 1813 287 1827
rect 113 1753 127 1767
rect 213 1753 227 1767
rect 93 1692 107 1706
rect 413 1793 427 1807
rect 313 1753 327 1767
rect 413 1753 427 1767
rect 773 2732 787 2746
rect 733 2713 747 2727
rect 733 2653 747 2667
rect 673 2513 687 2527
rect 693 2474 707 2488
rect 593 2433 607 2447
rect 573 2293 587 2307
rect 653 2413 667 2427
rect 693 2393 707 2407
rect 853 2913 867 2927
rect 833 2853 847 2867
rect 933 2993 947 3007
rect 1053 2994 1067 3008
rect 913 2813 927 2827
rect 993 2952 1007 2966
rect 993 2913 1007 2927
rect 1033 2873 1047 2887
rect 993 2833 1007 2847
rect 853 2774 867 2788
rect 893 2774 907 2788
rect 893 2732 907 2746
rect 793 2553 807 2567
rect 833 2474 847 2488
rect 773 2393 787 2407
rect 733 2353 747 2367
rect 773 2313 787 2327
rect 573 2254 587 2268
rect 753 2273 767 2287
rect 553 2212 567 2226
rect 493 2173 507 2187
rect 572 2173 586 2187
rect 593 2173 607 2187
rect 573 2133 587 2147
rect 453 1912 467 1926
rect 453 1813 467 1827
rect 433 1733 447 1747
rect 213 1673 227 1687
rect 253 1673 267 1687
rect 153 1613 167 1627
rect 33 1493 47 1507
rect 173 1493 187 1507
rect 13 1433 27 1447
rect 13 1392 27 1406
rect 93 1392 107 1406
rect 153 1353 167 1367
rect 113 1214 127 1228
rect 93 1172 107 1186
rect 213 1453 227 1467
rect 193 1213 207 1227
rect 273 1434 287 1448
rect 353 1692 367 1706
rect 413 1673 427 1687
rect 453 1673 467 1687
rect 373 1493 387 1507
rect 293 1433 307 1447
rect 413 1434 427 1448
rect 253 1373 267 1387
rect 353 1373 367 1387
rect 273 1214 287 1228
rect 213 1172 227 1186
rect 253 1172 267 1186
rect 293 1133 307 1147
rect 193 1073 207 1087
rect 133 1033 147 1047
rect 173 1033 187 1047
rect 133 973 147 987
rect 333 993 347 1007
rect 313 973 327 987
rect 233 913 247 927
rect 273 914 287 928
rect 333 953 347 967
rect 313 913 327 927
rect 153 853 167 867
rect 393 1353 407 1367
rect 393 1233 407 1247
rect 493 1912 507 1926
rect 533 1853 547 1867
rect 533 1734 547 1748
rect 553 1693 567 1707
rect 513 1553 527 1567
rect 493 1434 507 1448
rect 493 1373 507 1387
rect 493 1313 507 1327
rect 473 1293 487 1307
rect 413 1172 427 1186
rect 453 1172 467 1186
rect 493 1172 507 1186
rect 533 1493 547 1507
rect 533 1453 547 1467
rect 713 2212 727 2226
rect 653 2093 667 2107
rect 593 2033 607 2047
rect 573 1673 587 1687
rect 553 1434 567 1448
rect 633 1993 647 2007
rect 833 2254 847 2268
rect 773 2013 787 2027
rect 853 1954 867 1968
rect 613 1853 627 1867
rect 713 1912 727 1926
rect 753 1913 767 1927
rect 633 1833 647 1847
rect 833 1912 847 1926
rect 833 1873 847 1887
rect 653 1793 667 1807
rect 793 1793 807 1807
rect 813 1773 827 1787
rect 693 1734 707 1748
rect 753 1734 767 1748
rect 653 1673 667 1687
rect 613 1553 627 1567
rect 713 1692 727 1706
rect 813 1734 827 1748
rect 933 2773 947 2787
rect 1013 2774 1027 2788
rect 1053 2774 1067 2788
rect 913 2693 927 2707
rect 993 2732 1007 2746
rect 1073 2733 1087 2747
rect 933 2633 947 2647
rect 1033 2533 1047 2547
rect 1013 2473 1027 2487
rect 933 2432 947 2446
rect 1013 2432 1027 2446
rect 913 2393 927 2407
rect 973 2393 987 2407
rect 953 2254 967 2268
rect 1013 2254 1027 2268
rect 1013 2213 1027 2227
rect 973 2173 987 2187
rect 973 2113 987 2127
rect 1153 3252 1167 3266
rect 1153 3213 1167 3227
rect 1273 3353 1287 3367
rect 1213 3333 1227 3347
rect 1593 4034 1607 4048
rect 1632 4033 1646 4047
rect 1653 4034 1667 4048
rect 1693 4034 1707 4048
rect 1773 4034 1787 4048
rect 1573 3992 1587 4006
rect 1633 3992 1647 4006
rect 1713 3992 1727 4006
rect 1753 3992 1767 4006
rect 1653 3953 1667 3967
rect 1653 3932 1667 3946
rect 1633 3913 1647 3927
rect 1533 3853 1547 3867
rect 1493 3833 1507 3847
rect 1493 3772 1507 3786
rect 1493 3593 1507 3607
rect 1453 3533 1467 3547
rect 1333 3453 1347 3467
rect 1313 3353 1327 3367
rect 1333 3333 1347 3347
rect 1293 3313 1307 3327
rect 1393 3313 1407 3327
rect 1473 3353 1487 3367
rect 1213 3252 1227 3266
rect 1253 3252 1267 3266
rect 1213 3113 1227 3127
rect 1133 3093 1147 3107
rect 1153 3053 1167 3067
rect 1153 3013 1167 3027
rect 1393 3013 1407 3027
rect 1273 2994 1287 3008
rect 1313 2994 1327 3008
rect 1473 3193 1487 3207
rect 1453 3173 1467 3187
rect 1893 4353 1907 4367
rect 1993 4512 2007 4526
rect 2253 4513 2267 4527
rect 2153 4493 2167 4507
rect 2253 4453 2267 4467
rect 2033 4433 2047 4447
rect 2233 4433 2247 4447
rect 1973 4334 1987 4348
rect 2213 4334 2227 4348
rect 2193 4313 2207 4327
rect 1833 4293 1847 4307
rect 1913 4292 1927 4306
rect 2093 4292 2107 4306
rect 2213 4292 2227 4306
rect 2033 4253 2047 4267
rect 2153 4253 2167 4267
rect 1833 4213 1847 4227
rect 1933 4073 1947 4087
rect 1873 4034 1887 4048
rect 1833 3992 1847 4006
rect 1813 3853 1827 3867
rect 1853 3853 1867 3867
rect 1593 3814 1607 3828
rect 1692 3814 1706 3828
rect 1613 3772 1627 3786
rect 1653 3772 1667 3786
rect 1553 3673 1567 3687
rect 1533 3533 1547 3547
rect 1713 3813 1727 3827
rect 1793 3814 1807 3828
rect 1873 3813 1887 3827
rect 1713 3772 1727 3786
rect 1813 3772 1827 3786
rect 1853 3772 1867 3786
rect 1693 3753 1707 3767
rect 1773 3753 1787 3767
rect 1733 3633 1747 3647
rect 1733 3573 1747 3587
rect 1973 3913 1987 3927
rect 2053 4033 2067 4047
rect 2093 4034 2107 4048
rect 2053 3933 2067 3947
rect 2133 3913 2147 3927
rect 2213 3913 2227 3927
rect 1993 3893 2007 3907
rect 2033 3893 2047 3907
rect 1953 3814 1967 3828
rect 1993 3813 2007 3827
rect 1893 3753 1907 3767
rect 1933 3753 1947 3767
rect 2013 3772 2027 3786
rect 2073 3772 2087 3786
rect 2193 3814 2207 3828
rect 1973 3733 1987 3747
rect 2133 3733 2147 3747
rect 2553 5013 2567 5027
rect 2553 4953 2567 4967
rect 2633 5032 2647 5046
rect 2633 4953 2647 4967
rect 2613 4913 2627 4927
rect 2553 4853 2567 4867
rect 2693 5074 2707 5088
rect 2713 5032 2727 5046
rect 2953 5813 2967 5827
rect 2953 5673 2967 5687
rect 2873 5594 2887 5608
rect 2913 5594 2927 5608
rect 2933 5552 2947 5566
rect 3113 5852 3127 5866
rect 3073 5813 3087 5827
rect 3153 5813 3167 5827
rect 3013 5713 3027 5727
rect 2993 5493 3007 5507
rect 2933 5473 2947 5487
rect 2973 5433 2987 5447
rect 2873 5393 2887 5407
rect 2933 5374 2947 5388
rect 2893 5293 2907 5307
rect 2853 5233 2867 5247
rect 2893 5173 2907 5187
rect 2833 5153 2847 5167
rect 2773 5093 2787 5107
rect 2813 5093 2827 5107
rect 2673 4993 2687 5007
rect 2653 4853 2667 4867
rect 2513 4593 2527 4607
rect 2473 4573 2487 4587
rect 2513 4554 2527 4568
rect 2393 4512 2407 4526
rect 2333 4473 2347 4487
rect 2373 4473 2387 4487
rect 2313 4453 2327 4467
rect 2453 4512 2467 4526
rect 2673 4833 2687 4847
rect 2613 4812 2627 4826
rect 2673 4812 2687 4826
rect 2573 4553 2587 4567
rect 2613 4554 2627 4568
rect 2553 4493 2567 4507
rect 2573 4433 2587 4447
rect 2413 4413 2427 4427
rect 2473 4413 2487 4427
rect 2553 4413 2567 4427
rect 2633 4413 2647 4427
rect 2873 5074 2887 5088
rect 2833 5032 2847 5046
rect 2913 5074 2927 5088
rect 2893 4993 2907 5007
rect 2973 5333 2987 5347
rect 3193 5893 3207 5907
rect 3253 5894 3267 5908
rect 3213 5852 3227 5866
rect 3293 5852 3307 5866
rect 3353 5833 3367 5847
rect 3173 5793 3187 5807
rect 3133 5773 3147 5787
rect 3373 5713 3387 5727
rect 3153 5673 3167 5687
rect 3133 5594 3147 5608
rect 3053 5552 3067 5566
rect 3093 5552 3107 5566
rect 3233 5653 3247 5667
rect 3333 5653 3347 5667
rect 3193 5613 3207 5627
rect 3193 5594 3207 5608
rect 3313 5613 3327 5627
rect 3273 5593 3287 5607
rect 3393 5693 3407 5707
rect 3373 5613 3387 5627
rect 3073 5493 3087 5507
rect 3153 5374 3167 5388
rect 3053 5233 3067 5247
rect 3273 5552 3287 5566
rect 3313 5552 3327 5566
rect 3373 5552 3387 5566
rect 3373 5513 3387 5527
rect 3213 5493 3227 5507
rect 3233 5413 3247 5427
rect 3333 5413 3347 5427
rect 3273 5374 3287 5388
rect 3333 5374 3347 5388
rect 3173 5273 3187 5287
rect 3093 5193 3107 5207
rect 3013 5133 3027 5147
rect 3093 5133 3107 5147
rect 3073 5074 3087 5088
rect 2953 5032 2967 5046
rect 2913 4973 2927 4987
rect 2793 4953 2807 4967
rect 2773 4913 2787 4927
rect 2833 4913 2847 4927
rect 2773 4854 2787 4868
rect 2873 4893 2887 4907
rect 3073 4973 3087 4987
rect 2913 4854 2927 4868
rect 2973 4854 2987 4868
rect 2833 4812 2847 4826
rect 2893 4812 2907 4826
rect 2933 4812 2947 4826
rect 2753 4793 2767 4807
rect 2973 4713 2987 4727
rect 3013 4873 3027 4887
rect 2753 4653 2767 4667
rect 2993 4653 3007 4667
rect 2713 4633 2727 4647
rect 2793 4554 2807 4568
rect 2873 4554 2887 4568
rect 2733 4473 2747 4487
rect 2693 4453 2707 4467
rect 2673 4353 2687 4367
rect 2713 4413 2727 4427
rect 2693 4333 2707 4347
rect 2293 4292 2307 4306
rect 2433 4292 2447 4306
rect 2473 4292 2487 4306
rect 2673 4292 2687 4306
rect 2373 4253 2387 4267
rect 2493 4253 2507 4267
rect 2613 4253 2627 4267
rect 2333 4193 2347 4207
rect 2393 4173 2407 4187
rect 2293 4053 2307 4067
rect 2273 3992 2287 4006
rect 2333 3992 2347 4006
rect 2273 3853 2287 3867
rect 2333 3853 2347 3867
rect 2273 3813 2287 3827
rect 2313 3814 2327 3828
rect 2253 3772 2267 3786
rect 2233 3693 2247 3707
rect 2253 3673 2267 3687
rect 2233 3653 2247 3667
rect 1933 3633 1947 3647
rect 1613 3514 1627 3528
rect 1693 3514 1707 3528
rect 1533 3433 1547 3447
rect 1633 3473 1647 3487
rect 1713 3472 1727 3486
rect 1853 3514 1867 3528
rect 1993 3514 2007 3528
rect 2093 3514 2107 3528
rect 2133 3514 2147 3528
rect 2173 3514 2187 3528
rect 1833 3472 1847 3486
rect 1733 3433 1747 3447
rect 1773 3433 1787 3447
rect 1533 3353 1547 3367
rect 1573 3373 1587 3387
rect 1553 3313 1567 3327
rect 1553 3252 1567 3266
rect 1593 3252 1607 3266
rect 1813 3373 1827 3387
rect 1813 3333 1827 3347
rect 1933 3472 1947 3486
rect 2013 3393 2027 3407
rect 2053 3393 2067 3407
rect 1873 3313 1887 3327
rect 1753 3252 1767 3266
rect 1633 3173 1647 3187
rect 1493 3133 1507 3147
rect 1713 3133 1727 3147
rect 1453 3113 1467 3127
rect 1193 2953 1207 2967
rect 1173 2893 1187 2907
rect 1113 2853 1127 2867
rect 1293 2933 1307 2947
rect 1293 2893 1307 2907
rect 1172 2833 1186 2847
rect 1193 2833 1207 2847
rect 1413 2993 1427 3007
rect 1693 3093 1707 3107
rect 1673 3053 1687 3067
rect 1513 3013 1527 3027
rect 1573 3013 1587 3027
rect 1553 2973 1567 2987
rect 1373 2953 1387 2967
rect 1313 2873 1327 2887
rect 1353 2873 1367 2887
rect 1393 2873 1407 2887
rect 1213 2732 1227 2746
rect 1293 2732 1307 2746
rect 1373 2732 1387 2746
rect 1373 2653 1387 2667
rect 1633 2933 1647 2947
rect 1573 2893 1587 2907
rect 1933 3252 1947 3266
rect 1993 3193 2007 3207
rect 1873 3173 1887 3187
rect 1753 3113 1767 3127
rect 1773 2994 1787 3008
rect 1813 2994 1827 3008
rect 1853 2993 1867 3007
rect 1713 2952 1727 2966
rect 1753 2952 1767 2966
rect 1853 2933 1867 2947
rect 1953 3133 1967 3147
rect 1913 2994 1927 3008
rect 2173 3433 2187 3447
rect 2133 3393 2147 3407
rect 2113 3293 2127 3307
rect 2093 3073 2107 3087
rect 2253 3413 2267 3427
rect 2213 3294 2227 3308
rect 2333 3772 2347 3786
rect 2453 4034 2467 4048
rect 2553 4034 2567 4048
rect 2553 3993 2567 4007
rect 2513 3913 2527 3927
rect 2433 3873 2447 3887
rect 2473 3853 2487 3867
rect 2673 4053 2687 4067
rect 2773 4453 2787 4467
rect 2833 4433 2847 4447
rect 2793 4334 2807 4348
rect 2733 4193 2747 4207
rect 2773 4093 2787 4107
rect 2753 4033 2767 4047
rect 2633 3893 2647 3907
rect 2513 3813 2527 3827
rect 2613 3813 2627 3827
rect 2453 3772 2467 3786
rect 2493 3772 2507 3786
rect 2533 3772 2547 3786
rect 2593 3772 2607 3786
rect 2633 3772 2647 3786
rect 2693 3992 2707 4006
rect 2853 4373 2867 4387
rect 2873 4353 2887 4367
rect 2933 4512 2947 4526
rect 2993 4473 3007 4487
rect 2933 4413 2947 4427
rect 2893 4333 2907 4347
rect 2973 4393 2987 4407
rect 2873 4313 2887 4327
rect 2873 4253 2887 4267
rect 2853 4233 2867 4247
rect 2953 4292 2967 4306
rect 3153 5093 3167 5107
rect 3133 5033 3147 5047
rect 3093 4873 3107 4887
rect 3053 4812 3067 4826
rect 3153 4793 3167 4807
rect 3253 5332 3267 5346
rect 3293 5332 3307 5346
rect 3193 5173 3207 5187
rect 3213 5173 3227 5187
rect 3253 5153 3267 5167
rect 3253 5113 3267 5127
rect 3313 5133 3327 5147
rect 3293 5093 3307 5107
rect 3273 5073 3287 5087
rect 3233 5032 3247 5046
rect 3233 4893 3247 4907
rect 3193 4793 3207 4807
rect 3173 4733 3187 4747
rect 3093 4713 3107 4727
rect 3033 4633 3047 4647
rect 3093 4573 3107 4587
rect 3173 4573 3187 4587
rect 3033 4512 3047 4526
rect 3073 4512 3087 4526
rect 3153 4493 3167 4507
rect 3113 4473 3127 4487
rect 3093 4353 3107 4367
rect 3073 4253 3087 4267
rect 3173 4393 3187 4407
rect 3013 4213 3027 4227
rect 3033 4193 3047 4207
rect 2913 4133 2927 4147
rect 2913 4093 2927 4107
rect 3113 4213 3127 4227
rect 3073 4173 3087 4187
rect 2873 4053 2887 4067
rect 2913 4053 2927 4067
rect 3033 4053 3047 4067
rect 2993 4034 3007 4048
rect 2813 3953 2827 3967
rect 2773 3873 2787 3887
rect 2713 3814 2727 3828
rect 2753 3814 2767 3828
rect 2653 3753 2667 3767
rect 2753 3753 2767 3767
rect 2513 3693 2527 3707
rect 2393 3613 2407 3627
rect 2493 3613 2507 3627
rect 2433 3593 2447 3607
rect 2393 3514 2407 3528
rect 2413 3413 2427 3427
rect 2353 3373 2367 3387
rect 2273 3333 2287 3347
rect 2393 3333 2407 3347
rect 2453 3333 2467 3347
rect 2253 3293 2267 3307
rect 2353 3293 2367 3307
rect 2133 3252 2147 3266
rect 2193 3252 2207 3266
rect 2233 3252 2247 3266
rect 2333 3252 2347 3266
rect 2393 3233 2407 3247
rect 2273 3173 2287 3187
rect 2273 3113 2287 3127
rect 2133 3033 2147 3047
rect 2233 3013 2247 3027
rect 2173 2994 2187 3008
rect 2233 2994 2247 3008
rect 2373 3093 2387 3107
rect 2313 2994 2327 3008
rect 1933 2952 1947 2966
rect 1993 2952 2007 2966
rect 2073 2952 2087 2966
rect 1873 2913 1887 2927
rect 1933 2913 1947 2927
rect 1793 2893 1807 2907
rect 1433 2853 1447 2867
rect 1493 2833 1507 2847
rect 1533 2813 1547 2827
rect 1433 2732 1447 2746
rect 1513 2732 1527 2746
rect 1593 2873 1607 2887
rect 1672 2873 1686 2887
rect 1693 2873 1707 2887
rect 1773 2853 1787 2867
rect 1613 2774 1627 2788
rect 1653 2774 1667 2788
rect 1693 2774 1707 2788
rect 1413 2633 1427 2647
rect 1473 2633 1487 2647
rect 1333 2573 1347 2587
rect 1093 2553 1107 2567
rect 1073 2474 1087 2488
rect 1273 2513 1287 2527
rect 1173 2473 1187 2487
rect 1213 2474 1227 2488
rect 1273 2474 1287 2488
rect 1333 2474 1347 2488
rect 1393 2474 1407 2488
rect 1513 2474 1527 2488
rect 1173 2353 1187 2367
rect 1093 2273 1107 2287
rect 1133 2254 1147 2268
rect 1253 2293 1267 2307
rect 1333 2293 1347 2307
rect 1433 2353 1447 2367
rect 1113 2212 1127 2226
rect 1173 2212 1187 2226
rect 1073 2193 1087 2207
rect 1053 2013 1067 2027
rect 1033 1993 1047 2007
rect 953 1954 967 1968
rect 913 1873 927 1887
rect 973 1873 987 1887
rect 893 1733 907 1747
rect 773 1692 787 1706
rect 833 1692 847 1706
rect 873 1692 887 1706
rect 813 1673 827 1687
rect 753 1613 767 1627
rect 673 1573 687 1587
rect 753 1553 767 1567
rect 653 1433 667 1447
rect 713 1434 727 1448
rect 573 1313 587 1327
rect 613 1293 627 1307
rect 573 1233 587 1247
rect 613 1214 627 1228
rect 633 1173 647 1187
rect 553 1133 567 1147
rect 493 1073 507 1087
rect 453 1033 467 1047
rect 413 953 427 967
rect 353 913 367 927
rect 413 914 427 928
rect 293 872 307 886
rect 333 872 347 886
rect 233 833 247 847
rect 293 813 307 827
rect 193 713 207 727
rect 253 713 267 727
rect 113 694 127 708
rect 173 693 187 707
rect 133 652 147 666
rect 133 513 147 527
rect 173 513 187 527
rect 253 694 267 708
rect 233 652 247 666
rect 273 613 287 627
rect 233 593 247 607
rect 353 833 367 847
rect 433 853 447 867
rect 573 993 587 1007
rect 733 1373 747 1387
rect 773 1313 787 1327
rect 673 1273 687 1287
rect 653 1133 667 1147
rect 633 953 647 967
rect 613 914 627 928
rect 553 813 567 827
rect 593 773 607 787
rect 653 773 667 787
rect 533 753 547 767
rect 493 733 507 747
rect 413 694 427 708
rect 453 694 467 708
rect 353 652 367 666
rect 393 652 407 666
rect 353 613 367 627
rect 433 593 447 607
rect 353 513 367 527
rect 333 413 347 427
rect 333 373 347 387
rect 453 413 467 427
rect 113 352 127 366
rect 113 313 127 327
rect 213 352 227 366
rect 273 352 287 366
rect 353 352 367 366
rect 393 352 407 366
rect 433 352 447 366
rect 593 752 607 766
rect 532 693 546 707
rect 553 694 567 708
rect 633 653 647 667
rect 513 453 527 467
rect 573 453 587 467
rect 793 1253 807 1267
rect 713 1214 727 1228
rect 773 1214 787 1228
rect 733 1113 747 1127
rect 733 914 747 928
rect 793 853 807 867
rect 713 813 727 827
rect 733 753 747 767
rect 833 1453 847 1467
rect 1053 1853 1067 1867
rect 1053 1813 1067 1827
rect 992 1773 1006 1787
rect 1013 1773 1027 1787
rect 933 1692 947 1706
rect 973 1692 987 1706
rect 1013 1673 1027 1687
rect 933 1593 947 1607
rect 913 1453 927 1467
rect 1273 2212 1287 2226
rect 1333 2212 1347 2226
rect 1373 2212 1387 2226
rect 1593 2732 1607 2746
rect 1753 2773 1767 2787
rect 1673 2732 1687 2746
rect 1813 2813 1827 2827
rect 1853 2774 1867 2788
rect 1913 2773 1927 2787
rect 1773 2732 1787 2746
rect 1833 2732 1847 2746
rect 1873 2732 1887 2746
rect 1613 2693 1627 2707
rect 1713 2693 1727 2707
rect 2113 2873 2127 2887
rect 1993 2853 2007 2867
rect 1953 2773 1967 2787
rect 2033 2813 2047 2827
rect 1953 2732 1967 2746
rect 1993 2713 2007 2727
rect 1913 2693 1927 2707
rect 1973 2692 1987 2706
rect 2073 2713 2087 2727
rect 1793 2653 1807 2667
rect 2013 2653 2027 2667
rect 1773 2553 1787 2567
rect 1593 2474 1607 2488
rect 1633 2474 1647 2488
rect 1713 2474 1727 2488
rect 1553 2433 1567 2447
rect 1613 2432 1627 2446
rect 1573 2254 1587 2268
rect 1633 2253 1647 2267
rect 1473 2193 1487 2207
rect 1413 2153 1427 2167
rect 1233 2073 1247 2087
rect 1173 2013 1187 2027
rect 1093 1953 1107 1967
rect 1133 1954 1147 1968
rect 1233 1954 1247 1968
rect 1073 1692 1087 1706
rect 1053 1573 1067 1587
rect 1073 1513 1087 1527
rect 1153 1873 1167 1887
rect 1153 1852 1167 1866
rect 1293 1793 1307 1807
rect 1273 1773 1287 1787
rect 1273 1734 1287 1748
rect 1433 1912 1447 1926
rect 1493 1912 1507 1926
rect 1473 1893 1487 1907
rect 1433 1853 1447 1867
rect 1353 1793 1367 1807
rect 1393 1793 1407 1807
rect 1333 1733 1347 1747
rect 1293 1692 1307 1706
rect 1113 1673 1127 1687
rect 973 1433 987 1447
rect 1053 1434 1067 1448
rect 1093 1434 1107 1448
rect 833 1373 847 1387
rect 873 1273 887 1287
rect 953 1313 967 1327
rect 913 1253 927 1267
rect 853 1214 867 1228
rect 893 1214 907 1228
rect 913 1172 927 1186
rect 873 1153 887 1167
rect 873 993 887 1007
rect 913 953 927 967
rect 1033 1392 1047 1406
rect 1093 1393 1107 1407
rect 993 1253 1007 1267
rect 1073 1253 1087 1267
rect 993 1213 1007 1227
rect 1033 1214 1047 1228
rect 973 1172 987 1186
rect 1053 1172 1067 1186
rect 1013 1113 1027 1127
rect 973 953 987 967
rect 953 914 967 928
rect 1013 914 1027 928
rect 913 893 927 907
rect 853 872 867 886
rect 1033 872 1047 886
rect 1173 1633 1187 1647
rect 1213 1493 1227 1507
rect 1173 1434 1187 1448
rect 1213 1434 1227 1448
rect 1593 2212 1607 2226
rect 1673 2212 1687 2226
rect 1633 2173 1647 2187
rect 1533 1954 1547 1968
rect 1633 1954 1647 1968
rect 1733 2173 1747 2187
rect 2153 2693 2167 2707
rect 2193 2973 2207 2987
rect 2253 2893 2267 2907
rect 2193 2813 2207 2827
rect 2493 3073 2507 3087
rect 2453 3033 2467 3047
rect 2413 2994 2427 3008
rect 2493 3013 2507 3027
rect 2753 3633 2767 3647
rect 2553 3514 2567 3528
rect 2593 3514 2607 3528
rect 2653 3513 2667 3527
rect 2693 3514 2707 3528
rect 2633 3493 2647 3507
rect 2533 3353 2547 3367
rect 2633 3433 2647 3447
rect 2593 3353 2607 3367
rect 2573 3313 2587 3327
rect 2713 3453 2727 3467
rect 2653 3413 2667 3427
rect 2573 3252 2587 3266
rect 2793 3813 2807 3827
rect 2773 3553 2787 3567
rect 2913 3993 2927 4007
rect 3013 3992 3027 4006
rect 2853 3893 2867 3907
rect 3013 3893 3027 3907
rect 2873 3814 2887 3828
rect 2933 3814 2947 3828
rect 2993 3814 3007 3828
rect 2813 3653 2827 3667
rect 2913 3773 2927 3787
rect 2893 3713 2907 3727
rect 2893 3593 2907 3607
rect 2853 3553 2867 3567
rect 2893 3553 2907 3567
rect 3133 4193 3147 4207
rect 3253 4773 3267 4787
rect 3293 4973 3307 4987
rect 3473 6414 3487 6428
rect 3753 6433 3767 6447
rect 3913 6433 3927 6447
rect 3613 6414 3627 6428
rect 3493 6372 3507 6386
rect 3573 6372 3587 6386
rect 3533 6333 3547 6347
rect 3693 6414 3707 6428
rect 3773 6414 3787 6428
rect 3833 6414 3847 6428
rect 3673 6372 3687 6386
rect 3713 6372 3727 6386
rect 3753 6372 3767 6386
rect 4153 6473 4167 6487
rect 4893 6473 4907 6487
rect 4933 6473 4947 6487
rect 5213 6473 5227 6487
rect 4013 6414 4027 6428
rect 4053 6413 4067 6427
rect 4113 6414 4127 6428
rect 4433 6453 4447 6467
rect 4293 6414 4307 6428
rect 4913 6453 4927 6467
rect 4473 6433 4487 6447
rect 4613 6433 4627 6447
rect 4513 6413 4527 6427
rect 4573 6414 4587 6428
rect 4793 6433 4807 6447
rect 4893 6433 4907 6447
rect 3773 6353 3787 6367
rect 3733 6273 3747 6287
rect 3613 6253 3627 6267
rect 3573 6213 3587 6227
rect 3553 6193 3567 6207
rect 3493 6153 3507 6167
rect 3513 6072 3527 6086
rect 3553 6073 3567 6087
rect 3633 6153 3647 6167
rect 3673 6153 3687 6167
rect 3593 6013 3607 6027
rect 3693 6033 3707 6047
rect 3653 5993 3667 6007
rect 3593 5973 3607 5987
rect 3553 5953 3567 5967
rect 3433 5773 3447 5787
rect 3433 5713 3447 5727
rect 3493 5633 3507 5647
rect 3653 5953 3667 5967
rect 3673 5852 3687 5866
rect 3553 5813 3567 5827
rect 3613 5773 3627 5787
rect 3573 5653 3587 5667
rect 3453 5594 3467 5608
rect 3493 5594 3507 5608
rect 3533 5594 3547 5608
rect 3433 5553 3447 5567
rect 3513 5552 3527 5566
rect 3453 5493 3467 5507
rect 3593 5594 3607 5608
rect 3533 5453 3547 5467
rect 3573 5453 3587 5467
rect 3493 5413 3507 5427
rect 3413 5374 3427 5388
rect 3473 5373 3487 5387
rect 3453 5332 3467 5346
rect 3353 5293 3367 5307
rect 3333 5093 3347 5107
rect 3513 5393 3527 5407
rect 3493 5253 3507 5267
rect 3473 5233 3487 5247
rect 3433 5173 3447 5187
rect 3353 5074 3367 5088
rect 3333 5032 3347 5046
rect 3333 4993 3347 5007
rect 3493 5153 3507 5167
rect 3553 5413 3567 5427
rect 3753 6253 3767 6267
rect 3753 6213 3767 6227
rect 3813 6372 3827 6386
rect 3913 6372 3927 6386
rect 3993 6372 4007 6386
rect 4833 6414 4847 6428
rect 5093 6433 5107 6447
rect 5053 6414 5067 6428
rect 5453 6453 5467 6467
rect 5233 6433 5247 6447
rect 5273 6433 5287 6447
rect 5393 6433 5407 6447
rect 5253 6414 5267 6428
rect 5293 6413 5307 6427
rect 5353 6414 5367 6428
rect 4133 6372 4147 6386
rect 4193 6353 4207 6367
rect 4173 6293 4187 6307
rect 4053 6273 4067 6287
rect 4053 6233 4067 6247
rect 3833 6114 3847 6128
rect 3873 6114 3887 6128
rect 3953 6114 3967 6128
rect 3993 6114 4007 6128
rect 4033 6114 4047 6128
rect 3753 6093 3767 6107
rect 3813 6072 3827 6086
rect 3873 6073 3887 6087
rect 3933 6072 3947 6086
rect 3993 6053 4007 6067
rect 3973 6033 3987 6047
rect 3913 5993 3927 6007
rect 3813 5953 3827 5967
rect 3873 5953 3887 5967
rect 3893 5933 3907 5947
rect 3853 5894 3867 5908
rect 3753 5852 3767 5866
rect 3793 5852 3807 5866
rect 3833 5852 3847 5866
rect 3893 5852 3907 5866
rect 3733 5653 3747 5667
rect 3673 5633 3687 5647
rect 3713 5594 3727 5608
rect 3653 5552 3667 5566
rect 3793 5793 3807 5807
rect 3873 5693 3887 5707
rect 3793 5653 3807 5667
rect 3793 5632 3807 5646
rect 3773 5594 3787 5608
rect 3833 5594 3847 5608
rect 3933 5933 3947 5947
rect 3953 5894 3967 5908
rect 4093 6153 4107 6167
rect 4073 6133 4087 6147
rect 4173 6114 4187 6128
rect 4073 6072 4087 6086
rect 4113 6072 4127 6086
rect 4173 6053 4187 6067
rect 4313 6372 4327 6386
rect 4413 6372 4427 6386
rect 4453 6372 4467 6386
rect 4513 6372 4527 6386
rect 4273 6233 4287 6247
rect 4713 6372 4727 6386
rect 4753 6372 4767 6386
rect 4793 6372 4807 6386
rect 4833 6373 4847 6387
rect 4873 6372 4887 6386
rect 4913 6372 4927 6386
rect 5033 6372 5047 6386
rect 4653 6333 4667 6347
rect 4593 6253 4607 6267
rect 4313 6193 4327 6207
rect 4493 6193 4507 6207
rect 4273 6153 4287 6167
rect 4273 6114 4287 6128
rect 4313 6114 4327 6128
rect 4373 6114 4387 6128
rect 4453 6114 4467 6128
rect 4593 6173 4607 6187
rect 4613 6114 4627 6128
rect 4853 6233 4867 6247
rect 4673 6173 4687 6187
rect 4293 6072 4307 6086
rect 4273 6053 4287 6067
rect 4193 6033 4207 6047
rect 4073 6013 4087 6027
rect 4053 5993 4067 6007
rect 4033 5973 4047 5987
rect 4053 5894 4067 5908
rect 3973 5852 3987 5866
rect 4233 5933 4247 5947
rect 4133 5894 4147 5908
rect 4173 5894 4187 5908
rect 4073 5852 4087 5866
rect 4113 5852 4127 5866
rect 4153 5833 4167 5847
rect 4653 6113 4667 6127
rect 4693 6114 4707 6128
rect 4753 6114 4767 6128
rect 4633 6072 4647 6086
rect 4673 6072 4687 6086
rect 4433 6033 4447 6047
rect 4473 6033 4487 6047
rect 4373 6013 4387 6027
rect 4333 5993 4347 6007
rect 4313 5894 4327 5908
rect 4253 5833 4267 5847
rect 4053 5813 4067 5827
rect 4233 5813 4247 5827
rect 3933 5793 3947 5807
rect 3913 5633 3927 5647
rect 4033 5713 4047 5727
rect 4153 5713 4167 5727
rect 3953 5594 3967 5608
rect 3993 5594 4007 5608
rect 4193 5693 4207 5707
rect 4193 5653 4207 5667
rect 4153 5613 4167 5627
rect 3793 5553 3807 5567
rect 3773 5493 3787 5507
rect 3653 5413 3667 5427
rect 3613 5393 3627 5407
rect 3693 5453 3707 5467
rect 3693 5413 3707 5427
rect 3692 5373 3706 5387
rect 3713 5374 3727 5388
rect 3653 5333 3667 5347
rect 3733 5332 3747 5346
rect 3573 5273 3587 5287
rect 3933 5553 3947 5567
rect 4013 5552 4027 5566
rect 4173 5552 4187 5566
rect 4093 5533 4107 5547
rect 3873 5493 3887 5507
rect 3853 5453 3867 5467
rect 3813 5373 3827 5387
rect 4013 5393 4027 5407
rect 4053 5393 4067 5407
rect 3813 5332 3827 5346
rect 3853 5332 3867 5346
rect 3893 5332 3907 5346
rect 3993 5332 4007 5346
rect 4033 5332 4047 5346
rect 3733 5253 3747 5267
rect 3773 5253 3787 5267
rect 3533 5153 3547 5167
rect 3513 5133 3527 5147
rect 3573 5113 3587 5127
rect 3673 5113 3687 5127
rect 3433 4933 3447 4947
rect 3473 4873 3487 4887
rect 3413 4854 3427 4868
rect 3313 4812 3327 4826
rect 3353 4812 3367 4826
rect 3393 4812 3407 4826
rect 3453 4813 3467 4827
rect 3293 4773 3307 4787
rect 3353 4633 3367 4647
rect 3233 4593 3247 4607
rect 3273 4593 3287 4607
rect 3273 4554 3287 4568
rect 3333 4533 3347 4547
rect 3293 4493 3307 4507
rect 3253 4473 3267 4487
rect 3433 4713 3447 4727
rect 3453 4693 3467 4707
rect 3593 5074 3607 5088
rect 3633 5074 3647 5088
rect 3713 5074 3727 5088
rect 3573 5013 3587 5027
rect 3993 5313 4007 5327
rect 4033 5273 4047 5287
rect 4073 5273 4087 5287
rect 3813 5213 3827 5227
rect 3893 5193 3907 5207
rect 3773 5173 3787 5187
rect 3873 5093 3887 5107
rect 3773 5074 3787 5088
rect 3813 5074 3827 5088
rect 3653 5032 3667 5046
rect 3712 5033 3726 5047
rect 3733 5033 3747 5047
rect 3793 5032 3807 5046
rect 3633 5013 3647 5027
rect 3593 4973 3607 4987
rect 3613 4893 3627 4907
rect 3533 4873 3547 4887
rect 3573 4854 3587 4868
rect 3513 4812 3527 4826
rect 3513 4733 3527 4747
rect 3493 4633 3507 4647
rect 3473 4593 3487 4607
rect 3413 4554 3427 4568
rect 3493 4553 3507 4567
rect 3353 4512 3367 4526
rect 3393 4512 3407 4526
rect 3473 4513 3487 4527
rect 3433 4493 3447 4507
rect 3493 4493 3507 4507
rect 3333 4453 3347 4467
rect 3293 4433 3307 4447
rect 3253 4334 3267 4348
rect 3353 4373 3367 4387
rect 3333 4334 3347 4348
rect 3273 4292 3287 4306
rect 3153 4173 3167 4187
rect 3193 4173 3207 4187
rect 3233 4173 3247 4187
rect 3193 4133 3207 4147
rect 3173 3913 3187 3927
rect 3253 3913 3267 3927
rect 3113 3833 3127 3847
rect 3253 3813 3267 3827
rect 3013 3772 3027 3786
rect 3053 3772 3067 3786
rect 3113 3772 3127 3786
rect 3173 3772 3187 3786
rect 3233 3772 3247 3786
rect 2993 3713 3007 3727
rect 3093 3673 3107 3687
rect 3113 3673 3127 3687
rect 2873 3533 2887 3547
rect 2913 3533 2927 3547
rect 2833 3514 2847 3528
rect 3153 3653 3167 3667
rect 3033 3514 3047 3528
rect 3093 3514 3107 3528
rect 3133 3513 3147 3527
rect 2773 3473 2787 3487
rect 2753 3453 2767 3467
rect 2733 3353 2747 3367
rect 2773 3333 2787 3347
rect 2813 3472 2827 3486
rect 2853 3472 2867 3486
rect 2833 3453 2847 3467
rect 2873 3433 2887 3447
rect 2833 3413 2847 3427
rect 2813 3373 2827 3387
rect 2793 3293 2807 3307
rect 2613 3233 2627 3247
rect 2553 3193 2567 3207
rect 2533 3013 2547 3027
rect 2373 2933 2387 2947
rect 2433 2913 2447 2927
rect 2993 3433 3007 3447
rect 2913 3353 2927 3367
rect 2973 3313 2987 3327
rect 2913 3294 2927 3308
rect 2813 3252 2827 3266
rect 2893 3252 2907 3266
rect 2933 3252 2947 3266
rect 2973 3252 2987 3266
rect 3093 3333 3107 3347
rect 3133 3333 3147 3347
rect 3053 3313 3067 3327
rect 3093 3294 3107 3308
rect 3073 3153 3087 3167
rect 3433 4413 3447 4427
rect 3453 4334 3467 4348
rect 3373 4292 3387 4306
rect 3433 4292 3447 4306
rect 3373 4233 3387 4247
rect 3333 4153 3347 4167
rect 3373 4133 3387 4147
rect 3313 4053 3327 4067
rect 3353 3992 3367 4006
rect 3873 5013 3887 5027
rect 3713 4973 3727 4987
rect 3793 4973 3807 4987
rect 3833 4973 3847 4987
rect 3653 4933 3667 4947
rect 3593 4793 3607 4807
rect 3633 4793 3647 4807
rect 3553 4713 3567 4727
rect 3573 4613 3587 4627
rect 3533 4593 3547 4607
rect 3533 4553 3547 4567
rect 3533 4513 3547 4527
rect 3593 4493 3607 4507
rect 3553 4453 3567 4467
rect 3533 4333 3547 4347
rect 3473 4113 3487 4127
rect 3513 4193 3527 4207
rect 3513 4073 3527 4087
rect 3393 4053 3407 4067
rect 3493 4053 3507 4067
rect 3373 3853 3387 3867
rect 3293 3833 3307 3847
rect 3353 3833 3367 3847
rect 3273 3633 3287 3647
rect 3353 3753 3367 3767
rect 3353 3613 3367 3627
rect 3613 4413 3627 4427
rect 3553 4292 3567 4306
rect 3553 4253 3567 4267
rect 3573 4213 3587 4227
rect 3553 4153 3567 4167
rect 3473 3992 3487 4006
rect 3533 3992 3547 4006
rect 3413 3853 3427 3867
rect 3393 3573 3407 3587
rect 3233 3553 3247 3567
rect 3273 3514 3287 3528
rect 3313 3514 3327 3528
rect 3213 3472 3227 3486
rect 3213 3433 3227 3447
rect 2613 3013 2627 3027
rect 2653 2994 2667 3008
rect 2693 2994 2707 3008
rect 2893 3033 2907 3047
rect 3013 3033 3027 3047
rect 2873 2994 2887 3008
rect 2553 2952 2567 2966
rect 2593 2952 2607 2966
rect 2633 2933 2647 2947
rect 2673 2933 2687 2947
rect 2573 2893 2587 2907
rect 2533 2853 2547 2867
rect 2493 2833 2507 2847
rect 2293 2793 2307 2807
rect 2493 2793 2507 2807
rect 2193 2774 2207 2788
rect 2253 2774 2267 2788
rect 2173 2653 2187 2667
rect 2073 2513 2087 2527
rect 1893 2474 1907 2488
rect 1953 2474 1967 2488
rect 2013 2474 2027 2488
rect 2133 2432 2147 2446
rect 2133 2353 2147 2367
rect 1913 2293 1927 2307
rect 1973 2293 1987 2307
rect 1873 2254 1887 2268
rect 1913 2254 1927 2268
rect 1953 2254 1967 2268
rect 1833 2173 1847 2187
rect 1793 2013 1807 2027
rect 1693 1954 1707 1968
rect 1733 1954 1747 1968
rect 1853 2113 1867 2127
rect 2033 2254 2047 2268
rect 2093 2253 2107 2267
rect 2053 2212 2067 2226
rect 2093 2212 2107 2226
rect 2013 2193 2027 2207
rect 1973 2173 1987 2187
rect 2053 2173 2067 2187
rect 1953 2153 1967 2167
rect 1933 2093 1947 2107
rect 1893 2073 1907 2087
rect 1893 2033 1907 2047
rect 1893 1954 1907 1968
rect 1613 1912 1627 1926
rect 1673 1913 1687 1927
rect 1553 1893 1567 1907
rect 1753 1912 1767 1926
rect 1693 1873 1707 1887
rect 1533 1853 1547 1867
rect 1753 1853 1767 1867
rect 1513 1753 1527 1767
rect 1673 1753 1687 1767
rect 1573 1734 1587 1748
rect 1613 1734 1627 1748
rect 1413 1692 1427 1706
rect 1493 1693 1507 1707
rect 1553 1692 1567 1706
rect 1953 1973 1967 1987
rect 1933 1853 1947 1867
rect 1873 1833 1887 1847
rect 1793 1813 1807 1827
rect 1813 1734 1827 1748
rect 1453 1673 1467 1687
rect 1613 1673 1627 1687
rect 1573 1533 1587 1547
rect 1533 1513 1547 1527
rect 1493 1434 1507 1448
rect 1753 1692 1767 1706
rect 1753 1633 1767 1647
rect 1733 1553 1747 1567
rect 1633 1453 1647 1467
rect 1693 1453 1707 1467
rect 1573 1433 1587 1447
rect 1673 1434 1687 1448
rect 1193 1392 1207 1406
rect 1393 1392 1407 1406
rect 1453 1393 1467 1407
rect 1513 1392 1527 1406
rect 1513 1313 1527 1327
rect 1153 1273 1167 1287
rect 1253 1273 1267 1287
rect 1353 1273 1367 1287
rect 1113 1253 1127 1267
rect 1133 1214 1147 1228
rect 1233 1193 1247 1207
rect 1173 1172 1187 1186
rect 1153 993 1167 1007
rect 1093 914 1107 928
rect 1313 1214 1327 1228
rect 1393 1213 1407 1227
rect 1473 1214 1487 1228
rect 1593 1392 1607 1406
rect 1653 1392 1667 1406
rect 1573 1273 1587 1287
rect 1693 1353 1707 1367
rect 1693 1313 1707 1327
rect 1672 1273 1686 1287
rect 1693 1273 1707 1287
rect 1593 1233 1607 1247
rect 1293 1172 1307 1186
rect 1333 1153 1347 1167
rect 1393 1153 1407 1167
rect 1493 1172 1507 1186
rect 1453 1113 1467 1127
rect 1413 1093 1427 1107
rect 1293 973 1307 987
rect 1513 973 1527 987
rect 1493 933 1507 947
rect 1193 914 1207 928
rect 1253 914 1267 928
rect 1333 914 1347 928
rect 1473 913 1487 927
rect 1633 1172 1647 1186
rect 1653 1093 1667 1107
rect 1693 953 1707 967
rect 1673 933 1687 947
rect 1733 1353 1747 1367
rect 1833 1692 1847 1706
rect 2013 1833 2027 1847
rect 1913 1793 1927 1807
rect 1953 1793 1967 1807
rect 1893 1734 1907 1748
rect 2313 2713 2327 2727
rect 2273 2673 2287 2687
rect 2273 2633 2287 2647
rect 2233 2473 2247 2487
rect 2273 2474 2287 2488
rect 2313 2474 2327 2488
rect 2352 2474 2366 2488
rect 2373 2474 2387 2488
rect 2533 2713 2547 2727
rect 2453 2573 2467 2587
rect 2293 2413 2307 2427
rect 2333 2413 2347 2427
rect 2233 2373 2247 2387
rect 2193 2333 2207 2347
rect 2173 2293 2187 2307
rect 2213 2254 2227 2268
rect 2513 2533 2527 2547
rect 2373 2433 2387 2447
rect 2393 2413 2407 2427
rect 2473 2432 2487 2446
rect 2433 2413 2447 2427
rect 2373 2333 2387 2347
rect 2353 2253 2367 2267
rect 2193 2212 2207 2226
rect 2332 2212 2346 2226
rect 2353 2213 2367 2227
rect 2273 2173 2287 2187
rect 2133 2153 2147 2167
rect 2233 2153 2247 2167
rect 2313 2093 2327 2107
rect 2233 2053 2247 2067
rect 2293 2053 2307 2067
rect 2093 1954 2107 1968
rect 2153 1954 2167 1968
rect 2313 1973 2327 1987
rect 2333 1954 2347 1968
rect 2393 2293 2407 2307
rect 2453 2254 2467 2268
rect 2633 2793 2647 2807
rect 2613 2573 2627 2587
rect 2573 2474 2587 2488
rect 2613 2474 2627 2488
rect 2653 2474 2667 2488
rect 2593 2413 2607 2427
rect 2653 2413 2667 2427
rect 2593 2353 2607 2367
rect 2533 2293 2547 2307
rect 2513 2273 2527 2287
rect 2613 2313 2627 2327
rect 2613 2273 2627 2287
rect 2573 2212 2587 2226
rect 2613 2193 2627 2207
rect 2552 2173 2566 2187
rect 2573 2173 2587 2187
rect 2493 2153 2507 2167
rect 2453 2133 2467 2147
rect 2493 2113 2507 2127
rect 2453 2073 2467 2087
rect 2393 2053 2407 2067
rect 2373 1973 2387 1987
rect 2433 1954 2447 1968
rect 2233 1933 2247 1947
rect 2133 1912 2147 1926
rect 2173 1873 2187 1887
rect 2253 1913 2267 1927
rect 2313 1912 2327 1926
rect 2373 1912 2387 1926
rect 2433 1873 2447 1887
rect 2233 1853 2247 1867
rect 2313 1853 2327 1867
rect 2153 1833 2167 1847
rect 2113 1793 2127 1807
rect 2053 1753 2067 1767
rect 1953 1734 1967 1748
rect 1993 1734 2007 1748
rect 1873 1613 1887 1627
rect 1873 1573 1887 1587
rect 1793 1553 1807 1567
rect 1773 1473 1787 1487
rect 1753 1333 1767 1347
rect 1833 1453 1847 1467
rect 1873 1434 1887 1448
rect 1973 1692 1987 1706
rect 2113 1692 2127 1706
rect 2053 1673 2067 1687
rect 2013 1653 2027 1667
rect 2013 1553 2027 1567
rect 1933 1493 1947 1507
rect 1813 1392 1827 1406
rect 1833 1293 1847 1307
rect 1753 1093 1767 1107
rect 1093 872 1107 886
rect 1173 872 1187 886
rect 1313 872 1327 886
rect 1353 872 1367 886
rect 1433 873 1447 887
rect 1073 853 1087 867
rect 1133 853 1147 867
rect 1313 853 1327 867
rect 1493 853 1507 867
rect 1593 873 1607 887
rect 1633 872 1647 886
rect 1533 853 1547 867
rect 853 813 867 827
rect 993 813 1007 827
rect 773 694 787 708
rect 813 693 827 707
rect 673 633 687 647
rect 653 493 667 507
rect 653 433 667 447
rect 633 413 647 427
rect 593 394 607 408
rect 512 353 526 367
rect 533 353 547 367
rect 313 313 327 327
rect 493 313 507 327
rect 153 253 167 267
rect 213 233 227 247
rect 573 352 587 366
rect 753 652 767 666
rect 1553 773 1567 787
rect 933 753 947 767
rect 893 733 907 747
rect 1233 713 1247 727
rect 1353 713 1367 727
rect 1433 713 1447 727
rect 1493 713 1507 727
rect 1033 694 1047 708
rect 1073 694 1087 708
rect 1133 694 1147 708
rect 1193 694 1207 708
rect 1333 694 1347 708
rect 1393 694 1407 708
rect 853 673 867 687
rect 833 652 847 666
rect 813 613 827 627
rect 813 453 827 467
rect 953 652 967 666
rect 913 633 927 647
rect 973 473 987 487
rect 913 453 927 467
rect 713 433 727 447
rect 833 433 847 447
rect 873 413 887 427
rect 753 394 767 408
rect 813 393 827 407
rect 673 352 687 366
rect 733 313 747 327
rect 773 273 787 287
rect 652 233 666 247
rect 673 233 687 247
rect 573 213 587 227
rect 633 213 647 227
rect 413 193 427 207
rect 533 193 547 207
rect 373 174 387 188
rect 493 173 507 187
rect 633 174 647 188
rect 313 132 327 146
rect 353 132 367 146
rect 493 113 507 127
rect 233 93 247 107
rect 393 93 407 107
rect 613 113 627 127
rect 713 174 727 188
rect 753 174 767 188
rect 1093 652 1107 666
rect 1213 652 1227 666
rect 1253 652 1267 666
rect 1133 613 1147 627
rect 1213 613 1227 627
rect 1293 593 1307 607
rect 1233 493 1247 507
rect 1053 473 1067 487
rect 1193 473 1207 487
rect 1033 413 1047 427
rect 1113 453 1127 467
rect 1153 413 1167 427
rect 1373 652 1387 666
rect 1333 493 1347 507
rect 1413 613 1427 627
rect 1393 493 1407 507
rect 1353 453 1367 467
rect 1373 453 1387 467
rect 1313 413 1327 427
rect 1153 352 1167 366
rect 1213 352 1227 366
rect 1253 352 1267 366
rect 1292 353 1306 367
rect 1493 652 1507 666
rect 1573 652 1587 666
rect 1553 613 1567 627
rect 1533 593 1547 607
rect 1673 853 1687 867
rect 1753 914 1767 928
rect 1913 1393 1927 1407
rect 1973 1473 1987 1487
rect 2293 1813 2307 1827
rect 2273 1793 2287 1807
rect 2173 1753 2187 1767
rect 2233 1734 2247 1748
rect 2173 1673 2187 1687
rect 2153 1653 2167 1667
rect 2393 1833 2407 1847
rect 2333 1734 2347 1748
rect 2753 2952 2767 2966
rect 2793 2952 2807 2966
rect 2833 2952 2847 2966
rect 2813 2913 2827 2927
rect 2793 2813 2807 2827
rect 2693 2773 2707 2787
rect 2793 2732 2807 2746
rect 2753 2553 2767 2567
rect 2713 2474 2727 2488
rect 2753 2474 2767 2488
rect 2693 2433 2707 2447
rect 2693 2373 2707 2387
rect 2753 2413 2767 2427
rect 2733 2353 2747 2367
rect 2793 2433 2807 2447
rect 2773 2373 2787 2387
rect 2873 2813 2887 2827
rect 2933 2994 2947 3008
rect 2953 2893 2967 2907
rect 2973 2873 2987 2887
rect 2973 2833 2987 2847
rect 3133 3093 3147 3107
rect 3173 2994 3187 3008
rect 3373 3514 3387 3528
rect 3433 3813 3447 3827
rect 3473 3814 3487 3828
rect 3533 3773 3547 3787
rect 3773 4853 3787 4867
rect 3693 4812 3707 4826
rect 3693 4753 3707 4767
rect 3673 4633 3687 4647
rect 3673 4573 3687 4587
rect 3833 4933 3847 4947
rect 3853 4854 3867 4868
rect 3913 5113 3927 5127
rect 3973 5074 3987 5088
rect 3933 5013 3947 5027
rect 3793 4812 3807 4826
rect 3833 4812 3847 4826
rect 3913 4753 3927 4767
rect 3913 4713 3927 4727
rect 3753 4693 3767 4707
rect 3733 4673 3747 4687
rect 3713 4593 3727 4607
rect 3713 4553 3727 4567
rect 3793 4613 3807 4627
rect 3853 4613 3867 4627
rect 3793 4554 3807 4568
rect 3833 4554 3847 4568
rect 3713 4513 3727 4527
rect 3672 4413 3686 4427
rect 3693 4413 3707 4427
rect 3773 4512 3787 4526
rect 3793 4473 3807 4487
rect 3733 4453 3747 4467
rect 3713 4373 3727 4387
rect 3693 4253 3707 4267
rect 3653 4213 3667 4227
rect 3773 4233 3787 4247
rect 3693 4193 3707 4207
rect 3733 4193 3747 4207
rect 3653 4073 3667 4087
rect 3713 4133 3727 4147
rect 3753 4133 3767 4147
rect 3733 4093 3747 4107
rect 3713 4073 3727 4087
rect 3693 4033 3707 4047
rect 3613 3992 3627 4006
rect 3693 3993 3707 4007
rect 3713 3973 3727 3987
rect 3653 3913 3667 3927
rect 3613 3893 3627 3907
rect 3653 3873 3667 3887
rect 3613 3853 3627 3867
rect 3613 3814 3627 3828
rect 3693 3814 3707 3828
rect 3493 3733 3507 3747
rect 3433 3613 3447 3627
rect 3453 3593 3467 3607
rect 3433 3473 3447 3487
rect 3253 3393 3267 3407
rect 3333 3433 3347 3447
rect 3393 3433 3407 3447
rect 3333 3294 3347 3308
rect 3373 3252 3387 3266
rect 3313 3213 3327 3227
rect 3373 3213 3387 3227
rect 3233 2994 3247 3008
rect 3153 2952 3167 2966
rect 3213 2953 3227 2967
rect 3093 2813 3107 2827
rect 2893 2653 2907 2667
rect 2873 2593 2887 2607
rect 2873 2474 2887 2488
rect 3053 2774 3067 2788
rect 2993 2732 3007 2746
rect 3033 2732 3047 2746
rect 2973 2653 2987 2667
rect 3073 2653 3087 2667
rect 2953 2473 2967 2487
rect 2693 2193 2707 2207
rect 2773 2212 2787 2226
rect 2733 2173 2747 2187
rect 2713 2153 2727 2167
rect 2493 1954 2507 1968
rect 2553 1954 2567 1968
rect 2613 1954 2627 1968
rect 2673 1954 2687 1968
rect 2473 1913 2487 1927
rect 2553 1873 2567 1887
rect 2473 1833 2487 1847
rect 2453 1793 2467 1807
rect 2313 1692 2327 1706
rect 2293 1633 2307 1647
rect 2193 1593 2207 1607
rect 2273 1593 2287 1607
rect 2173 1573 2187 1587
rect 2073 1453 2087 1467
rect 2133 1434 2147 1448
rect 1993 1392 2007 1406
rect 2153 1393 2167 1407
rect 1933 1373 1947 1387
rect 2033 1373 2047 1387
rect 2073 1373 2087 1387
rect 2013 1293 2027 1307
rect 2073 1293 2087 1307
rect 1873 1253 1887 1267
rect 1853 1233 1867 1247
rect 1933 1214 1947 1228
rect 1993 1213 2007 1227
rect 1873 1172 1887 1186
rect 1913 1172 1927 1186
rect 2053 1253 2067 1267
rect 2073 1233 2087 1247
rect 2053 1214 2067 1228
rect 2013 1172 2027 1186
rect 2073 1172 2087 1186
rect 2493 1733 2507 1747
rect 2613 1853 2627 1867
rect 2633 1813 2647 1827
rect 2613 1793 2627 1807
rect 2613 1753 2627 1767
rect 2413 1692 2427 1706
rect 2493 1692 2507 1706
rect 2533 1692 2547 1706
rect 2573 1692 2587 1706
rect 2613 1692 2627 1706
rect 2333 1673 2347 1687
rect 2373 1673 2387 1687
rect 2773 2153 2787 2167
rect 2813 2153 2827 2167
rect 2793 1893 2807 1907
rect 2833 1893 2847 1907
rect 2813 1853 2827 1867
rect 2713 1753 2727 1767
rect 2693 1734 2707 1748
rect 2893 2353 2907 2367
rect 2873 2254 2887 2268
rect 2913 2212 2927 2226
rect 3293 2952 3307 2966
rect 3233 2913 3247 2927
rect 3293 2913 3307 2927
rect 3253 2853 3267 2867
rect 3133 2813 3147 2827
rect 3113 2633 3127 2647
rect 3153 2774 3167 2788
rect 3213 2774 3227 2788
rect 3173 2732 3187 2746
rect 3153 2693 3167 2707
rect 3213 2673 3227 2687
rect 3173 2633 3187 2647
rect 2993 2573 3007 2587
rect 3133 2573 3147 2587
rect 3153 2533 3167 2547
rect 3053 2432 3067 2446
rect 3093 2432 3107 2446
rect 3033 2393 3047 2407
rect 3153 2393 3167 2407
rect 2993 2254 3007 2268
rect 3153 2353 3167 2367
rect 3093 2313 3107 2327
rect 3313 2813 3327 2827
rect 3413 3353 3427 3367
rect 3413 3294 3427 3308
rect 3413 3253 3427 3267
rect 3413 3193 3427 3207
rect 3393 3133 3407 3147
rect 3373 2774 3387 2788
rect 3293 2733 3307 2747
rect 3353 2732 3367 2746
rect 3413 3073 3427 3087
rect 3473 3573 3487 3587
rect 3553 3693 3567 3707
rect 3553 3653 3567 3667
rect 3633 3772 3647 3786
rect 3593 3753 3607 3767
rect 3673 3773 3687 3787
rect 3593 3713 3607 3727
rect 3573 3613 3587 3627
rect 3513 3553 3527 3567
rect 3493 3513 3507 3527
rect 3953 4893 3967 4907
rect 3933 4673 3947 4687
rect 3993 4953 4007 4967
rect 4073 5213 4087 5227
rect 4173 5513 4187 5527
rect 4213 5374 4227 5388
rect 4113 5332 4127 5346
rect 4233 5313 4247 5327
rect 4193 5253 4207 5267
rect 4133 5213 4147 5227
rect 4133 5173 4147 5187
rect 4153 5153 4167 5167
rect 4153 5113 4167 5127
rect 4053 5033 4067 5047
rect 4053 4933 4067 4947
rect 4093 5074 4107 5088
rect 4213 5133 4227 5147
rect 4193 5013 4207 5027
rect 4133 4993 4147 5007
rect 4113 4953 4127 4967
rect 4133 4913 4147 4927
rect 4033 4893 4047 4907
rect 4073 4893 4087 4907
rect 4113 4893 4127 4907
rect 4033 4854 4047 4868
rect 4073 4854 4087 4868
rect 3973 4812 3987 4826
rect 4013 4812 4027 4826
rect 4033 4713 4047 4727
rect 3953 4613 3967 4627
rect 3913 4554 3927 4568
rect 3953 4554 3967 4568
rect 4013 4554 4027 4568
rect 3873 4513 3887 4527
rect 3853 4433 3867 4447
rect 3853 4412 3867 4426
rect 3933 4512 3947 4526
rect 3973 4433 3987 4447
rect 3893 4373 3907 4387
rect 3933 4334 3947 4348
rect 3953 4292 3967 4306
rect 3933 4253 3947 4267
rect 3913 4213 3927 4227
rect 3873 4193 3887 4207
rect 3933 4173 3947 4187
rect 3853 4153 3867 4167
rect 3893 4113 3907 4127
rect 3833 4072 3847 4086
rect 3793 4034 3807 4048
rect 3873 4053 3887 4067
rect 3733 3933 3747 3947
rect 3813 3973 3827 3987
rect 3913 4073 3927 4087
rect 3953 4073 3967 4087
rect 3993 4413 4007 4427
rect 3993 4334 4007 4348
rect 3993 4093 4007 4107
rect 3933 4053 3947 4067
rect 3973 4034 3987 4048
rect 3893 3993 3907 4007
rect 3953 3992 3967 4006
rect 3833 3933 3847 3947
rect 3793 3772 3807 3786
rect 3733 3713 3747 3727
rect 3693 3693 3707 3707
rect 3753 3673 3767 3687
rect 3733 3613 3747 3627
rect 3793 3633 3807 3647
rect 3753 3593 3767 3607
rect 3793 3593 3807 3607
rect 3793 3553 3807 3567
rect 3653 3513 3667 3527
rect 3693 3514 3707 3528
rect 3473 3433 3487 3447
rect 3553 3433 3567 3447
rect 3633 3433 3647 3447
rect 3533 3294 3547 3308
rect 3493 3213 3507 3227
rect 3453 3113 3467 3127
rect 3433 3053 3447 3067
rect 3473 3053 3487 3067
rect 3473 2993 3487 3007
rect 3413 2953 3427 2967
rect 3393 2713 3407 2727
rect 3253 2653 3267 2667
rect 3453 2952 3467 2966
rect 3493 2952 3507 2966
rect 3453 2893 3467 2907
rect 3513 2833 3527 2847
rect 3453 2774 3467 2788
rect 3453 2713 3467 2727
rect 3413 2613 3427 2627
rect 3273 2593 3287 2607
rect 3213 2573 3227 2587
rect 3213 2493 3227 2507
rect 3413 2573 3427 2587
rect 3433 2553 3447 2567
rect 3413 2533 3427 2547
rect 3273 2474 3287 2488
rect 3333 2474 3347 2488
rect 3433 2473 3447 2487
rect 3413 2433 3427 2447
rect 3213 2413 3227 2427
rect 3173 2333 3187 2347
rect 3293 2333 3307 2347
rect 3353 2333 3367 2347
rect 3413 2333 3427 2347
rect 3073 2293 3087 2307
rect 3173 2273 3187 2287
rect 3093 2253 3107 2267
rect 2973 2212 2987 2226
rect 2993 2133 3007 2147
rect 2993 2093 3007 2107
rect 3053 2212 3067 2226
rect 3213 2212 3227 2226
rect 3013 2033 3027 2047
rect 2933 1993 2947 2007
rect 3013 1993 3027 2007
rect 3113 2113 3127 2127
rect 3133 2093 3147 2107
rect 3113 2073 3127 2087
rect 2873 1954 2887 1968
rect 2913 1954 2927 1968
rect 2953 1954 2967 1968
rect 2933 1912 2947 1926
rect 2873 1873 2887 1887
rect 2973 1873 2987 1887
rect 3013 1873 3027 1887
rect 2893 1853 2907 1867
rect 2853 1813 2867 1827
rect 2853 1773 2867 1787
rect 2793 1733 2807 1747
rect 2953 1793 2967 1807
rect 2933 1773 2947 1787
rect 2893 1734 2907 1748
rect 2773 1713 2787 1727
rect 2513 1653 2527 1667
rect 2633 1653 2647 1667
rect 2333 1573 2347 1587
rect 2292 1513 2306 1527
rect 2313 1513 2327 1527
rect 2193 1393 2207 1407
rect 2293 1392 2307 1406
rect 2253 1333 2267 1347
rect 2233 1273 2247 1287
rect 2293 1273 2307 1287
rect 2273 1213 2287 1227
rect 1953 1133 1967 1147
rect 2173 1133 2187 1147
rect 1833 1093 1847 1107
rect 1973 953 1987 967
rect 1793 913 1807 927
rect 1813 914 1827 928
rect 2053 914 2067 928
rect 2093 914 2107 928
rect 2133 914 2147 928
rect 1753 853 1767 867
rect 1733 733 1747 747
rect 1653 694 1667 708
rect 1713 694 1727 708
rect 1873 872 1887 886
rect 1993 872 2007 886
rect 1913 773 1927 787
rect 1993 773 2007 787
rect 1833 694 1847 708
rect 1873 694 1887 708
rect 1953 733 1967 747
rect 1693 652 1707 666
rect 1733 652 1747 666
rect 1653 613 1667 627
rect 1973 694 1987 708
rect 2013 694 2027 708
rect 2113 872 2127 886
rect 2213 1172 2227 1186
rect 2253 1172 2267 1186
rect 2253 1013 2267 1027
rect 2413 1473 2427 1487
rect 2473 1433 2487 1447
rect 2393 1392 2407 1406
rect 2413 1253 2427 1267
rect 2453 1253 2467 1267
rect 2333 1233 2347 1247
rect 2373 1214 2387 1228
rect 2333 1173 2347 1187
rect 2253 914 2267 928
rect 2313 914 2327 928
rect 2193 873 2207 887
rect 2273 793 2287 807
rect 2273 733 2287 747
rect 2313 733 2327 747
rect 2193 694 2207 708
rect 1973 653 1987 667
rect 2033 652 2047 666
rect 2113 653 2127 667
rect 1893 633 1907 647
rect 2033 631 2047 645
rect 2073 633 2087 647
rect 1633 573 1647 587
rect 1773 573 1787 587
rect 1553 493 1567 507
rect 1473 473 1487 487
rect 1513 413 1527 427
rect 1733 473 1747 487
rect 1793 473 1807 487
rect 1653 433 1667 447
rect 1593 394 1607 408
rect 1633 394 1647 408
rect 1313 352 1327 366
rect 1373 352 1387 366
rect 1413 352 1427 366
rect 1533 352 1547 366
rect 893 313 907 327
rect 1693 394 1707 408
rect 2033 433 2047 447
rect 1813 394 1827 408
rect 1873 394 1887 408
rect 1913 394 1927 408
rect 2073 394 2087 408
rect 1713 352 1727 366
rect 1753 352 1767 366
rect 1793 353 1807 367
rect 1653 313 1667 327
rect 1253 273 1267 287
rect 1393 273 1407 287
rect 1573 273 1587 287
rect 1633 273 1647 287
rect 973 253 987 267
rect 1173 253 1187 267
rect 913 233 927 247
rect 873 174 887 188
rect 1033 174 1047 188
rect 1073 174 1087 188
rect 1313 213 1327 227
rect 1353 174 1367 188
rect 1753 313 1767 327
rect 1473 213 1487 227
rect 1673 213 1687 227
rect 1713 213 1727 227
rect 1413 173 1427 187
rect 1513 193 1527 207
rect 1633 174 1647 188
rect 1733 193 1747 207
rect 653 132 667 146
rect 693 132 707 146
rect 733 132 747 146
rect 813 132 827 146
rect 853 113 867 127
rect 973 132 987 146
rect 1053 132 1067 146
rect 1253 132 1267 146
rect 1293 132 1307 146
rect 1193 113 1207 127
rect 1413 132 1427 146
rect 1653 132 1667 146
rect 1793 273 1807 287
rect 1973 373 1987 387
rect 1833 253 1847 267
rect 1813 193 1827 207
rect 1933 352 1947 366
rect 2053 352 2067 366
rect 1973 313 1987 327
rect 2093 293 2107 307
rect 2073 253 2087 267
rect 1893 233 1907 247
rect 2013 233 2027 247
rect 1733 132 1747 146
rect 1913 173 1927 187
rect 1973 174 1987 188
rect 2053 213 2067 227
rect 1813 132 1827 146
rect 1853 132 1867 146
rect 1893 132 1907 146
rect 1333 113 1347 127
rect 1373 113 1387 127
rect 733 93 747 107
rect 893 93 907 107
rect 1013 93 1027 107
rect 1953 132 1967 146
rect 1993 132 2007 146
rect 2013 113 2027 127
rect 1913 93 1927 107
rect 1993 93 2007 107
rect 93 73 107 87
rect 593 73 607 87
rect 633 73 647 87
rect 1653 73 1667 87
rect 1973 73 1987 87
rect 2233 633 2247 647
rect 2253 433 2267 447
rect 2153 394 2167 408
rect 2213 394 2227 408
rect 2133 213 2147 227
rect 2073 173 2087 187
rect 2113 174 2127 188
rect 2233 352 2247 366
rect 2273 352 2287 366
rect 2213 233 2227 247
rect 2393 1172 2407 1186
rect 2453 1172 2467 1186
rect 2433 953 2447 967
rect 2393 914 2407 928
rect 2713 1633 2727 1647
rect 2673 1593 2687 1607
rect 2713 1513 2727 1527
rect 2613 1453 2627 1467
rect 2533 1434 2547 1448
rect 2673 1434 2687 1448
rect 2513 1393 2527 1407
rect 2573 1392 2587 1406
rect 2693 1393 2707 1407
rect 2493 1373 2507 1387
rect 2553 1214 2567 1228
rect 2613 1213 2627 1227
rect 2793 1692 2807 1706
rect 2833 1692 2847 1706
rect 2792 1653 2806 1667
rect 2813 1653 2827 1667
rect 2853 1653 2867 1667
rect 2773 1593 2787 1607
rect 2833 1593 2847 1607
rect 2793 1513 2807 1527
rect 2793 1373 2807 1387
rect 2733 1313 2747 1327
rect 2773 1313 2787 1327
rect 2733 1214 2747 1228
rect 2493 1173 2507 1187
rect 2533 1172 2547 1186
rect 2573 1172 2587 1186
rect 2693 1153 2707 1167
rect 2553 1073 2567 1087
rect 2673 1033 2687 1047
rect 2553 1013 2567 1027
rect 2513 953 2527 967
rect 2473 913 2487 927
rect 2413 773 2427 787
rect 2413 733 2427 747
rect 2473 733 2487 747
rect 2393 533 2407 547
rect 2373 473 2387 487
rect 2353 433 2367 447
rect 2373 394 2387 408
rect 2473 473 2487 487
rect 2433 453 2447 467
rect 2433 394 2447 408
rect 2633 933 2647 947
rect 2593 914 2607 928
rect 2653 873 2667 887
rect 2593 833 2607 847
rect 2633 833 2647 847
rect 2533 793 2547 807
rect 2593 793 2607 807
rect 2553 773 2567 787
rect 2533 733 2547 747
rect 2513 713 2527 727
rect 2513 533 2527 547
rect 2573 533 2587 547
rect 2493 413 2507 427
rect 2353 353 2367 367
rect 2393 313 2407 327
rect 2333 213 2347 227
rect 2313 193 2327 207
rect 2353 174 2367 188
rect 2413 293 2427 307
rect 2453 293 2467 307
rect 2453 213 2467 227
rect 2433 173 2447 187
rect 2613 493 2627 507
rect 2533 413 2547 427
rect 2513 352 2527 366
rect 2493 193 2507 207
rect 2293 132 2307 146
rect 2133 113 2147 127
rect 2393 132 2407 146
rect 2333 93 2347 107
rect 2433 93 2447 107
rect 1933 13 1947 27
rect 2053 13 2067 27
rect 2433 13 2447 27
rect 2573 394 2587 408
rect 2693 873 2707 887
rect 2893 1673 2907 1687
rect 2873 1633 2887 1647
rect 2873 1434 2887 1448
rect 3073 1954 3087 1968
rect 3153 2033 3167 2047
rect 3093 1893 3107 1907
rect 3133 1912 3147 1926
rect 3113 1813 3127 1827
rect 3033 1753 3047 1767
rect 3013 1734 3027 1748
rect 3233 2013 3247 2027
rect 3333 2212 3347 2226
rect 3313 2173 3327 2187
rect 3213 1912 3227 1926
rect 3253 1912 3267 1926
rect 3293 1913 3307 1927
rect 3193 1793 3207 1807
rect 3253 1793 3267 1807
rect 3173 1753 3187 1767
rect 3153 1733 3167 1747
rect 2953 1673 2967 1687
rect 2933 1653 2947 1667
rect 2993 1633 3007 1647
rect 2973 1613 2987 1627
rect 2933 1434 2947 1448
rect 3073 1692 3087 1706
rect 3132 1673 3146 1687
rect 3153 1673 3167 1687
rect 3253 1734 3267 1748
rect 3273 1693 3287 1707
rect 3353 2013 3367 2027
rect 3333 1953 3347 1967
rect 3513 2593 3527 2607
rect 3513 2493 3527 2507
rect 3533 2473 3547 2487
rect 3453 2393 3467 2407
rect 3573 3413 3587 3427
rect 3873 3953 3887 3967
rect 3853 3753 3867 3767
rect 3933 3913 3947 3927
rect 3933 3814 3947 3828
rect 4073 4613 4087 4627
rect 4053 4553 4067 4567
rect 4133 4854 4147 4868
rect 4173 4854 4187 4868
rect 4333 5852 4347 5866
rect 4293 5813 4307 5827
rect 4733 6072 4747 6086
rect 4893 6213 4907 6227
rect 4953 6293 4967 6307
rect 4913 6153 4927 6167
rect 4873 6133 4887 6147
rect 4913 6114 4927 6128
rect 4993 6173 5007 6187
rect 4893 6072 4907 6086
rect 4953 6053 4967 6067
rect 4773 6033 4787 6047
rect 4853 6033 4867 6047
rect 4933 6033 4947 6047
rect 4693 5993 4707 6007
rect 4433 5973 4447 5987
rect 4853 5953 4867 5967
rect 4433 5933 4447 5947
rect 4753 5933 4767 5947
rect 4393 5893 4407 5907
rect 4573 5894 4587 5908
rect 4633 5894 4647 5908
rect 4673 5894 4687 5908
rect 4793 5894 4807 5908
rect 4373 5793 4387 5807
rect 4453 5852 4467 5866
rect 4533 5833 4547 5847
rect 4393 5693 4407 5707
rect 4273 5653 4287 5667
rect 4333 5594 4347 5608
rect 4433 5594 4447 5608
rect 4473 5594 4487 5608
rect 4513 5594 4527 5608
rect 4273 5553 4287 5567
rect 4273 5513 4287 5527
rect 4313 5513 4327 5527
rect 4433 5513 4447 5527
rect 4373 5493 4387 5507
rect 4373 5453 4387 5467
rect 4333 5374 4347 5388
rect 4413 5374 4427 5388
rect 4273 5332 4287 5346
rect 4313 5332 4327 5346
rect 4353 5332 4367 5346
rect 4253 5253 4267 5267
rect 4333 5213 4347 5227
rect 4413 5253 4427 5267
rect 4353 5193 4367 5207
rect 4393 5193 4407 5207
rect 4333 5113 4347 5127
rect 4393 5093 4407 5107
rect 4293 5074 4307 5088
rect 4333 5074 4347 5088
rect 4313 5032 4327 5046
rect 4493 5553 4507 5567
rect 4453 5453 4467 5467
rect 4553 5753 4567 5767
rect 4633 5753 4647 5767
rect 4573 5713 4587 5727
rect 4613 5713 4627 5727
rect 4553 5633 4567 5647
rect 4633 5653 4647 5667
rect 4733 5833 4747 5847
rect 4733 5793 4747 5807
rect 4733 5693 4747 5707
rect 4673 5633 4687 5647
rect 4512 5513 4526 5527
rect 4533 5513 4547 5527
rect 4473 5332 4487 5346
rect 4513 5253 4527 5267
rect 4593 5594 4607 5608
rect 4633 5593 4647 5607
rect 4593 5533 4607 5547
rect 4613 5513 4627 5527
rect 4833 5753 4847 5767
rect 4813 5693 4827 5707
rect 4773 5673 4787 5687
rect 4773 5594 4787 5608
rect 4693 5533 4707 5547
rect 4693 5493 4707 5507
rect 4633 5473 4647 5487
rect 4673 5473 4687 5487
rect 4593 5433 4607 5447
rect 4573 5413 4587 5427
rect 4573 5332 4587 5346
rect 4613 5332 4627 5346
rect 4673 5273 4687 5287
rect 4713 5473 4727 5487
rect 4813 5473 4827 5487
rect 4753 5433 4767 5447
rect 4893 5894 4907 5908
rect 4913 5833 4927 5847
rect 4993 6033 5007 6047
rect 5233 6372 5247 6386
rect 5293 6372 5307 6386
rect 5133 6333 5147 6347
rect 5193 6333 5207 6347
rect 5053 6114 5067 6128
rect 5113 6113 5127 6127
rect 5073 6053 5087 6067
rect 5013 6013 5027 6027
rect 5473 6413 5487 6427
rect 5533 6413 5547 6427
rect 5413 6353 5427 6367
rect 5453 6353 5467 6367
rect 5373 6293 5387 6307
rect 5173 6273 5187 6287
rect 5193 6253 5207 6267
rect 5173 6233 5187 6247
rect 5213 6193 5227 6207
rect 5373 6193 5387 6207
rect 5193 6173 5207 6187
rect 5213 6153 5227 6167
rect 5513 6372 5527 6386
rect 5713 6473 5727 6487
rect 5893 6473 5907 6487
rect 5693 6433 5707 6447
rect 5673 6414 5687 6428
rect 5913 6453 5927 6467
rect 5953 6453 5967 6467
rect 5793 6433 5807 6447
rect 5813 6414 5827 6428
rect 5853 6414 5867 6428
rect 6073 6433 6087 6447
rect 5993 6414 6007 6428
rect 6033 6414 6047 6428
rect 5633 6373 5647 6387
rect 5693 6372 5707 6386
rect 5753 6372 5767 6386
rect 5653 6353 5667 6367
rect 5873 6372 5887 6386
rect 5913 6373 5927 6387
rect 5973 6372 5987 6386
rect 5793 6353 5807 6367
rect 5833 6293 5847 6307
rect 5753 6273 5767 6287
rect 5573 6193 5587 6207
rect 5773 6173 5787 6187
rect 5473 6153 5487 6167
rect 5673 6153 5687 6167
rect 5413 6114 5427 6128
rect 5453 6114 5467 6128
rect 5133 6072 5147 6086
rect 5193 6072 5207 6086
rect 5233 6072 5247 6086
rect 5353 6072 5367 6086
rect 5153 5993 5167 6007
rect 5053 5913 5067 5927
rect 5113 5913 5127 5927
rect 5033 5852 5047 5866
rect 5073 5793 5087 5807
rect 5133 5773 5147 5787
rect 5393 5953 5407 5967
rect 5213 5913 5227 5927
rect 5253 5894 5267 5908
rect 5313 5893 5327 5907
rect 5373 5894 5387 5908
rect 5413 5894 5427 5908
rect 5233 5852 5247 5866
rect 5193 5793 5207 5807
rect 5153 5693 5167 5707
rect 4953 5673 4967 5687
rect 4853 5594 4867 5608
rect 4893 5594 4907 5608
rect 4773 5413 4787 5427
rect 4833 5413 4847 5427
rect 4813 5374 4827 5388
rect 4733 5333 4747 5347
rect 4713 5293 4727 5307
rect 4713 5272 4727 5286
rect 4613 5253 4627 5267
rect 4653 5253 4667 5267
rect 4693 5253 4707 5267
rect 4553 5233 4567 5247
rect 4573 5213 4587 5227
rect 4433 5173 4447 5187
rect 4473 5113 4487 5127
rect 4553 5093 4567 5107
rect 4513 5074 4527 5088
rect 4493 5032 4507 5046
rect 4273 5013 4287 5027
rect 4273 4913 4287 4927
rect 4233 4873 4247 4887
rect 4173 4773 4187 4787
rect 4113 4574 4127 4588
rect 4113 4553 4127 4567
rect 4033 4513 4047 4527
rect 4093 4493 4107 4507
rect 4233 4812 4247 4826
rect 4293 4812 4307 4826
rect 4193 4753 4207 4767
rect 4453 4993 4467 5007
rect 4513 4993 4527 5007
rect 4373 4933 4387 4947
rect 4373 4854 4387 4868
rect 4433 4854 4447 4868
rect 4393 4812 4407 4826
rect 4293 4733 4307 4747
rect 4253 4713 4267 4727
rect 4193 4673 4207 4687
rect 4253 4554 4267 4568
rect 4293 4553 4307 4567
rect 4373 4593 4387 4607
rect 4533 4973 4547 4987
rect 4473 4873 4487 4887
rect 4553 4933 4567 4947
rect 4533 4854 4547 4868
rect 4493 4812 4507 4826
rect 4473 4753 4487 4767
rect 4453 4693 4467 4707
rect 4413 4633 4427 4647
rect 4413 4593 4427 4607
rect 4173 4493 4187 4507
rect 4213 4493 4227 4507
rect 4233 4473 4247 4487
rect 4153 4413 4167 4427
rect 4193 4413 4207 4427
rect 4173 4393 4187 4407
rect 4113 4373 4127 4387
rect 4033 4333 4047 4347
rect 4153 4334 4167 4348
rect 4053 4292 4067 4306
rect 4273 4393 4287 4407
rect 4213 4373 4227 4387
rect 4193 4334 4207 4348
rect 4033 4233 4047 4247
rect 4173 4233 4187 4247
rect 4013 3953 4027 3967
rect 4073 4213 4087 4227
rect 4173 4193 4187 4207
rect 4133 4113 4147 4127
rect 4073 4093 4087 4107
rect 4093 4053 4107 4067
rect 4073 3992 4087 4006
rect 4033 3893 4047 3907
rect 4073 3893 4087 3907
rect 4313 4433 4327 4447
rect 4373 4493 4387 4507
rect 4353 4413 4367 4427
rect 4353 4373 4367 4387
rect 4293 4353 4307 4367
rect 4313 4334 4327 4348
rect 4273 4273 4287 4287
rect 4213 4053 4227 4067
rect 4453 4513 4467 4526
rect 4453 4512 4467 4513
rect 4433 4433 4447 4447
rect 4453 4393 4467 4407
rect 4393 4333 4407 4347
rect 4593 5173 4607 5187
rect 4653 5094 4667 5108
rect 4653 5073 4667 5087
rect 4693 5074 4707 5088
rect 4593 4853 4607 4867
rect 4573 4793 4587 4807
rect 4553 4733 4567 4747
rect 4593 4733 4607 4747
rect 4633 5013 4647 5027
rect 4673 4873 4687 4887
rect 4733 5213 4747 5227
rect 4773 5293 4787 5307
rect 4833 5233 4847 5247
rect 4773 5133 4787 5147
rect 4753 5113 4767 5127
rect 4753 5074 4767 5088
rect 4793 5074 4807 5088
rect 4813 5032 4827 5046
rect 4913 5533 4927 5547
rect 5173 5653 5187 5667
rect 5073 5633 5087 5647
rect 5113 5633 5127 5647
rect 5033 5594 5047 5608
rect 5013 5552 5027 5566
rect 5053 5552 5067 5566
rect 5153 5593 5167 5607
rect 5313 5633 5327 5647
rect 5253 5594 5267 5608
rect 5313 5594 5327 5608
rect 5173 5553 5187 5567
rect 4893 5493 4907 5507
rect 4953 5493 4967 5507
rect 5013 5493 5027 5507
rect 5213 5492 5227 5506
rect 4953 5433 4967 5447
rect 4993 5413 5007 5427
rect 4953 5374 4967 5388
rect 4933 5233 4947 5247
rect 4953 5193 4967 5207
rect 4913 5113 4927 5127
rect 4993 5113 5007 5127
rect 4893 5073 4907 5087
rect 4893 5033 4907 5047
rect 4873 5013 4887 5027
rect 4773 4973 4787 4987
rect 4833 4973 4847 4987
rect 4893 4953 4907 4967
rect 4733 4933 4747 4947
rect 4833 4933 4847 4947
rect 4873 4913 4887 4927
rect 4833 4893 4847 4907
rect 4733 4873 4747 4887
rect 4713 4853 4727 4867
rect 4713 4813 4727 4827
rect 4673 4793 4687 4807
rect 4653 4733 4667 4747
rect 4493 4653 4507 4667
rect 4613 4653 4627 4667
rect 4653 4653 4667 4667
rect 4473 4353 4487 4367
rect 4633 4593 4647 4607
rect 4613 4554 4627 4568
rect 4653 4554 4667 4568
rect 4513 4512 4527 4526
rect 4513 4433 4527 4447
rect 4313 4253 4327 4267
rect 4373 4253 4387 4267
rect 4113 3873 4127 3887
rect 4093 3853 4107 3867
rect 4093 3832 4107 3846
rect 3973 3813 3987 3827
rect 4073 3813 4087 3827
rect 3873 3733 3887 3747
rect 3933 3733 3947 3747
rect 3913 3693 3927 3707
rect 3833 3653 3847 3667
rect 3913 3633 3927 3647
rect 3833 3514 3847 3528
rect 3873 3514 3887 3528
rect 3813 3433 3827 3447
rect 3913 3513 3927 3527
rect 3973 3773 3987 3787
rect 3953 3713 3967 3727
rect 3953 3692 3967 3706
rect 3893 3472 3907 3486
rect 3933 3473 3947 3487
rect 3653 3393 3667 3407
rect 3733 3393 3747 3407
rect 3773 3393 3787 3407
rect 3793 3373 3807 3387
rect 3633 3333 3647 3347
rect 3733 3333 3747 3347
rect 3693 3294 3707 3308
rect 3733 3294 3747 3308
rect 3673 3153 3687 3167
rect 3633 3073 3647 3087
rect 3673 3073 3687 3087
rect 3613 3013 3627 3027
rect 3973 3633 3987 3647
rect 3973 3593 3987 3607
rect 4053 3772 4067 3786
rect 4273 4034 4287 4048
rect 4253 3992 4267 4006
rect 4213 3973 4227 3987
rect 4113 3733 4127 3747
rect 4093 3713 4107 3727
rect 4033 3593 4047 3607
rect 4213 3593 4227 3607
rect 3993 3553 4007 3567
rect 3993 3532 4007 3546
rect 3973 3513 3987 3527
rect 4093 3553 4107 3567
rect 4073 3533 4087 3547
rect 3953 3413 3967 3427
rect 4133 3514 4147 3528
rect 4173 3514 4187 3528
rect 4213 3514 4227 3528
rect 4093 3473 4107 3487
rect 4153 3472 4167 3486
rect 4192 3473 4206 3487
rect 4213 3473 4227 3487
rect 4153 3413 4167 3427
rect 4073 3373 4087 3387
rect 4113 3373 4127 3387
rect 3853 3252 3867 3266
rect 3813 3213 3827 3227
rect 3913 3073 3927 3087
rect 3813 2993 3827 3007
rect 3853 2994 3867 3008
rect 3693 2953 3707 2967
rect 3573 2913 3587 2927
rect 3673 2913 3687 2927
rect 3613 2793 3627 2807
rect 3653 2774 3667 2788
rect 3793 2953 3807 2967
rect 3733 2913 3747 2927
rect 3733 2873 3747 2887
rect 3913 2913 3927 2927
rect 3873 2873 3887 2887
rect 3813 2813 3827 2827
rect 3713 2793 3727 2807
rect 3693 2774 3707 2788
rect 3773 2774 3787 2788
rect 3813 2774 3827 2788
rect 3713 2752 3727 2766
rect 3573 2713 3587 2727
rect 3553 2413 3567 2427
rect 3513 2353 3527 2367
rect 3493 2273 3507 2287
rect 3533 2273 3547 2287
rect 3433 2173 3447 2187
rect 3393 2113 3407 2127
rect 3533 2213 3547 2227
rect 3513 2093 3527 2107
rect 3473 2073 3487 2087
rect 3473 2032 3487 2046
rect 3393 1993 3407 2007
rect 3373 1973 3387 1987
rect 3373 1912 3387 1926
rect 3413 1912 3427 1926
rect 3393 1893 3407 1907
rect 3393 1853 3407 1867
rect 3353 1813 3367 1827
rect 3333 1773 3347 1787
rect 3333 1734 3347 1748
rect 3193 1673 3207 1687
rect 3172 1633 3186 1647
rect 3193 1633 3207 1647
rect 3153 1613 3167 1627
rect 2993 1593 3007 1607
rect 3033 1593 3047 1607
rect 3093 1593 3107 1607
rect 3073 1553 3087 1567
rect 2993 1473 3007 1487
rect 2893 1393 2907 1407
rect 2953 1392 2967 1406
rect 2873 1373 2887 1387
rect 2853 1313 2867 1327
rect 3013 1313 3027 1327
rect 3073 1313 3087 1327
rect 3073 1273 3087 1287
rect 2833 1253 2847 1267
rect 2792 1213 2806 1227
rect 2813 1213 2827 1227
rect 2873 1214 2887 1228
rect 3013 1214 3027 1228
rect 2772 1153 2786 1167
rect 2793 1153 2807 1167
rect 2853 1153 2867 1167
rect 3193 1513 3207 1527
rect 3253 1473 3267 1487
rect 3133 1434 3147 1448
rect 3193 1434 3207 1448
rect 3113 1393 3127 1407
rect 3313 1692 3327 1706
rect 3493 1973 3507 1987
rect 3693 2733 3707 2747
rect 3673 2713 3687 2727
rect 3733 2713 3747 2727
rect 3713 2693 3727 2707
rect 3633 2673 3647 2687
rect 3753 2673 3767 2687
rect 3613 2653 3627 2667
rect 3593 2613 3607 2627
rect 3713 2593 3727 2607
rect 3673 2513 3687 2527
rect 3693 2493 3707 2507
rect 3613 2453 3627 2467
rect 3593 2353 3607 2367
rect 3613 2313 3627 2327
rect 3652 2413 3666 2427
rect 3673 2413 3687 2427
rect 3593 2273 3607 2287
rect 3633 2273 3647 2287
rect 3593 2254 3607 2268
rect 3633 2212 3647 2226
rect 3593 2173 3607 2187
rect 3573 2093 3587 2107
rect 3533 2033 3547 2047
rect 3633 2053 3647 2067
rect 3633 1893 3647 1907
rect 3613 1853 3627 1867
rect 3513 1833 3527 1847
rect 3593 1833 3607 1847
rect 3493 1813 3507 1827
rect 3413 1793 3427 1807
rect 3473 1793 3487 1807
rect 3593 1793 3607 1807
rect 3613 1773 3627 1787
rect 3513 1753 3527 1767
rect 3573 1753 3587 1767
rect 3453 1734 3467 1748
rect 3493 1733 3507 1747
rect 3433 1692 3447 1706
rect 3353 1653 3367 1667
rect 3393 1652 3407 1666
rect 3373 1593 3387 1607
rect 3313 1573 3327 1587
rect 3293 1493 3307 1507
rect 3353 1533 3367 1547
rect 3313 1473 3327 1487
rect 3293 1453 3307 1467
rect 3273 1434 3287 1448
rect 3413 1633 3427 1647
rect 3413 1593 3427 1607
rect 3233 1353 3247 1367
rect 3113 1293 3127 1307
rect 3173 1293 3187 1307
rect 3113 1213 3127 1227
rect 3213 1273 3227 1287
rect 3113 1172 3127 1186
rect 3153 1172 3167 1186
rect 3193 1172 3207 1186
rect 2993 1133 3007 1147
rect 2893 1013 2907 1027
rect 2813 953 2827 967
rect 2753 914 2767 928
rect 2793 914 2807 928
rect 2853 914 2867 928
rect 2913 914 2927 928
rect 2953 914 2967 928
rect 2773 853 2787 867
rect 2713 773 2727 787
rect 2873 872 2887 886
rect 2933 872 2947 886
rect 2773 733 2787 747
rect 2813 733 2827 747
rect 2693 713 2707 727
rect 2813 694 2827 708
rect 2773 673 2787 687
rect 2633 473 2647 487
rect 2593 352 2607 366
rect 2553 193 2567 207
rect 2533 13 2547 27
rect 2633 174 2647 188
rect 2693 493 2707 507
rect 2833 652 2847 666
rect 2973 833 2987 847
rect 2773 573 2787 587
rect 2753 453 2767 467
rect 2713 394 2727 408
rect 2833 413 2847 427
rect 2793 394 2807 408
rect 2693 352 2707 366
rect 2733 352 2747 366
rect 2773 333 2787 347
rect 2673 173 2687 187
rect 2933 652 2947 666
rect 2973 613 2987 627
rect 2873 533 2887 547
rect 2913 453 2927 467
rect 2953 394 2967 408
rect 2993 394 3007 408
rect 2893 352 2907 366
rect 2933 352 2947 366
rect 2873 313 2887 327
rect 2913 313 2927 327
rect 2833 293 2847 307
rect 2993 273 3007 287
rect 3093 1133 3107 1147
rect 3033 1053 3047 1067
rect 3233 1053 3247 1067
rect 3133 953 3147 967
rect 3093 914 3107 928
rect 3172 914 3186 928
rect 3193 914 3207 928
rect 3373 1393 3387 1407
rect 3333 1373 3347 1387
rect 3313 1214 3327 1228
rect 3433 1533 3447 1547
rect 3433 1473 3447 1487
rect 3453 1434 3467 1448
rect 3633 1733 3647 1747
rect 3513 1693 3527 1707
rect 3593 1692 3607 1706
rect 3613 1673 3627 1687
rect 3513 1653 3527 1667
rect 3553 1613 3567 1627
rect 3613 1573 3627 1587
rect 3553 1533 3567 1547
rect 3613 1513 3627 1527
rect 3713 2474 3727 2488
rect 3813 2474 3827 2488
rect 3693 2373 3707 2387
rect 3693 2333 3707 2347
rect 3693 2133 3707 2147
rect 3673 2093 3687 2107
rect 3673 1933 3687 1947
rect 3753 2453 3767 2467
rect 3893 2853 3907 2867
rect 3793 2413 3807 2427
rect 3873 2413 3887 2427
rect 4013 3333 4027 3347
rect 3993 3252 4007 3266
rect 3973 3113 3987 3127
rect 3993 3073 4007 3087
rect 3973 3033 3987 3047
rect 3973 2893 3987 2907
rect 3953 2853 3967 2867
rect 4073 3294 4087 3308
rect 4053 3252 4067 3266
rect 4073 3213 4087 3227
rect 4033 3193 4047 3207
rect 4033 3113 4047 3127
rect 4133 3253 4147 3267
rect 4113 3173 4127 3187
rect 4093 3153 4107 3167
rect 4113 3113 4127 3127
rect 4073 3013 4087 3027
rect 4073 2952 4087 2966
rect 4113 2933 4127 2947
rect 4073 2913 4087 2927
rect 4033 2833 4047 2847
rect 3993 2793 4007 2807
rect 4033 2793 4047 2807
rect 3913 2773 3927 2787
rect 3933 2732 3947 2746
rect 3993 2732 4007 2746
rect 4033 2732 4047 2746
rect 3913 2673 3927 2687
rect 4053 2673 4067 2687
rect 4053 2593 4067 2607
rect 4053 2572 4067 2586
rect 3973 2553 3987 2567
rect 4013 2493 4027 2507
rect 3973 2433 3987 2447
rect 3953 2413 3967 2427
rect 3893 2393 3907 2407
rect 3953 2392 3967 2406
rect 3793 2254 3807 2268
rect 3753 2153 3767 2167
rect 3753 2093 3767 2107
rect 3713 2053 3727 2067
rect 3813 2212 3827 2226
rect 3913 2212 3927 2226
rect 3853 2173 3867 2187
rect 3773 2073 3787 2087
rect 4113 2873 4127 2887
rect 4093 2853 4107 2867
rect 4093 2813 4107 2827
rect 4253 3953 4267 3967
rect 4413 4213 4427 4227
rect 4413 4073 4427 4087
rect 4333 4034 4347 4048
rect 4373 4034 4387 4048
rect 4273 3913 4287 3927
rect 4313 3913 4327 3927
rect 4393 3992 4407 4006
rect 4433 3992 4447 4006
rect 4393 3953 4407 3967
rect 4413 3933 4427 3947
rect 4393 3913 4407 3927
rect 4333 3853 4347 3867
rect 4373 3853 4387 3867
rect 4273 3813 4287 3827
rect 4313 3814 4327 3828
rect 4293 3772 4307 3786
rect 4373 3773 4387 3787
rect 4313 3673 4327 3687
rect 4293 3514 4307 3528
rect 4333 3514 4347 3528
rect 4273 3473 4287 3487
rect 4253 3413 4267 3427
rect 4213 3333 4227 3347
rect 4233 3294 4247 3308
rect 4173 3093 4187 3107
rect 4253 3253 4267 3267
rect 4213 3173 4227 3187
rect 4213 3133 4227 3147
rect 4213 3073 4227 3087
rect 4193 3013 4207 3027
rect 4293 3453 4307 3467
rect 4373 3473 4387 3487
rect 4353 3393 4367 3407
rect 4293 3373 4307 3387
rect 4493 4093 4507 4107
rect 4613 4453 4627 4467
rect 4573 4353 4587 4367
rect 4553 4333 4567 4347
rect 4533 4253 4547 4267
rect 4533 4213 4547 4227
rect 4593 4213 4607 4227
rect 4573 4073 4587 4087
rect 4533 4034 4547 4048
rect 4573 4034 4587 4048
rect 4633 4034 4647 4048
rect 4493 3993 4507 4007
rect 4553 3992 4567 4006
rect 4573 3973 4587 3987
rect 4473 3913 4487 3927
rect 4473 3873 4487 3887
rect 4473 3814 4487 3828
rect 4513 3814 4527 3828
rect 4553 3913 4567 3927
rect 4433 3773 4447 3787
rect 4413 3473 4427 3487
rect 4293 3333 4307 3347
rect 4373 3333 4387 3347
rect 4333 3294 4347 3308
rect 4373 3294 4387 3308
rect 4293 3253 4307 3267
rect 4353 3252 4367 3266
rect 4453 3733 4467 3747
rect 4533 3733 4547 3747
rect 4493 3693 4507 3707
rect 4633 3973 4647 3987
rect 4593 3913 4607 3927
rect 4633 3873 4647 3887
rect 4693 4733 4707 4747
rect 4693 4612 4707 4626
rect 4693 4573 4707 4587
rect 4753 4853 4767 4867
rect 4773 4813 4787 4827
rect 4813 4812 4827 4826
rect 4732 4753 4746 4767
rect 4753 4753 4767 4767
rect 4813 4753 4827 4767
rect 4673 4413 4687 4427
rect 4673 4273 4687 4287
rect 4673 4153 4687 4167
rect 4793 4554 4807 4568
rect 4853 4733 4867 4747
rect 4833 4653 4847 4667
rect 4773 4512 4787 4526
rect 4733 4453 4747 4467
rect 4753 4334 4767 4348
rect 4733 4273 4747 4287
rect 4773 4253 4787 4267
rect 4713 4173 4727 4187
rect 4693 4113 4707 4127
rect 4753 4113 4767 4127
rect 4833 4473 4847 4487
rect 4833 4333 4847 4347
rect 4933 5013 4947 5027
rect 4993 4993 5007 5007
rect 4973 4973 4987 4987
rect 5093 5374 5107 5388
rect 5133 5374 5147 5388
rect 5193 5374 5207 5388
rect 5033 5353 5047 5367
rect 5253 5433 5267 5447
rect 5213 5353 5227 5367
rect 5433 5853 5447 5867
rect 5353 5773 5367 5787
rect 5473 6073 5487 6087
rect 5573 6114 5587 6128
rect 5613 6114 5627 6128
rect 5713 6114 5727 6128
rect 5553 6072 5567 6086
rect 5653 6053 5667 6067
rect 5693 6053 5707 6067
rect 5753 6053 5767 6067
rect 5593 6033 5607 6047
rect 5493 5893 5507 5907
rect 5553 5894 5567 5908
rect 5453 5713 5467 5727
rect 5433 5653 5447 5667
rect 5373 5633 5387 5647
rect 5393 5593 5407 5607
rect 5453 5594 5467 5608
rect 5493 5594 5507 5608
rect 5373 5552 5387 5566
rect 5433 5552 5447 5566
rect 5473 5552 5487 5566
rect 5393 5413 5407 5427
rect 5393 5374 5407 5388
rect 5793 6153 5807 6167
rect 5793 6113 5807 6127
rect 5873 6133 5887 6147
rect 5933 6333 5947 6347
rect 6013 6333 6027 6347
rect 6613 6473 6627 6487
rect 6693 6473 6707 6487
rect 6493 6453 6507 6467
rect 6173 6433 6187 6447
rect 6233 6413 6247 6427
rect 6293 6414 6307 6428
rect 6333 6414 6347 6428
rect 6373 6414 6387 6428
rect 6412 6413 6426 6427
rect 6433 6413 6447 6427
rect 6533 6414 6547 6428
rect 6573 6413 6587 6427
rect 6193 6372 6207 6386
rect 6233 6372 6247 6386
rect 6153 6353 6167 6367
rect 6313 6353 6327 6367
rect 6413 6372 6427 6386
rect 6073 6273 6087 6287
rect 6113 6273 6127 6287
rect 5933 6233 5947 6247
rect 5993 6173 6007 6187
rect 6093 6173 6107 6187
rect 6073 6133 6087 6147
rect 5753 5993 5767 6007
rect 5713 5933 5727 5947
rect 5753 5894 5767 5908
rect 5853 6072 5867 6086
rect 5912 6073 5926 6087
rect 5933 6073 5947 6087
rect 5973 6072 5987 6086
rect 6013 6072 6027 6086
rect 5813 5993 5827 6007
rect 5953 5973 5967 5987
rect 5933 5933 5947 5947
rect 5813 5894 5827 5908
rect 5853 5894 5867 5908
rect 5893 5894 5907 5908
rect 5653 5833 5667 5847
rect 5693 5833 5707 5847
rect 5772 5853 5786 5867
rect 5793 5853 5807 5867
rect 5613 5773 5627 5787
rect 5573 5594 5587 5608
rect 5693 5693 5707 5707
rect 5653 5653 5667 5667
rect 5553 5553 5567 5567
rect 5553 5532 5567 5546
rect 5493 5513 5507 5527
rect 5533 5513 5547 5527
rect 5473 5413 5487 5427
rect 5053 5293 5067 5307
rect 5113 5332 5127 5346
rect 5093 5313 5107 5327
rect 5073 5273 5087 5287
rect 5053 5233 5067 5247
rect 5033 5153 5047 5167
rect 5193 5333 5207 5347
rect 5273 5332 5287 5346
rect 5333 5333 5347 5347
rect 5373 5332 5387 5346
rect 5413 5332 5427 5346
rect 5473 5332 5487 5346
rect 5153 5233 5167 5247
rect 5252 5113 5266 5127
rect 5273 5113 5287 5127
rect 5213 5093 5227 5107
rect 5093 5074 5107 5088
rect 5313 5074 5327 5088
rect 5353 5074 5367 5088
rect 5153 5032 5167 5046
rect 5213 5033 5227 5047
rect 5253 5032 5267 5046
rect 5293 5032 5307 5046
rect 5333 5013 5347 5027
rect 5693 5593 5707 5607
rect 5593 5553 5607 5567
rect 5573 5493 5587 5507
rect 5673 5533 5687 5547
rect 5633 5493 5647 5507
rect 5633 5453 5647 5467
rect 5673 5413 5687 5427
rect 5653 5393 5667 5407
rect 5573 5332 5587 5346
rect 5633 5332 5647 5346
rect 5493 5293 5507 5307
rect 5533 5293 5547 5307
rect 5393 5233 5407 5247
rect 5433 5113 5447 5127
rect 5473 5074 5487 5088
rect 5393 5032 5407 5046
rect 5453 5032 5467 5046
rect 5493 5032 5507 5046
rect 5353 4993 5367 5007
rect 5373 4973 5387 4987
rect 5113 4953 5127 4967
rect 5053 4913 5067 4927
rect 5153 4913 5167 4927
rect 5033 4853 5047 4867
rect 4973 4812 4987 4826
rect 5013 4753 5027 4767
rect 4933 4733 4947 4747
rect 5093 4853 5107 4867
rect 5273 4893 5287 4907
rect 5212 4853 5226 4867
rect 5233 4854 5247 4868
rect 5273 4854 5287 4868
rect 5313 4854 5327 4868
rect 5353 4854 5367 4868
rect 5173 4812 5187 4826
rect 5093 4773 5107 4787
rect 5133 4773 5147 4787
rect 4873 4653 4887 4667
rect 4913 4653 4927 4667
rect 5013 4653 5027 4667
rect 4913 4613 4927 4627
rect 4953 4554 4967 4568
rect 4993 4513 5007 4527
rect 4973 4473 4987 4487
rect 4893 4393 4907 4407
rect 4933 4393 4947 4407
rect 4973 4393 4987 4407
rect 4873 4353 4887 4367
rect 4953 4353 4967 4367
rect 4673 3973 4687 3987
rect 4713 3973 4727 3987
rect 4653 3853 4667 3867
rect 4673 3814 4687 3828
rect 4573 3653 4587 3667
rect 4573 3593 4587 3607
rect 4553 3573 4567 3587
rect 4493 3514 4507 3528
rect 4573 3514 4587 3528
rect 4453 3473 4467 3487
rect 4433 3433 4447 3447
rect 4433 3333 4447 3347
rect 4432 3294 4446 3308
rect 4513 3472 4527 3486
rect 4533 3333 4547 3347
rect 4473 3313 4487 3327
rect 4513 3313 4527 3327
rect 4413 3213 4427 3227
rect 4373 3193 4387 3207
rect 4333 3173 4347 3187
rect 4313 3133 4327 3147
rect 4273 3113 4287 3127
rect 4313 3033 4327 3047
rect 4293 3013 4307 3027
rect 4313 2994 4327 3008
rect 4233 2952 4247 2966
rect 4193 2933 4207 2947
rect 4153 2913 4167 2927
rect 4133 2833 4147 2847
rect 4313 2953 4327 2967
rect 4273 2893 4287 2907
rect 4233 2873 4247 2887
rect 4273 2853 4287 2867
rect 4193 2813 4207 2827
rect 4133 2774 4147 2788
rect 4213 2773 4227 2787
rect 4313 2774 4327 2788
rect 4413 3073 4427 3087
rect 4373 2994 4387 3008
rect 4453 3293 4467 3307
rect 4533 3294 4547 3308
rect 4453 3253 4467 3267
rect 4433 2993 4447 3007
rect 4473 3133 4487 3147
rect 4393 2952 4407 2966
rect 4453 2953 4467 2967
rect 4533 3213 4547 3227
rect 4573 3433 4587 3447
rect 4613 3753 4627 3767
rect 4633 3713 4647 3727
rect 4613 3693 4627 3707
rect 4733 3853 4747 3867
rect 4813 4034 4827 4048
rect 4873 4273 4887 4287
rect 5153 4713 5167 4727
rect 5133 4653 5147 4667
rect 5073 4554 5087 4568
rect 5093 4512 5107 4526
rect 5233 4773 5247 4787
rect 5353 4813 5367 4827
rect 5293 4753 5307 4767
rect 5433 4893 5447 4907
rect 5513 4873 5527 4887
rect 5473 4854 5487 4868
rect 5453 4812 5467 4826
rect 5373 4713 5387 4727
rect 5213 4633 5227 4647
rect 5313 4633 5327 4647
rect 5213 4612 5227 4626
rect 5253 4573 5267 4587
rect 5213 4553 5227 4567
rect 5293 4553 5307 4567
rect 5173 4533 5187 4547
rect 5093 4433 5107 4447
rect 5033 4413 5047 4427
rect 5053 4353 5067 4367
rect 5013 4333 5027 4347
rect 5133 4512 5147 4526
rect 5153 4413 5167 4427
rect 5193 4513 5207 4527
rect 5233 4493 5247 4507
rect 5273 4453 5287 4467
rect 5193 4433 5207 4447
rect 5233 4353 5247 4367
rect 5113 4333 5127 4347
rect 4973 4273 4987 4287
rect 4953 4253 4967 4267
rect 4893 4213 4907 4227
rect 4893 4173 4907 4187
rect 5073 4292 5087 4306
rect 5073 4173 5087 4187
rect 5033 4093 5047 4107
rect 5073 4093 5087 4107
rect 4893 4034 4907 4048
rect 4953 4034 4967 4048
rect 4793 3893 4807 3907
rect 4833 3893 4847 3907
rect 4793 3872 4807 3886
rect 4833 3813 4847 3827
rect 4733 3753 4747 3767
rect 4713 3713 4727 3727
rect 4833 3773 4847 3787
rect 4773 3653 4787 3667
rect 4753 3593 4767 3607
rect 4693 3573 4707 3587
rect 4653 3533 4667 3547
rect 4613 3353 4627 3367
rect 4673 3472 4687 3486
rect 4673 3453 4687 3467
rect 4753 3453 4767 3467
rect 4713 3413 4727 3427
rect 4693 3393 4707 3407
rect 4733 3393 4747 3407
rect 4633 3333 4647 3347
rect 4613 3313 4627 3327
rect 4713 3313 4727 3327
rect 4673 3294 4687 3308
rect 4633 3233 4647 3247
rect 4573 3193 4587 3207
rect 4553 3173 4567 3187
rect 4513 3073 4527 3087
rect 4613 3113 4627 3127
rect 4593 3073 4607 3087
rect 4513 2994 4527 3008
rect 4553 2994 4567 3008
rect 4493 2953 4507 2967
rect 4533 2952 4547 2966
rect 4493 2893 4507 2907
rect 4353 2793 4367 2807
rect 4353 2772 4367 2786
rect 4433 2774 4447 2788
rect 4113 2713 4127 2727
rect 4213 2732 4227 2746
rect 4253 2732 4267 2746
rect 4153 2693 4167 2707
rect 4113 2653 4127 2667
rect 4073 2513 4087 2527
rect 4073 2432 4087 2446
rect 4053 2413 4067 2427
rect 4013 2373 4027 2387
rect 4093 2373 4107 2387
rect 4053 2353 4067 2367
rect 3973 2273 3987 2287
rect 4033 2273 4047 2287
rect 4053 2212 4067 2226
rect 3953 2153 3967 2167
rect 4033 2153 4047 2167
rect 4013 2113 4027 2127
rect 3873 2073 3887 2087
rect 3853 2013 3867 2027
rect 3853 1933 3867 1947
rect 3733 1912 3747 1926
rect 3793 1912 3807 1926
rect 3693 1853 3707 1867
rect 3773 1853 3787 1867
rect 3733 1833 3747 1847
rect 3713 1813 3727 1827
rect 3832 1833 3846 1847
rect 3853 1833 3867 1847
rect 3713 1773 3727 1787
rect 3773 1773 3787 1787
rect 3813 1753 3827 1767
rect 3753 1734 3767 1748
rect 3793 1713 3807 1727
rect 3733 1692 3747 1706
rect 3993 2033 4007 2047
rect 3973 2013 3987 2027
rect 3913 1954 3927 1968
rect 3993 1993 4007 2007
rect 4013 1853 4027 1867
rect 3893 1773 3907 1787
rect 3933 1773 3947 1787
rect 3873 1753 3887 1767
rect 4053 2053 4067 2067
rect 4053 2032 4067 2046
rect 4073 2013 4087 2027
rect 4053 1993 4067 2007
rect 4133 2513 4147 2527
rect 4353 2693 4367 2707
rect 4293 2653 4307 2667
rect 4173 2613 4187 2627
rect 4413 2732 4427 2746
rect 4473 2733 4487 2747
rect 4453 2713 4467 2727
rect 4453 2692 4467 2706
rect 4313 2593 4327 2607
rect 4373 2593 4387 2607
rect 4213 2573 4227 2587
rect 4173 2533 4187 2547
rect 4153 2493 4167 2507
rect 4133 2432 4147 2446
rect 4193 2432 4207 2446
rect 4133 2313 4147 2327
rect 4113 2213 4127 2227
rect 4353 2533 4367 2547
rect 4393 2474 4407 2488
rect 4353 2393 4367 2407
rect 4353 2353 4367 2367
rect 4313 2313 4327 2327
rect 4393 2393 4407 2407
rect 4373 2293 4387 2307
rect 4173 2273 4187 2287
rect 4253 2253 4267 2267
rect 4353 2254 4367 2268
rect 4193 2212 4207 2226
rect 4193 2173 4207 2187
rect 4153 2153 4167 2167
rect 4133 2113 4147 2127
rect 4113 2093 4127 2107
rect 4193 2053 4207 2067
rect 4233 2053 4247 2067
rect 4153 1993 4167 2007
rect 4133 1954 4147 1968
rect 4213 1993 4227 2007
rect 4193 1953 4207 1967
rect 4293 2212 4307 2226
rect 4373 2213 4387 2227
rect 4293 2173 4307 2187
rect 4153 1873 4167 1887
rect 4093 1853 4107 1867
rect 3973 1753 3987 1767
rect 4033 1753 4047 1767
rect 3953 1733 3967 1747
rect 3813 1693 3827 1707
rect 3873 1692 3887 1706
rect 3913 1692 3927 1706
rect 3813 1672 3827 1686
rect 3793 1653 3807 1667
rect 3872 1613 3886 1627
rect 3893 1613 3907 1627
rect 3773 1593 3787 1607
rect 3813 1593 3827 1607
rect 3693 1573 3707 1587
rect 3793 1572 3807 1586
rect 3833 1573 3847 1587
rect 3653 1553 3667 1567
rect 3713 1533 3727 1547
rect 3633 1493 3647 1507
rect 3693 1493 3707 1507
rect 3413 1393 3427 1407
rect 3613 1433 3627 1447
rect 3653 1434 3667 1448
rect 3793 1493 3807 1507
rect 3713 1473 3727 1487
rect 3773 1473 3787 1487
rect 3733 1433 3747 1447
rect 3693 1413 3707 1427
rect 3453 1333 3467 1347
rect 3513 1333 3527 1347
rect 3493 1214 3507 1228
rect 3553 1253 3567 1267
rect 3593 1253 3607 1267
rect 3433 1172 3447 1186
rect 3533 1172 3547 1186
rect 3393 1053 3407 1067
rect 3373 1013 3387 1027
rect 3413 1013 3427 1027
rect 3333 993 3347 1007
rect 3273 953 3287 967
rect 3313 953 3327 967
rect 3273 914 3287 928
rect 3373 914 3387 928
rect 3173 873 3187 887
rect 3113 853 3127 867
rect 3073 833 3087 847
rect 3133 773 3147 787
rect 3073 733 3087 747
rect 3253 872 3267 886
rect 3433 914 3447 928
rect 3433 853 3447 867
rect 3653 1353 3667 1367
rect 3673 1313 3687 1327
rect 3653 1293 3667 1307
rect 3613 1093 3627 1107
rect 3633 1073 3647 1087
rect 3613 1033 3627 1047
rect 3893 1493 3907 1507
rect 3933 1533 3947 1547
rect 3913 1453 3927 1467
rect 4013 1734 4027 1748
rect 4113 1833 4127 1847
rect 4053 1733 4067 1747
rect 4093 1733 4107 1747
rect 4153 1793 4167 1807
rect 4133 1713 4147 1727
rect 4033 1692 4047 1706
rect 4113 1693 4127 1707
rect 4053 1653 4067 1667
rect 4033 1613 4047 1627
rect 4073 1613 4087 1627
rect 4053 1593 4067 1607
rect 3973 1533 3987 1547
rect 3993 1493 4007 1507
rect 3953 1473 3967 1487
rect 3973 1453 3987 1467
rect 3873 1413 3887 1427
rect 3793 1392 3807 1406
rect 3793 1353 3807 1367
rect 3793 1293 3807 1307
rect 3833 1293 3847 1307
rect 3733 1253 3747 1267
rect 3913 1253 3927 1267
rect 3753 1233 3767 1247
rect 3713 1214 3727 1228
rect 3833 1213 3847 1227
rect 3873 1214 3887 1228
rect 3993 1313 4007 1327
rect 3673 1053 3687 1067
rect 3733 1053 3747 1067
rect 3753 993 3767 1007
rect 3653 953 3667 967
rect 3733 953 3747 967
rect 3613 914 3627 928
rect 3533 853 3547 867
rect 3413 833 3427 847
rect 3493 833 3507 847
rect 3633 793 3647 807
rect 3813 1093 3827 1107
rect 3813 1013 3827 1027
rect 3773 973 3787 987
rect 3933 1172 3947 1186
rect 3973 1172 3987 1186
rect 3933 1113 3947 1127
rect 3973 1113 3987 1127
rect 4073 1453 4087 1467
rect 4033 1434 4047 1448
rect 4133 1533 4147 1547
rect 4133 1473 4147 1487
rect 4113 1434 4127 1448
rect 4053 1393 4067 1407
rect 4033 1313 4047 1327
rect 4033 1233 4047 1247
rect 4093 1373 4107 1387
rect 4133 1293 4147 1307
rect 4093 1214 4107 1228
rect 4013 1153 4027 1167
rect 4073 1153 4087 1167
rect 4013 1093 4027 1107
rect 3993 1073 4007 1087
rect 3933 1013 3947 1027
rect 4113 1013 4127 1027
rect 3833 953 3847 967
rect 3873 953 3887 967
rect 3793 872 3807 886
rect 3793 853 3807 867
rect 3753 813 3767 827
rect 3733 773 3747 787
rect 3713 753 3727 767
rect 3193 733 3207 747
rect 3513 733 3527 747
rect 3253 694 3267 708
rect 3293 694 3307 708
rect 3373 694 3387 708
rect 3413 694 3427 708
rect 3453 694 3467 708
rect 3493 694 3507 708
rect 3213 673 3227 687
rect 3353 673 3367 687
rect 3313 652 3327 666
rect 3373 653 3387 667
rect 3353 633 3367 647
rect 3433 633 3447 647
rect 3153 613 3167 627
rect 3253 613 3267 627
rect 3113 573 3127 587
rect 3033 533 3047 547
rect 3113 513 3127 527
rect 3033 493 3047 507
rect 3073 453 3087 467
rect 3073 413 3087 427
rect 3033 393 3047 407
rect 3093 352 3107 366
rect 3713 713 3727 727
rect 3553 694 3567 708
rect 3593 694 3607 708
rect 3673 693 3687 707
rect 3773 773 3787 787
rect 3813 773 3827 787
rect 3753 693 3767 707
rect 3513 652 3527 666
rect 3573 652 3587 666
rect 3733 652 3747 666
rect 3973 993 3987 1007
rect 4253 1953 4267 1967
rect 4373 2153 4387 2167
rect 4413 2353 4427 2367
rect 4573 2833 4587 2847
rect 4613 3033 4627 3047
rect 4613 2994 4627 3008
rect 4613 2953 4627 2967
rect 4593 2793 4607 2807
rect 4693 3193 4707 3207
rect 4873 3973 4887 3987
rect 4933 3973 4947 3987
rect 4913 3933 4927 3947
rect 4873 3893 4887 3907
rect 4853 3713 4867 3727
rect 5193 4334 5207 4348
rect 5233 4334 5247 4348
rect 5293 4334 5307 4348
rect 5253 4292 5267 4306
rect 5153 4233 5167 4247
rect 5213 4233 5227 4247
rect 5473 4573 5487 4587
rect 5333 4554 5347 4568
rect 5373 4554 5387 4568
rect 5333 4493 5347 4507
rect 5393 4493 5407 4507
rect 5653 5193 5667 5207
rect 5733 5833 5747 5847
rect 5733 5613 5747 5627
rect 5873 5852 5887 5866
rect 5933 5773 5947 5787
rect 6093 6013 6107 6027
rect 6073 5894 6087 5908
rect 6293 6213 6307 6227
rect 6153 6113 6167 6127
rect 6253 6113 6267 6127
rect 6233 6073 6247 6087
rect 6153 6033 6167 6047
rect 6193 6033 6207 6047
rect 5873 5753 5887 5767
rect 5953 5753 5967 5767
rect 5813 5633 5827 5647
rect 5793 5613 5807 5627
rect 5753 5593 5767 5607
rect 5833 5594 5847 5608
rect 5773 5552 5787 5566
rect 5813 5552 5827 5566
rect 5733 5493 5747 5507
rect 5733 5413 5747 5427
rect 5713 5393 5727 5407
rect 5833 5533 5847 5547
rect 5813 5493 5827 5507
rect 5793 5374 5807 5388
rect 5753 5332 5767 5346
rect 5693 5293 5707 5307
rect 5793 5293 5807 5307
rect 5693 5253 5707 5267
rect 5673 5133 5687 5147
rect 5593 5093 5607 5107
rect 5693 5093 5707 5107
rect 5733 5093 5747 5107
rect 5793 5093 5807 5107
rect 5633 5074 5647 5088
rect 5693 5032 5707 5046
rect 5753 5032 5767 5046
rect 6033 5852 6047 5866
rect 5913 5633 5927 5647
rect 5993 5633 6007 5647
rect 5893 5594 5907 5608
rect 5873 5533 5887 5547
rect 5933 5594 5947 5608
rect 5953 5552 5967 5566
rect 5993 5552 6007 5566
rect 5973 5493 5987 5507
rect 5893 5453 5907 5467
rect 5953 5453 5967 5467
rect 5853 5413 5867 5427
rect 5873 5374 5887 5388
rect 5913 5374 5927 5388
rect 5673 4913 5687 4927
rect 5713 4913 5727 4927
rect 5613 4874 5627 4888
rect 5573 4854 5587 4868
rect 5613 4853 5627 4867
rect 5753 4873 5767 4887
rect 5853 5332 5867 5346
rect 5893 5332 5907 5346
rect 5953 5333 5967 5347
rect 5853 5293 5867 5307
rect 5673 4812 5687 4826
rect 5553 4793 5567 4807
rect 5593 4793 5607 4807
rect 5633 4793 5647 4807
rect 5813 4812 5827 4826
rect 5513 4573 5527 4587
rect 5593 4633 5607 4647
rect 5473 4493 5487 4507
rect 5433 4413 5447 4427
rect 5413 4373 5427 4387
rect 5373 4334 5387 4348
rect 5353 4292 5367 4306
rect 5433 4293 5447 4307
rect 5293 4232 5307 4246
rect 5253 4093 5267 4107
rect 5173 4034 5187 4048
rect 5053 3992 5067 4006
rect 5133 3993 5147 4007
rect 5173 3973 5187 3987
rect 4993 3953 5007 3967
rect 4973 3913 4987 3927
rect 4953 3893 4967 3907
rect 5013 3873 5027 3887
rect 4913 3814 4927 3828
rect 4993 3853 5007 3867
rect 4993 3813 5007 3827
rect 5033 3814 5047 3828
rect 5093 3814 5107 3828
rect 5133 3814 5147 3828
rect 4973 3772 4987 3786
rect 5013 3772 5027 3786
rect 4933 3633 4947 3647
rect 4993 3633 5007 3647
rect 5033 3633 5047 3647
rect 4873 3613 4887 3627
rect 4913 3613 4927 3627
rect 4833 3593 4847 3607
rect 4793 3513 4807 3527
rect 4853 3533 4867 3547
rect 4793 3473 4807 3487
rect 4773 3294 4787 3308
rect 4753 3273 4767 3287
rect 4673 3113 4687 3127
rect 4653 3093 4667 3107
rect 4653 3013 4667 3027
rect 4713 3053 4727 3067
rect 4713 2994 4727 3008
rect 4753 2993 4767 3007
rect 4733 2952 4747 2966
rect 4713 2933 4727 2947
rect 4693 2873 4707 2887
rect 4633 2853 4647 2867
rect 4693 2852 4707 2866
rect 4613 2774 4627 2788
rect 4533 2733 4547 2747
rect 4493 2693 4507 2707
rect 4473 2573 4487 2587
rect 4513 2533 4527 2547
rect 4473 2473 4487 2487
rect 4553 2693 4567 2707
rect 4693 2733 4707 2747
rect 4873 3453 4887 3467
rect 4833 3353 4847 3367
rect 4833 3294 4847 3308
rect 4873 3233 4887 3247
rect 4873 3193 4887 3207
rect 4813 3073 4827 3087
rect 4793 3053 4807 3067
rect 4813 2993 4827 3007
rect 4853 3073 4867 3087
rect 4933 3533 4947 3547
rect 5033 3593 5047 3607
rect 4933 3472 4947 3486
rect 4973 3472 4987 3486
rect 5113 3772 5127 3786
rect 5093 3753 5107 3767
rect 5073 3713 5087 3727
rect 5053 3573 5067 3587
rect 5353 4034 5367 4048
rect 5253 3973 5267 3987
rect 5273 3873 5287 3887
rect 5213 3813 5227 3827
rect 5193 3772 5207 3786
rect 5413 4033 5427 4047
rect 5413 3992 5427 4006
rect 5533 4512 5547 4526
rect 5573 4512 5587 4526
rect 5473 4413 5487 4427
rect 5573 4473 5587 4487
rect 5513 4453 5527 4467
rect 5533 4433 5547 4447
rect 5493 4333 5507 4347
rect 6193 5894 6207 5908
rect 6233 5893 6247 5907
rect 6133 5813 6147 5827
rect 6133 5693 6147 5707
rect 6113 5633 6127 5647
rect 6073 5593 6087 5607
rect 6113 5594 6127 5608
rect 6153 5594 6167 5608
rect 6213 5852 6227 5866
rect 6473 6372 6487 6386
rect 6433 6173 6447 6187
rect 6453 6153 6467 6167
rect 6313 6133 6327 6147
rect 6353 6072 6367 6086
rect 6293 5973 6307 5987
rect 6653 6414 6667 6428
rect 6633 6372 6647 6386
rect 6673 6372 6687 6386
rect 6613 6273 6627 6287
rect 6713 6293 6727 6307
rect 6773 6293 6787 6307
rect 6633 6213 6647 6227
rect 6573 6153 6587 6167
rect 6533 6133 6547 6147
rect 6513 6114 6527 6128
rect 6413 6053 6427 6067
rect 6453 6053 6467 6067
rect 6353 5913 6367 5927
rect 6273 5893 6287 5907
rect 6313 5894 6327 5908
rect 6393 5893 6407 5907
rect 6253 5813 6267 5827
rect 6293 5852 6307 5866
rect 6333 5852 6347 5866
rect 6373 5852 6387 5866
rect 6193 5594 6207 5608
rect 6373 5653 6387 5667
rect 6313 5633 6327 5647
rect 6073 5553 6087 5567
rect 6033 5493 6047 5507
rect 6013 5453 6027 5467
rect 6293 5593 6307 5607
rect 6333 5613 6347 5627
rect 6533 6072 6547 6086
rect 6453 6032 6467 6046
rect 6493 6033 6507 6047
rect 6533 6033 6547 6047
rect 6453 5893 6467 5907
rect 6493 5894 6507 5908
rect 6573 6013 6587 6027
rect 6453 5853 6467 5867
rect 6433 5793 6447 5807
rect 6413 5613 6427 5627
rect 6233 5533 6247 5547
rect 6273 5533 6287 5547
rect 6313 5533 6327 5547
rect 6193 5493 6207 5507
rect 6133 5473 6147 5487
rect 6273 5493 6287 5507
rect 6093 5433 6107 5447
rect 6233 5433 6247 5447
rect 6033 5374 6047 5388
rect 6073 5374 6087 5388
rect 6112 5373 6126 5387
rect 6133 5373 6147 5387
rect 6193 5374 6207 5388
rect 5973 5293 5987 5307
rect 5893 5073 5907 5087
rect 5973 5074 5987 5088
rect 5913 5032 5927 5046
rect 5993 5033 6007 5047
rect 6113 5332 6127 5346
rect 6053 5193 6067 5207
rect 6093 5133 6107 5147
rect 6213 5332 6227 5346
rect 6233 5313 6247 5327
rect 6173 5273 6187 5287
rect 6213 5153 6227 5167
rect 6133 5073 6147 5087
rect 6053 5053 6067 5067
rect 6033 5033 6047 5047
rect 6013 4973 6027 4987
rect 6013 4913 6027 4927
rect 5873 4854 5887 4868
rect 5933 4854 5947 4868
rect 5973 4854 5987 4868
rect 5853 4773 5867 4787
rect 5753 4753 5767 4767
rect 5773 4733 5787 4747
rect 5593 4373 5607 4387
rect 5693 4554 5707 4568
rect 5793 4713 5807 4727
rect 5773 4554 5787 4568
rect 6033 4853 6047 4867
rect 5873 4633 5887 4647
rect 5833 4593 5847 4607
rect 5753 4513 5767 4527
rect 5872 4554 5886 4568
rect 5913 4812 5927 4826
rect 5953 4812 5967 4826
rect 6013 4812 6027 4826
rect 5933 4793 5947 4807
rect 5913 4773 5927 4787
rect 5893 4553 5907 4567
rect 5813 4512 5827 4526
rect 5833 4493 5847 4507
rect 5813 4453 5827 4467
rect 5793 4433 5807 4447
rect 5633 4393 5647 4407
rect 5613 4334 5627 4348
rect 5473 4292 5487 4306
rect 5513 4292 5527 4306
rect 5553 4292 5567 4306
rect 5613 4292 5627 4306
rect 5673 4413 5687 4427
rect 5713 4334 5727 4348
rect 5753 4334 5767 4348
rect 5653 4292 5667 4306
rect 5693 4292 5707 4306
rect 5733 4292 5747 4306
rect 5753 4273 5767 4287
rect 5453 4233 5467 4247
rect 5633 4233 5647 4247
rect 5733 4153 5747 4167
rect 5513 4133 5527 4147
rect 5633 4133 5647 4147
rect 5473 4093 5487 4107
rect 5613 4093 5627 4107
rect 5673 4034 5687 4048
rect 5393 3973 5407 3987
rect 5333 3953 5347 3967
rect 5413 3814 5427 3828
rect 5493 3992 5507 4006
rect 5593 3992 5607 4006
rect 5653 3992 5667 4006
rect 5533 3973 5547 3987
rect 5673 3973 5687 3987
rect 5513 3814 5527 3828
rect 5433 3772 5447 3786
rect 5493 3772 5507 3786
rect 5493 3733 5507 3747
rect 5233 3693 5247 3707
rect 5433 3693 5447 3707
rect 5473 3693 5487 3707
rect 5173 3653 5187 3667
rect 5233 3613 5247 3627
rect 5093 3553 5107 3567
rect 5133 3533 5147 3547
rect 5193 3533 5207 3547
rect 5073 3514 5087 3528
rect 5133 3514 5147 3528
rect 5153 3472 5167 3486
rect 5073 3453 5087 3467
rect 4953 3433 4967 3447
rect 5033 3433 5047 3447
rect 4933 3353 4947 3367
rect 4853 3013 4867 3027
rect 4873 2994 4887 3008
rect 5333 3593 5347 3607
rect 5253 3573 5267 3587
rect 5333 3553 5347 3567
rect 5373 3553 5387 3567
rect 5253 3513 5267 3527
rect 5333 3514 5347 3528
rect 5233 3473 5247 3487
rect 5273 3472 5287 3486
rect 5293 3453 5307 3467
rect 5213 3393 5227 3407
rect 5193 3373 5207 3387
rect 5193 3333 5207 3347
rect 5013 3294 5027 3308
rect 5093 3294 5107 3308
rect 5133 3294 5147 3308
rect 5073 3273 5087 3287
rect 4993 3252 5007 3266
rect 5073 3233 5087 3247
rect 4953 3213 4967 3227
rect 5033 3213 5047 3227
rect 5253 3294 5267 3308
rect 5393 3514 5407 3528
rect 5473 3514 5487 3528
rect 5573 3833 5587 3847
rect 5613 3814 5627 3828
rect 5593 3772 5607 3786
rect 5633 3733 5647 3747
rect 5533 3713 5547 3727
rect 5593 3693 5607 3707
rect 5533 3633 5547 3647
rect 5313 3433 5327 3447
rect 5373 3433 5387 3447
rect 5453 3472 5467 3486
rect 5453 3413 5467 3427
rect 5493 3413 5507 3427
rect 5393 3393 5407 3407
rect 5373 3333 5387 3347
rect 5473 3333 5487 3347
rect 5353 3294 5367 3308
rect 5433 3294 5447 3308
rect 5053 3193 5067 3207
rect 5313 3233 5327 3247
rect 5273 3193 5287 3207
rect 5313 3153 5327 3167
rect 5073 3113 5087 3127
rect 5033 3053 5047 3067
rect 4953 2994 4967 3008
rect 4773 2833 4787 2847
rect 4753 2774 4767 2788
rect 4853 2952 4867 2966
rect 4933 2953 4947 2967
rect 5133 3033 5147 3047
rect 5213 3033 5227 3047
rect 5093 2994 5107 3008
rect 5173 2994 5187 3008
rect 4713 2713 4727 2727
rect 4753 2713 4767 2727
rect 4633 2693 4647 2707
rect 4613 2613 4627 2627
rect 4593 2553 4607 2567
rect 4573 2513 4587 2527
rect 4613 2513 4627 2527
rect 4553 2493 4567 2507
rect 4473 2413 4487 2427
rect 4513 2373 4527 2387
rect 4413 2253 4427 2267
rect 4453 2254 4467 2268
rect 4493 2254 4507 2268
rect 4393 2133 4407 2147
rect 4313 2073 4327 2087
rect 4313 2013 4327 2027
rect 4453 2193 4467 2207
rect 4313 1912 4327 1926
rect 4413 1953 4427 1967
rect 4293 1893 4307 1907
rect 4273 1653 4287 1667
rect 4233 1553 4247 1567
rect 4193 1533 4207 1547
rect 4173 1453 4187 1467
rect 4233 1493 4247 1507
rect 4273 1493 4287 1507
rect 4193 1433 4207 1447
rect 4313 1813 4327 1827
rect 4293 1453 4307 1467
rect 4173 1273 4187 1287
rect 4153 1133 4167 1147
rect 4173 933 4187 947
rect 4033 913 4047 927
rect 3953 872 3967 886
rect 3953 833 3967 847
rect 3873 773 3887 787
rect 3873 733 3887 747
rect 3793 713 3807 727
rect 3913 694 3927 708
rect 3793 652 3807 666
rect 3613 613 3627 627
rect 3673 613 3687 627
rect 3513 513 3527 527
rect 3193 473 3207 487
rect 3253 473 3267 487
rect 3493 473 3507 487
rect 3093 333 3107 347
rect 3153 333 3167 347
rect 3053 313 3067 327
rect 3053 213 3067 227
rect 2653 132 2667 146
rect 2893 73 2907 87
rect 3093 174 3107 188
rect 3133 174 3147 188
rect 3273 453 3287 467
rect 3393 453 3407 467
rect 3233 394 3247 408
rect 3313 394 3327 408
rect 3453 394 3467 408
rect 3593 473 3607 487
rect 3553 394 3567 408
rect 3893 652 3907 666
rect 4033 853 4047 867
rect 3972 813 3986 827
rect 3993 813 4007 827
rect 3973 773 3987 787
rect 4033 733 4047 747
rect 4253 1392 4267 1406
rect 4353 1793 4367 1807
rect 4393 1853 4407 1867
rect 4393 1793 4407 1807
rect 4413 1733 4427 1747
rect 4353 1653 4367 1667
rect 4413 1693 4427 1707
rect 4493 2193 4507 2207
rect 4473 2173 4487 2187
rect 4473 2073 4487 2087
rect 4473 1973 4487 1987
rect 4453 1953 4467 1967
rect 4553 2413 4567 2427
rect 4533 2293 4547 2307
rect 4533 2272 4547 2286
rect 4593 2353 4607 2367
rect 4593 2313 4607 2327
rect 4693 2513 4707 2527
rect 4633 2353 4647 2367
rect 4613 2293 4627 2307
rect 4573 2273 4587 2287
rect 4633 2273 4647 2287
rect 4613 2254 4627 2268
rect 4553 2173 4567 2187
rect 4553 2152 4567 2166
rect 4533 2073 4547 2087
rect 4633 2193 4647 2207
rect 4713 2432 4727 2446
rect 4693 2373 4707 2387
rect 4673 2333 4687 2347
rect 4673 2273 4687 2287
rect 4653 2153 4667 2167
rect 4653 2132 4667 2146
rect 4573 2113 4587 2127
rect 4613 2033 4627 2047
rect 4593 1993 4607 2007
rect 4493 1912 4507 1926
rect 4553 1913 4567 1927
rect 4473 1873 4487 1887
rect 4453 1733 4467 1747
rect 4433 1673 4447 1687
rect 4453 1653 4467 1667
rect 4413 1633 4427 1647
rect 4653 1993 4667 2007
rect 4773 2673 4787 2687
rect 4773 2432 4787 2446
rect 5013 2952 5027 2966
rect 5073 2953 5087 2967
rect 4973 2913 4987 2927
rect 4913 2853 4927 2867
rect 4913 2774 4927 2788
rect 4873 2713 4887 2727
rect 4953 2732 4967 2746
rect 4933 2713 4947 2727
rect 4893 2653 4907 2667
rect 4853 2593 4867 2607
rect 4813 2433 4827 2447
rect 4813 2393 4827 2407
rect 4753 2373 4767 2387
rect 4773 2353 4787 2367
rect 4713 2233 4727 2247
rect 4713 2212 4727 2226
rect 4693 2193 4707 2207
rect 4693 1993 4707 2007
rect 4653 1972 4667 1986
rect 4613 1953 4627 1967
rect 4593 1913 4607 1927
rect 4673 1912 4687 1926
rect 4573 1873 4587 1887
rect 4633 1873 4647 1887
rect 4573 1833 4587 1847
rect 4533 1813 4547 1827
rect 4593 1813 4607 1827
rect 4513 1692 4527 1706
rect 4573 1692 4587 1706
rect 4513 1671 4527 1685
rect 4473 1613 4487 1627
rect 4353 1593 4367 1607
rect 4393 1593 4407 1607
rect 4493 1593 4507 1607
rect 4333 1513 4347 1527
rect 4333 1373 4347 1387
rect 4313 1353 4327 1367
rect 4453 1513 4467 1527
rect 4413 1434 4427 1448
rect 4373 1353 4387 1367
rect 4353 1333 4367 1347
rect 4333 1273 4347 1287
rect 4273 1253 4287 1267
rect 4233 1214 4247 1228
rect 4353 1253 4367 1267
rect 4333 1233 4347 1247
rect 4313 1214 4327 1228
rect 4253 1153 4267 1167
rect 4333 1093 4347 1107
rect 4433 1392 4447 1406
rect 4493 1373 4507 1387
rect 4453 1353 4467 1367
rect 4393 1313 4407 1327
rect 4393 1273 4407 1287
rect 4373 1214 4387 1228
rect 4373 1172 4387 1186
rect 4573 1553 4587 1567
rect 4533 1513 4547 1527
rect 4453 1233 4467 1247
rect 4513 1253 4527 1267
rect 4693 1813 4707 1827
rect 4653 1734 4667 1748
rect 4673 1693 4687 1707
rect 4653 1653 4667 1667
rect 4653 1593 4667 1607
rect 4793 2212 4807 2226
rect 4753 2193 4767 2207
rect 4873 2373 4887 2387
rect 4913 2313 4927 2327
rect 4853 2293 4867 2307
rect 4793 2173 4807 2187
rect 4833 2173 4847 2187
rect 5153 2952 5167 2966
rect 5253 3013 5267 3027
rect 5373 3252 5387 3266
rect 5413 3252 5427 3266
rect 5513 3153 5527 3167
rect 5553 3593 5567 3607
rect 5633 3633 5647 3647
rect 5633 3514 5647 3528
rect 5733 3953 5747 3967
rect 6113 5032 6127 5046
rect 6133 4993 6147 5007
rect 6093 4854 6107 4868
rect 6193 5032 6207 5046
rect 6173 4993 6187 5007
rect 6153 4973 6167 4987
rect 6173 4933 6187 4947
rect 6213 4893 6227 4907
rect 6053 4733 6067 4747
rect 6113 4713 6127 4727
rect 5993 4633 6007 4647
rect 6033 4633 6047 4647
rect 5993 4593 6007 4607
rect 6293 5413 6307 5427
rect 6393 5552 6407 5566
rect 6373 5513 6387 5527
rect 6333 5493 6347 5507
rect 6333 5374 6347 5388
rect 6373 5374 6387 5388
rect 6293 5333 6307 5347
rect 6353 5332 6367 5346
rect 6273 5313 6287 5327
rect 6373 5273 6387 5287
rect 6253 5113 6267 5127
rect 6313 5074 6327 5088
rect 6373 5074 6387 5088
rect 6293 5032 6307 5046
rect 6293 5013 6307 5027
rect 6333 4993 6347 5007
rect 6353 4953 6367 4967
rect 6333 4933 6347 4947
rect 6253 4913 6267 4927
rect 6233 4853 6247 4867
rect 6333 4893 6347 4907
rect 6293 4854 6307 4868
rect 6233 4813 6247 4827
rect 6253 4793 6267 4807
rect 6273 4753 6287 4767
rect 6373 4913 6387 4927
rect 6353 4773 6367 4787
rect 6313 4733 6327 4747
rect 6413 5513 6427 5527
rect 6553 5853 6567 5867
rect 6513 5793 6527 5807
rect 6473 5773 6487 5787
rect 6633 6114 6647 6128
rect 6673 6114 6687 6128
rect 6633 6053 6647 6067
rect 6613 6013 6627 6027
rect 6693 6013 6707 6027
rect 6653 5894 6667 5908
rect 6733 6053 6747 6067
rect 6713 5893 6727 5907
rect 6773 5893 6787 5907
rect 6473 5752 6487 5766
rect 6552 5753 6566 5767
rect 6573 5753 6587 5767
rect 6593 5713 6607 5727
rect 6493 5653 6507 5667
rect 6513 5614 6527 5628
rect 6493 5593 6507 5607
rect 6533 5593 6547 5607
rect 6633 5793 6647 5807
rect 6733 5833 6747 5847
rect 6673 5773 6687 5787
rect 6653 5753 6667 5767
rect 6633 5673 6647 5687
rect 6473 5513 6487 5527
rect 6613 5553 6627 5567
rect 6573 5513 6587 5527
rect 6613 5513 6627 5527
rect 6553 5473 6567 5487
rect 6493 5433 6507 5447
rect 6453 5413 6467 5427
rect 6513 5393 6527 5407
rect 6473 5332 6487 5346
rect 6513 5332 6527 5346
rect 6413 5293 6427 5307
rect 6413 5173 6427 5187
rect 6453 5113 6467 5127
rect 6493 5313 6507 5327
rect 6493 5173 6507 5187
rect 6553 5153 6567 5167
rect 6473 5013 6487 5027
rect 6433 4993 6447 5007
rect 6513 4993 6527 5007
rect 6413 4913 6427 4927
rect 6393 4893 6407 4907
rect 6493 4953 6507 4967
rect 6553 4953 6567 4967
rect 6433 4873 6447 4887
rect 6453 4854 6467 4868
rect 6513 4913 6527 4927
rect 6532 4893 6546 4907
rect 6553 4893 6567 4907
rect 6433 4812 6447 4826
rect 6453 4773 6467 4787
rect 6433 4713 6447 4727
rect 6273 4693 6287 4707
rect 6373 4693 6387 4707
rect 6253 4673 6267 4687
rect 6233 4593 6247 4607
rect 6153 4573 6167 4587
rect 6373 4613 6387 4627
rect 6453 4613 6467 4627
rect 6393 4593 6407 4607
rect 6093 4553 6107 4567
rect 6133 4554 6147 4568
rect 6193 4554 6207 4568
rect 5853 4373 5867 4387
rect 5933 4372 5947 4386
rect 5813 4333 5827 4347
rect 5873 4334 5887 4348
rect 5913 4334 5927 4348
rect 5813 4292 5827 4306
rect 5793 4273 5807 4287
rect 5813 4113 5827 4127
rect 5793 4073 5807 4087
rect 5773 4033 5787 4047
rect 5893 4273 5907 4287
rect 5853 4213 5867 4227
rect 5873 4073 5887 4087
rect 5833 4033 5847 4047
rect 5813 3992 5827 4006
rect 5813 3953 5827 3967
rect 5753 3893 5767 3907
rect 5693 3833 5707 3847
rect 5733 3833 5747 3847
rect 5773 3814 5787 3828
rect 5853 3893 5867 3907
rect 5833 3813 5847 3827
rect 5693 3793 5707 3807
rect 5673 3513 5687 3527
rect 5613 3472 5627 3486
rect 5553 3393 5567 3407
rect 5673 3473 5687 3487
rect 5653 3373 5667 3387
rect 5613 3294 5627 3308
rect 5653 3253 5667 3267
rect 5633 3233 5647 3247
rect 5593 3193 5607 3207
rect 5613 3153 5627 3167
rect 5593 3093 5607 3107
rect 5333 3073 5347 3087
rect 5533 3073 5547 3087
rect 5493 3033 5507 3047
rect 5553 3033 5567 3047
rect 5453 2994 5467 3008
rect 5393 2973 5407 2987
rect 5253 2953 5267 2967
rect 5173 2933 5187 2947
rect 5213 2933 5227 2947
rect 5133 2853 5147 2867
rect 5093 2833 5107 2847
rect 4973 2673 4987 2687
rect 4953 2513 4967 2527
rect 5113 2732 5127 2746
rect 5053 2613 5067 2627
rect 4973 2473 4987 2487
rect 5013 2474 5027 2488
rect 4953 2413 4967 2427
rect 4993 2393 5007 2407
rect 4933 2273 4947 2287
rect 4973 2273 4987 2287
rect 4933 2212 4947 2226
rect 4853 2113 4867 2127
rect 4833 2093 4847 2107
rect 4833 2053 4847 2067
rect 4753 1973 4767 1987
rect 4733 1954 4747 1968
rect 4733 1873 4747 1887
rect 4853 1972 4867 1986
rect 4813 1954 4827 1968
rect 4893 2172 4907 2186
rect 4793 1912 4807 1926
rect 4913 2153 4927 2167
rect 4913 2053 4927 2067
rect 4973 2053 4987 2067
rect 4913 1973 4927 1987
rect 4933 1953 4947 1967
rect 5073 2433 5087 2447
rect 5033 2393 5047 2407
rect 5033 2313 5047 2327
rect 5013 2253 5027 2267
rect 5013 2213 5027 2227
rect 5053 2133 5067 2147
rect 5013 2093 5027 2107
rect 5113 2432 5127 2446
rect 5113 2373 5127 2387
rect 5233 2833 5247 2847
rect 5213 2732 5227 2746
rect 5173 2613 5187 2627
rect 5173 2513 5187 2527
rect 5633 3133 5647 3147
rect 5753 3772 5767 3786
rect 5793 3693 5807 3707
rect 5793 3553 5807 3567
rect 5833 3553 5847 3567
rect 5713 3514 5727 3528
rect 5753 3514 5767 3528
rect 5833 3473 5847 3487
rect 5793 3433 5807 3447
rect 5773 3413 5787 3427
rect 5813 3393 5827 3407
rect 5793 3373 5807 3387
rect 5973 4453 5987 4467
rect 5953 4273 5967 4287
rect 5933 4213 5947 4227
rect 6033 4393 6047 4407
rect 6013 4373 6027 4387
rect 5993 4333 6007 4347
rect 6153 4512 6167 4526
rect 6113 4473 6127 4487
rect 6073 4373 6087 4387
rect 6053 4353 6067 4367
rect 6153 4473 6167 4487
rect 6273 4554 6287 4568
rect 6233 4512 6247 4526
rect 6133 4433 6147 4447
rect 6193 4433 6207 4447
rect 6113 4333 6127 4347
rect 6093 4292 6107 4306
rect 6153 4393 6167 4407
rect 6053 4252 6067 4266
rect 5993 4193 6007 4207
rect 5973 4153 5987 4167
rect 5933 4054 5947 4068
rect 5973 4053 5987 4067
rect 5893 4033 5907 4047
rect 5933 4033 5947 4047
rect 6033 4013 6047 4027
rect 5893 3993 5907 4007
rect 5913 3973 5927 3987
rect 5953 3973 5967 3987
rect 5993 3973 6007 3987
rect 5933 3853 5947 3867
rect 6033 3973 6047 3987
rect 6013 3913 6027 3927
rect 6073 4213 6087 4227
rect 6093 4113 6107 4127
rect 6233 4393 6247 4407
rect 6213 4373 6227 4387
rect 6193 4353 6207 4367
rect 6293 4373 6307 4387
rect 6253 4334 6267 4348
rect 6193 4292 6207 4306
rect 6273 4293 6287 4307
rect 6253 4273 6267 4287
rect 6173 4253 6187 4267
rect 6213 4173 6227 4187
rect 6153 4093 6167 4107
rect 6193 4093 6207 4107
rect 6173 4073 6187 4087
rect 6073 3933 6087 3947
rect 6013 3873 6027 3887
rect 6053 3873 6067 3887
rect 5913 3772 5927 3786
rect 5933 3593 5947 3607
rect 5913 3533 5927 3547
rect 5993 3773 6007 3787
rect 6073 3814 6087 3828
rect 6093 3773 6107 3787
rect 6093 3733 6107 3747
rect 6053 3693 6067 3707
rect 6133 3973 6147 3987
rect 6193 3953 6207 3967
rect 6133 3933 6147 3947
rect 6153 3913 6167 3927
rect 6153 3813 6167 3827
rect 6353 4453 6367 4467
rect 6333 4433 6347 4447
rect 6313 4293 6327 4307
rect 6293 4233 6307 4247
rect 6273 4173 6287 4187
rect 6253 4093 6267 4107
rect 6393 4512 6407 4526
rect 6393 4433 6407 4447
rect 6373 4393 6387 4407
rect 6433 4413 6447 4427
rect 6473 4413 6487 4427
rect 6453 4372 6467 4386
rect 6433 4353 6447 4367
rect 6453 4333 6467 4347
rect 6353 4293 6367 4307
rect 6393 4273 6407 4287
rect 6333 4253 6347 4267
rect 6333 4213 6347 4227
rect 6273 4034 6287 4048
rect 6313 4033 6327 4047
rect 6413 4213 6427 4227
rect 6393 4193 6407 4207
rect 6253 3993 6267 4007
rect 6272 3953 6286 3967
rect 6293 3953 6307 3967
rect 6253 3913 6267 3927
rect 6212 3853 6226 3867
rect 6233 3853 6247 3867
rect 6273 3853 6287 3867
rect 6233 3814 6247 3828
rect 6173 3772 6187 3786
rect 6173 3713 6187 3727
rect 6213 3713 6227 3727
rect 6113 3673 6127 3687
rect 6053 3593 6067 3607
rect 6093 3593 6107 3607
rect 5953 3533 5967 3547
rect 5973 3514 5987 3528
rect 6013 3514 6027 3528
rect 6133 3514 6147 3528
rect 5873 3473 5887 3487
rect 5913 3472 5927 3486
rect 5953 3472 5967 3486
rect 5953 3453 5967 3467
rect 5873 3413 5887 3427
rect 5733 3333 5747 3347
rect 5813 3333 5827 3347
rect 5853 3333 5867 3347
rect 5733 3253 5747 3267
rect 5713 3233 5727 3247
rect 5773 3233 5787 3247
rect 5693 3033 5707 3047
rect 5653 2994 5667 3008
rect 5693 2994 5707 3008
rect 5393 2913 5407 2927
rect 5413 2893 5427 2907
rect 5433 2893 5447 2907
rect 5373 2774 5387 2788
rect 5553 2952 5567 2966
rect 5593 2952 5607 2966
rect 5633 2952 5647 2966
rect 5753 3113 5767 3127
rect 5593 2873 5607 2887
rect 5653 2873 5667 2887
rect 5693 2873 5707 2887
rect 5733 2873 5747 2887
rect 5473 2853 5487 2867
rect 5573 2833 5587 2847
rect 5433 2773 5447 2787
rect 5473 2774 5487 2788
rect 5513 2774 5527 2788
rect 5353 2732 5367 2746
rect 5393 2673 5407 2687
rect 5253 2653 5267 2667
rect 5293 2653 5307 2667
rect 5253 2613 5267 2627
rect 5313 2573 5327 2587
rect 5273 2513 5287 2527
rect 5413 2553 5427 2567
rect 5353 2474 5367 2488
rect 5133 2353 5147 2367
rect 5113 2253 5127 2267
rect 5273 2433 5287 2447
rect 5213 2373 5227 2387
rect 5193 2353 5207 2367
rect 5153 2253 5167 2267
rect 5233 2313 5247 2327
rect 5273 2273 5287 2287
rect 5233 2254 5247 2268
rect 5133 2212 5147 2226
rect 5113 2153 5127 2167
rect 5033 2073 5047 2087
rect 5093 2073 5107 2087
rect 5013 1953 5027 1967
rect 4773 1873 4787 1887
rect 4813 1873 4827 1887
rect 4753 1853 4767 1867
rect 4733 1733 4747 1747
rect 4773 1734 4787 1748
rect 4753 1692 4767 1706
rect 4713 1673 4727 1687
rect 4693 1573 4707 1587
rect 4633 1533 4647 1547
rect 4733 1653 4747 1667
rect 4753 1573 4767 1587
rect 4652 1493 4666 1507
rect 4673 1493 4687 1507
rect 4593 1434 4607 1448
rect 4613 1392 4627 1406
rect 4733 1453 4747 1467
rect 4693 1433 4707 1447
rect 4833 1793 4847 1807
rect 4833 1734 4847 1748
rect 4813 1493 4827 1507
rect 4673 1353 4687 1367
rect 4633 1313 4647 1327
rect 4533 1214 4547 1228
rect 4573 1214 4587 1228
rect 4493 1193 4507 1207
rect 4373 1132 4387 1146
rect 4293 1053 4307 1067
rect 4353 1053 4367 1067
rect 4413 1073 4427 1087
rect 4373 1033 4387 1047
rect 4333 973 4347 987
rect 4213 914 4227 928
rect 4312 914 4326 928
rect 4333 913 4347 927
rect 4593 1093 4607 1107
rect 4773 1373 4787 1387
rect 4893 1873 4907 1887
rect 5013 1932 5027 1946
rect 4953 1912 4967 1926
rect 4913 1753 4927 1767
rect 4933 1692 4947 1706
rect 4873 1673 4887 1687
rect 4853 1553 4867 1567
rect 4973 1692 4987 1706
rect 4953 1613 4967 1627
rect 4973 1553 4987 1567
rect 4953 1453 4967 1467
rect 4913 1434 4927 1448
rect 4833 1353 4847 1367
rect 4653 1293 4667 1307
rect 4693 1293 4707 1307
rect 4693 1253 4707 1267
rect 4973 1353 4987 1367
rect 4953 1273 4967 1287
rect 4893 1233 4907 1247
rect 4733 1214 4747 1228
rect 4813 1214 4827 1228
rect 4873 1214 4887 1228
rect 4913 1214 4927 1228
rect 4653 1172 4667 1186
rect 4713 1172 4727 1186
rect 4753 1132 4767 1146
rect 4473 1013 4487 1027
rect 4633 1013 4647 1027
rect 4473 953 4487 967
rect 4633 953 4647 967
rect 4473 914 4487 928
rect 4593 914 4607 928
rect 4693 933 4707 947
rect 4193 853 4207 867
rect 4193 832 4207 846
rect 4153 813 4167 827
rect 4153 773 4167 787
rect 4113 753 4127 767
rect 4053 713 4067 727
rect 3973 693 3987 707
rect 4033 694 4047 708
rect 4153 693 4167 707
rect 4253 813 4267 827
rect 4233 773 4247 787
rect 4273 753 4287 767
rect 4233 694 4247 708
rect 4013 652 4027 666
rect 3853 593 3867 607
rect 3933 593 3947 607
rect 3973 593 3987 607
rect 4013 553 4027 567
rect 3833 533 3847 547
rect 3953 533 3967 547
rect 3513 373 3527 387
rect 3313 353 3327 367
rect 3433 352 3447 366
rect 3573 352 3587 366
rect 3613 352 3627 366
rect 3253 333 3267 347
rect 3233 313 3247 327
rect 3813 394 3827 408
rect 3873 473 3887 487
rect 3853 433 3867 447
rect 3753 352 3767 366
rect 3833 352 3847 366
rect 3673 313 3687 327
rect 3613 293 3627 307
rect 3313 273 3327 287
rect 3673 273 3687 287
rect 3833 273 3847 287
rect 3233 213 3247 227
rect 3033 132 3047 146
rect 3073 113 3087 127
rect 3293 173 3307 187
rect 3572 253 3586 267
rect 3593 253 3607 267
rect 3573 193 3587 207
rect 3353 174 3367 188
rect 3393 174 3407 188
rect 3553 174 3567 188
rect 3653 193 3667 207
rect 3753 193 3767 207
rect 3633 173 3647 187
rect 3293 113 3307 127
rect 3413 132 3427 146
rect 3573 132 3587 146
rect 3713 174 3727 188
rect 3913 394 3927 408
rect 3993 373 4007 387
rect 3913 333 3927 347
rect 3873 273 3887 287
rect 3853 253 3867 267
rect 3873 193 3887 207
rect 3933 233 3947 247
rect 4173 652 4187 666
rect 4213 652 4227 666
rect 4253 613 4267 627
rect 4233 592 4247 606
rect 4153 513 4167 527
rect 4093 493 4107 507
rect 4053 433 4067 447
rect 4613 872 4627 886
rect 4713 914 4727 928
rect 4953 1213 4967 1227
rect 4893 1172 4907 1186
rect 4853 1093 4867 1107
rect 4813 1053 4827 1067
rect 4793 914 4807 928
rect 4853 913 4867 927
rect 4713 873 4727 887
rect 4773 872 4787 886
rect 4453 833 4467 847
rect 4653 833 4667 847
rect 4693 833 4707 847
rect 4733 833 4747 847
rect 4373 753 4387 767
rect 4573 753 4587 767
rect 4493 733 4507 747
rect 4293 692 4307 706
rect 4413 694 4427 708
rect 4452 693 4466 707
rect 4473 693 4487 707
rect 4233 394 4247 408
rect 4313 593 4327 607
rect 4393 652 4407 666
rect 4353 633 4367 647
rect 4373 613 4387 627
rect 4353 593 4367 607
rect 4393 593 4407 607
rect 4373 573 4387 587
rect 4333 513 4347 527
rect 4013 352 4027 366
rect 4073 352 4087 366
rect 4213 352 4227 366
rect 4453 473 4467 487
rect 4413 433 4427 447
rect 4533 694 4547 708
rect 4493 652 4507 666
rect 4553 652 4567 666
rect 4593 633 4607 647
rect 4693 694 4707 708
rect 4793 694 4807 708
rect 4673 652 4687 666
rect 4713 652 4727 666
rect 4573 613 4587 627
rect 4373 394 4387 408
rect 4353 352 4367 366
rect 4393 352 4407 366
rect 4293 333 4307 347
rect 4333 333 4347 347
rect 4113 313 4127 327
rect 4133 273 4147 287
rect 4113 253 4127 267
rect 4093 213 4107 227
rect 3993 193 4007 207
rect 4073 193 4087 207
rect 4033 174 4047 188
rect 4233 233 4247 247
rect 4133 193 4147 207
rect 4113 173 4127 187
rect 4153 173 4167 187
rect 4193 174 4207 188
rect 4133 153 4147 167
rect 3653 132 3667 146
rect 3693 132 3707 146
rect 3733 132 3747 146
rect 3833 132 3847 146
rect 3893 132 3907 146
rect 3573 113 3587 127
rect 3633 113 3647 127
rect 4093 132 4107 146
rect 3933 93 3947 107
rect 4053 93 4067 107
rect 3213 73 3227 87
rect 3373 73 3387 87
rect 3533 73 3547 87
rect 4213 132 4227 146
rect 4392 273 4406 287
rect 4413 273 4427 287
rect 4393 213 4407 227
rect 4313 193 4327 207
rect 4353 193 4367 207
rect 4373 132 4387 146
rect 4493 394 4507 408
rect 4533 394 4547 408
rect 4473 273 4487 287
rect 4433 253 4447 267
rect 4493 253 4507 267
rect 4433 213 4447 227
rect 4413 132 4427 146
rect 4453 173 4467 187
rect 4553 213 4567 227
rect 4533 174 4547 188
rect 4473 132 4487 146
rect 4393 113 4407 127
rect 4313 73 4327 87
rect 3133 33 3147 47
rect 4153 33 4167 47
rect 4753 633 4767 647
rect 4673 593 4687 607
rect 4713 593 4727 607
rect 4853 872 4867 886
rect 4893 1113 4907 1127
rect 5013 1873 5027 1887
rect 5073 2033 5087 2047
rect 5133 1873 5147 1887
rect 5113 1853 5127 1867
rect 5093 1753 5107 1767
rect 5033 1692 5047 1706
rect 5073 1653 5087 1667
rect 5073 1613 5087 1627
rect 5073 1453 5087 1467
rect 5013 1434 5027 1448
rect 5093 1433 5107 1447
rect 5013 1333 5027 1347
rect 4993 1213 5007 1227
rect 5053 1353 5067 1367
rect 5033 1253 5047 1267
rect 5173 2212 5187 2226
rect 5213 2173 5227 2187
rect 5273 2133 5287 2147
rect 5273 2093 5287 2107
rect 5253 1973 5267 1987
rect 5173 1953 5187 1967
rect 5213 1954 5227 1968
rect 5153 1853 5167 1867
rect 5133 1833 5147 1847
rect 5233 1912 5247 1926
rect 5173 1773 5187 1787
rect 5253 1773 5267 1787
rect 5193 1734 5207 1748
rect 5173 1692 5187 1706
rect 5213 1692 5227 1706
rect 5253 1692 5267 1706
rect 5133 1633 5147 1647
rect 5333 2432 5347 2446
rect 5373 2353 5387 2367
rect 5573 2732 5587 2746
rect 5533 2693 5547 2707
rect 5613 2774 5627 2788
rect 5693 2774 5707 2788
rect 5673 2732 5687 2746
rect 5713 2732 5727 2746
rect 5613 2693 5627 2707
rect 5593 2593 5607 2607
rect 5473 2573 5487 2587
rect 5513 2573 5527 2587
rect 5473 2513 5487 2527
rect 5453 2474 5467 2488
rect 5573 2553 5587 2567
rect 5433 2432 5447 2446
rect 5493 2432 5507 2446
rect 5533 2413 5547 2427
rect 5673 2474 5687 2488
rect 5733 2473 5747 2487
rect 5613 2433 5627 2447
rect 5613 2373 5627 2387
rect 5693 2432 5707 2446
rect 5853 3253 5867 3267
rect 5833 3193 5847 3207
rect 5813 3153 5827 3167
rect 5833 2994 5847 3008
rect 5773 2853 5787 2867
rect 5933 3393 5947 3407
rect 5893 3373 5907 3387
rect 6013 3413 6027 3427
rect 6053 3413 6067 3427
rect 5973 3294 5987 3308
rect 6033 3333 6047 3347
rect 6013 3273 6027 3287
rect 5913 3252 5927 3266
rect 5893 3233 5907 3247
rect 5873 2953 5887 2967
rect 5913 3193 5927 3207
rect 5953 3173 5967 3187
rect 5973 3133 5987 3147
rect 5953 3113 5967 3127
rect 5913 3073 5927 3087
rect 5933 3033 5947 3047
rect 5913 2993 5927 3007
rect 6013 3073 6027 3087
rect 5973 2994 5987 3008
rect 5913 2953 5927 2967
rect 6113 3472 6127 3486
rect 6193 3613 6207 3627
rect 6113 3373 6127 3387
rect 6073 3333 6087 3347
rect 6073 3294 6087 3308
rect 6173 3472 6187 3486
rect 6173 3393 6187 3407
rect 6173 3353 6187 3367
rect 6173 3313 6187 3327
rect 6053 3253 6067 3267
rect 6133 3252 6147 3266
rect 6173 3253 6187 3267
rect 6093 3233 6107 3247
rect 6053 3133 6067 3147
rect 6133 3133 6147 3147
rect 6053 3073 6067 3087
rect 5833 2853 5847 2867
rect 5893 2853 5907 2867
rect 5793 2833 5807 2847
rect 5873 2774 5887 2788
rect 5773 2732 5787 2746
rect 5953 2933 5967 2947
rect 5853 2693 5867 2707
rect 5793 2593 5807 2607
rect 5773 2533 5787 2547
rect 5773 2493 5787 2507
rect 5833 2553 5847 2567
rect 5813 2493 5827 2507
rect 5773 2413 5787 2427
rect 5753 2393 5767 2407
rect 5653 2353 5667 2367
rect 5573 2313 5587 2327
rect 5733 2313 5747 2327
rect 5413 2293 5427 2307
rect 5353 2273 5367 2287
rect 5393 2254 5407 2268
rect 5473 2253 5487 2267
rect 5533 2254 5547 2268
rect 5613 2254 5627 2268
rect 5373 2212 5387 2226
rect 5333 2053 5347 2067
rect 5453 2053 5467 2067
rect 5373 1993 5387 2007
rect 5413 1954 5427 1968
rect 5513 2212 5527 2226
rect 5513 2173 5527 2187
rect 5593 2213 5607 2227
rect 5513 2133 5527 2147
rect 5553 2133 5567 2147
rect 5473 2033 5487 2047
rect 5573 2093 5587 2107
rect 5693 2254 5707 2268
rect 5813 2353 5827 2367
rect 5813 2332 5827 2346
rect 5773 2293 5787 2307
rect 5873 2373 5887 2387
rect 5913 2713 5927 2727
rect 5953 2873 5967 2887
rect 6033 2952 6047 2966
rect 6133 3033 6147 3047
rect 6093 2994 6107 3008
rect 6113 2952 6127 2966
rect 6153 2952 6167 2966
rect 6213 3514 6227 3528
rect 6353 3993 6367 4007
rect 6333 3893 6347 3907
rect 6393 3992 6407 4006
rect 6453 4253 6467 4267
rect 6433 4193 6447 4207
rect 6473 4213 6487 4227
rect 6593 5413 6607 5427
rect 6693 5673 6707 5687
rect 6733 5593 6747 5607
rect 6733 5553 6747 5567
rect 6713 5513 6727 5527
rect 6653 5433 6667 5447
rect 6633 5413 6647 5427
rect 6633 5374 6647 5388
rect 6733 5473 6747 5487
rect 6713 5373 6727 5387
rect 6613 5333 6627 5347
rect 6593 5133 6607 5147
rect 6713 5333 6727 5347
rect 6693 5313 6707 5327
rect 6733 5313 6747 5327
rect 6653 5273 6667 5287
rect 6713 5133 6727 5147
rect 6613 5113 6627 5127
rect 6653 5113 6667 5127
rect 6613 5074 6627 5088
rect 6693 5033 6707 5047
rect 6673 4993 6687 5007
rect 6673 4953 6687 4967
rect 6633 4893 6647 4907
rect 6653 4873 6667 4887
rect 6613 4854 6627 4868
rect 6553 4812 6567 4826
rect 6533 4713 6547 4727
rect 6632 4812 6646 4826
rect 6653 4813 6667 4827
rect 6593 4793 6607 4807
rect 6633 4753 6647 4767
rect 6593 4733 6607 4747
rect 6533 4673 6547 4687
rect 6573 4673 6587 4687
rect 6593 4613 6607 4627
rect 6532 4553 6546 4567
rect 6553 4554 6567 4568
rect 6573 4512 6587 4526
rect 6573 4491 6587 4505
rect 6613 4493 6627 4507
rect 6513 4453 6527 4467
rect 6513 4393 6527 4407
rect 6553 4373 6567 4387
rect 6513 4333 6527 4347
rect 6593 4433 6607 4447
rect 6633 4473 6647 4487
rect 6613 4393 6627 4407
rect 6573 4353 6587 4367
rect 6593 4334 6607 4348
rect 6533 4292 6547 4306
rect 6553 4273 6567 4287
rect 6493 4193 6507 4207
rect 6453 4153 6467 4167
rect 6473 4133 6487 4147
rect 6533 4133 6547 4147
rect 6533 4093 6547 4107
rect 6513 4034 6527 4048
rect 6453 3992 6467 4006
rect 6473 3973 6487 3987
rect 6433 3953 6447 3967
rect 6453 3933 6467 3947
rect 6413 3893 6427 3907
rect 6393 3833 6407 3847
rect 6313 3813 6327 3827
rect 6353 3814 6367 3828
rect 6313 3753 6327 3767
rect 6313 3673 6327 3687
rect 6273 3613 6287 3627
rect 6293 3573 6307 3587
rect 6273 3553 6287 3567
rect 6293 3513 6307 3527
rect 6293 3473 6307 3487
rect 6253 3353 6267 3367
rect 6213 3293 6227 3307
rect 6353 3673 6367 3687
rect 6413 3772 6427 3786
rect 6413 3753 6427 3767
rect 6453 3733 6467 3747
rect 6453 3712 6467 3726
rect 6373 3653 6387 3667
rect 6393 3553 6407 3567
rect 6433 3553 6447 3567
rect 6353 3513 6367 3527
rect 6453 3513 6467 3527
rect 6373 3453 6387 3467
rect 6333 3413 6347 3427
rect 6333 3373 6347 3387
rect 6293 3333 6307 3347
rect 6273 3313 6287 3327
rect 6353 3313 6367 3327
rect 6273 3252 6287 3266
rect 6333 3253 6347 3267
rect 6273 3193 6287 3207
rect 6233 3173 6247 3187
rect 6693 4813 6707 4827
rect 6693 4693 6707 4707
rect 6753 4593 6767 4607
rect 6733 4473 6747 4487
rect 6733 4433 6747 4447
rect 6713 4353 6727 4367
rect 6693 4334 6707 4348
rect 6773 4333 6787 4347
rect 6573 4193 6587 4207
rect 6633 4253 6647 4267
rect 6573 4172 6587 4186
rect 6613 4173 6627 4187
rect 6553 3973 6567 3987
rect 6713 4292 6727 4306
rect 6673 4233 6687 4247
rect 6653 4153 6667 4167
rect 6613 4073 6627 4087
rect 6613 4034 6627 4048
rect 6733 4273 6747 4287
rect 6713 4233 6727 4247
rect 6693 4073 6707 4087
rect 6693 4033 6707 4047
rect 6573 3933 6587 3947
rect 6593 3913 6607 3927
rect 6513 3873 6527 3887
rect 6493 3833 6507 3847
rect 6553 3833 6567 3847
rect 6533 3772 6547 3786
rect 6653 3973 6667 3987
rect 6633 3893 6647 3907
rect 6493 3733 6507 3747
rect 6473 3453 6487 3467
rect 6413 3333 6427 3347
rect 6433 3333 6447 3347
rect 6393 3313 6407 3327
rect 6373 3253 6387 3267
rect 6353 3073 6367 3087
rect 6253 3033 6267 3047
rect 6313 3033 6327 3047
rect 6213 2953 6227 2967
rect 6253 2993 6267 3007
rect 6313 2994 6327 3008
rect 6453 3252 6467 3266
rect 6413 3153 6427 3167
rect 6613 3693 6627 3707
rect 6593 3673 6607 3687
rect 6553 3653 6567 3667
rect 6513 3533 6527 3547
rect 6453 3133 6467 3147
rect 6473 3113 6487 3127
rect 6393 3053 6407 3067
rect 6433 3053 6447 3067
rect 6233 2933 6247 2947
rect 6153 2913 6167 2927
rect 6192 2913 6206 2927
rect 6213 2913 6227 2927
rect 6073 2893 6087 2907
rect 6133 2893 6147 2907
rect 6053 2813 6067 2827
rect 5993 2793 6007 2807
rect 6033 2774 6047 2788
rect 6133 2853 6147 2867
rect 6093 2813 6107 2827
rect 5973 2733 5987 2747
rect 5953 2713 5967 2727
rect 5933 2633 5947 2647
rect 6273 2933 6287 2947
rect 6253 2833 6267 2847
rect 6153 2793 6167 2807
rect 6113 2773 6127 2787
rect 6193 2793 6207 2807
rect 6053 2713 6067 2727
rect 6013 2673 6027 2687
rect 6033 2633 6047 2647
rect 5973 2493 5987 2507
rect 5993 2474 6007 2488
rect 6093 2732 6107 2746
rect 6093 2673 6107 2687
rect 6253 2753 6267 2767
rect 6173 2732 6187 2746
rect 6333 2952 6347 2966
rect 6373 2953 6387 2967
rect 6573 3633 6587 3647
rect 6613 3553 6627 3567
rect 6573 3533 6587 3547
rect 6573 3472 6587 3486
rect 6693 3993 6707 4007
rect 6693 3913 6707 3927
rect 6693 3873 6707 3887
rect 6773 4293 6787 4307
rect 6753 4253 6767 4267
rect 6733 4193 6747 4207
rect 6733 3853 6747 3867
rect 6753 3813 6767 3827
rect 6653 3772 6667 3786
rect 6713 3772 6727 3786
rect 6753 3773 6767 3787
rect 6733 3693 6747 3707
rect 6693 3553 6707 3567
rect 6653 3513 6667 3527
rect 6732 3514 6746 3528
rect 6773 3633 6787 3647
rect 6773 3553 6787 3567
rect 6753 3513 6767 3527
rect 6633 3473 6647 3487
rect 6653 3453 6667 3467
rect 6713 3472 6727 3486
rect 6693 3453 6707 3467
rect 6732 3453 6746 3467
rect 6673 3373 6687 3387
rect 6693 3353 6707 3367
rect 6613 3333 6627 3347
rect 6673 3333 6687 3347
rect 6593 3313 6607 3327
rect 6633 3294 6647 3308
rect 6533 3273 6547 3287
rect 6513 3073 6527 3087
rect 6533 3053 6547 3067
rect 6513 3033 6527 3047
rect 6533 3013 6547 3027
rect 6473 2993 6487 3007
rect 6513 2994 6527 3008
rect 6293 2893 6307 2907
rect 6353 2893 6367 2907
rect 6393 2893 6407 2907
rect 6233 2713 6247 2727
rect 6273 2713 6287 2727
rect 6133 2693 6147 2707
rect 6073 2573 6087 2587
rect 6053 2553 6067 2567
rect 6053 2513 6067 2527
rect 5913 2413 5927 2427
rect 5893 2333 5907 2347
rect 5833 2293 5847 2307
rect 5633 2193 5647 2207
rect 5693 2193 5707 2207
rect 5633 2073 5647 2087
rect 5613 2053 5627 2067
rect 5593 1993 5607 2007
rect 5573 1954 5587 1968
rect 5533 1912 5547 1926
rect 5393 1893 5407 1907
rect 5453 1893 5467 1907
rect 5353 1873 5367 1887
rect 5333 1853 5347 1867
rect 5453 1773 5467 1787
rect 5393 1733 5407 1747
rect 5713 1912 5727 1926
rect 5813 2273 5827 2287
rect 6013 2432 6027 2446
rect 6113 2593 6127 2607
rect 6213 2533 6227 2547
rect 6173 2513 6187 2527
rect 6073 2393 6087 2407
rect 5993 2373 6007 2387
rect 6053 2373 6067 2387
rect 5913 2254 5927 2268
rect 5813 2212 5827 2226
rect 5853 2212 5867 2226
rect 5893 2193 5907 2207
rect 5833 2033 5847 2047
rect 5873 1993 5887 2007
rect 5833 1954 5847 1968
rect 5553 1733 5567 1747
rect 5593 1734 5607 1748
rect 5633 1734 5647 1748
rect 5353 1692 5367 1706
rect 5533 1713 5547 1727
rect 5473 1673 5487 1687
rect 5533 1653 5547 1667
rect 5293 1613 5307 1627
rect 5393 1613 5407 1627
rect 5353 1593 5367 1607
rect 5313 1493 5327 1507
rect 5193 1434 5207 1448
rect 5433 1553 5447 1567
rect 5413 1473 5427 1487
rect 5153 1373 5167 1387
rect 5133 1353 5147 1367
rect 5113 1333 5127 1347
rect 5133 1253 5147 1267
rect 5073 1172 5087 1186
rect 5053 1153 5067 1167
rect 4973 1093 4987 1107
rect 5033 1093 5047 1107
rect 5093 1053 5107 1067
rect 5093 1013 5107 1027
rect 5053 993 5067 1007
rect 4933 914 4947 928
rect 4893 872 4907 886
rect 4953 872 4967 886
rect 4953 813 4967 827
rect 4873 793 4887 807
rect 4913 793 4927 807
rect 4873 694 4887 708
rect 4833 653 4847 667
rect 4973 713 4987 727
rect 4813 633 4827 647
rect 4793 573 4807 587
rect 4653 553 4667 567
rect 4813 533 4827 547
rect 4893 652 4907 666
rect 4953 652 4967 666
rect 4853 633 4867 647
rect 4973 613 4987 627
rect 4833 453 4847 467
rect 4713 433 4727 447
rect 4713 394 4727 408
rect 4753 394 4767 408
rect 5013 913 5027 927
rect 5053 914 5067 928
rect 5213 1313 5227 1327
rect 5273 1313 5287 1327
rect 5153 1213 5167 1227
rect 5213 1214 5227 1228
rect 5193 1172 5207 1186
rect 5253 1172 5267 1186
rect 5293 1214 5307 1228
rect 5373 1373 5387 1387
rect 5373 1333 5387 1347
rect 5273 1113 5287 1127
rect 5273 1053 5287 1067
rect 5133 933 5147 947
rect 5013 872 5027 886
rect 5033 713 5047 727
rect 5173 753 5187 767
rect 5113 733 5127 747
rect 5233 872 5247 886
rect 5213 694 5227 708
rect 5353 1172 5367 1186
rect 5333 1093 5347 1107
rect 5313 1053 5327 1067
rect 5313 1013 5327 1027
rect 5253 693 5267 707
rect 5293 693 5307 707
rect 5393 1113 5407 1127
rect 5353 1073 5367 1087
rect 5393 933 5407 947
rect 5613 1673 5627 1687
rect 5653 1653 5667 1667
rect 5613 1533 5627 1547
rect 5453 1513 5467 1527
rect 5553 1513 5567 1527
rect 5593 1493 5607 1507
rect 5553 1434 5567 1448
rect 5453 1353 5467 1367
rect 5493 1353 5507 1367
rect 5593 1293 5607 1307
rect 5553 1253 5567 1267
rect 5533 1233 5547 1247
rect 5533 1153 5547 1167
rect 5493 1133 5507 1147
rect 6113 2432 6127 2446
rect 6193 2433 6207 2447
rect 6153 2393 6167 2407
rect 6113 2333 6127 2347
rect 6013 2293 6027 2307
rect 5973 2253 5987 2267
rect 6053 2254 6067 2268
rect 6093 2293 6107 2307
rect 5953 2193 5967 2207
rect 6033 2173 6047 2187
rect 5973 2133 5987 2147
rect 5973 1993 5987 2007
rect 6033 1993 6047 2007
rect 5953 1953 5967 1967
rect 5953 1912 5967 1926
rect 6013 1912 6027 1926
rect 5933 1873 5947 1887
rect 6013 1873 6027 1887
rect 5853 1833 5867 1847
rect 5853 1773 5867 1787
rect 5773 1734 5787 1748
rect 5813 1734 5827 1748
rect 5713 1553 5727 1567
rect 5693 1473 5707 1487
rect 5673 1434 5687 1448
rect 5673 1333 5687 1347
rect 5673 1233 5687 1247
rect 5713 1214 5727 1228
rect 5753 1673 5767 1687
rect 5833 1693 5847 1707
rect 5793 1434 5807 1448
rect 5853 1553 5867 1567
rect 5813 1392 5827 1406
rect 5773 1353 5787 1367
rect 5613 1172 5627 1186
rect 5693 1172 5707 1186
rect 5653 1133 5667 1147
rect 5593 1113 5607 1127
rect 5973 1813 5987 1827
rect 5973 1773 5987 1787
rect 5933 1734 5947 1748
rect 5913 1673 5927 1687
rect 5893 1613 5907 1627
rect 5953 1613 5967 1627
rect 6153 2273 6167 2287
rect 6213 2413 6227 2427
rect 6193 2253 6207 2267
rect 6113 2033 6127 2047
rect 6173 2212 6187 2226
rect 6213 2213 6227 2227
rect 6333 2732 6347 2746
rect 6393 2733 6407 2747
rect 6353 2693 6367 2707
rect 6333 2573 6347 2587
rect 6293 2513 6307 2527
rect 6293 2474 6307 2488
rect 6313 2413 6327 2427
rect 6313 2353 6327 2367
rect 6293 2333 6307 2347
rect 6433 2933 6447 2947
rect 6573 3252 6587 3266
rect 6553 2933 6567 2947
rect 6493 2913 6507 2927
rect 6533 2913 6547 2927
rect 6453 2893 6467 2907
rect 6533 2892 6547 2906
rect 6473 2853 6487 2867
rect 6493 2813 6507 2827
rect 6473 2793 6487 2807
rect 6493 2774 6507 2788
rect 6433 2733 6447 2747
rect 6473 2732 6487 2746
rect 6433 2673 6447 2687
rect 6413 2653 6427 2667
rect 6413 2593 6427 2607
rect 6473 2513 6487 2527
rect 6613 3153 6627 3167
rect 6673 3153 6687 3167
rect 6653 3033 6667 3047
rect 6613 2994 6627 3008
rect 6693 2993 6707 3007
rect 6593 2953 6607 2967
rect 6733 3373 6747 3387
rect 6473 2474 6487 2488
rect 6433 2433 6447 2447
rect 6413 2413 6427 2427
rect 6393 2353 6407 2367
rect 6373 2333 6387 2347
rect 6313 2293 6327 2307
rect 6353 2313 6367 2327
rect 6433 2293 6447 2307
rect 6493 2413 6507 2427
rect 6533 2433 6547 2447
rect 6333 2253 6347 2267
rect 6253 2213 6267 2227
rect 6373 2253 6387 2267
rect 6413 2254 6427 2268
rect 6453 2253 6467 2267
rect 6493 2253 6507 2267
rect 6233 2153 6247 2167
rect 6213 2133 6227 2147
rect 6133 2013 6147 2027
rect 6113 1954 6127 1968
rect 6173 1954 6187 1968
rect 6213 1954 6227 1968
rect 6093 1793 6107 1807
rect 6013 1593 6027 1607
rect 6093 1734 6107 1748
rect 6193 1912 6207 1926
rect 6313 2212 6327 2226
rect 6353 2212 6367 2226
rect 6293 2173 6307 2187
rect 6273 2153 6287 2167
rect 6273 1913 6287 1927
rect 6153 1833 6167 1847
rect 6193 1793 6207 1807
rect 6173 1733 6187 1747
rect 6113 1673 6127 1687
rect 6073 1613 6087 1627
rect 6073 1553 6087 1567
rect 6033 1533 6047 1547
rect 5913 1493 5927 1507
rect 5973 1493 5987 1507
rect 6053 1473 6067 1487
rect 6013 1434 6027 1448
rect 5893 1413 5907 1427
rect 5913 1353 5927 1367
rect 5833 1293 5847 1307
rect 5873 1293 5887 1307
rect 5773 1253 5787 1267
rect 5753 1133 5767 1147
rect 5733 1093 5747 1107
rect 5733 1013 5747 1027
rect 5613 973 5627 987
rect 5453 913 5467 927
rect 5493 914 5507 928
rect 5413 872 5427 886
rect 5493 873 5507 887
rect 5693 914 5707 928
rect 5573 872 5587 886
rect 5613 872 5627 886
rect 5593 833 5607 847
rect 5513 813 5527 827
rect 5333 773 5347 787
rect 5533 773 5547 787
rect 5353 694 5367 708
rect 5413 694 5427 708
rect 5493 694 5507 708
rect 5113 652 5127 666
rect 5153 652 5167 666
rect 5233 652 5247 666
rect 5333 652 5347 666
rect 5713 872 5727 886
rect 5733 853 5747 867
rect 5673 813 5687 827
rect 5693 773 5707 787
rect 5653 694 5667 708
rect 5413 633 5427 647
rect 5473 633 5487 647
rect 5593 652 5607 666
rect 5633 652 5647 666
rect 5673 652 5687 666
rect 5253 613 5267 627
rect 5233 593 5247 607
rect 5093 573 5107 587
rect 5393 593 5407 607
rect 5373 553 5387 567
rect 5513 612 5527 626
rect 5433 553 5447 567
rect 5273 513 5287 527
rect 5413 513 5427 527
rect 5173 453 5187 467
rect 4993 394 5007 408
rect 4833 373 4847 387
rect 4673 333 4687 347
rect 4593 213 4607 227
rect 4613 173 4627 187
rect 4713 233 4727 247
rect 4773 233 4787 247
rect 4733 173 4747 187
rect 4653 132 4667 146
rect 4693 132 4707 146
rect 5213 394 5227 408
rect 4993 352 5007 366
rect 5073 352 5087 366
rect 4833 213 4847 227
rect 4893 213 4907 227
rect 5133 313 5147 327
rect 4993 213 5007 227
rect 4913 174 4927 188
rect 4953 174 4967 188
rect 5293 394 5307 408
rect 5333 394 5347 408
rect 5393 352 5407 366
rect 5353 333 5367 347
rect 5293 313 5307 327
rect 5633 413 5647 427
rect 5513 394 5527 408
rect 5633 394 5647 408
rect 5673 394 5687 408
rect 5433 333 5447 347
rect 5313 293 5327 307
rect 5273 273 5287 287
rect 5193 253 5207 267
rect 5213 213 5227 227
rect 4813 132 4827 146
rect 4893 132 4907 146
rect 5013 132 5027 146
rect 5153 132 5167 146
rect 4973 113 4987 127
rect 4613 93 4627 107
rect 4773 93 4787 107
rect 5333 273 5347 287
rect 5393 253 5407 267
rect 5373 213 5387 227
rect 5613 352 5627 366
rect 5692 353 5706 367
rect 5713 353 5727 367
rect 5653 333 5667 347
rect 5693 313 5707 327
rect 5873 1233 5887 1247
rect 5793 1172 5807 1186
rect 5793 953 5807 967
rect 5793 873 5807 887
rect 5933 1293 5947 1307
rect 5913 993 5927 1007
rect 5873 914 5887 928
rect 5993 1392 6007 1406
rect 6053 1392 6067 1406
rect 6433 2212 6447 2226
rect 6513 2213 6527 2227
rect 6473 2073 6487 2087
rect 6433 2033 6447 2047
rect 6413 2013 6427 2027
rect 6333 1993 6347 2007
rect 6373 1993 6387 2007
rect 6433 1993 6447 2007
rect 6413 1973 6427 1987
rect 6373 1954 6387 1968
rect 6313 1912 6327 1926
rect 6313 1833 6327 1847
rect 6293 1753 6307 1767
rect 6333 1753 6347 1767
rect 6253 1734 6267 1748
rect 6273 1692 6287 1706
rect 6273 1593 6287 1607
rect 6233 1513 6247 1527
rect 6193 1493 6207 1507
rect 6093 1473 6107 1487
rect 6173 1473 6187 1487
rect 6233 1473 6247 1487
rect 6153 1434 6167 1448
rect 6193 1434 6207 1448
rect 6093 1373 6107 1387
rect 6073 1333 6087 1347
rect 6173 1373 6187 1387
rect 6153 1333 6167 1347
rect 6073 1273 6087 1287
rect 6133 1273 6147 1287
rect 6013 1253 6027 1267
rect 5972 1233 5986 1247
rect 5993 1233 6007 1247
rect 6053 1213 6067 1227
rect 5973 1172 5987 1186
rect 6033 1173 6047 1187
rect 6013 1153 6027 1167
rect 5953 1093 5967 1107
rect 5933 914 5947 928
rect 5813 853 5827 867
rect 5893 872 5907 886
rect 5973 993 5987 1007
rect 6113 1214 6127 1228
rect 6193 1253 6207 1267
rect 6073 1172 6087 1186
rect 6133 1172 6147 1186
rect 6253 1434 6267 1448
rect 6573 2853 6587 2867
rect 6653 2933 6667 2947
rect 6673 2893 6687 2907
rect 6633 2853 6647 2867
rect 6613 2833 6627 2847
rect 6593 2813 6607 2827
rect 6713 2933 6727 2947
rect 6613 2732 6627 2746
rect 6673 2733 6687 2747
rect 6653 2693 6667 2707
rect 6633 2673 6647 2687
rect 6653 2553 6667 2567
rect 6653 2532 6667 2546
rect 6633 2493 6647 2507
rect 6673 2473 6687 2487
rect 6573 2333 6587 2347
rect 6673 2433 6687 2447
rect 6633 2413 6647 2427
rect 6613 2313 6627 2327
rect 6653 2293 6667 2307
rect 6633 2212 6647 2226
rect 6573 2133 6587 2147
rect 6553 1972 6567 1986
rect 6493 1954 6507 1968
rect 6513 1912 6527 1926
rect 6553 1893 6567 1907
rect 6553 1872 6567 1886
rect 6453 1853 6467 1867
rect 6513 1853 6527 1867
rect 6373 1833 6387 1847
rect 6433 1833 6447 1847
rect 6433 1793 6447 1807
rect 6393 1753 6407 1767
rect 6473 1734 6487 1748
rect 6373 1692 6387 1706
rect 6373 1593 6387 1607
rect 6353 1553 6367 1567
rect 6333 1473 6347 1487
rect 6453 1692 6467 1706
rect 6533 1753 6547 1767
rect 6613 2013 6627 2027
rect 6653 2073 6667 2087
rect 6713 2693 6727 2707
rect 6713 2653 6727 2667
rect 6693 2413 6707 2427
rect 6693 2392 6707 2406
rect 6673 2013 6687 2027
rect 6633 1973 6647 1987
rect 6633 1912 6647 1926
rect 6653 1893 6667 1907
rect 6633 1833 6647 1847
rect 6593 1793 6607 1807
rect 6573 1753 6587 1767
rect 6553 1733 6567 1747
rect 6613 1773 6627 1787
rect 6673 1873 6687 1887
rect 6673 1793 6687 1807
rect 6553 1693 6567 1707
rect 6533 1593 6547 1607
rect 6513 1573 6527 1587
rect 6433 1553 6447 1567
rect 6493 1513 6507 1527
rect 6373 1434 6387 1448
rect 6273 1333 6287 1347
rect 6273 1293 6287 1307
rect 6253 1273 6267 1287
rect 6313 1392 6327 1406
rect 6533 1493 6547 1507
rect 6433 1432 6447 1446
rect 6493 1434 6507 1448
rect 6613 1692 6627 1706
rect 6593 1613 6607 1627
rect 6673 1613 6687 1627
rect 6573 1593 6587 1607
rect 6353 1333 6367 1347
rect 6293 1253 6307 1267
rect 6373 1253 6387 1267
rect 6253 1233 6267 1247
rect 6313 1214 6327 1228
rect 6053 1073 6067 1087
rect 6073 1053 6087 1067
rect 5993 973 6007 987
rect 6033 973 6047 987
rect 5793 773 5807 787
rect 5853 773 5867 787
rect 5973 872 5987 886
rect 5953 753 5967 767
rect 5833 733 5847 747
rect 5933 733 5947 747
rect 5913 693 5927 707
rect 6033 914 6047 928
rect 6133 914 6147 928
rect 6053 872 6067 886
rect 6093 872 6107 886
rect 5993 694 6007 708
rect 6053 693 6067 707
rect 6233 1153 6247 1167
rect 6333 1172 6347 1186
rect 6313 1153 6327 1167
rect 6293 1073 6307 1087
rect 6193 973 6207 987
rect 6433 1313 6447 1327
rect 6433 1292 6447 1306
rect 6513 1392 6527 1406
rect 6533 1313 6547 1327
rect 6473 1214 6487 1228
rect 6453 1172 6467 1186
rect 6393 1113 6407 1127
rect 6513 1153 6527 1167
rect 6493 1073 6507 1087
rect 6373 1013 6387 1027
rect 6473 1013 6487 1027
rect 6333 953 6347 967
rect 6233 914 6247 928
rect 6313 914 6327 928
rect 6213 872 6227 886
rect 6453 914 6467 928
rect 6133 833 6147 847
rect 6213 753 6227 767
rect 5753 652 5767 666
rect 5813 652 5827 666
rect 5853 613 5867 627
rect 6013 652 6027 666
rect 6173 694 6187 708
rect 6073 652 6087 666
rect 6113 652 6127 666
rect 5973 613 5987 627
rect 5913 453 5927 467
rect 6173 453 6187 467
rect 5853 413 5867 427
rect 5753 394 5767 408
rect 5813 394 5827 408
rect 6013 413 6027 427
rect 5913 394 5927 408
rect 5973 394 5987 408
rect 6133 394 6147 408
rect 5753 333 5767 347
rect 5633 293 5647 307
rect 5733 293 5747 307
rect 5513 273 5527 287
rect 5593 273 5607 287
rect 5493 253 5507 267
rect 5513 213 5527 227
rect 5553 213 5567 227
rect 5473 174 5487 188
rect 5693 253 5707 267
rect 5633 174 5647 188
rect 5273 132 5287 146
rect 5313 132 5327 146
rect 5372 132 5386 146
rect 5393 132 5407 146
rect 5453 132 5467 146
rect 5493 132 5507 146
rect 5553 132 5567 146
rect 5613 132 5627 146
rect 6353 872 6367 886
rect 6313 833 6327 847
rect 6373 693 6387 707
rect 6233 613 6247 627
rect 6333 652 6347 666
rect 6373 652 6387 666
rect 6293 593 6307 607
rect 6313 453 6327 467
rect 6273 394 6287 408
rect 5953 352 5967 366
rect 5993 333 6007 347
rect 5833 313 5847 327
rect 5913 313 5927 327
rect 6073 313 6087 327
rect 5793 293 5807 307
rect 5953 273 5967 287
rect 5773 233 5787 247
rect 5813 233 5827 247
rect 5913 174 5927 188
rect 5993 233 6007 247
rect 6153 352 6167 366
rect 6213 352 6227 366
rect 6293 352 6307 366
rect 6113 273 6127 287
rect 6233 273 6247 287
rect 6093 233 6107 247
rect 6233 233 6247 247
rect 6213 213 6227 227
rect 6253 174 6267 188
rect 6433 694 6447 708
rect 6573 1373 6587 1387
rect 6573 1333 6587 1347
rect 6613 1593 6627 1607
rect 6733 1833 6747 1847
rect 6713 1733 6727 1747
rect 6693 1553 6707 1567
rect 6673 1513 6687 1527
rect 6653 1493 6667 1507
rect 6653 1453 6667 1467
rect 6713 1453 6727 1467
rect 6773 3453 6787 3467
rect 6773 3113 6787 3127
rect 6773 3073 6787 3087
rect 6773 1753 6787 1767
rect 6773 1573 6787 1587
rect 6653 1392 6667 1406
rect 6753 1393 6767 1407
rect 6693 1373 6707 1387
rect 6593 1253 6607 1267
rect 6573 1213 6587 1227
rect 6553 1153 6567 1167
rect 6613 1153 6627 1167
rect 6553 1113 6567 1127
rect 6533 833 6547 847
rect 6673 914 6687 928
rect 6573 872 6587 886
rect 6533 733 6547 747
rect 6473 693 6487 707
rect 6473 652 6487 666
rect 6393 593 6407 607
rect 6393 394 6407 408
rect 6433 394 6447 408
rect 6613 753 6627 767
rect 6673 753 6687 767
rect 6593 733 6607 747
rect 6593 652 6607 666
rect 6553 613 6567 627
rect 6533 394 6547 408
rect 6653 394 6667 408
rect 6453 352 6467 366
rect 6393 333 6407 347
rect 6373 293 6387 307
rect 6553 353 6567 367
rect 6493 253 6507 267
rect 6433 174 6447 188
rect 6633 293 6647 307
rect 6593 233 6607 247
rect 6773 753 6787 767
rect 6613 174 6627 188
rect 6733 174 6747 188
rect 5773 132 5787 146
rect 5813 133 5827 147
rect 5933 132 5947 146
rect 5993 133 6007 147
rect 6032 133 6046 147
rect 6053 132 6067 146
rect 6233 132 6247 146
rect 6333 133 6347 146
rect 6333 132 6347 133
rect 6413 132 6427 146
rect 5993 93 6007 107
rect 6033 93 6047 107
rect 6093 93 6107 107
rect 6633 132 6647 146
rect 5213 33 5227 47
rect 5893 33 5907 47
rect 6453 33 6467 47
rect 6593 33 6607 47
rect 4453 13 4467 27
rect 4573 13 4587 27
<< metal3 >>
rect 2807 6516 2833 6524
rect 3007 6516 3093 6524
rect 547 6496 1273 6504
rect 1287 6496 2333 6504
rect 3707 6496 3973 6504
rect 5587 6496 6133 6504
rect 2707 6476 2853 6484
rect 2907 6476 3193 6484
rect 3447 6476 3513 6484
rect 3536 6476 3944 6484
rect 187 6456 573 6464
rect 587 6456 1393 6464
rect 1407 6456 1473 6464
rect 1527 6456 1733 6464
rect 2747 6456 3264 6464
rect 3256 6444 3264 6456
rect 3536 6464 3544 6476
rect 3287 6456 3544 6464
rect 3936 6464 3944 6476
rect 4167 6476 4893 6484
rect 4947 6476 5213 6484
rect 5727 6476 5893 6484
rect 6627 6476 6693 6484
rect 3936 6456 4433 6464
rect 4927 6456 5453 6464
rect 5467 6456 5913 6464
rect 5967 6456 6493 6464
rect 3256 6436 3753 6444
rect 3767 6436 3913 6444
rect 4487 6436 4613 6444
rect 4627 6436 4793 6444
rect 4807 6436 4893 6444
rect 5107 6436 5233 6444
rect 5287 6436 5393 6444
rect 5707 6436 5793 6444
rect 6087 6436 6173 6444
rect 127 6417 213 6425
rect 287 6416 373 6424
rect 447 6416 533 6424
rect 627 6416 733 6424
rect 747 6416 793 6424
rect 907 6416 924 6424
rect 387 6375 413 6383
rect 467 6376 553 6384
rect 767 6376 873 6384
rect 916 6384 924 6416
rect 967 6416 1033 6424
rect 1047 6416 1153 6424
rect 1347 6416 1433 6424
rect 1447 6416 1573 6424
rect 1627 6417 1673 6425
rect 1787 6417 1833 6425
rect 1847 6416 1913 6424
rect 1967 6416 2033 6424
rect 2147 6416 2233 6424
rect 2287 6416 2344 6424
rect 2096 6404 2104 6414
rect 2027 6396 2104 6404
rect 2336 6404 2344 6416
rect 2367 6417 2393 6425
rect 2467 6416 2533 6424
rect 2647 6417 2693 6425
rect 3047 6416 3184 6424
rect 2336 6396 2564 6404
rect 916 6376 1053 6384
rect 1307 6376 1413 6384
rect 1467 6375 1513 6383
rect 1647 6375 1693 6383
rect 1807 6376 1933 6384
rect 1947 6375 1973 6383
rect 2127 6375 2173 6383
rect 2227 6375 2253 6383
rect 2556 6386 2564 6396
rect 3176 6386 3184 6416
rect 3207 6416 3333 6424
rect 3387 6416 3473 6424
rect 3627 6417 3693 6425
rect 3787 6417 3833 6425
rect 4016 6404 4024 6414
rect 4067 6416 4113 6424
rect 4307 6416 4513 6424
rect 4527 6416 4573 6424
rect 4847 6417 5053 6425
rect 5256 6404 5264 6414
rect 5307 6416 5353 6424
rect 5487 6416 5533 6424
rect 5547 6416 5673 6424
rect 5776 6416 5813 6424
rect 3676 6396 3784 6404
rect 4016 6396 4124 6404
rect 5256 6396 5324 6404
rect 3676 6386 3684 6396
rect 2327 6376 2413 6384
rect 2567 6376 2673 6384
rect 2687 6376 2833 6384
rect 3507 6375 3573 6383
rect 3727 6375 3753 6383
rect 3776 6384 3784 6396
rect 3776 6376 3813 6384
rect 3927 6375 3993 6383
rect 4116 6384 4124 6396
rect 4116 6376 4133 6384
rect 4327 6376 4413 6384
rect 4467 6375 4513 6383
rect 4527 6376 4713 6384
rect 4767 6375 4793 6383
rect 4847 6376 4873 6384
rect 4927 6376 5033 6384
rect 5247 6375 5293 6383
rect 5316 6384 5324 6396
rect 5316 6376 5513 6384
rect 5527 6376 5633 6384
rect 5707 6375 5753 6383
rect 87 6356 293 6364
rect 927 6356 1013 6364
rect 1187 6356 1333 6364
rect 2296 6364 2304 6372
rect 1547 6356 2284 6364
rect 2296 6356 2333 6364
rect 1147 6336 1673 6344
rect 1687 6336 1933 6344
rect 1947 6336 2013 6344
rect 2276 6344 2284 6356
rect 3227 6356 3353 6364
rect 3367 6356 3773 6364
rect 4156 6356 4193 6364
rect 2276 6336 2513 6344
rect 2527 6336 2633 6344
rect 2887 6336 3273 6344
rect 4156 6344 4164 6356
rect 5427 6356 5453 6364
rect 5776 6364 5784 6416
rect 5867 6416 5993 6424
rect 6047 6416 6233 6424
rect 6307 6417 6333 6425
rect 6387 6416 6412 6424
rect 6447 6416 6533 6424
rect 6587 6416 6653 6424
rect 5887 6375 5913 6383
rect 5927 6376 5973 6384
rect 6207 6375 6233 6383
rect 6427 6375 6473 6383
rect 6647 6375 6673 6383
rect 5667 6356 5784 6364
rect 5807 6356 6153 6364
rect 6167 6356 6313 6364
rect 3547 6336 4164 6344
rect 4667 6336 5133 6344
rect 5147 6336 5193 6344
rect 5656 6344 5664 6353
rect 5207 6336 5664 6344
rect 5947 6336 6013 6344
rect 167 6316 453 6324
rect 2047 6316 2213 6324
rect 2467 6316 3053 6324
rect 1787 6296 1833 6304
rect 3127 6296 4173 6304
rect 4967 6296 5373 6304
rect 5387 6296 5833 6304
rect 6727 6296 6773 6304
rect 1607 6276 1733 6284
rect 2127 6276 2173 6284
rect 2187 6276 2353 6284
rect 3747 6276 4053 6284
rect 5187 6276 5753 6284
rect 5916 6276 6073 6284
rect 2427 6256 3113 6264
rect 3287 6256 3613 6264
rect 3767 6256 4593 6264
rect 5916 6264 5924 6276
rect 6127 6276 6613 6284
rect 5207 6256 5924 6264
rect 1487 6236 1753 6244
rect 3367 6236 3604 6244
rect 567 6216 593 6224
rect 1707 6216 2113 6224
rect 3356 6216 3573 6224
rect 1067 6196 1233 6204
rect 1307 6196 1573 6204
rect 1687 6196 2133 6204
rect 2527 6196 2713 6204
rect 2727 6196 3013 6204
rect 3356 6204 3364 6216
rect 3596 6224 3604 6236
rect 4067 6236 4273 6244
rect 4867 6236 5173 6244
rect 5196 6236 5933 6244
rect 3596 6216 3753 6224
rect 5196 6224 5204 6236
rect 4907 6216 5204 6224
rect 6307 6216 6633 6224
rect 3027 6196 3364 6204
rect 3567 6196 4313 6204
rect 4507 6196 5213 6204
rect 5387 6196 5573 6204
rect 607 6176 813 6184
rect 827 6176 933 6184
rect 1207 6176 1593 6184
rect 1667 6176 2213 6184
rect 2767 6176 2993 6184
rect 3067 6176 3313 6184
rect 4607 6176 4673 6184
rect 5007 6176 5193 6184
rect 5787 6176 5993 6184
rect 6107 6176 6433 6184
rect 307 6156 464 6164
rect 456 6147 464 6156
rect 747 6156 853 6164
rect 867 6156 953 6164
rect 1387 6156 1533 6164
rect 1547 6156 1613 6164
rect 1747 6156 2073 6164
rect 2887 6156 2913 6164
rect 2927 6156 3153 6164
rect 3427 6156 3493 6164
rect 3507 6156 3633 6164
rect 3687 6156 4093 6164
rect 4287 6156 4913 6164
rect 5227 6156 5473 6164
rect 5687 6156 5793 6164
rect 6467 6156 6573 6164
rect 467 6136 653 6144
rect 147 6117 213 6125
rect 227 6116 253 6124
rect 787 6116 893 6124
rect 1027 6117 1093 6125
rect 1427 6117 1453 6125
rect 1587 6116 1673 6124
rect 1687 6116 1753 6124
rect 336 6104 344 6114
rect 1916 6116 1964 6124
rect 336 6096 533 6104
rect 1836 6104 1844 6114
rect 1916 6104 1924 6116
rect 1836 6096 1924 6104
rect 1956 6104 1964 6116
rect 2187 6116 2293 6124
rect 2627 6117 2813 6125
rect 3027 6116 3113 6124
rect 1996 6104 2004 6114
rect 1956 6096 2093 6104
rect 2576 6087 2584 6114
rect 3173 6124 3187 6133
rect 3876 6136 4073 6144
rect 3876 6128 3884 6136
rect 4087 6136 4873 6144
rect 3173 6120 3193 6124
rect 3176 6116 3193 6120
rect 3847 6117 3873 6125
rect 4007 6117 4033 6125
rect 4187 6117 4273 6125
rect 3767 6096 3804 6104
rect 167 6076 313 6084
rect 487 6076 553 6084
rect 596 6076 613 6084
rect 596 6064 604 6076
rect 627 6076 753 6084
rect 867 6075 913 6083
rect 1407 6076 1473 6084
rect 1567 6076 1733 6084
rect 1787 6076 1813 6084
rect 1947 6076 1973 6084
rect 2227 6076 2313 6084
rect 2327 6076 2433 6084
rect 2567 6076 2584 6087
rect 2567 6073 2580 6076
rect 2927 6075 2993 6083
rect 3127 6075 3173 6083
rect 3287 6076 3333 6084
rect 3387 6075 3413 6083
rect 3527 6076 3553 6084
rect 3796 6084 3804 6096
rect 3796 6076 3813 6084
rect 3887 6076 3933 6084
rect 940 6064 953 6067
rect 367 6056 604 6064
rect 936 6056 953 6064
rect 940 6053 953 6056
rect 967 6056 1013 6064
rect 1027 6056 1213 6064
rect 1767 6056 1853 6064
rect 2647 6056 2733 6064
rect 2747 6056 2993 6064
rect 3956 6064 3964 6114
rect 4296 6086 4304 6136
rect 5887 6136 6073 6144
rect 6087 6136 6313 6144
rect 4327 6117 4373 6125
rect 4467 6116 4613 6124
rect 4640 6124 4653 6127
rect 4636 6113 4653 6124
rect 4707 6117 4753 6125
rect 4767 6116 4913 6124
rect 5067 6116 5113 6124
rect 5427 6117 5453 6125
rect 5587 6117 5613 6125
rect 5627 6116 5713 6124
rect 5807 6116 6153 6124
rect 6167 6116 6253 6124
rect 4636 6086 4644 6113
rect 4087 6075 4113 6083
rect 4687 6075 4733 6083
rect 4747 6076 4893 6084
rect 5147 6075 5193 6083
rect 5247 6076 5353 6084
rect 5487 6076 5553 6084
rect 5867 6076 5912 6084
rect 5947 6076 5973 6084
rect 6027 6076 6233 6084
rect 6247 6076 6353 6084
rect 3956 6056 3993 6064
rect 4187 6056 4273 6064
rect 4967 6056 5073 6064
rect 5667 6056 5693 6064
rect 5707 6056 5753 6064
rect 6427 6056 6453 6064
rect 6516 6047 6524 6114
rect 6536 6086 6544 6133
rect 6647 6117 6673 6125
rect 6647 6056 6733 6064
rect 1087 6036 1293 6044
rect 2167 6036 2533 6044
rect 2827 6036 2853 6044
rect 2867 6036 3053 6044
rect 3707 6036 3973 6044
rect 4207 6036 4433 6044
rect 4487 6036 4773 6044
rect 4787 6036 4853 6044
rect 4947 6036 4993 6044
rect 5607 6036 6153 6044
rect 6167 6036 6193 6044
rect 6467 6036 6493 6044
rect 6516 6036 6533 6047
rect 6520 6033 6533 6036
rect 87 6016 113 6024
rect 127 6016 353 6024
rect 2567 6016 2744 6024
rect 2736 6007 2744 6016
rect 3267 6016 3413 6024
rect 3607 6016 4073 6024
rect 4387 6016 5013 6024
rect 5616 6016 6093 6024
rect 1367 5996 1513 6004
rect 1927 5996 2013 6004
rect 2027 5996 2313 6004
rect 2747 5996 2933 6004
rect 2947 5996 3073 6004
rect 3667 5996 3913 6004
rect 3927 5996 4053 6004
rect 4347 5996 4693 6004
rect 5616 6004 5624 6016
rect 6587 6016 6613 6024
rect 6627 6016 6693 6024
rect 5167 5996 5624 6004
rect 5767 5996 5813 6004
rect 547 5976 573 5984
rect 1627 5976 1913 5984
rect 2367 5976 2593 5984
rect 3247 5976 3593 5984
rect 4047 5976 4433 5984
rect 5967 5976 6293 5984
rect 667 5956 833 5964
rect 1707 5956 2073 5964
rect 2087 5956 2393 5964
rect 3067 5956 3213 5964
rect 3267 5956 3553 5964
rect 3567 5956 3653 5964
rect 3827 5956 3873 5964
rect 4867 5956 5393 5964
rect 447 5936 513 5944
rect 527 5936 713 5944
rect 1067 5936 1233 5944
rect 1247 5936 1413 5944
rect 1696 5944 1704 5953
rect 1467 5936 1704 5944
rect 2507 5936 2944 5944
rect 2936 5927 2944 5936
rect 3047 5936 3893 5944
rect 3947 5936 4233 5944
rect 4447 5936 4753 5944
rect 5727 5936 5933 5944
rect 5947 5936 6084 5944
rect 807 5916 873 5924
rect 1487 5916 1533 5924
rect 1547 5924 1560 5927
rect 1547 5916 1564 5924
rect 1547 5913 1560 5916
rect 1747 5916 1793 5924
rect 2027 5916 2133 5924
rect 2147 5916 2373 5924
rect 2947 5916 3093 5924
rect 3107 5916 3173 5924
rect 5067 5916 5113 5924
rect 5127 5916 5213 5924
rect 6076 5924 6084 5936
rect 6076 5916 6353 5924
rect 167 5897 233 5905
rect 307 5896 373 5904
rect 627 5897 1093 5905
rect 1167 5897 1193 5905
rect 1307 5896 1353 5904
rect 1487 5897 1573 5905
rect 1667 5896 1753 5904
rect 1887 5897 1953 5905
rect 2247 5897 2273 5905
rect 2336 5896 2453 5904
rect 1756 5884 1764 5894
rect 2336 5884 2344 5896
rect 2467 5896 2593 5904
rect 2807 5896 2833 5904
rect 2847 5897 2893 5905
rect 2936 5896 3053 5904
rect 1756 5876 2344 5884
rect 187 5856 313 5864
rect 387 5855 413 5863
rect 527 5855 553 5863
rect 747 5856 793 5864
rect 867 5856 1013 5864
rect 1107 5856 1213 5864
rect 1387 5856 1513 5864
rect 2336 5866 2344 5876
rect 1527 5856 1533 5864
rect 1987 5856 2113 5864
rect 2187 5855 2293 5863
rect 2387 5856 2433 5864
rect 2807 5855 2873 5863
rect 2936 5864 2944 5896
rect 3107 5896 3193 5904
rect 3867 5896 3953 5904
rect 4067 5897 4133 5905
rect 4187 5896 4313 5904
rect 3256 5884 3264 5894
rect 3856 5884 3864 5894
rect 4407 5896 4573 5904
rect 4587 5897 4633 5905
rect 4687 5897 4793 5905
rect 4807 5896 4893 5904
rect 5267 5896 5313 5904
rect 5427 5896 5493 5904
rect 3196 5876 3264 5884
rect 3816 5876 3864 5884
rect 2927 5856 2944 5864
rect 3007 5855 3113 5863
rect 3196 5864 3204 5876
rect 3127 5856 3204 5864
rect 3227 5855 3293 5863
rect 3687 5856 3753 5864
rect 3767 5855 3793 5863
rect 847 5836 893 5844
rect 907 5836 953 5844
rect 967 5836 1293 5844
rect 2847 5836 2873 5844
rect 3816 5844 3824 5876
rect 3847 5855 3893 5863
rect 3907 5856 3973 5864
rect 4087 5855 4113 5863
rect 4347 5856 4453 5864
rect 5016 5856 5033 5864
rect 3367 5836 3824 5844
rect 4167 5836 4253 5844
rect 4547 5836 4733 5844
rect 5016 5844 5024 5856
rect 5047 5856 5233 5864
rect 5376 5864 5384 5894
rect 5507 5896 5553 5904
rect 5827 5897 5853 5905
rect 6087 5897 6193 5905
rect 6220 5904 6233 5907
rect 5756 5867 5764 5894
rect 5896 5884 5904 5894
rect 6216 5893 6233 5904
rect 6287 5896 6313 5904
rect 6380 5904 6393 5907
rect 6376 5893 6393 5904
rect 6507 5896 6653 5904
rect 6760 5904 6773 5907
rect 6756 5893 6773 5904
rect 5896 5876 5964 5884
rect 5376 5856 5433 5864
rect 5756 5856 5772 5867
rect 5760 5853 5772 5856
rect 5807 5856 5873 5864
rect 4927 5836 5024 5844
rect 5667 5836 5693 5844
rect 5796 5844 5804 5853
rect 5956 5864 5964 5876
rect 6216 5866 6224 5893
rect 6376 5866 6384 5893
rect 6456 5867 6464 5893
rect 5956 5856 6033 5864
rect 6307 5855 6333 5863
rect 6716 5864 6724 5893
rect 6567 5856 6724 5864
rect 6756 5847 6764 5893
rect 5747 5836 5804 5844
rect 6747 5836 6764 5847
rect 6747 5833 6760 5836
rect 127 5816 453 5824
rect 607 5816 773 5824
rect 1827 5816 1973 5824
rect 2587 5816 2953 5824
rect 3087 5816 3153 5824
rect 3567 5816 4053 5824
rect 4247 5816 4293 5824
rect 6147 5816 6253 5824
rect 1087 5796 1153 5804
rect 1167 5796 1333 5804
rect 1487 5796 2173 5804
rect 2627 5796 2673 5804
rect 2687 5796 2853 5804
rect 3187 5796 3793 5804
rect 3947 5796 4373 5804
rect 4747 5796 5073 5804
rect 5087 5796 5193 5804
rect 6447 5796 6513 5804
rect 6527 5796 6633 5804
rect 1787 5776 1873 5784
rect 1887 5776 2153 5784
rect 2267 5776 3133 5784
rect 3447 5776 3613 5784
rect 5147 5776 5353 5784
rect 5367 5776 5613 5784
rect 5947 5776 6473 5784
rect 6487 5776 6673 5784
rect 2027 5756 2053 5764
rect 2767 5756 4553 5764
rect 4647 5756 4833 5764
rect 5887 5756 5953 5764
rect 6487 5756 6552 5764
rect 6587 5756 6653 5764
rect 1727 5736 1793 5744
rect 1807 5736 2233 5744
rect 2407 5736 2473 5744
rect 2487 5736 2753 5744
rect 367 5716 1533 5724
rect 1547 5716 2013 5724
rect 2067 5716 2253 5724
rect 2307 5716 2493 5724
rect 3027 5716 3373 5724
rect 3447 5716 4033 5724
rect 4167 5716 4573 5724
rect 4587 5716 4613 5724
rect 5467 5716 6593 5724
rect 287 5696 313 5704
rect 2036 5696 2713 5704
rect 2036 5687 2044 5696
rect 3407 5696 3873 5704
rect 4207 5696 4393 5704
rect 4747 5696 4813 5704
rect 4827 5696 5153 5704
rect 5707 5696 6133 5704
rect 1147 5676 1233 5684
rect 1647 5676 1892 5684
rect 1927 5676 2032 5684
rect 2067 5676 2373 5684
rect 2807 5676 2953 5684
rect 2967 5676 3153 5684
rect 4787 5676 4953 5684
rect 6647 5676 6693 5684
rect 427 5656 453 5664
rect 467 5656 613 5664
rect 1267 5656 2693 5664
rect 2896 5656 3233 5664
rect 1427 5636 1473 5644
rect 1487 5636 2433 5644
rect 2896 5644 2904 5656
rect 3247 5656 3333 5664
rect 3587 5656 3733 5664
rect 3807 5656 4193 5664
rect 4287 5656 4633 5664
rect 5187 5656 5433 5664
rect 5447 5656 5653 5664
rect 6387 5656 6493 5664
rect 2567 5636 2904 5644
rect 3507 5636 3673 5644
rect 3807 5636 3913 5644
rect 4567 5636 4624 5644
rect 220 5624 233 5627
rect 216 5613 233 5624
rect 467 5616 653 5624
rect 1907 5616 2053 5624
rect 3207 5616 3313 5624
rect 3387 5616 4153 5624
rect 216 5584 224 5613
rect 196 5576 224 5584
rect 236 5596 313 5604
rect 67 5555 113 5563
rect 196 5544 204 5576
rect 236 5547 244 5596
rect 507 5597 553 5605
rect 747 5596 773 5604
rect 927 5596 1073 5604
rect 1567 5597 1593 5605
rect 1196 5584 1204 5594
rect 1176 5576 1204 5584
rect 1876 5584 1884 5594
rect 2267 5596 2293 5604
rect 2347 5597 2393 5605
rect 2667 5596 2813 5604
rect 2887 5597 2913 5605
rect 3147 5597 3193 5605
rect 1876 5576 1993 5584
rect 287 5556 333 5564
rect 427 5555 473 5563
rect 1176 5564 1184 5576
rect 2616 5584 2624 5594
rect 3287 5596 3424 5604
rect 2616 5576 2713 5584
rect 3416 5584 3424 5596
rect 3467 5597 3493 5605
rect 3547 5597 3593 5605
rect 3727 5596 3773 5604
rect 3787 5597 3833 5605
rect 3967 5597 3993 5605
rect 4347 5596 4433 5604
rect 4527 5597 4593 5605
rect 4616 5604 4624 5636
rect 4687 5636 5073 5644
rect 5087 5636 5113 5644
rect 5327 5636 5373 5644
rect 5827 5636 5913 5644
rect 5927 5636 5993 5644
rect 6127 5636 6313 5644
rect 5747 5616 5793 5624
rect 6320 5624 6333 5627
rect 6316 5613 6333 5624
rect 6427 5616 6513 5624
rect 4616 5596 4633 5604
rect 3416 5576 4044 5584
rect 1127 5556 1184 5564
rect 1327 5556 1453 5564
rect 1467 5556 1553 5564
rect 1727 5555 1753 5563
rect 1907 5556 1973 5564
rect 2067 5556 2153 5564
rect 2207 5556 2313 5564
rect 2467 5556 2553 5564
rect 2947 5556 3053 5564
rect 3107 5555 3273 5563
rect 3327 5555 3373 5563
rect 3447 5556 3513 5564
rect 3667 5556 3793 5564
rect 3947 5556 4013 5564
rect 4036 5564 4044 5576
rect 4476 5567 4484 5594
rect 4787 5597 4853 5605
rect 4907 5596 5033 5604
rect 5047 5596 5153 5604
rect 5327 5596 5393 5604
rect 5256 5584 5264 5594
rect 5407 5596 5453 5604
rect 5507 5597 5573 5605
rect 5847 5596 5893 5604
rect 5907 5597 5933 5605
rect 6060 5604 6073 5607
rect 6056 5593 6073 5604
rect 6167 5597 6193 5605
rect 6207 5596 6293 5604
rect 5036 5576 5264 5584
rect 4036 5556 4173 5564
rect 4187 5556 4273 5564
rect 4476 5556 4493 5567
rect 4480 5553 4493 5556
rect 5036 5564 5044 5576
rect 5027 5556 5044 5564
rect 5067 5556 5173 5564
rect 5387 5555 5433 5563
rect 5487 5556 5553 5564
rect 5696 5564 5704 5593
rect 5607 5556 5704 5564
rect 5756 5564 5764 5593
rect 5756 5556 5773 5564
rect 5827 5556 5953 5564
rect 6056 5564 6064 5593
rect 6007 5556 6064 5564
rect 6116 5564 6124 5594
rect 6087 5556 6124 5564
rect 6316 5547 6324 5613
rect 6507 5596 6533 5604
rect 6736 5567 6744 5593
rect 6407 5556 6613 5564
rect 156 5540 204 5544
rect 153 5536 204 5540
rect 153 5527 167 5536
rect 227 5536 244 5547
rect 227 5533 240 5536
rect 527 5536 893 5544
rect 1207 5536 1233 5544
rect 1547 5536 1613 5544
rect 4107 5536 4593 5544
rect 4707 5536 4913 5544
rect 5567 5536 5673 5544
rect 5847 5536 5873 5544
rect 6247 5536 6273 5544
rect 1007 5516 1653 5524
rect 1667 5516 2173 5524
rect 2227 5516 2333 5524
rect 2387 5516 2593 5524
rect 2647 5516 2773 5524
rect 2787 5516 3373 5524
rect 4187 5516 4273 5524
rect 4287 5516 4313 5524
rect 4447 5516 4512 5524
rect 4547 5516 4613 5524
rect 5507 5516 5533 5524
rect 6387 5516 6413 5524
rect 6487 5516 6573 5524
rect 6627 5516 6713 5524
rect 247 5496 393 5504
rect 2636 5504 2644 5513
rect 407 5496 2644 5504
rect 3007 5496 3073 5504
rect 3227 5496 3453 5504
rect 3787 5496 3873 5504
rect 4387 5496 4693 5504
rect 4907 5496 4953 5504
rect 4967 5496 5013 5504
rect 5227 5496 5573 5504
rect 5587 5496 5633 5504
rect 5747 5496 5813 5504
rect 5987 5496 6033 5504
rect 6207 5496 6273 5504
rect 6287 5496 6333 5504
rect 547 5476 633 5484
rect 1327 5476 2132 5484
rect 2167 5476 2613 5484
rect 2667 5476 2933 5484
rect 4647 5476 4673 5484
rect 4727 5476 4813 5484
rect 6147 5476 6553 5484
rect 6567 5476 6733 5484
rect 807 5456 1093 5464
rect 1367 5456 1873 5464
rect 2347 5456 2513 5464
rect 3547 5456 3573 5464
rect 3707 5456 3853 5464
rect 3867 5456 4373 5464
rect 4467 5456 5633 5464
rect 5647 5456 5893 5464
rect 5967 5456 6013 5464
rect 2267 5436 2293 5444
rect 2507 5436 2713 5444
rect 2727 5436 2973 5444
rect 4607 5436 4753 5444
rect 4967 5436 5253 5444
rect 6107 5436 6233 5444
rect 6507 5436 6653 5444
rect 1147 5416 1413 5424
rect 2207 5416 2233 5424
rect 2667 5416 2733 5424
rect 3247 5416 3333 5424
rect 3507 5416 3553 5424
rect 3567 5416 3653 5424
rect 3707 5416 4573 5424
rect 4787 5416 4833 5424
rect 4847 5416 4993 5424
rect 5407 5416 5473 5424
rect 5687 5416 5733 5424
rect 5747 5416 5853 5424
rect 6307 5416 6453 5424
rect 6607 5416 6633 5424
rect 627 5396 673 5404
rect 687 5396 793 5404
rect 907 5396 933 5404
rect 127 5376 153 5384
rect 167 5376 213 5384
rect 847 5376 944 5384
rect 936 5364 944 5376
rect 967 5376 1013 5384
rect 1287 5376 1453 5384
rect 1547 5377 1573 5385
rect 1627 5376 1693 5384
rect 2096 5384 2104 5413
rect 2267 5396 2393 5404
rect 2407 5396 2873 5404
rect 3527 5396 3613 5404
rect 4027 5396 4053 5404
rect 5667 5396 5713 5404
rect 6500 5404 6513 5407
rect 6496 5393 6513 5404
rect 2096 5376 2124 5384
rect 936 5356 1033 5364
rect 2116 5364 2124 5376
rect 2147 5377 2173 5385
rect 2387 5376 2453 5384
rect 2627 5377 2693 5385
rect 2787 5376 2813 5384
rect 3167 5377 3273 5385
rect 3347 5377 3413 5385
rect 2116 5356 2153 5364
rect 67 5336 93 5344
rect 227 5335 273 5343
rect 607 5336 733 5344
rect 747 5335 773 5343
rect 827 5335 872 5343
rect 907 5335 933 5343
rect 1127 5336 1293 5344
rect 1427 5335 1453 5343
rect 1767 5335 1813 5343
rect 2207 5336 2273 5344
rect 2487 5336 2593 5344
rect 2687 5335 2713 5343
rect 2936 5344 2944 5374
rect 3487 5376 3692 5384
rect 3727 5376 3813 5384
rect 3827 5376 4213 5384
rect 4347 5377 4413 5385
rect 4967 5376 5004 5384
rect 2727 5336 2944 5344
rect 2987 5336 3253 5344
rect 3307 5336 3453 5344
rect 3667 5336 3733 5344
rect 3827 5335 3853 5343
rect 3907 5336 3993 5344
rect 4047 5335 4113 5343
rect 4287 5335 4313 5343
rect 4367 5336 4473 5344
rect 4587 5335 4613 5343
rect 4816 5344 4824 5374
rect 4747 5336 4824 5344
rect 4996 5344 5004 5376
rect 5147 5377 5193 5385
rect 5407 5376 5584 5384
rect 5096 5364 5104 5374
rect 5047 5356 5104 5364
rect 5176 5356 5213 5364
rect 4996 5336 5024 5344
rect 4007 5316 4233 5324
rect 5016 5324 5024 5336
rect 5176 5344 5184 5356
rect 5127 5336 5184 5344
rect 5207 5336 5273 5344
rect 5576 5346 5584 5376
rect 5807 5377 5873 5385
rect 5927 5376 6033 5384
rect 6087 5376 6112 5384
rect 6147 5376 6193 5384
rect 6347 5377 6373 5385
rect 5756 5356 5864 5364
rect 5756 5346 5764 5356
rect 5856 5346 5864 5356
rect 5347 5336 5373 5344
rect 5427 5335 5473 5343
rect 5647 5335 5753 5343
rect 5907 5336 5953 5344
rect 6127 5335 6213 5343
rect 6307 5336 6353 5344
rect 6367 5336 6473 5344
rect 6496 5327 6504 5393
rect 6616 5376 6633 5384
rect 6616 5347 6624 5376
rect 6716 5347 6724 5373
rect 6527 5336 6544 5344
rect 5016 5316 5093 5324
rect 6247 5316 6273 5324
rect 6536 5324 6544 5336
rect 6536 5316 6693 5324
rect 6707 5316 6733 5324
rect 707 5296 973 5304
rect 2407 5296 2473 5304
rect 2547 5296 2753 5304
rect 2767 5296 2893 5304
rect 3367 5296 4713 5304
rect 4787 5296 5053 5304
rect 5507 5296 5533 5304
rect 5707 5296 5793 5304
rect 5867 5296 5973 5304
rect 6356 5296 6413 5304
rect 1027 5276 1673 5284
rect 1687 5276 2013 5284
rect 2327 5276 2393 5284
rect 2407 5276 3173 5284
rect 3587 5276 4033 5284
rect 4087 5276 4673 5284
rect 4727 5276 5073 5284
rect 6356 5284 6364 5296
rect 6187 5276 6364 5284
rect 6387 5276 6653 5284
rect 247 5256 293 5264
rect 2067 5256 2173 5264
rect 2227 5256 2353 5264
rect 2527 5256 3493 5264
rect 3747 5256 3773 5264
rect 4207 5256 4253 5264
rect 4427 5256 4513 5264
rect 4627 5256 4653 5264
rect 4707 5256 5693 5264
rect 347 5236 1193 5244
rect 1207 5236 1353 5244
rect 2207 5236 2333 5244
rect 2667 5236 2853 5244
rect 2867 5236 3053 5244
rect 3067 5236 3473 5244
rect 4567 5236 4833 5244
rect 4847 5236 4933 5244
rect 5067 5236 5153 5244
rect 5167 5236 5393 5244
rect 1727 5216 2373 5224
rect 2687 5216 3813 5224
rect 3876 5216 4073 5224
rect 247 5196 1073 5204
rect 2167 5196 2433 5204
rect 2447 5196 2633 5204
rect 2767 5196 3093 5204
rect 3876 5204 3884 5216
rect 4147 5216 4333 5224
rect 4587 5216 4733 5224
rect 3107 5196 3884 5204
rect 3907 5196 4353 5204
rect 4407 5196 4953 5204
rect 5667 5196 6053 5204
rect 1947 5176 2033 5184
rect 2047 5176 2333 5184
rect 2907 5176 3193 5184
rect 3207 5176 3213 5184
rect 3227 5176 3433 5184
rect 3787 5176 4133 5184
rect 4447 5176 4593 5184
rect 6427 5176 6493 5184
rect 1187 5156 1253 5164
rect 1587 5156 2673 5164
rect 2847 5156 3253 5164
rect 3507 5156 3533 5164
rect 4167 5156 5033 5164
rect 6227 5156 6553 5164
rect 127 5136 1093 5144
rect 3027 5136 3093 5144
rect 3327 5136 3513 5144
rect 4227 5136 4773 5144
rect 5687 5136 6093 5144
rect 6607 5136 6713 5144
rect 1627 5116 1693 5124
rect 2187 5116 2253 5124
rect 3267 5116 3573 5124
rect 3587 5116 3673 5124
rect 3687 5116 3913 5124
rect 3927 5116 4153 5124
rect 4347 5116 4473 5124
rect 4767 5116 4913 5124
rect 5007 5116 5252 5124
rect 5287 5116 5433 5124
rect 6267 5116 6453 5124
rect 6627 5116 6653 5124
rect 1287 5096 1373 5104
rect 1387 5096 1813 5104
rect 2447 5096 2653 5104
rect 2787 5096 2813 5104
rect 3167 5096 3293 5104
rect 3347 5096 3873 5104
rect 3887 5096 4393 5104
rect 4567 5096 4653 5104
rect 5227 5096 5593 5104
rect 5607 5096 5693 5104
rect 5747 5096 5793 5104
rect 87 5084 100 5087
rect 87 5073 104 5084
rect 167 5077 193 5085
rect 367 5077 393 5085
rect 447 5076 633 5084
rect 687 5076 813 5084
rect 827 5076 933 5084
rect 1147 5077 1193 5085
rect 1627 5076 1673 5084
rect 96 5046 104 5073
rect 147 5036 213 5044
rect 327 5036 353 5044
rect 367 5036 533 5044
rect 976 5044 984 5074
rect 1236 5064 1244 5074
rect 1867 5077 1913 5085
rect 1967 5077 1993 5085
rect 2127 5077 2153 5085
rect 2167 5077 2213 5085
rect 2307 5077 2353 5085
rect 2607 5076 2693 5084
rect 2887 5077 2913 5085
rect 2927 5076 3073 5084
rect 1236 5056 1513 5064
rect 787 5036 984 5044
rect 1127 5036 1173 5044
rect 1607 5035 1653 5043
rect 1667 5035 1693 5043
rect 1907 5035 2032 5043
rect 2056 5040 2093 5044
rect 2053 5036 2093 5040
rect 2053 5027 2067 5036
rect 2256 5044 2264 5073
rect 2227 5036 2264 5044
rect 2347 5036 2413 5044
rect 2507 5035 2533 5043
rect 2556 5027 2564 5074
rect 3287 5076 3353 5084
rect 3607 5077 3633 5085
rect 3727 5077 3773 5085
rect 3827 5076 3973 5084
rect 4107 5076 4293 5084
rect 4347 5076 4513 5084
rect 4527 5076 4653 5084
rect 4707 5077 4753 5085
rect 4807 5076 4893 5084
rect 5107 5076 5264 5084
rect 2647 5035 2713 5043
rect 2847 5035 2953 5043
rect 3147 5036 3233 5044
rect 3247 5035 3333 5043
rect 3667 5036 3712 5044
rect 3747 5036 3793 5044
rect 4067 5036 4304 5044
rect 127 5016 233 5024
rect 307 5016 333 5024
rect 3587 5016 3633 5024
rect 3887 5016 3933 5024
rect 4207 5016 4273 5024
rect 4296 5024 4304 5036
rect 4327 5036 4493 5044
rect 4827 5036 4893 5044
rect 5167 5036 5213 5044
rect 5256 5046 5264 5076
rect 5327 5077 5353 5085
rect 5367 5076 5473 5084
rect 5636 5064 5644 5074
rect 5496 5056 5644 5064
rect 5496 5046 5504 5056
rect 5307 5040 5344 5044
rect 5307 5036 5347 5040
rect 5333 5027 5347 5036
rect 5407 5035 5453 5043
rect 5707 5035 5753 5043
rect 5896 5044 5904 5073
rect 5976 5047 5984 5074
rect 6327 5077 6373 5085
rect 6136 5064 6144 5073
rect 6067 5056 6144 5064
rect 5896 5036 5913 5044
rect 5976 5036 5993 5047
rect 5980 5033 5993 5036
rect 6047 5036 6113 5044
rect 6207 5035 6293 5043
rect 6616 5044 6624 5074
rect 6616 5036 6693 5044
rect 4296 5016 4633 5024
rect 4887 5016 4933 5024
rect 6307 5016 6473 5024
rect 527 4996 573 5004
rect 667 4996 1433 5004
rect 1787 4996 1853 5004
rect 1867 4996 2233 5004
rect 2367 4996 2473 5004
rect 2687 4996 2893 5004
rect 3347 4996 4133 5004
rect 4467 4996 4513 5004
rect 5007 4996 5353 5004
rect 6147 4996 6173 5004
rect 6347 4996 6433 5004
rect 6527 4996 6673 5004
rect 707 4976 1193 4984
rect 1827 4976 1933 4984
rect 2027 4976 2213 4984
rect 2927 4976 3073 4984
rect 3307 4976 3593 4984
rect 3727 4976 3793 4984
rect 3807 4976 3833 4984
rect 4547 4976 4773 4984
rect 4847 4976 4973 4984
rect 5387 4976 6013 4984
rect 6027 4976 6153 4984
rect 2567 4956 2633 4964
rect 2647 4956 2793 4964
rect 3596 4964 3604 4973
rect 3596 4956 3993 4964
rect 4007 4956 4113 4964
rect 4907 4956 5113 4964
rect 6367 4956 6493 4964
rect 6567 4956 6673 4964
rect 267 4936 692 4944
rect 727 4936 853 4944
rect 867 4936 993 4944
rect 1007 4936 1253 4944
rect 1527 4936 1873 4944
rect 2007 4936 2313 4944
rect 3447 4936 3653 4944
rect 3847 4936 4053 4944
rect 4387 4936 4553 4944
rect 4747 4936 4833 4944
rect 6187 4936 6333 4944
rect 427 4916 733 4924
rect 1007 4916 1473 4924
rect 1747 4916 1893 4924
rect 2467 4916 2613 4924
rect 2787 4916 2833 4924
rect 4147 4916 4273 4924
rect 4287 4916 4824 4924
rect 4816 4907 4824 4916
rect 4887 4916 5053 4924
rect 5167 4916 5673 4924
rect 5727 4916 6013 4924
rect 6267 4916 6373 4924
rect 6427 4916 6513 4924
rect 587 4896 673 4904
rect 1247 4896 1313 4904
rect 1747 4896 1813 4904
rect 1987 4896 2292 4904
rect 2327 4896 2873 4904
rect 3247 4896 3613 4904
rect 3967 4896 4033 4904
rect 4087 4896 4113 4904
rect 4816 4896 4833 4907
rect 4820 4893 4833 4896
rect 5287 4896 5433 4904
rect 6227 4896 6333 4904
rect 6407 4896 6532 4904
rect 6567 4896 6633 4904
rect 967 4876 1053 4884
rect 1647 4876 1993 4884
rect 3027 4876 3093 4884
rect 3256 4876 3473 4884
rect -24 4856 153 4864
rect 387 4856 453 4864
rect 527 4856 613 4864
rect 700 4864 713 4867
rect 696 4853 713 4864
rect 827 4856 933 4864
rect 1047 4857 1073 4865
rect 1087 4857 1133 4865
rect 1147 4856 1273 4864
rect 1407 4856 1613 4864
rect 696 4826 704 4853
rect 1636 4826 1644 4873
rect 1747 4857 1853 4865
rect 2027 4857 2093 4865
rect 2567 4856 2653 4864
rect 2927 4857 2973 4865
rect 3256 4864 3264 4876
rect 3487 4876 3533 4884
rect 4247 4876 4473 4884
rect 4687 4876 4733 4884
rect 5527 4876 5613 4884
rect 5627 4876 5753 4884
rect 2996 4856 3264 4864
rect 2316 4836 2673 4844
rect 467 4815 493 4823
rect 547 4815 573 4823
rect 987 4815 1073 4823
rect 1127 4816 1293 4824
rect 1347 4815 1393 4823
rect 1507 4816 1593 4824
rect 1707 4815 1753 4823
rect 1907 4816 1993 4824
rect 2316 4826 2324 4836
rect 2776 4844 2784 4854
rect 2996 4844 3004 4856
rect 3587 4856 3773 4864
rect 2716 4836 3004 4844
rect 3056 4836 3384 4844
rect 2207 4816 2313 4824
rect 2487 4816 2613 4824
rect 2716 4824 2724 4836
rect 3056 4826 3064 4836
rect 2687 4816 2724 4824
rect 2847 4815 2893 4823
rect 2947 4816 3053 4824
rect 3327 4815 3353 4823
rect 3376 4824 3384 4836
rect 3376 4816 3393 4824
rect 3416 4824 3424 4854
rect 3867 4856 4033 4864
rect 4087 4856 4133 4864
rect 4147 4857 4173 4865
rect 4236 4856 4373 4864
rect 3416 4816 3453 4824
rect 4236 4826 4244 4856
rect 4447 4857 4533 4865
rect 4607 4856 4713 4864
rect 4727 4856 4753 4864
rect 4976 4856 5033 4864
rect 4676 4836 4824 4844
rect 3527 4815 3693 4823
rect 3807 4815 3833 4823
rect 3987 4815 4013 4823
rect 4307 4815 4393 4823
rect 4407 4816 4493 4824
rect 4676 4824 4684 4836
rect 4507 4816 4684 4824
rect 4727 4816 4773 4824
rect 4816 4826 4824 4836
rect 4976 4826 4984 4856
rect 5107 4856 5212 4864
rect 5247 4857 5273 4865
rect 5327 4857 5353 4865
rect 5367 4856 5473 4864
rect 5187 4816 5353 4824
rect 5576 4824 5584 4854
rect 5627 4856 5644 4864
rect 5467 4816 5584 4824
rect 5636 4807 5644 4856
rect 5887 4857 5933 4865
rect 5987 4856 6033 4864
rect 6096 4844 6104 4854
rect 6276 4856 6293 4864
rect 5936 4836 6104 4844
rect 5687 4815 5813 4823
rect 5827 4816 5913 4824
rect 5936 4807 5944 4836
rect 6236 4827 6244 4853
rect 5967 4815 6013 4823
rect 6276 4807 6284 4856
rect 6436 4826 6444 4873
rect 6467 4856 6524 4864
rect 627 4796 653 4804
rect 767 4796 833 4804
rect 2387 4796 2753 4804
rect 2767 4796 3153 4804
rect 3167 4796 3193 4804
rect 3607 4796 3633 4804
rect 4587 4796 4673 4804
rect 5567 4796 5593 4804
rect 6267 4796 6284 4807
rect 6516 4804 6524 4856
rect 6653 4864 6667 4873
rect 6627 4860 6667 4864
rect 6627 4856 6664 4860
rect 6567 4815 6632 4823
rect 6667 4816 6693 4824
rect 6516 4796 6593 4804
rect 6267 4793 6280 4796
rect 947 4776 1013 4784
rect 1027 4776 1113 4784
rect 1187 4776 1353 4784
rect 1367 4776 1433 4784
rect 1607 4776 1733 4784
rect 2127 4776 2213 4784
rect 3267 4776 3293 4784
rect 4187 4776 5093 4784
rect 5147 4776 5233 4784
rect 5867 4776 5913 4784
rect 6367 4776 6453 4784
rect 207 4756 253 4764
rect 367 4756 753 4764
rect 2287 4756 2353 4764
rect 2367 4756 3693 4764
rect 3927 4756 4193 4764
rect 4487 4756 4732 4764
rect 4767 4756 4813 4764
rect 4827 4756 5013 4764
rect 5307 4756 5753 4764
rect 6287 4756 6633 4764
rect 3187 4736 3513 4744
rect 3527 4736 4293 4744
rect 4567 4736 4593 4744
rect 4667 4736 4693 4744
rect 4867 4736 4933 4744
rect 5787 4736 6053 4744
rect 6327 4736 6593 4744
rect 1527 4716 2353 4724
rect 2987 4716 3093 4724
rect 3107 4716 3433 4724
rect 3567 4716 3913 4724
rect 4047 4716 4253 4724
rect 5167 4716 5373 4724
rect 5807 4716 6113 4724
rect 6447 4716 6533 4724
rect 67 4696 133 4704
rect 147 4696 453 4704
rect 1487 4696 2373 4704
rect 3467 4696 3753 4704
rect 3767 4696 4224 4704
rect 847 4676 1453 4684
rect 3747 4676 3933 4684
rect 3947 4676 4193 4684
rect 4216 4684 4224 4696
rect 4467 4696 6273 4704
rect 6387 4696 6693 4704
rect 4216 4676 6253 4684
rect 6547 4676 6573 4684
rect 227 4656 293 4664
rect 307 4656 593 4664
rect 1547 4656 1713 4664
rect 1727 4656 2113 4664
rect 2387 4656 2433 4664
rect 2767 4656 2993 4664
rect 4507 4656 4613 4664
rect 4667 4656 4833 4664
rect 4887 4656 4913 4664
rect 5027 4656 5133 4664
rect 127 4636 173 4644
rect 1327 4636 1513 4644
rect 2367 4636 2713 4644
rect 3047 4636 3353 4644
rect 3367 4636 3493 4644
rect 3687 4636 4413 4644
rect 5227 4636 5313 4644
rect 5607 4636 5873 4644
rect 6007 4636 6033 4644
rect 327 4616 513 4624
rect 1747 4616 2313 4624
rect 3587 4616 3793 4624
rect 3867 4616 3953 4624
rect 3967 4616 4073 4624
rect 4707 4616 4913 4624
rect 5227 4616 6373 4624
rect 6467 4616 6593 4624
rect 2407 4596 2513 4604
rect 3247 4596 3273 4604
rect 3487 4596 3533 4604
rect 3727 4596 4373 4604
rect 4427 4596 4633 4604
rect 5847 4596 5993 4604
rect 6247 4596 6393 4604
rect 6767 4604 6780 4607
rect 6767 4593 6784 4604
rect 367 4576 484 4584
rect 476 4568 484 4576
rect 1987 4576 2093 4584
rect 2367 4576 2473 4584
rect 3107 4576 3173 4584
rect 3687 4576 4113 4584
rect 4596 4576 4693 4584
rect -24 4556 93 4564
rect 407 4557 433 4565
rect 487 4557 553 4565
rect 687 4557 1053 4565
rect 1107 4556 1193 4564
rect 1587 4556 1633 4564
rect 1647 4557 1673 4565
rect 156 4544 164 4554
rect 1947 4556 2013 4564
rect 2027 4556 2133 4564
rect 2387 4557 2513 4565
rect 156 4536 324 4544
rect 47 4515 293 4523
rect 316 4524 324 4536
rect 1007 4536 1564 4544
rect 316 4516 373 4524
rect 1556 4526 1564 4536
rect 2276 4527 2284 4554
rect 2587 4556 2613 4564
rect 2807 4557 2873 4565
rect 3427 4556 3493 4564
rect 3276 4544 3284 4554
rect 3547 4556 3664 4564
rect 3276 4536 3333 4544
rect 3656 4544 3664 4556
rect 3727 4556 3784 4564
rect 3656 4536 3704 4544
rect 3696 4527 3704 4536
rect 447 4516 533 4524
rect 1707 4516 1793 4524
rect 1867 4516 1993 4524
rect 2267 4516 2284 4527
rect 2267 4513 2280 4516
rect 2407 4515 2453 4523
rect 2947 4516 3033 4524
rect 3047 4515 3073 4523
rect 3367 4515 3393 4523
rect 3487 4516 3533 4524
rect 3696 4516 3713 4527
rect 3700 4513 3713 4516
rect 3776 4526 3784 4556
rect 3807 4557 3833 4565
rect 3967 4557 4013 4565
rect 4027 4556 4053 4564
rect 3916 4524 3924 4554
rect 4127 4556 4253 4564
rect 4596 4564 4604 4576
rect 5267 4576 5473 4584
rect 5487 4576 5513 4584
rect 4307 4556 4604 4564
rect 4627 4557 4653 4565
rect 4967 4556 5073 4564
rect 4796 4544 4804 4554
rect 5347 4557 5373 4565
rect 5707 4557 5773 4565
rect 5787 4556 5872 4564
rect 4796 4536 5173 4544
rect 5216 4544 5224 4553
rect 5293 4544 5307 4553
rect 5196 4540 5307 4544
rect 5336 4544 5344 4554
rect 6107 4556 6133 4564
rect 5193 4536 5304 4540
rect 5336 4536 5544 4544
rect 5193 4527 5207 4536
rect 3887 4516 3924 4524
rect 3947 4516 4033 4524
rect 4467 4515 4513 4523
rect 4787 4516 4984 4524
rect 167 4496 253 4504
rect 1467 4496 1533 4504
rect 2167 4496 2553 4504
rect 2567 4496 3153 4504
rect 3307 4496 3433 4504
rect 3507 4496 3593 4504
rect 4107 4496 4173 4504
rect 4227 4496 4373 4504
rect 4976 4504 4984 4516
rect 5007 4516 5093 4524
rect 5107 4515 5133 4523
rect 5536 4526 5544 4536
rect 5587 4515 5753 4523
rect 5767 4515 5813 4523
rect 4976 4496 5233 4504
rect 5247 4496 5333 4504
rect 5407 4496 5473 4504
rect 5896 4504 5904 4553
rect 6156 4526 6164 4573
rect 6207 4557 6273 4565
rect 6546 4553 6547 4560
rect 6533 4544 6547 4553
rect 6376 4540 6547 4544
rect 6556 4544 6564 4554
rect 6376 4536 6543 4540
rect 6556 4536 6604 4544
rect 6376 4524 6384 4536
rect 6247 4516 6384 4524
rect 6407 4515 6573 4523
rect 6596 4507 6604 4536
rect 6580 4505 6604 4507
rect 5847 4496 5904 4504
rect 6587 4496 6604 4505
rect 6587 4493 6600 4496
rect 6776 4504 6784 4593
rect 6627 4496 6784 4504
rect 287 4476 333 4484
rect 407 4476 453 4484
rect 807 4476 913 4484
rect 2347 4476 2373 4484
rect 2387 4476 2733 4484
rect 3007 4476 3113 4484
rect 3127 4476 3253 4484
rect 3807 4476 4233 4484
rect 4847 4476 4973 4484
rect 5587 4476 6113 4484
rect 6127 4476 6153 4484
rect 6647 4476 6733 4484
rect 747 4456 1073 4464
rect 1087 4456 1373 4464
rect 1467 4456 1513 4464
rect 2267 4456 2313 4464
rect 2707 4456 2773 4464
rect 3347 4456 3553 4464
rect 3567 4456 3733 4464
rect 4236 4464 4244 4473
rect 4236 4456 4613 4464
rect 4627 4456 4733 4464
rect 5287 4456 5513 4464
rect 5827 4456 5973 4464
rect 6367 4456 6513 4464
rect 347 4436 693 4444
rect 1787 4436 2033 4444
rect 2047 4436 2233 4444
rect 2587 4436 2833 4444
rect 3307 4436 3853 4444
rect 3987 4436 4313 4444
rect 4447 4436 4513 4444
rect 5107 4436 5193 4444
rect 5547 4436 5793 4444
rect 6147 4436 6193 4444
rect 6347 4436 6393 4444
rect 6607 4436 6733 4444
rect 667 4416 833 4424
rect 1227 4416 1413 4424
rect 2427 4416 2473 4424
rect 2567 4416 2633 4424
rect 2727 4416 2933 4424
rect 3447 4416 3613 4424
rect 3627 4416 3672 4424
rect 3707 4416 3853 4424
rect 4007 4416 4153 4424
rect 4207 4416 4353 4424
rect 4536 4416 4673 4424
rect 347 4396 473 4404
rect 1647 4396 1673 4404
rect 1687 4396 1833 4404
rect 2987 4396 3173 4404
rect 4187 4396 4273 4404
rect 4536 4404 4544 4416
rect 5047 4416 5153 4424
rect 5447 4416 5473 4424
rect 5487 4416 5673 4424
rect 6447 4416 6473 4424
rect 4467 4396 4544 4404
rect 4556 4396 4893 4404
rect 987 4376 1293 4384
rect 2867 4376 3353 4384
rect 3727 4376 3893 4384
rect 4127 4376 4213 4384
rect 4556 4384 4564 4396
rect 4947 4396 4973 4404
rect 4987 4396 5633 4404
rect 6047 4396 6153 4404
rect 6247 4396 6373 4404
rect 6527 4396 6613 4404
rect 4367 4376 4564 4384
rect 5427 4376 5593 4384
rect 5867 4376 5933 4384
rect 6027 4376 6073 4384
rect 6087 4376 6213 4384
rect 6227 4376 6293 4384
rect 6467 4376 6553 4384
rect 47 4356 113 4364
rect 127 4356 193 4364
rect 907 4356 933 4364
rect 1827 4356 1893 4364
rect 1907 4356 2673 4364
rect 2887 4356 3093 4364
rect 4136 4356 4293 4364
rect 267 4336 313 4344
rect 447 4336 573 4344
rect 396 4324 404 4334
rect 727 4337 793 4345
rect 847 4337 873 4345
rect 716 4324 724 4334
rect 1047 4336 1133 4344
rect 1156 4336 1373 4344
rect 396 4316 724 4324
rect 207 4295 233 4303
rect 287 4296 333 4304
rect 1156 4306 1164 4336
rect 1387 4336 1453 4344
rect 1467 4336 1493 4344
rect 1627 4336 1733 4344
rect 1987 4337 2213 4345
rect 2680 4344 2693 4347
rect 2676 4333 2693 4344
rect 2096 4316 2193 4324
rect 547 4295 573 4303
rect 596 4296 813 4304
rect 107 4276 153 4284
rect 596 4284 604 4296
rect 1007 4295 1033 4303
rect 1267 4295 1293 4303
rect 1687 4295 1713 4303
rect 2096 4306 2104 4316
rect 2676 4306 2684 4333
rect 2796 4324 2804 4334
rect 3267 4337 3333 4345
rect 3467 4336 3533 4344
rect 3947 4337 3993 4345
rect 4136 4344 4144 4356
rect 4487 4356 4573 4364
rect 4887 4356 4953 4364
rect 5067 4356 5233 4364
rect 6396 4356 6433 4364
rect 4047 4336 4144 4344
rect 4167 4337 4193 4345
rect 2796 4316 2873 4324
rect 2893 4324 2907 4333
rect 2893 4320 2964 4324
rect 2896 4316 2964 4320
rect 2956 4306 2964 4316
rect 1847 4296 1913 4304
rect 2227 4295 2293 4303
rect 2447 4295 2473 4303
rect 3287 4295 3373 4303
rect 3447 4295 3553 4303
rect 3967 4295 4053 4303
rect 427 4276 604 4284
rect 967 4276 1113 4284
rect 4316 4284 4324 4334
rect 4407 4336 4553 4344
rect 4767 4336 4833 4344
rect 5127 4336 5193 4344
rect 5247 4337 5293 4345
rect 5307 4336 5373 4344
rect 5627 4337 5713 4345
rect 5767 4336 5813 4344
rect 5827 4336 5873 4344
rect 5927 4336 5993 4344
rect 5016 4304 5024 4333
rect 5493 4324 5507 4333
rect 5436 4320 5507 4324
rect 5433 4316 5504 4320
rect 5433 4307 5447 4316
rect 5016 4296 5073 4304
rect 5267 4296 5353 4304
rect 5487 4295 5513 4303
rect 5567 4295 5613 4303
rect 5667 4295 5693 4303
rect 5747 4295 5813 4303
rect 6056 4304 6064 4353
rect 6100 4344 6113 4347
rect 6096 4333 6113 4344
rect 6096 4306 6104 4333
rect 6196 4324 6204 4353
rect 6396 4344 6404 4356
rect 6267 4336 6404 4344
rect 6416 4336 6453 4344
rect 6416 4324 6424 4336
rect 6196 4316 6224 4324
rect 6356 4320 6424 4324
rect 5827 4296 6064 4304
rect 6107 4296 6193 4304
rect 4287 4276 4324 4284
rect 4687 4276 4733 4284
rect 4887 4276 4973 4284
rect 5767 4276 5793 4284
rect 5907 4276 5953 4284
rect 6216 4284 6224 4316
rect 6353 4316 6424 4320
rect 6353 4307 6367 4316
rect 6287 4296 6313 4304
rect 6516 4304 6524 4333
rect 6436 4296 6524 4304
rect 6216 4276 6253 4284
rect 6436 4284 6444 4296
rect 6576 4304 6584 4353
rect 6607 4336 6693 4344
rect 6713 4344 6727 4353
rect 6713 4340 6744 4344
rect 6716 4336 6744 4340
rect 6576 4296 6713 4304
rect 6407 4276 6444 4284
rect 6536 4287 6544 4292
rect 6736 4287 6744 4336
rect 6776 4307 6784 4333
rect 6536 4276 6553 4287
rect 6540 4273 6553 4276
rect 1287 4256 2033 4264
rect 2047 4256 2153 4264
rect 2167 4256 2373 4264
rect 2387 4256 2493 4264
rect 2507 4256 2613 4264
rect 2887 4256 3073 4264
rect 3567 4256 3693 4264
rect 3707 4256 3933 4264
rect 4327 4256 4373 4264
rect 4547 4256 4773 4264
rect 4787 4256 4953 4264
rect 6067 4256 6173 4264
rect 6347 4256 6453 4264
rect 6647 4256 6753 4264
rect 127 4236 833 4244
rect 887 4236 2853 4244
rect 3387 4236 3773 4244
rect 4047 4236 4173 4244
rect 5167 4236 5213 4244
rect 5307 4236 5453 4244
rect 5647 4236 6293 4244
rect 6687 4236 6713 4244
rect 307 4216 373 4224
rect 487 4216 593 4224
rect 607 4216 1193 4224
rect 1427 4216 1833 4224
rect 3027 4216 3113 4224
rect 3587 4216 3653 4224
rect 3667 4216 3913 4224
rect 3927 4216 4073 4224
rect 4427 4216 4533 4224
rect 4607 4216 4893 4224
rect 5867 4216 5933 4224
rect 6087 4216 6333 4224
rect 6427 4216 6473 4224
rect 2347 4196 2733 4204
rect 2747 4196 3033 4204
rect 3147 4196 3513 4204
rect 3707 4196 3733 4204
rect 3887 4196 4173 4204
rect 6007 4196 6393 4204
rect 6407 4196 6433 4204
rect 6507 4196 6573 4204
rect 6587 4196 6733 4204
rect 1767 4176 2393 4184
rect 3087 4176 3153 4184
rect 3207 4176 3233 4184
rect 3696 4184 3704 4193
rect 3247 4176 3704 4184
rect 3947 4176 4713 4184
rect 4907 4176 5073 4184
rect 6227 4176 6273 4184
rect 6587 4176 6613 4184
rect 3347 4156 3553 4164
rect 3867 4156 4673 4164
rect 5747 4156 5973 4164
rect 6467 4156 6653 4164
rect 447 4136 1313 4144
rect 2927 4136 3193 4144
rect 3387 4136 3713 4144
rect 3767 4136 5513 4144
rect 5527 4136 5633 4144
rect 6487 4136 6533 4144
rect 287 4116 353 4124
rect 1367 4116 1733 4124
rect 3196 4124 3204 4133
rect 3196 4116 3473 4124
rect 3907 4116 4133 4124
rect 4396 4116 4693 4124
rect 567 4096 873 4104
rect 2787 4096 2913 4104
rect 3747 4096 3993 4104
rect 4396 4104 4404 4116
rect 4707 4116 4753 4124
rect 5827 4116 6093 4124
rect 4087 4096 4404 4104
rect 4507 4096 5033 4104
rect 5047 4096 5073 4104
rect 5087 4096 5253 4104
rect 5267 4096 5473 4104
rect 5487 4096 5613 4104
rect 6167 4096 6193 4104
rect 6267 4096 6533 4104
rect 327 4076 393 4084
rect 1467 4076 1933 4084
rect 3527 4076 3653 4084
rect 3727 4076 3833 4084
rect 3927 4076 3953 4084
rect 4427 4076 4573 4084
rect 5807 4076 5873 4084
rect 5887 4076 6173 4084
rect 6627 4076 6693 4084
rect 256 4056 473 4064
rect 36 4006 44 4053
rect 256 4048 264 4056
rect 487 4056 593 4064
rect 616 4056 944 4064
rect 127 4037 153 4045
rect 227 4037 253 4045
rect 367 4036 513 4044
rect 616 4044 624 4056
rect 527 4036 624 4044
rect 107 3996 133 4004
rect 307 3996 333 4004
rect 656 4004 664 4034
rect 847 4036 913 4044
rect 936 4044 944 4056
rect 2307 4056 2673 4064
rect 2887 4056 2913 4064
rect 3047 4056 3313 4064
rect 3407 4056 3493 4064
rect 3887 4056 3933 4064
rect 4107 4056 4213 4064
rect 5947 4056 5973 4064
rect 936 4036 953 4044
rect 967 4037 993 4045
rect 1047 4036 1093 4044
rect 1107 4036 1273 4044
rect 1607 4036 1632 4044
rect 1667 4037 1693 4045
rect 1787 4036 1873 4044
rect 2067 4036 2093 4044
rect 2467 4037 2553 4045
rect 2767 4036 2993 4044
rect 3807 4036 3973 4044
rect 3987 4036 4273 4044
rect 3696 4007 3704 4033
rect 547 3996 664 4004
rect 787 3995 833 4003
rect 887 3996 933 4004
rect 1467 3996 1573 4004
rect 1647 3995 1713 4003
rect 1767 3995 1833 4003
rect 2287 3996 2333 4004
rect 2567 3996 2693 4004
rect 2927 3996 3013 4004
rect 3367 3996 3473 4004
rect 3547 3995 3613 4003
rect 4076 4006 4084 4036
rect 4347 4037 4373 4045
rect 4387 4036 4533 4044
rect 4587 4037 4633 4045
rect 4827 4037 4893 4045
rect 4967 4037 5173 4045
rect 5367 4036 5413 4044
rect 5427 4036 5673 4044
rect 5847 4036 5864 4044
rect 4416 4016 4564 4024
rect 3907 3996 3953 4004
rect 4216 4000 4253 4004
rect 4213 3996 4253 4000
rect 4213 3987 4227 3996
rect 4416 4004 4424 4016
rect 4407 3996 4424 4004
rect 4447 3996 4493 4004
rect 4556 4006 4564 4016
rect 5067 3996 5133 4004
rect 5427 3995 5493 4003
rect 5607 3995 5653 4003
rect 607 3976 713 3984
rect 3727 3976 3813 3984
rect 4587 3976 4633 3984
rect 4687 3976 4713 3984
rect 4887 3976 4933 3984
rect 5187 3976 5253 3984
rect 5407 3976 5533 3984
rect 5776 3984 5784 4033
rect 5856 4024 5864 4036
rect 5907 4036 5933 4044
rect 5856 4016 6033 4024
rect 6276 4007 6284 4034
rect 5827 3996 5893 4004
rect 6267 3996 6284 4007
rect 6316 4024 6324 4033
rect 6516 4024 6524 4034
rect 6316 4016 6524 4024
rect 6316 4004 6324 4016
rect 6316 3996 6353 4004
rect 6267 3993 6280 3996
rect 6407 3995 6453 4003
rect 5687 3976 5784 3984
rect 5927 3976 5953 3984
rect 6007 3976 6033 3984
rect 6047 3976 6133 3984
rect 6487 3976 6553 3984
rect 6616 3984 6624 4034
rect 6696 4007 6704 4033
rect 6616 3976 6653 3984
rect 127 3956 373 3964
rect 967 3956 993 3964
rect 1387 3956 1653 3964
rect 1667 3956 2813 3964
rect 3887 3956 4013 3964
rect 4267 3956 4393 3964
rect 5007 3956 5333 3964
rect 5747 3956 5813 3964
rect 6207 3956 6272 3964
rect 6307 3956 6433 3964
rect 407 3936 493 3944
rect 1667 3936 2053 3944
rect 3747 3936 3833 3944
rect 4427 3936 4913 3944
rect 6087 3936 6133 3944
rect 6467 3936 6573 3944
rect 727 3916 1093 3924
rect 1427 3916 1633 3924
rect 1656 3916 1973 3924
rect 947 3896 1033 3904
rect 1656 3904 1664 3916
rect 2147 3916 2213 3924
rect 2527 3916 3173 3924
rect 3267 3916 3653 3924
rect 3947 3916 4273 3924
rect 4327 3916 4393 3924
rect 4487 3916 4553 3924
rect 4607 3916 4973 3924
rect 6027 3916 6153 3924
rect 6167 3916 6253 3924
rect 6607 3916 6693 3924
rect 1487 3896 1664 3904
rect 2007 3896 2033 3904
rect 2647 3896 2853 3904
rect 3027 3896 3613 3904
rect 4047 3896 4073 3904
rect 4807 3896 4833 3904
rect 4887 3896 4953 3904
rect 5767 3896 5853 3904
rect 6347 3896 6413 3904
rect 6427 3896 6633 3904
rect 987 3876 1333 3884
rect 2447 3876 2773 3884
rect 3667 3876 4113 3884
rect 4487 3876 4633 3884
rect 4807 3876 5013 3884
rect 5027 3876 5273 3884
rect 6027 3876 6053 3884
rect 6527 3876 6693 3884
rect 587 3856 1193 3864
rect 1547 3856 1813 3864
rect 1867 3856 2273 3864
rect 2347 3856 2473 3864
rect 3387 3856 3413 3864
rect 3627 3856 4093 3864
rect 4256 3856 4333 3864
rect 367 3836 433 3844
rect 1267 3836 1373 3844
rect 1447 3836 1493 3844
rect 3127 3836 3284 3844
rect 167 3775 193 3783
rect 656 3784 664 3814
rect 707 3816 773 3824
rect 1067 3816 1133 3824
rect 656 3776 693 3784
rect 847 3775 973 3783
rect 1016 3767 1024 3814
rect 1207 3816 1273 3824
rect 1607 3817 1692 3825
rect 1727 3816 1793 3824
rect 1887 3816 1953 3824
rect 2007 3824 2020 3827
rect 2007 3813 2024 3824
rect 2207 3816 2273 3824
rect 2287 3816 2313 3824
rect 2500 3824 2513 3827
rect 2496 3813 2513 3824
rect 2536 3816 2613 3824
rect 2016 3786 2024 3813
rect 2496 3786 2504 3813
rect 2536 3786 2544 3816
rect 2727 3817 2753 3825
rect 2767 3816 2793 3824
rect 2887 3816 2924 3824
rect 2916 3787 2924 3816
rect 2947 3817 2993 3825
rect 3240 3824 3253 3827
rect 3236 3813 3253 3824
rect 1287 3775 1313 3783
rect 1367 3775 1413 3783
rect 1507 3776 1613 3784
rect 1667 3775 1713 3783
rect 1827 3775 1853 3783
rect 2087 3775 2253 3783
rect 2347 3776 2453 3784
rect 2607 3775 2633 3783
rect 3236 3786 3244 3813
rect 3027 3775 3053 3783
rect 3127 3776 3173 3784
rect 267 3756 293 3764
rect 307 3756 473 3764
rect 1707 3756 1773 3764
rect 1787 3756 1893 3764
rect 1907 3756 1933 3764
rect 2667 3756 2753 3764
rect 3276 3764 3284 3836
rect 3307 3836 3353 3844
rect 4256 3844 4264 3856
rect 4387 3856 4653 3864
rect 4747 3856 4993 3864
rect 5947 3856 6212 3864
rect 6247 3856 6273 3864
rect 4107 3836 4264 3844
rect 5587 3836 5693 3844
rect 5707 3836 5733 3844
rect 6407 3836 6493 3844
rect 6507 3836 6553 3844
rect 3447 3816 3473 3824
rect 3627 3817 3693 3825
rect 3796 3816 3933 3824
rect 3276 3756 3353 3764
rect 1987 3736 2133 3744
rect 3536 3744 3544 3773
rect 3647 3776 3673 3784
rect 3796 3786 3804 3816
rect 4060 3824 4073 3827
rect 4056 3813 4073 3824
rect 4327 3816 4473 3824
rect 4527 3816 4604 3824
rect 3976 3787 3984 3813
rect 4056 3786 4064 3813
rect 4276 3784 4284 3813
rect 4276 3776 4293 3784
rect 4387 3776 4433 3784
rect 3607 3756 3853 3764
rect 3507 3736 3544 3744
rect 3887 3736 3933 3744
rect 4127 3736 4453 3744
rect 4467 3736 4533 3744
rect 4596 3744 4604 3816
rect 4687 3816 4764 3824
rect 4756 3804 4764 3816
rect 4927 3816 4993 3824
rect 5047 3817 5093 3825
rect 5147 3816 5213 3824
rect 5427 3817 5513 3825
rect 5627 3820 5704 3824
rect 5627 3816 5707 3820
rect 4756 3796 4824 3804
rect 4627 3756 4733 3764
rect 4816 3764 4824 3796
rect 4836 3787 4844 3813
rect 5693 3807 5707 3816
rect 5787 3816 5833 3824
rect 6076 3787 6084 3814
rect 6167 3824 6180 3827
rect 6167 3813 6184 3824
rect 6247 3816 6313 3824
rect 6736 3824 6744 3853
rect 6367 3816 6744 3824
rect 4987 3775 5013 3783
rect 5027 3776 5113 3784
rect 5207 3775 5433 3783
rect 5507 3775 5593 3783
rect 5607 3776 5753 3784
rect 5927 3776 5993 3784
rect 6076 3776 6093 3787
rect 6080 3773 6093 3776
rect 6176 3786 6184 3813
rect 6756 3787 6764 3813
rect 6427 3776 6533 3784
rect 6667 3775 6713 3783
rect 4816 3756 5093 3764
rect 6327 3756 6413 3764
rect 4596 3736 5493 3744
rect 5647 3736 6093 3744
rect 6467 3736 6493 3744
rect 127 3716 153 3724
rect 207 3716 593 3724
rect 607 3716 1033 3724
rect 2907 3716 2993 3724
rect 3007 3716 3593 3724
rect 3747 3716 3953 3724
rect 3967 3716 4093 3724
rect 4647 3716 4713 3724
rect 4867 3716 5073 3724
rect 5547 3716 6173 3724
rect 6227 3716 6453 3724
rect 2247 3696 2513 3704
rect 2527 3696 3553 3704
rect 3707 3696 3913 3704
rect 3927 3696 3953 3704
rect 4507 3696 4613 3704
rect 5247 3696 5433 3704
rect 5447 3696 5473 3704
rect 5487 3696 5593 3704
rect 5807 3696 6053 3704
rect 6627 3696 6733 3704
rect 207 3676 413 3684
rect 427 3676 573 3684
rect 1107 3676 1173 3684
rect 1187 3676 1553 3684
rect 2267 3676 3093 3684
rect 3107 3676 3113 3684
rect 3767 3676 4313 3684
rect 6127 3676 6313 3684
rect 6367 3676 6593 3684
rect 947 3656 2233 3664
rect 2827 3656 3153 3664
rect 3567 3656 3833 3664
rect 4316 3664 4324 3673
rect 4316 3656 4573 3664
rect 4787 3656 5173 3664
rect 6387 3656 6553 3664
rect 707 3636 833 3644
rect 847 3636 1733 3644
rect 1947 3636 2753 3644
rect 3287 3636 3793 3644
rect 3927 3636 3973 3644
rect 4947 3636 4993 3644
rect 5007 3636 5033 3644
rect 5547 3636 5633 3644
rect 6587 3636 6773 3644
rect 2407 3616 2493 3624
rect 3367 3616 3433 3624
rect 3587 3616 3733 3624
rect 4887 3616 4913 3624
rect 5247 3616 5924 3624
rect 5916 3607 5924 3616
rect 6207 3616 6273 3624
rect 1267 3596 1493 3604
rect 2447 3596 2893 3604
rect 3036 3596 3453 3604
rect 1147 3576 1313 3584
rect 3036 3584 3044 3596
rect 3467 3596 3753 3604
rect 3807 3596 3973 3604
rect 4047 3596 4213 3604
rect 4587 3596 4753 3604
rect 4847 3596 5033 3604
rect 5347 3596 5553 3604
rect 5916 3596 5933 3607
rect 5920 3593 5933 3596
rect 6067 3596 6093 3604
rect 1747 3576 3044 3584
rect 3407 3576 3473 3584
rect 4567 3576 4693 3584
rect 5067 3576 5253 3584
rect 6116 3576 6293 3584
rect 267 3556 393 3564
rect 407 3556 453 3564
rect 587 3556 1464 3564
rect 1456 3547 1464 3556
rect 2787 3556 2853 3564
rect 2907 3556 3233 3564
rect 3247 3556 3513 3564
rect 3807 3556 3993 3564
rect 4107 3556 4644 3564
rect 4636 3547 4644 3556
rect 5107 3556 5333 3564
rect 5387 3556 5793 3564
rect 6116 3564 6124 3576
rect 5847 3556 6124 3564
rect 6287 3556 6393 3564
rect 6447 3556 6613 3564
rect 6707 3556 6773 3564
rect 1467 3536 1533 3544
rect 2887 3536 2913 3544
rect 4007 3536 4073 3544
rect 4636 3536 4653 3547
rect 4640 3533 4653 3536
rect 4667 3536 4853 3544
rect 4867 3536 4933 3544
rect 5147 3536 5193 3544
rect 5927 3544 5940 3547
rect 5927 3533 5944 3544
rect 6527 3536 6573 3544
rect -24 3516 93 3524
rect 336 3516 353 3524
rect 336 3487 344 3516
rect 447 3517 493 3525
rect 547 3517 573 3525
rect 627 3517 673 3525
rect 727 3517 773 3525
rect 1027 3516 1053 3524
rect 396 3504 404 3514
rect 876 3504 884 3514
rect 1107 3516 1133 3524
rect 1287 3516 1304 3524
rect 396 3496 544 3504
rect 876 3496 1073 3504
rect 147 3476 293 3484
rect 387 3480 424 3484
rect 387 3476 427 3480
rect 413 3467 427 3476
rect 447 3475 513 3483
rect 536 3484 544 3496
rect 536 3476 553 3484
rect 607 3476 693 3484
rect 787 3476 853 3484
rect 967 3476 1113 3484
rect 167 3456 233 3464
rect 1176 3464 1184 3514
rect 1216 3487 1224 3514
rect 1296 3487 1304 3516
rect 1627 3517 1693 3525
rect 1867 3516 1993 3524
rect 2107 3517 2133 3525
rect 2187 3517 2393 3525
rect 2407 3516 2553 3524
rect 2607 3516 2653 3524
rect 2556 3504 2564 3514
rect 2667 3516 2693 3524
rect 2936 3516 3033 3524
rect 2556 3496 2633 3504
rect 1207 3476 1224 3487
rect 1207 3473 1220 3476
rect 1647 3476 1713 3484
rect 1847 3475 1933 3483
rect 2787 3476 2813 3484
rect 2836 3467 2844 3514
rect 2936 3504 2944 3516
rect 3107 3516 3133 3524
rect 3287 3517 3313 3525
rect 2856 3496 2944 3504
rect 2856 3486 2864 3496
rect 3376 3484 3384 3514
rect 3667 3516 3693 3524
rect 3847 3517 3873 3525
rect 3887 3516 3913 3524
rect 4187 3517 4213 3525
rect 4507 3517 4573 3525
rect 3227 3476 3384 3484
rect 3496 3484 3504 3513
rect 3973 3504 3987 3513
rect 4136 3504 4144 3514
rect 3973 3500 4184 3504
rect 3976 3496 4184 3500
rect 4176 3487 4184 3496
rect 3447 3476 3504 3484
rect 3907 3476 3933 3484
rect 4107 3476 4153 3484
rect 4176 3476 4192 3487
rect 4180 3473 4192 3476
rect 4227 3476 4273 3484
rect 4296 3467 4304 3514
rect 4336 3484 4344 3514
rect 5087 3517 5133 3525
rect 5267 3524 5280 3527
rect 5267 3513 5284 3524
rect 5407 3517 5473 3525
rect 4796 3487 4804 3513
rect 4336 3476 4373 3484
rect 4427 3476 4453 3484
rect 4527 3476 4673 3484
rect 4947 3475 4973 3483
rect 5167 3476 5233 3484
rect 5276 3486 5284 3513
rect 1176 3456 1333 3464
rect 2727 3456 2753 3464
rect 4687 3456 4753 3464
rect 4887 3456 5073 3464
rect 5336 3464 5344 3514
rect 5467 3476 5613 3484
rect 5636 3464 5644 3514
rect 5727 3517 5753 3525
rect 5676 3487 5684 3513
rect 5936 3504 5944 3533
rect 5916 3496 5944 3504
rect 5847 3476 5873 3484
rect 5916 3486 5924 3496
rect 5956 3486 5964 3533
rect 5987 3517 6013 3525
rect 6147 3517 6213 3525
rect 6280 3524 6293 3527
rect 6276 3513 6293 3524
rect 6667 3524 6680 3527
rect 6667 3513 6684 3524
rect 6276 3487 6284 3513
rect 6127 3475 6173 3483
rect 6276 3476 6293 3487
rect 6280 3473 6293 3476
rect 6356 3467 6364 3513
rect 6453 3504 6467 3513
rect 6676 3504 6684 3513
rect 6453 3500 6664 3504
rect 6456 3496 6664 3500
rect 6676 3496 6724 3504
rect 6587 3476 6633 3484
rect 6656 3484 6664 3496
rect 6716 3486 6724 3496
rect 6656 3476 6684 3484
rect 6676 3467 6684 3476
rect 6735 3467 6743 3514
rect 6767 3524 6780 3527
rect 6767 3513 6784 3524
rect 6776 3467 6784 3513
rect 5307 3456 5644 3464
rect 5856 3456 5953 3464
rect 307 3436 432 3444
rect 467 3436 653 3444
rect 1007 3436 1533 3444
rect 1547 3436 1733 3444
rect 1747 3436 1773 3444
rect 1787 3436 2173 3444
rect 2647 3436 2873 3444
rect 2887 3436 2993 3444
rect 3227 3436 3333 3444
rect 3407 3436 3473 3444
rect 3567 3436 3633 3444
rect 3676 3436 3813 3444
rect 347 3416 393 3424
rect 547 3416 613 3424
rect 2267 3416 2413 3424
rect 2667 3416 2833 3424
rect 3676 3424 3684 3436
rect 4447 3436 4573 3444
rect 4967 3436 5033 3444
rect 5327 3436 5373 3444
rect 5856 3444 5864 3456
rect 6356 3456 6373 3467
rect 6360 3453 6373 3456
rect 6487 3456 6653 3464
rect 6676 3456 6693 3467
rect 6680 3453 6693 3456
rect 5807 3436 5864 3444
rect 3587 3416 3684 3424
rect 3967 3416 4153 3424
rect 4167 3416 4253 3424
rect 4727 3416 5453 3424
rect 5507 3416 5773 3424
rect 5887 3416 6013 3424
rect 6067 3416 6333 3424
rect 567 3396 893 3404
rect 2027 3396 2053 3404
rect 2067 3396 2133 3404
rect 3267 3396 3653 3404
rect 3747 3396 3773 3404
rect 4367 3396 4693 3404
rect 4747 3396 5213 3404
rect 5227 3396 5393 3404
rect 5567 3396 5813 3404
rect 5947 3396 6173 3404
rect 147 3376 1573 3384
rect 1827 3376 2353 3384
rect 2827 3376 3164 3384
rect 1287 3356 1313 3364
rect 1327 3356 1473 3364
rect 1487 3356 1533 3364
rect 2547 3356 2593 3364
rect 2747 3356 2913 3364
rect 3156 3364 3164 3376
rect 3807 3376 4073 3384
rect 4087 3376 4113 3384
rect 4307 3376 5193 3384
rect 5667 3376 5793 3384
rect 5907 3376 6113 3384
rect 6347 3376 6673 3384
rect 3156 3356 3413 3364
rect 4627 3356 4833 3364
rect 4847 3356 4933 3364
rect 6187 3356 6253 3364
rect 6733 3364 6747 3373
rect 6707 3360 6747 3364
rect 6707 3356 6744 3360
rect 867 3336 993 3344
rect 1047 3336 1213 3344
rect 1347 3336 1813 3344
rect 2287 3336 2393 3344
rect 2467 3336 2773 3344
rect 2787 3336 3093 3344
rect 3147 3336 3633 3344
rect 3647 3336 3733 3344
rect 4027 3336 4213 3344
rect 4307 3336 4373 3344
rect 4447 3336 4533 3344
rect 4647 3336 4704 3344
rect 4696 3327 4704 3336
rect 5207 3336 5373 3344
rect 5487 3336 5733 3344
rect 5827 3336 5853 3344
rect 6047 3336 6073 3344
rect 6307 3336 6413 3344
rect 6427 3336 6433 3344
rect 6627 3336 6673 3344
rect 1307 3316 1393 3324
rect 1887 3316 1944 3324
rect -24 3296 193 3304
rect 207 3296 273 3304
rect 627 3296 664 3304
rect -24 3256 93 3264
rect 507 3255 553 3263
rect 656 3264 664 3296
rect 907 3297 993 3305
rect 1107 3297 1133 3305
rect 656 3256 733 3264
rect 1036 3264 1044 3294
rect 1556 3266 1564 3313
rect 1936 3266 1944 3316
rect 2987 3316 3053 3324
rect 4356 3316 4473 3324
rect 2127 3296 2213 3304
rect 2240 3304 2253 3307
rect 2236 3293 2253 3304
rect 2340 3304 2353 3307
rect 2336 3293 2353 3304
rect 2236 3266 2244 3293
rect 2336 3266 2344 3293
rect 2576 3266 2584 3313
rect 2807 3296 2913 3304
rect 3107 3297 3333 3305
rect 3427 3297 3533 3305
rect 3707 3296 3733 3304
rect 3996 3296 4073 3304
rect 3996 3284 4004 3296
rect 4356 3304 4364 3316
rect 4527 3316 4613 3324
rect 4696 3316 4713 3327
rect 4700 3313 4713 3316
rect 6187 3316 6273 3324
rect 6367 3316 6393 3324
rect 6436 3324 6444 3333
rect 6436 3316 6593 3324
rect 4347 3296 4364 3304
rect 4387 3297 4432 3305
rect 3916 3276 4004 3284
rect 1036 3256 1153 3264
rect 1227 3255 1253 3263
rect 1607 3255 1753 3263
rect 2147 3255 2193 3263
rect 2827 3255 2893 3263
rect 2947 3255 2973 3263
rect 3387 3256 3413 3264
rect 3916 3264 3924 3276
rect 3867 3256 3924 3264
rect 4007 3255 4053 3263
rect 4236 3264 4244 3294
rect 4336 3284 4344 3294
rect 4547 3297 4673 3305
rect 4787 3297 4833 3305
rect 5027 3296 5064 3304
rect 4256 3280 4344 3284
rect 4147 3256 4244 3264
rect 4253 3276 4344 3280
rect 4253 3267 4267 3276
rect 4456 3267 4464 3293
rect 5056 3287 5064 3296
rect 5107 3297 5133 3305
rect 5147 3296 5253 3304
rect 5367 3297 5433 3305
rect 5987 3296 6044 3304
rect 4767 3276 5004 3284
rect 5056 3276 5073 3287
rect 4307 3256 4353 3264
rect 4996 3266 5004 3276
rect 5060 3273 5073 3276
rect 5387 3255 5413 3263
rect 5616 3264 5624 3294
rect 5616 3260 5644 3264
rect 5616 3256 5647 3260
rect 5633 3247 5647 3256
rect 5667 3256 5733 3264
rect 5867 3255 5913 3263
rect 387 3236 433 3244
rect 1027 3236 1073 3244
rect 2407 3236 2613 3244
rect 4647 3236 4873 3244
rect 5087 3236 5313 3244
rect 5727 3236 5773 3244
rect 6016 3244 6024 3273
rect 5907 3236 6024 3244
rect 6036 3244 6044 3296
rect 6076 3267 6084 3294
rect 6227 3304 6240 3307
rect 6227 3293 6244 3304
rect 6067 3256 6084 3267
rect 6067 3253 6080 3256
rect 6147 3255 6173 3263
rect 6236 3264 6244 3293
rect 6616 3296 6633 3304
rect 6616 3284 6624 3296
rect 6547 3276 6624 3284
rect 6236 3256 6273 3264
rect 6347 3256 6373 3264
rect 6467 3256 6573 3264
rect 6036 3236 6093 3244
rect 767 3216 1153 3224
rect 3327 3216 3373 3224
rect 3387 3216 3493 3224
rect 3827 3216 4073 3224
rect 4427 3216 4533 3224
rect 4967 3216 5033 3224
rect 447 3196 673 3204
rect 1487 3196 1993 3204
rect 2007 3196 2553 3204
rect 3427 3196 4033 3204
rect 4387 3196 4573 3204
rect 4707 3196 4873 3204
rect 5067 3196 5273 3204
rect 5607 3196 5833 3204
rect 5927 3196 6273 3204
rect 1467 3176 1633 3184
rect 1647 3176 1873 3184
rect 1887 3176 2273 3184
rect 4127 3176 4213 3184
rect 4227 3176 4333 3184
rect 4347 3176 4553 3184
rect 5967 3176 6233 3184
rect 3087 3156 3673 3164
rect 3687 3156 4093 3164
rect 5327 3156 5513 3164
rect 5527 3156 5613 3164
rect 5827 3156 6413 3164
rect 6427 3156 6613 3164
rect 6627 3156 6673 3164
rect 547 3136 833 3144
rect 1507 3136 1713 3144
rect 1727 3136 1953 3144
rect 3407 3136 4213 3144
rect 4327 3136 4473 3144
rect 5647 3136 5973 3144
rect 5987 3136 6053 3144
rect 6147 3136 6453 3144
rect 267 3116 1093 3124
rect 1227 3116 1453 3124
rect 1767 3116 2273 3124
rect 3467 3116 3973 3124
rect 4047 3116 4113 3124
rect 4287 3116 4613 3124
rect 4687 3116 5073 3124
rect 5767 3116 5953 3124
rect 6487 3116 6773 3124
rect 667 3096 1053 3104
rect 1147 3096 1693 3104
rect 2387 3096 3133 3104
rect 4187 3096 4653 3104
rect 4836 3096 5593 3104
rect 4836 3087 4844 3096
rect 5756 3104 5764 3113
rect 5636 3096 5764 3104
rect 567 3076 813 3084
rect 1107 3076 2093 3084
rect 2507 3076 3413 3084
rect 3647 3076 3673 3084
rect 3687 3076 3913 3084
rect 3927 3076 3993 3084
rect 4227 3076 4413 3084
rect 4527 3076 4593 3084
rect 4827 3076 4844 3087
rect 4827 3073 4840 3076
rect 4867 3076 5333 3084
rect 5636 3084 5644 3096
rect 5547 3076 5644 3084
rect 5927 3076 6013 3084
rect 6067 3076 6353 3084
rect 6527 3076 6773 3084
rect 747 3056 933 3064
rect 1167 3056 1673 3064
rect 3447 3056 3473 3064
rect 4727 3056 4793 3064
rect 4807 3056 5033 3064
rect 6407 3056 6433 3064
rect 6447 3056 6533 3064
rect -24 3024 -16 3044
rect 427 3036 553 3044
rect 2147 3036 2453 3044
rect 2907 3036 3013 3044
rect 3987 3036 4313 3044
rect 4627 3036 5133 3044
rect 5147 3036 5213 3044
rect 5436 3036 5493 3044
rect -24 3016 113 3024
rect 527 3016 693 3024
rect 847 3016 1013 3024
rect 1027 3016 1153 3024
rect 1527 3016 1573 3024
rect 2247 3016 2493 3024
rect 2547 3016 2613 3024
rect 3296 3016 3613 3024
rect -24 2996 253 3004
rect 607 2997 633 3005
rect 787 2996 933 3004
rect 1067 2996 1124 3004
rect 1116 2984 1124 2996
rect 1287 2997 1313 3005
rect 1393 3004 1407 3013
rect 1376 3000 1407 3004
rect 1376 2996 1404 3000
rect 276 2976 724 2984
rect 1116 2976 1144 2984
rect 276 2964 284 2976
rect 167 2956 284 2964
rect 307 2956 653 2964
rect 716 2966 724 2976
rect 807 2955 993 2963
rect 1136 2964 1144 2976
rect 1376 2967 1384 2996
rect 1736 2996 1773 3004
rect 1136 2956 1193 2964
rect 527 2936 573 2944
rect 1416 2944 1424 2993
rect 1736 2984 1744 2996
rect 1567 2976 1744 2984
rect 1727 2955 1753 2963
rect 1816 2964 1824 2994
rect 1867 2996 1913 3004
rect 2187 2997 2233 3005
rect 2327 2996 2413 3004
rect 2667 2997 2693 3005
rect 2887 2997 2933 3005
rect 3187 2997 3233 3005
rect 2316 2984 2324 2994
rect 2207 2976 2324 2984
rect 1816 2956 1933 2964
rect 2007 2955 2073 2963
rect 2567 2955 2593 2963
rect 2607 2956 2753 2964
rect 2807 2955 2833 2963
rect 3167 2956 3213 2964
rect 3296 2966 3304 3016
rect 4087 3024 4100 3027
rect 4087 3013 4104 3024
rect 4207 3016 4293 3024
rect 4667 3016 4853 3024
rect 5436 3024 5444 3036
rect 5507 3036 5553 3044
rect 5707 3036 5933 3044
rect 5947 3036 6133 3044
rect 6267 3036 6313 3044
rect 6327 3036 6513 3044
rect 6596 3036 6653 3044
rect 5267 3016 5444 3024
rect 6596 3024 6604 3036
rect 6547 3016 6604 3024
rect 3827 2996 3853 3004
rect 3473 2984 3487 2993
rect 3416 2980 3487 2984
rect 4096 2984 4104 3013
rect 4327 2997 4373 3005
rect 4447 2996 4513 3004
rect 4476 2984 4484 2996
rect 4627 2997 4713 3005
rect 3413 2976 3484 2980
rect 4096 2976 4144 2984
rect 3413 2967 3427 2976
rect 3467 2956 3493 2964
rect 3707 2956 3793 2964
rect 4087 2960 4124 2964
rect 4087 2956 4127 2960
rect 4113 2947 4127 2956
rect 1307 2936 1424 2944
rect 1647 2936 1853 2944
rect 1867 2936 2373 2944
rect 2647 2936 2673 2944
rect 4136 2944 4144 2976
rect 4436 2976 4484 2984
rect 4556 2984 4564 2994
rect 4887 2997 4953 3005
rect 5107 2997 5173 3005
rect 5667 2997 5693 3005
rect 5707 2996 5833 3004
rect 4753 2984 4767 2993
rect 4556 2980 4767 2984
rect 4556 2976 4764 2980
rect 4247 2956 4313 2964
rect 4436 2964 4444 2976
rect 4407 2956 4444 2964
rect 4467 2956 4493 2964
rect 4547 2956 4613 2964
rect 4136 2936 4193 2944
rect 4636 2944 4644 2976
rect 4816 2964 4824 2993
rect 5456 2984 5464 2994
rect 5987 2996 6093 3004
rect 6327 2996 6473 3004
rect 6527 2997 6613 3005
rect 5407 2976 5464 2984
rect 5916 2967 5924 2993
rect 4747 2956 4824 2964
rect 4867 2956 4933 2964
rect 5027 2956 5073 2964
rect 5167 2956 5253 2964
rect 5567 2955 5593 2963
rect 5647 2956 5873 2964
rect 6047 2955 6113 2963
rect 6167 2956 6213 2964
rect 6256 2964 6264 2993
rect 6596 2967 6604 2997
rect 6256 2956 6333 2964
rect 6387 2964 6400 2967
rect 6387 2953 6404 2964
rect 4636 2936 4713 2944
rect 5187 2936 5213 2944
rect 6036 2944 6044 2952
rect 5967 2936 6044 2944
rect 6247 2936 6273 2944
rect 6396 2944 6404 2953
rect 6696 2947 6704 2993
rect 6396 2936 6433 2944
rect 6567 2936 6653 2944
rect 6696 2936 6713 2947
rect 6700 2933 6713 2936
rect 456 2916 853 2924
rect 456 2907 464 2916
rect 867 2916 993 2924
rect 1887 2916 1933 2924
rect 2447 2916 2813 2924
rect 3247 2916 3293 2924
rect 3587 2916 3673 2924
rect 3747 2916 3913 2924
rect 4087 2916 4153 2924
rect 4987 2916 5393 2924
rect 6167 2916 6192 2924
rect 6227 2916 6424 2924
rect 227 2896 453 2904
rect 1187 2896 1293 2904
rect 1587 2896 1793 2904
rect 2267 2896 2573 2904
rect 2967 2896 3453 2904
rect 3936 2896 3973 2904
rect 1047 2876 1313 2884
rect 1367 2876 1393 2884
rect 1607 2876 1672 2884
rect 1707 2876 2113 2884
rect 2987 2876 3733 2884
rect 3936 2884 3944 2896
rect 4287 2896 4484 2904
rect 3887 2876 3944 2884
rect 4127 2876 4233 2884
rect 4476 2884 4484 2896
rect 4507 2896 5413 2904
rect 5427 2896 5433 2904
rect 6087 2896 6133 2904
rect 6307 2896 6353 2904
rect 6367 2896 6393 2904
rect 6416 2904 6424 2916
rect 6507 2916 6533 2924
rect 6416 2896 6453 2904
rect 6547 2896 6673 2904
rect 4476 2876 4693 2884
rect 5607 2876 5653 2884
rect 5667 2876 5693 2884
rect 5747 2876 5953 2884
rect 147 2856 313 2864
rect 327 2856 573 2864
rect 787 2856 833 2864
rect 1127 2856 1433 2864
rect 1447 2856 1773 2864
rect 1787 2856 1993 2864
rect 2547 2856 3253 2864
rect 3907 2856 3953 2864
rect 4107 2856 4273 2864
rect 4647 2856 4693 2864
rect 4927 2856 5133 2864
rect 5487 2856 5773 2864
rect 5787 2856 5833 2864
rect 5907 2856 6133 2864
rect 6487 2856 6573 2864
rect 6587 2856 6633 2864
rect 1007 2836 1172 2844
rect 1207 2836 1493 2844
rect 2507 2836 2973 2844
rect 3527 2836 4033 2844
rect 4147 2836 4573 2844
rect 4587 2836 4773 2844
rect 4787 2836 5093 2844
rect 5247 2836 5573 2844
rect 5587 2836 5793 2844
rect 6267 2836 6613 2844
rect 527 2816 633 2824
rect 927 2816 1533 2824
rect 1547 2816 1813 2824
rect 1827 2816 2033 2824
rect 2047 2816 2193 2824
rect 2207 2816 2793 2824
rect 2807 2816 2873 2824
rect 3107 2816 3133 2824
rect 3147 2816 3313 2824
rect 3827 2816 4093 2824
rect 4207 2816 4604 2824
rect 4596 2807 4604 2816
rect 6067 2816 6093 2824
rect 6507 2816 6593 2824
rect 2307 2796 2493 2804
rect 2507 2796 2633 2804
rect 3627 2796 3713 2804
rect 4007 2796 4033 2804
rect 4367 2804 4380 2807
rect 4367 2793 4384 2804
rect 6007 2796 6153 2804
rect 6207 2796 6473 2804
rect 227 2776 364 2784
rect 356 2747 364 2776
rect 407 2777 453 2785
rect 507 2776 613 2784
rect 867 2777 893 2785
rect 947 2776 1013 2784
rect 1627 2777 1653 2785
rect 1707 2776 1753 2784
rect -24 2736 93 2744
rect 607 2735 773 2743
rect 907 2735 993 2743
rect 1056 2744 1064 2774
rect 1867 2776 1913 2784
rect 1967 2776 2193 2784
rect 2207 2777 2253 2785
rect 2707 2776 2824 2784
rect 2816 2764 2824 2776
rect 2976 2776 3024 2784
rect 2976 2764 2984 2776
rect 2816 2756 2984 2764
rect 1056 2736 1073 2744
rect 1087 2736 1213 2744
rect 1307 2735 1373 2743
rect 1447 2735 1513 2743
rect 1607 2735 1673 2743
rect 1787 2735 1833 2743
rect 1887 2735 1953 2743
rect 2807 2735 2993 2743
rect 3016 2744 3024 2776
rect 3067 2777 3153 2785
rect 3227 2776 3373 2784
rect 3387 2777 3453 2785
rect 3667 2777 3693 2785
rect 3736 2776 3773 2784
rect 3736 2767 3744 2776
rect 3787 2776 3813 2784
rect 3720 2766 3744 2767
rect 3727 2756 3744 2766
rect 4147 2776 4213 2784
rect 4327 2777 4353 2785
rect 3913 2764 3927 2773
rect 3913 2760 3984 2764
rect 3916 2756 3984 2760
rect 3727 2753 3740 2756
rect 3016 2736 3033 2744
rect 3056 2736 3173 2744
rect 227 2716 333 2724
rect 2007 2716 2073 2724
rect 2087 2716 2313 2724
rect 3056 2724 3064 2736
rect 3307 2736 3353 2744
rect 3367 2736 3693 2744
rect 3736 2740 3933 2744
rect 3733 2736 3933 2740
rect 3733 2727 3747 2736
rect 2547 2716 3064 2724
rect 3407 2716 3453 2724
rect 3587 2716 3673 2724
rect 3976 2724 3984 2756
rect 4007 2735 4033 2743
rect 4227 2735 4253 2743
rect 4376 2744 4384 2793
rect 4447 2776 4484 2784
rect 4476 2747 4484 2776
rect 4596 2764 4604 2793
rect 4627 2776 4753 2784
rect 4767 2776 4913 2784
rect 5387 2776 5433 2784
rect 5487 2777 5513 2785
rect 5627 2777 5693 2785
rect 5887 2776 5984 2784
rect 4536 2760 4604 2764
rect 4533 2756 4604 2760
rect 4533 2747 4547 2756
rect 5976 2747 5984 2776
rect 6047 2776 6113 2784
rect 6507 2776 6644 2784
rect 6267 2756 6344 2764
rect 4376 2736 4413 2744
rect 4707 2736 4953 2744
rect 5127 2736 5213 2744
rect 5227 2736 5353 2744
rect 5587 2735 5673 2743
rect 5727 2735 5773 2743
rect 6336 2746 6344 2756
rect 6107 2735 6173 2743
rect 6407 2736 6433 2744
rect 6487 2736 6613 2744
rect 6636 2744 6644 2776
rect 6636 2736 6673 2744
rect 3976 2716 4113 2724
rect 4467 2716 4564 2724
rect 733 2704 747 2713
rect 4556 2707 4564 2716
rect 4727 2716 4753 2724
rect 4887 2716 4933 2724
rect 5927 2716 5953 2724
rect 6067 2716 6233 2724
rect 6247 2716 6273 2724
rect 507 2700 747 2704
rect 507 2696 744 2700
rect 927 2696 1613 2704
rect 1727 2696 1913 2704
rect 1987 2696 2153 2704
rect 3167 2696 3713 2704
rect 4167 2696 4353 2704
rect 4467 2696 4493 2704
rect 4567 2696 4633 2704
rect 5547 2696 5613 2704
rect 5627 2696 5853 2704
rect 6147 2696 6353 2704
rect 6667 2696 6713 2704
rect 47 2676 273 2684
rect 287 2676 373 2684
rect 2287 2676 3213 2684
rect 3647 2676 3753 2684
rect 3927 2676 4053 2684
rect 4787 2676 4973 2684
rect 4987 2676 5393 2684
rect 6027 2676 6093 2684
rect 6447 2676 6633 2684
rect 527 2656 733 2664
rect 1387 2656 1793 2664
rect 1807 2656 2013 2664
rect 2027 2656 2173 2664
rect 2187 2656 2893 2664
rect 2907 2656 2973 2664
rect 2987 2656 3073 2664
rect 3267 2656 3613 2664
rect 4127 2656 4293 2664
rect 4907 2656 5253 2664
rect 5267 2656 5293 2664
rect 6427 2656 6713 2664
rect 27 2636 393 2644
rect 647 2636 933 2644
rect 1427 2636 1473 2644
rect 1487 2636 2273 2644
rect 3127 2636 3173 2644
rect 5947 2636 6033 2644
rect 447 2616 593 2624
rect 3427 2616 3593 2624
rect 3607 2616 4173 2624
rect 4627 2616 5053 2624
rect 5067 2616 5173 2624
rect 5187 2616 5253 2624
rect 2887 2596 3273 2604
rect 3527 2596 3713 2604
rect 4067 2596 4313 2604
rect 4387 2596 4853 2604
rect 5607 2596 5793 2604
rect 6127 2596 6413 2604
rect 67 2576 393 2584
rect 407 2576 1333 2584
rect 2467 2576 2613 2584
rect 3007 2576 3133 2584
rect 3227 2576 3413 2584
rect 4067 2576 4213 2584
rect 4487 2576 5313 2584
rect 5327 2576 5473 2584
rect 5487 2576 5513 2584
rect 6087 2576 6333 2584
rect 587 2556 793 2564
rect 1107 2556 1773 2564
rect 1787 2556 2753 2564
rect 3447 2556 3973 2564
rect 4607 2556 5413 2564
rect 5587 2556 5833 2564
rect 5847 2556 6053 2564
rect 6667 2564 6680 2567
rect 6667 2553 6684 2564
rect 267 2536 333 2544
rect 1047 2536 2513 2544
rect 3167 2536 3413 2544
rect 4187 2536 4353 2544
rect 4367 2536 4513 2544
rect 5787 2536 6213 2544
rect 6227 2536 6653 2544
rect -24 2516 53 2524
rect -24 2476 -16 2516
rect 387 2516 473 2524
rect 487 2516 673 2524
rect 1287 2516 2073 2524
rect 3687 2516 4073 2524
rect 4087 2516 4133 2524
rect 4587 2516 4613 2524
rect 4707 2516 4953 2524
rect 4967 2516 5173 2524
rect 5287 2516 5473 2524
rect 6067 2516 6173 2524
rect 6307 2516 6473 2524
rect 3227 2504 3240 2507
rect 3227 2493 3244 2504
rect 3527 2496 3693 2504
rect 4027 2496 4153 2504
rect 4416 2496 4553 2504
rect 67 2476 153 2484
rect 547 2477 693 2485
rect 847 2477 1013 2485
rect 207 2436 273 2444
rect 296 2444 304 2474
rect 1027 2477 1073 2485
rect 1087 2476 1173 2484
rect 1227 2476 1273 2484
rect 1347 2477 1393 2485
rect 1527 2477 1593 2485
rect 1647 2477 1713 2485
rect 1907 2476 1953 2484
rect 2027 2476 2233 2484
rect 2327 2477 2352 2485
rect 2387 2477 2573 2485
rect 2667 2477 2713 2485
rect 2276 2464 2284 2474
rect 2276 2456 2404 2464
rect 296 2436 413 2444
rect 607 2436 933 2444
rect 947 2435 1013 2443
rect 1567 2436 1613 2444
rect 2147 2436 2373 2444
rect 2396 2444 2404 2456
rect 2396 2436 2473 2444
rect 2616 2444 2624 2474
rect 2756 2464 2764 2474
rect 2756 2456 2784 2464
rect 2776 2447 2784 2456
rect 2616 2436 2693 2444
rect 2776 2436 2793 2447
rect 2780 2433 2793 2436
rect 667 2416 924 2424
rect 916 2407 924 2416
rect 2307 2416 2333 2424
rect 2407 2416 2433 2424
rect 2607 2416 2653 2424
rect 2876 2424 2884 2474
rect 2967 2484 2980 2487
rect 2967 2473 2984 2484
rect 2976 2444 2984 2473
rect 2976 2436 3053 2444
rect 3067 2436 3093 2444
rect 3236 2427 3244 2493
rect 3287 2476 3333 2484
rect 3347 2476 3433 2484
rect 3727 2477 3813 2485
rect 4096 2476 4393 2484
rect 3536 2444 3544 2473
rect 3627 2456 3753 2464
rect 4096 2464 4104 2476
rect 4416 2484 4424 2496
rect 5716 2496 5773 2504
rect 4407 2476 4424 2484
rect 4487 2476 4973 2484
rect 5367 2477 5453 2485
rect 5016 2464 5024 2474
rect 4076 2456 4104 2464
rect 4816 2460 5084 2464
rect 4813 2456 5087 2460
rect 3427 2436 3544 2444
rect 4076 2446 4084 2456
rect 4813 2447 4827 2456
rect 3987 2436 4073 2444
rect 4147 2435 4193 2443
rect 4727 2435 4773 2443
rect 5073 2447 5087 2456
rect 5127 2435 5273 2443
rect 5287 2435 5333 2443
rect 5447 2435 5493 2443
rect 5676 2444 5684 2474
rect 5627 2436 5684 2444
rect 5716 2444 5724 2496
rect 5827 2496 5964 2504
rect 5956 2484 5964 2496
rect 5987 2496 6024 2504
rect 5956 2476 5993 2484
rect 5707 2436 5724 2444
rect 2767 2416 2884 2424
rect 3227 2416 3244 2427
rect 3227 2413 3240 2416
rect 3567 2416 3652 2424
rect 3687 2416 3793 2424
rect 3887 2416 3953 2424
rect 3967 2416 4053 2424
rect 4487 2416 4553 2424
rect 4967 2420 5004 2424
rect 4967 2416 5007 2420
rect 707 2396 773 2404
rect 927 2396 973 2404
rect 3047 2396 3153 2404
rect 3676 2404 3684 2413
rect 4993 2407 5007 2416
rect 5736 2424 5744 2473
rect 6016 2446 6024 2496
rect 6676 2504 6684 2553
rect 6676 2496 6724 2504
rect 6196 2476 6293 2484
rect 6196 2447 6204 2476
rect 6476 2464 6484 2474
rect 6636 2464 6644 2493
rect 6436 2460 6484 2464
rect 6536 2460 6644 2464
rect 6433 2456 6484 2460
rect 6533 2456 6644 2460
rect 6433 2447 6447 2456
rect 6027 2436 6113 2444
rect 6533 2447 6547 2456
rect 6676 2447 6684 2473
rect 5547 2416 5744 2424
rect 5787 2416 5913 2424
rect 6227 2416 6313 2424
rect 6427 2416 6493 2424
rect 6647 2416 6693 2424
rect 6716 2407 6724 2496
rect 3467 2396 3684 2404
rect 3907 2396 3953 2404
rect 4367 2396 4393 2404
rect 4636 2396 4813 2404
rect 2247 2376 2684 2384
rect 507 2356 733 2364
rect 1187 2356 1433 2364
rect 2147 2356 2593 2364
rect 2676 2364 2684 2376
rect 2707 2376 2773 2384
rect 2787 2376 3693 2384
rect 3707 2376 4013 2384
rect 4027 2376 4093 2384
rect 4107 2376 4513 2384
rect 4636 2384 4644 2396
rect 5047 2396 5753 2404
rect 6087 2396 6153 2404
rect 6700 2406 6724 2407
rect 6707 2396 6724 2406
rect 6707 2393 6720 2396
rect 4576 2376 4644 2384
rect 2676 2356 2733 2364
rect 2907 2356 3153 2364
rect 3527 2356 3593 2364
rect 4067 2356 4353 2364
rect 4576 2364 4584 2376
rect 4707 2376 4753 2384
rect 4887 2376 5113 2384
rect 5227 2376 5613 2384
rect 5627 2376 5873 2384
rect 6007 2376 6053 2384
rect 4427 2356 4584 2364
rect 4607 2356 4633 2364
rect 4787 2356 5133 2364
rect 5207 2356 5344 2364
rect 47 2336 173 2344
rect 2207 2336 2373 2344
rect 3187 2336 3293 2344
rect 3367 2336 3413 2344
rect 3707 2336 4673 2344
rect 5336 2344 5344 2356
rect 5387 2356 5653 2364
rect 5667 2356 5813 2364
rect 6327 2356 6393 2364
rect 5336 2336 5813 2344
rect 5907 2336 6113 2344
rect 6307 2336 6373 2344
rect 6387 2336 6573 2344
rect 356 2316 773 2324
rect 356 2307 364 2316
rect 2627 2316 3093 2324
rect 3436 2316 3613 2324
rect 47 2296 113 2304
rect 287 2296 353 2304
rect 427 2296 573 2304
rect 1267 2296 1333 2304
rect 1927 2296 1973 2304
rect 2187 2296 2393 2304
rect 2407 2296 2533 2304
rect 3436 2304 3444 2316
rect 4147 2316 4304 2324
rect 3087 2296 3444 2304
rect 4296 2304 4304 2316
rect 4327 2316 4593 2324
rect 4927 2316 5033 2324
rect 5047 2316 5233 2324
rect 5587 2316 5733 2324
rect 6367 2316 6613 2324
rect 4296 2296 4373 2304
rect 4387 2296 4533 2304
rect 4627 2296 4853 2304
rect 5427 2296 5773 2304
rect 5847 2296 6013 2304
rect 6107 2296 6313 2304
rect 6447 2296 6653 2304
rect 307 2276 373 2284
rect 767 2276 1093 2284
rect 2527 2276 2613 2284
rect 2996 2276 3173 2284
rect 2996 2268 3004 2276
rect 3507 2276 3533 2284
rect 3607 2276 3633 2284
rect 3776 2276 3973 2284
rect 127 2256 473 2264
rect 587 2256 724 2264
rect -24 2216 33 2224
rect 716 2226 724 2256
rect 847 2256 953 2264
rect 967 2257 1013 2265
rect 1147 2256 1573 2264
rect 1587 2256 1633 2264
rect 1927 2257 1953 2265
rect 2047 2256 2093 2264
rect 1876 2244 1884 2254
rect 2227 2256 2344 2264
rect 1876 2236 1944 2244
rect 36 2204 44 2213
rect 147 2216 233 2224
rect 247 2216 324 2224
rect 36 2196 93 2204
rect 316 2204 324 2216
rect 487 2215 553 2223
rect 1027 2216 1113 2224
rect 1187 2215 1273 2223
rect 1347 2215 1373 2223
rect 1607 2215 1673 2223
rect 1936 2224 1944 2236
rect 2336 2226 2344 2256
rect 2887 2257 2993 2265
rect 2356 2227 2364 2253
rect 1936 2216 2053 2224
rect 2107 2215 2193 2223
rect 2456 2224 2464 2254
rect 3107 2256 3593 2264
rect 3776 2244 3784 2276
rect 4047 2276 4173 2284
rect 4547 2276 4573 2284
rect 4647 2276 4673 2284
rect 4947 2276 4973 2284
rect 5287 2276 5353 2284
rect 5827 2276 6153 2284
rect 3807 2256 4244 2264
rect 4236 2244 4244 2256
rect 4267 2256 4353 2264
rect 4427 2256 4453 2264
rect 4507 2257 4613 2265
rect 5127 2256 5153 2264
rect 5247 2256 5384 2264
rect 3776 2236 3824 2244
rect 4236 2236 4304 2244
rect 2456 2216 2573 2224
rect 2787 2216 2913 2224
rect 2927 2216 2944 2224
rect 2987 2215 3053 2223
rect 3227 2216 3333 2224
rect 3816 2226 3824 2236
rect 3547 2216 3633 2224
rect 3927 2215 4053 2223
rect 4296 2226 4304 2236
rect 4576 2236 4713 2244
rect 4127 2216 4193 2224
rect 4576 2224 4584 2236
rect 4727 2236 4924 2244
rect 4387 2216 4584 2224
rect 4727 2215 4793 2223
rect 4916 2224 4924 2236
rect 5016 2227 5024 2253
rect 5376 2244 5384 2256
rect 5407 2256 5473 2264
rect 5547 2256 5604 2264
rect 5376 2236 5524 2244
rect 4916 2216 4933 2224
rect 5516 2226 5524 2236
rect 5596 2227 5604 2256
rect 5627 2257 5693 2265
rect 5927 2256 5973 2264
rect 6067 2256 6193 2264
rect 5147 2215 5173 2223
rect 5187 2216 5373 2224
rect 5827 2215 5853 2223
rect 6056 2224 6064 2254
rect 6320 2264 6333 2267
rect 6316 2253 6333 2264
rect 6387 2256 6413 2264
rect 6467 2256 6493 2264
rect 6056 2216 6173 2224
rect 6227 2216 6253 2224
rect 6316 2226 6324 2253
rect 6367 2215 6433 2223
rect 6527 2216 6633 2224
rect 316 2196 433 2204
rect 1087 2196 1473 2204
rect 1736 2196 2013 2204
rect 1736 2187 1744 2196
rect 2627 2196 2693 2204
rect 4467 2196 4493 2204
rect 4647 2196 4693 2204
rect 4707 2196 4753 2204
rect 5647 2196 5693 2204
rect 5907 2196 5953 2204
rect 347 2176 393 2184
rect 507 2176 572 2184
rect 607 2176 973 2184
rect 1647 2176 1733 2184
rect 1847 2176 1973 2184
rect 1987 2176 2053 2184
rect 2067 2176 2273 2184
rect 2287 2176 2552 2184
rect 2587 2176 2733 2184
rect 3327 2176 3433 2184
rect 3447 2176 3593 2184
rect 3607 2176 3853 2184
rect 4207 2176 4293 2184
rect 4487 2176 4553 2184
rect 4567 2176 4793 2184
rect 4847 2176 4893 2184
rect 5227 2176 5513 2184
rect 6047 2176 6293 2184
rect 1427 2156 1953 2164
rect 2147 2156 2233 2164
rect 2507 2156 2713 2164
rect 2727 2156 2773 2164
rect 2827 2156 3753 2164
rect 3967 2156 4033 2164
rect 4167 2156 4373 2164
rect 4567 2156 4653 2164
rect 4927 2156 5113 2164
rect 6247 2156 6273 2164
rect 587 2136 2124 2144
rect 987 2116 1853 2124
rect 2116 2124 2124 2136
rect 2236 2136 2453 2144
rect 2236 2124 2244 2136
rect 3007 2136 3693 2144
rect 4407 2136 4653 2144
rect 5067 2136 5273 2144
rect 5527 2136 5553 2144
rect 5987 2136 6213 2144
rect 6227 2136 6573 2144
rect 2116 2116 2244 2124
rect 2256 2116 2493 2124
rect 187 2096 433 2104
rect 447 2096 653 2104
rect 2256 2104 2264 2116
rect 3127 2116 3393 2124
rect 4027 2116 4133 2124
rect 4587 2116 4853 2124
rect 1947 2096 2264 2104
rect 2327 2096 2993 2104
rect 3147 2096 3513 2104
rect 3587 2096 3673 2104
rect 3767 2096 4113 2104
rect 4847 2096 5013 2104
rect 5287 2096 5573 2104
rect 196 2076 1233 2084
rect 196 2064 204 2076
rect 1907 2076 2424 2084
rect 87 2056 204 2064
rect 2247 2056 2293 2064
rect 2307 2056 2393 2064
rect 2416 2064 2424 2076
rect 2467 2076 3113 2084
rect 3487 2076 3773 2084
rect 3787 2076 3873 2084
rect 4327 2076 4473 2084
rect 4547 2076 5033 2084
rect 5047 2076 5093 2084
rect 5107 2076 5633 2084
rect 6487 2076 6653 2084
rect 3476 2064 3484 2073
rect 2416 2056 3484 2064
rect 3647 2056 3713 2064
rect 4067 2056 4193 2064
rect 4247 2056 4833 2064
rect 4927 2056 4973 2064
rect 5347 2056 5453 2064
rect 5467 2056 5613 2064
rect 607 2036 1893 2044
rect 3027 2036 3153 2044
rect 3487 2036 3533 2044
rect 4007 2036 4053 2044
rect 4627 2036 5073 2044
rect 5487 2036 5833 2044
rect 6127 2036 6433 2044
rect 787 2016 1053 2024
rect 1187 2016 1793 2024
rect 3247 2016 3353 2024
rect 3867 2016 3973 2024
rect 4087 2016 4313 2024
rect 6147 2016 6413 2024
rect 6627 2016 6673 2024
rect -24 1996 53 2004
rect 67 1996 93 2004
rect 647 1996 1033 2004
rect 2947 1996 3013 2004
rect 3407 1996 3624 2004
rect 1967 1976 2313 1984
rect 3387 1976 3493 1984
rect 3616 1984 3624 1996
rect 3896 1996 3993 2004
rect 3896 1984 3904 1996
rect 4067 1996 4153 2004
rect 4227 1996 4593 2004
rect 4667 1996 4693 2004
rect 4707 1996 5373 2004
rect 5607 1996 5873 2004
rect 5887 1996 5973 2004
rect 6047 1996 6333 2004
rect 6387 1996 6433 2004
rect 3616 1976 3904 1984
rect 4487 1976 4653 1984
rect -24 1956 73 1964
rect 247 1957 293 1965
rect 867 1956 953 1964
rect 967 1956 1093 1964
rect 1147 1957 1233 1965
rect 1547 1957 1633 1965
rect 1707 1957 1733 1965
rect 1776 1956 1893 1964
rect 427 1916 453 1924
rect 467 1915 493 1923
rect 727 1915 753 1923
rect 767 1915 833 1923
rect 1447 1915 1493 1923
rect 1627 1916 1673 1924
rect 1776 1924 1784 1956
rect 2107 1957 2153 1965
rect 2347 1956 2364 1964
rect 2136 1936 2233 1944
rect 2136 1926 2144 1936
rect 1767 1916 1784 1924
rect 2267 1916 2313 1924
rect 2356 1924 2364 1956
rect 2376 1944 2384 1973
rect 4767 1976 4853 1984
rect 4927 1976 5253 1984
rect 6427 1976 6553 1984
rect 2447 1957 2493 1965
rect 2567 1956 2613 1964
rect 2687 1956 2864 1964
rect 2856 1944 2864 1956
rect 2887 1957 2913 1965
rect 2967 1956 3073 1964
rect 3256 1956 3333 1964
rect 2376 1936 2404 1944
rect 2856 1936 2904 1944
rect 2356 1916 2373 1924
rect 2396 1924 2404 1936
rect 2396 1916 2473 1924
rect 2896 1924 2904 1936
rect 3256 1926 3264 1956
rect 4036 1956 4133 1964
rect 3316 1936 3384 1944
rect 3316 1927 3324 1936
rect 2896 1916 2933 1924
rect 3147 1915 3213 1923
rect 3307 1916 3324 1927
rect 3376 1926 3384 1936
rect 3687 1936 3853 1944
rect 3916 1944 3924 1954
rect 4036 1944 4044 1956
rect 4267 1956 4413 1964
rect 4496 1956 4613 1964
rect 3916 1936 4044 1944
rect 3307 1913 3320 1916
rect 3387 1916 3413 1924
rect 3747 1916 3793 1924
rect 4196 1924 4204 1953
rect 4196 1916 4313 1924
rect 1487 1896 1553 1904
rect 2807 1896 2833 1904
rect 2847 1896 3093 1904
rect 3407 1896 3633 1904
rect 4456 1904 4464 1953
rect 4496 1926 4504 1956
rect 4747 1957 4813 1965
rect 5027 1956 5173 1964
rect 5427 1956 5573 1964
rect 5847 1956 5953 1964
rect 4567 1916 4593 1924
rect 4687 1916 4793 1924
rect 4936 1924 4944 1953
rect 5216 1944 5224 1954
rect 6127 1957 6173 1965
rect 6387 1956 6493 1964
rect 6216 1944 6224 1954
rect 5027 1936 5224 1944
rect 5336 1936 5404 1944
rect 6216 1936 6304 1944
rect 4936 1916 4953 1924
rect 5336 1924 5344 1936
rect 5247 1916 5344 1924
rect 5396 1924 5404 1936
rect 5396 1916 5533 1924
rect 5547 1916 5713 1924
rect 5967 1915 6013 1923
rect 6207 1916 6273 1924
rect 6296 1924 6304 1936
rect 6636 1926 6644 1973
rect 6296 1916 6313 1924
rect 6327 1915 6513 1923
rect 4307 1896 4464 1904
rect 5407 1896 5453 1904
rect 6567 1896 6653 1904
rect 847 1876 913 1884
rect 927 1876 973 1884
rect 1167 1876 1693 1884
rect 2187 1876 2433 1884
rect 2567 1876 2873 1884
rect 2987 1876 3013 1884
rect 4167 1876 4204 1884
rect 367 1856 533 1864
rect 547 1856 613 1864
rect 1067 1856 1153 1864
rect 1447 1856 1533 1864
rect 1767 1856 1933 1864
rect 2247 1856 2313 1864
rect 2627 1856 2813 1864
rect 2907 1856 3393 1864
rect 3627 1856 3693 1864
rect 3787 1856 4013 1864
rect 4027 1856 4093 1864
rect 4196 1864 4204 1876
rect 4487 1876 4573 1884
rect 4647 1876 4733 1884
rect 4787 1876 4813 1884
rect 4827 1876 4893 1884
rect 4907 1876 5013 1884
rect 5147 1876 5353 1884
rect 5947 1876 6013 1884
rect 6567 1876 6673 1884
rect 4196 1856 4393 1864
rect 4767 1856 5113 1864
rect 5167 1856 5333 1864
rect 6467 1856 6513 1864
rect 27 1836 633 1844
rect 1887 1836 2013 1844
rect 2167 1836 2393 1844
rect 2487 1836 3513 1844
rect 3607 1836 3704 1844
rect 3696 1827 3704 1836
rect 3747 1836 3832 1844
rect 3867 1836 4113 1844
rect 4587 1836 5133 1844
rect 5867 1836 6153 1844
rect 6276 1836 6313 1844
rect 287 1816 453 1824
rect 1067 1816 1793 1824
rect 1807 1816 2293 1824
rect 2647 1816 2853 1824
rect 2976 1816 3113 1824
rect 2976 1807 2984 1816
rect 3367 1816 3493 1824
rect 3696 1816 3713 1827
rect 3700 1813 3713 1816
rect 4327 1816 4533 1824
rect 4607 1816 4693 1824
rect 6276 1824 6284 1836
rect 6387 1836 6433 1844
rect 6647 1836 6733 1844
rect 5987 1816 6284 1824
rect 427 1796 653 1804
rect 807 1796 1293 1804
rect 1307 1796 1353 1804
rect 1367 1796 1393 1804
rect 1927 1796 1953 1804
rect 2127 1796 2273 1804
rect 2467 1796 2613 1804
rect 2967 1796 2984 1807
rect 2967 1793 2980 1796
rect 3207 1796 3253 1804
rect 3427 1796 3473 1804
rect 3487 1796 3593 1804
rect 4167 1796 4353 1804
rect 4407 1796 4833 1804
rect 6107 1796 6193 1804
rect 6447 1796 6593 1804
rect 6607 1796 6673 1804
rect 827 1776 992 1784
rect 1027 1776 1273 1784
rect 2867 1776 2933 1784
rect 3347 1776 3613 1784
rect 3727 1776 3773 1784
rect 3907 1776 3933 1784
rect 5187 1776 5253 1784
rect 5267 1776 5453 1784
rect 5867 1776 5973 1784
rect 127 1756 213 1764
rect 327 1756 413 1764
rect 1527 1756 1673 1764
rect 2067 1756 2173 1764
rect 2627 1756 2713 1764
rect 3047 1756 3173 1764
rect 3527 1756 3573 1764
rect 3827 1756 3873 1764
rect 3987 1756 4033 1764
rect 4927 1756 5093 1764
rect 6307 1756 6333 1764
rect 6547 1756 6573 1764
rect 6613 1764 6627 1773
rect 6613 1760 6773 1764
rect 6616 1756 6773 1760
rect 356 1736 433 1744
rect 356 1706 364 1736
rect 707 1737 753 1745
rect 856 1736 893 1744
rect 536 1707 544 1734
rect -24 1696 93 1704
rect 536 1696 553 1707
rect 540 1693 553 1696
rect 727 1695 773 1703
rect 816 1687 824 1734
rect 856 1704 864 1736
rect 1287 1736 1333 1744
rect 1587 1737 1613 1745
rect 1827 1736 1884 1744
rect 1876 1724 1884 1736
rect 1907 1737 1953 1745
rect 2007 1736 2124 1744
rect 1876 1716 1984 1724
rect 847 1696 864 1704
rect 887 1695 933 1703
rect 987 1695 1073 1703
rect 1307 1696 1413 1704
rect 1976 1706 1984 1716
rect 2116 1706 2124 1736
rect 2247 1737 2333 1745
rect 2347 1736 2493 1744
rect 2707 1736 2793 1744
rect 2816 1736 2893 1744
rect 2816 1724 2824 1736
rect 3027 1736 3153 1744
rect 3267 1737 3333 1745
rect 3467 1736 3493 1744
rect 3647 1736 3753 1744
rect 3967 1736 4013 1744
rect 4067 1736 4093 1744
rect 4427 1736 4453 1744
rect 2787 1716 2824 1724
rect 3807 1716 3904 1724
rect 1507 1696 1553 1704
rect 1767 1695 1833 1703
rect 2327 1695 2413 1703
rect 2507 1695 2533 1703
rect 2587 1695 2613 1703
rect 2807 1695 2833 1703
rect 3087 1695 3273 1703
rect 3287 1695 3313 1703
rect 3447 1696 3513 1704
rect 3607 1696 3733 1704
rect 3827 1695 3873 1703
rect 3896 1704 3904 1716
rect 4656 1724 4664 1734
rect 4787 1737 4833 1745
rect 5207 1736 5393 1744
rect 5567 1736 5593 1744
rect 5647 1736 5773 1744
rect 5827 1736 5933 1744
rect 4147 1720 4684 1724
rect 4147 1716 4687 1720
rect 4673 1707 4687 1716
rect 3896 1696 3913 1704
rect 3927 1696 4033 1704
rect 4127 1696 4413 1704
rect 4527 1695 4573 1703
rect 4736 1704 4744 1733
rect 5456 1716 5533 1724
rect 4736 1696 4753 1704
rect 4947 1695 4973 1703
rect 5047 1696 5173 1704
rect 5227 1695 5253 1703
rect 5456 1704 5464 1716
rect 5836 1707 5844 1736
rect 5947 1736 6093 1744
rect 6187 1736 6253 1744
rect 6393 1744 6407 1753
rect 6393 1740 6473 1744
rect 6396 1736 6473 1740
rect 6616 1736 6713 1744
rect 6556 1707 6564 1733
rect 5367 1696 5464 1704
rect 6287 1696 6373 1704
rect 6387 1695 6453 1703
rect 6616 1706 6624 1736
rect 227 1676 253 1684
rect 427 1676 453 1684
rect 587 1676 653 1684
rect 1027 1676 1113 1684
rect 1467 1676 1613 1684
rect 2067 1676 2173 1684
rect 2347 1676 2373 1684
rect 2907 1676 2953 1684
rect 3096 1676 3132 1684
rect 2027 1656 2153 1664
rect 2527 1656 2633 1664
rect 2656 1656 2792 1664
rect 1187 1636 1753 1644
rect 2656 1644 2664 1656
rect 2827 1656 2853 1664
rect 3096 1664 3104 1676
rect 3167 1676 3193 1684
rect 3627 1676 3813 1684
rect 4447 1676 4513 1684
rect 4727 1676 4873 1684
rect 5487 1676 5613 1684
rect 5627 1676 5753 1684
rect 5927 1676 6113 1684
rect 2947 1656 3104 1664
rect 3367 1656 3393 1664
rect 3527 1656 3793 1664
rect 4067 1656 4273 1664
rect 4287 1656 4353 1664
rect 4467 1656 4653 1664
rect 4747 1656 5073 1664
rect 5547 1656 5653 1664
rect 2307 1636 2664 1644
rect 2727 1636 2873 1644
rect 2887 1636 2993 1644
rect 3007 1636 3172 1644
rect 3207 1636 3413 1644
rect 4427 1636 5133 1644
rect 167 1616 753 1624
rect 1887 1616 2944 1624
rect 947 1596 1384 1604
rect 687 1576 1053 1584
rect 1376 1584 1384 1596
rect 2207 1596 2273 1604
rect 2316 1596 2673 1604
rect 1376 1576 1873 1584
rect 2316 1584 2324 1596
rect 2787 1596 2833 1604
rect 2936 1604 2944 1616
rect 2987 1616 3153 1624
rect 3567 1616 3872 1624
rect 3907 1616 4033 1624
rect 4087 1616 4473 1624
rect 4516 1616 4953 1624
rect 2936 1596 2993 1604
rect 3047 1596 3093 1604
rect 3156 1604 3164 1613
rect 4516 1607 4524 1616
rect 5087 1616 5293 1624
rect 5407 1616 5893 1624
rect 5907 1616 5953 1624
rect 5967 1616 6073 1624
rect 6607 1616 6673 1624
rect 3156 1596 3373 1604
rect 3427 1596 3773 1604
rect 3827 1596 4053 1604
rect 4367 1596 4393 1604
rect 4507 1596 4524 1607
rect 4507 1593 4520 1596
rect 4667 1596 5353 1604
rect 6027 1596 6273 1604
rect 6387 1596 6533 1604
rect 6587 1596 6613 1604
rect 2187 1576 2324 1584
rect 2347 1576 3313 1584
rect 3376 1584 3384 1593
rect 3376 1576 3613 1584
rect 3707 1576 3793 1584
rect 3847 1576 4264 1584
rect 527 1556 613 1564
rect 627 1556 753 1564
rect 1747 1556 1793 1564
rect 2027 1556 3073 1564
rect 3356 1556 3653 1564
rect 3356 1547 3364 1556
rect 3667 1556 4233 1564
rect 4256 1564 4264 1576
rect 4707 1576 4753 1584
rect 6527 1576 6773 1584
rect 4256 1556 4573 1564
rect 4636 1556 4853 1564
rect 4636 1547 4644 1556
rect 4987 1556 5433 1564
rect 5727 1556 5853 1564
rect 6087 1556 6353 1564
rect 6447 1556 6693 1564
rect 1587 1536 3353 1544
rect 3447 1536 3553 1544
rect 3727 1536 3933 1544
rect 3947 1536 3973 1544
rect 3996 1536 4133 1544
rect 1087 1516 1533 1524
rect 1547 1516 2292 1524
rect 2327 1516 2713 1524
rect 2807 1516 3193 1524
rect 3996 1524 4004 1536
rect 4207 1536 4633 1544
rect 5627 1536 6033 1544
rect 3627 1516 4004 1524
rect 4347 1516 4453 1524
rect 4467 1516 4533 1524
rect 5467 1516 5553 1524
rect 6247 1516 6493 1524
rect 6507 1516 6673 1524
rect 47 1496 173 1504
rect 187 1496 373 1504
rect 547 1496 1213 1504
rect 2296 1504 2304 1513
rect 1947 1496 2004 1504
rect 2296 1496 3293 1504
rect 1787 1476 1973 1484
rect 1996 1484 2004 1496
rect 3647 1496 3693 1504
rect 3807 1496 3893 1504
rect 4007 1496 4233 1504
rect 4287 1496 4652 1504
rect 4687 1496 4813 1504
rect 5056 1496 5313 1504
rect 1996 1476 2413 1484
rect 3007 1476 3253 1484
rect 3327 1476 3433 1484
rect 3596 1476 3713 1484
rect 227 1456 533 1464
rect 847 1456 913 1464
rect 1647 1456 1693 1464
rect 1707 1456 1833 1464
rect 2087 1456 2613 1464
rect 3596 1464 3604 1476
rect 3787 1476 3953 1484
rect 5056 1484 5064 1496
rect 5327 1496 5593 1504
rect 5607 1496 5913 1504
rect 5987 1496 6193 1504
rect 6547 1496 6653 1504
rect 4147 1476 5064 1484
rect 5427 1476 5693 1484
rect 6067 1476 6093 1484
rect 6107 1476 6173 1484
rect 6247 1476 6333 1484
rect 3307 1456 3604 1464
rect 3796 1456 3913 1464
rect -24 1436 13 1444
rect 287 1436 293 1444
rect 307 1436 413 1444
rect 507 1437 553 1445
rect 667 1436 713 1444
rect 987 1436 1053 1444
rect 1107 1437 1173 1445
rect 1227 1436 1493 1444
rect 1507 1436 1573 1444
rect 1687 1436 1873 1444
rect 2116 1436 2133 1444
rect 1876 1424 1884 1434
rect 1876 1416 1964 1424
rect 27 1395 93 1403
rect 1047 1396 1093 1404
rect 1107 1396 1193 1404
rect 1407 1396 1453 1404
rect 1467 1396 1513 1404
rect 1607 1395 1653 1403
rect 1827 1396 1913 1404
rect 1956 1404 1964 1416
rect 1956 1396 1993 1404
rect 267 1376 353 1384
rect 367 1376 493 1384
rect 747 1376 833 1384
rect 1947 1376 2033 1384
rect 2116 1384 2124 1436
rect 2487 1436 2533 1444
rect 2887 1437 2933 1445
rect 3207 1437 3273 1445
rect 3467 1436 3613 1444
rect 2676 1407 2684 1434
rect 3136 1407 3144 1434
rect 2167 1396 2193 1404
rect 2307 1395 2393 1403
rect 2527 1396 2573 1404
rect 2676 1396 2693 1407
rect 2680 1393 2693 1396
rect 2907 1396 2953 1404
rect 3127 1396 3144 1407
rect 3127 1393 3140 1396
rect 3387 1396 3413 1404
rect 2087 1376 2124 1384
rect 2507 1376 2793 1384
rect 2807 1376 2873 1384
rect 3656 1384 3664 1434
rect 3796 1444 3804 1456
rect 3987 1456 4073 1464
rect 4187 1456 4293 1464
rect 4747 1456 4824 1464
rect 3747 1436 3804 1444
rect 4047 1437 4113 1445
rect 3707 1416 3784 1424
rect 3776 1404 3784 1416
rect 4193 1424 4207 1433
rect 3887 1420 4207 1424
rect 4276 1436 4413 1444
rect 3887 1416 4204 1420
rect 4053 1407 4067 1416
rect 3776 1396 3793 1404
rect 4276 1404 4284 1436
rect 4607 1436 4693 1444
rect 4816 1444 4824 1456
rect 4967 1456 5073 1464
rect 6667 1456 6713 1464
rect 4816 1436 4913 1444
rect 4927 1436 5013 1444
rect 5107 1436 5193 1444
rect 5567 1436 5673 1444
rect 5687 1436 5793 1444
rect 6027 1436 6153 1444
rect 6207 1437 6253 1445
rect 6387 1436 6404 1444
rect 5816 1416 5893 1424
rect 5816 1406 5824 1416
rect 4267 1396 4284 1404
rect 4447 1396 4613 1404
rect 6007 1395 6053 1403
rect 6156 1404 6164 1434
rect 6396 1424 6404 1436
rect 6447 1437 6493 1445
rect 6396 1416 6424 1424
rect 6156 1396 6313 1404
rect 6416 1404 6424 1416
rect 6416 1396 6513 1404
rect 6667 1396 6753 1404
rect 3347 1376 3664 1384
rect 4107 1376 4333 1384
rect 4416 1376 4493 1384
rect 167 1356 393 1364
rect 1707 1356 1733 1364
rect 3247 1356 3653 1364
rect 3807 1356 4313 1364
rect 4416 1364 4424 1376
rect 4787 1376 5153 1384
rect 5387 1376 5464 1384
rect 5456 1367 5464 1376
rect 6107 1376 6173 1384
rect 6587 1376 6693 1384
rect 4387 1356 4424 1364
rect 4467 1356 4673 1364
rect 4847 1356 4973 1364
rect 5067 1356 5133 1364
rect 5467 1356 5493 1364
rect 5787 1356 5913 1364
rect 1767 1336 2253 1344
rect 3467 1336 3513 1344
rect 4836 1344 4844 1353
rect 4367 1336 4844 1344
rect 5027 1336 5113 1344
rect 5127 1336 5373 1344
rect 5687 1336 6073 1344
rect 6167 1336 6273 1344
rect 6367 1336 6573 1344
rect 507 1316 573 1324
rect 787 1316 953 1324
rect 1527 1316 1693 1324
rect 2747 1316 2773 1324
rect 2867 1316 3013 1324
rect 3087 1316 3673 1324
rect 4007 1316 4033 1324
rect 4407 1316 4633 1324
rect 5227 1316 5273 1324
rect 6447 1316 6533 1324
rect 487 1296 613 1304
rect 627 1296 1833 1304
rect 2027 1296 2073 1304
rect 3127 1296 3173 1304
rect 3667 1296 3793 1304
rect 3847 1296 4133 1304
rect 4667 1296 4693 1304
rect 5607 1296 5833 1304
rect 5887 1296 5933 1304
rect 6287 1296 6433 1304
rect 687 1276 873 1284
rect 1167 1276 1253 1284
rect 1267 1276 1353 1284
rect 1587 1276 1672 1284
rect 2016 1284 2024 1293
rect 1707 1276 2024 1284
rect 2247 1276 2293 1284
rect 2416 1276 3073 1284
rect 2416 1267 2424 1276
rect 3087 1276 3213 1284
rect 4187 1276 4333 1284
rect 4407 1276 4953 1284
rect 6087 1276 6133 1284
rect 6267 1276 6584 1284
rect 6576 1267 6584 1276
rect 576 1256 793 1264
rect 576 1247 584 1256
rect 807 1256 913 1264
rect 1007 1256 1073 1264
rect 1127 1256 1873 1264
rect 1887 1256 2053 1264
rect 2067 1256 2413 1264
rect 2467 1256 2833 1264
rect 3567 1256 3593 1264
rect 3607 1256 3733 1264
rect 3856 1256 3913 1264
rect 407 1236 573 1244
rect 1607 1236 1853 1244
rect 2087 1236 2333 1244
rect 3856 1244 3864 1256
rect 4287 1256 4353 1264
rect 4527 1256 4693 1264
rect 5047 1256 5133 1264
rect 5567 1256 5773 1264
rect 6027 1256 6193 1264
rect 6307 1256 6373 1264
rect 6576 1256 6593 1267
rect 6580 1253 6593 1256
rect 3767 1236 3864 1244
rect 4347 1236 4453 1244
rect 5547 1236 5673 1244
rect 5887 1236 5972 1244
rect 6007 1236 6253 1244
rect 127 1216 193 1224
rect 287 1216 384 1224
rect -24 1176 93 1184
rect 107 1176 213 1184
rect 227 1175 253 1183
rect 376 1184 384 1216
rect 627 1216 644 1224
rect 636 1187 644 1216
rect 787 1217 853 1225
rect 907 1216 993 1224
rect 376 1176 413 1184
rect 467 1175 493 1183
rect 716 1164 724 1214
rect 1047 1216 1104 1224
rect 1096 1204 1104 1216
rect 1147 1217 1313 1225
rect 1407 1216 1473 1224
rect 1947 1216 1993 1224
rect 2067 1216 2224 1224
rect 1096 1196 1233 1204
rect 2216 1186 2224 1216
rect 2567 1216 2613 1224
rect 927 1175 973 1183
rect 987 1176 1053 1184
rect 1187 1176 1293 1184
rect 1507 1176 1633 1184
rect 1887 1175 1913 1183
rect 2027 1175 2073 1183
rect 2276 1184 2284 1213
rect 2267 1176 2284 1184
rect 2376 1184 2384 1214
rect 2747 1216 2792 1224
rect 2827 1216 2873 1224
rect 3027 1216 3113 1224
rect 3327 1216 3493 1224
rect 3716 1204 3724 1214
rect 3847 1216 3873 1224
rect 4033 1224 4047 1233
rect 4033 1220 4093 1224
rect 4036 1216 4093 1220
rect 4327 1217 4373 1225
rect 4547 1217 4573 1225
rect 4747 1216 4764 1224
rect 4236 1204 4244 1214
rect 3196 1196 4493 1204
rect 2347 1176 2384 1184
rect 2407 1175 2453 1183
rect 3196 1186 3204 1196
rect 2507 1176 2533 1184
rect 2587 1176 2804 1184
rect 2796 1167 2804 1176
rect 3127 1175 3153 1183
rect 3447 1175 3533 1183
rect 3947 1175 3973 1183
rect 4387 1176 4653 1184
rect 4667 1175 4713 1183
rect 716 1156 873 1164
rect 1347 1156 1393 1164
rect 2707 1156 2772 1164
rect 2807 1156 2853 1164
rect 4027 1156 4073 1164
rect 4087 1156 4253 1164
rect 307 1136 553 1144
rect 567 1136 653 1144
rect 1967 1136 2173 1144
rect 3007 1136 3093 1144
rect 4756 1146 4764 1216
rect 4827 1217 4873 1225
rect 4896 1186 4904 1233
rect 4927 1216 4944 1224
rect 4936 1164 4944 1216
rect 4967 1216 4993 1224
rect 5167 1216 5213 1224
rect 5227 1217 5293 1225
rect 5727 1216 5984 1224
rect 5976 1204 5984 1216
rect 6067 1216 6113 1224
rect 6327 1216 6473 1224
rect 6496 1216 6573 1224
rect 6496 1204 6504 1216
rect 5976 1200 6044 1204
rect 5976 1196 6047 1200
rect 6033 1187 6047 1196
rect 5087 1176 5193 1184
rect 5267 1176 5353 1184
rect 5627 1175 5693 1183
rect 5807 1175 5973 1183
rect 6456 1196 6504 1204
rect 6456 1186 6464 1196
rect 6087 1175 6133 1183
rect 6347 1176 6453 1184
rect 4936 1156 5053 1164
rect 5616 1164 5624 1172
rect 5547 1156 5624 1164
rect 6027 1156 6233 1164
rect 6247 1156 6313 1164
rect 6527 1156 6553 1164
rect 6567 1156 6613 1164
rect 4167 1136 4373 1144
rect 5507 1136 5653 1144
rect 5667 1136 5753 1144
rect 747 1116 1013 1124
rect 1027 1116 1453 1124
rect 2236 1116 3933 1124
rect 1427 1096 1653 1104
rect 1667 1096 1753 1104
rect 2236 1104 2244 1116
rect 3987 1116 4893 1124
rect 5287 1116 5393 1124
rect 5407 1116 5593 1124
rect 6407 1116 6553 1124
rect 1847 1096 2244 1104
rect 3627 1096 3813 1104
rect 4027 1096 4333 1104
rect 4607 1096 4853 1104
rect 4987 1096 5033 1104
rect 5047 1096 5333 1104
rect 5747 1096 5953 1104
rect 207 1076 493 1084
rect 2567 1076 3633 1084
rect 3647 1076 3993 1084
rect 4007 1076 4413 1084
rect 5367 1076 6053 1084
rect 6307 1076 6493 1084
rect 3047 1056 3233 1064
rect 3247 1056 3393 1064
rect 3687 1056 3733 1064
rect 3747 1056 4293 1064
rect 4367 1056 4813 1064
rect 5107 1056 5273 1064
rect 5327 1056 6073 1064
rect 147 1036 173 1044
rect 187 1036 453 1044
rect 2687 1036 3613 1044
rect 4387 1036 5124 1044
rect 2267 1016 2553 1024
rect 2907 1016 3373 1024
rect 3387 1016 3413 1024
rect 3827 1016 3933 1024
rect 4127 1016 4473 1024
rect 4647 1016 5093 1024
rect 5116 1024 5124 1036
rect 5116 1016 5313 1024
rect 5536 1016 5733 1024
rect 347 996 573 1004
rect 887 996 1153 1004
rect 3347 996 3753 1004
rect 3767 996 3973 1004
rect 5536 1004 5544 1016
rect 6387 1016 6473 1024
rect 5067 996 5544 1004
rect 5927 996 5973 1004
rect 147 976 313 984
rect 1307 976 1513 984
rect 3787 976 4333 984
rect 4636 976 5613 984
rect 4636 967 4644 976
rect 6007 976 6033 984
rect 6047 976 6193 984
rect 347 956 413 964
rect 647 956 913 964
rect 927 956 973 964
rect 1707 956 1973 964
rect 2447 956 2513 964
rect 2527 956 2784 964
rect 1507 936 1673 944
rect 2456 936 2633 944
rect 247 916 273 924
rect 327 916 353 924
rect 367 916 413 924
rect 627 916 733 924
rect 967 917 1013 925
rect 1107 917 1193 925
rect 1267 917 1333 925
rect 1347 916 1473 924
rect 1767 917 1793 925
rect 1807 917 1813 925
rect 2067 917 2093 925
rect 2147 916 2253 924
rect 2327 917 2393 925
rect 2456 924 2464 936
rect 2776 944 2784 956
rect 2827 956 3133 964
rect 3287 956 3313 964
rect 3667 956 3733 964
rect 3847 956 3873 964
rect 4487 956 4633 964
rect 5807 956 6333 964
rect 2776 936 4173 944
rect 4707 936 5133 944
rect 5147 936 5393 944
rect 2407 916 2464 924
rect 2487 916 2593 924
rect 2807 916 2853 924
rect 2867 917 2913 925
rect 3107 917 3172 925
rect 3207 917 3273 925
rect 3387 917 3433 925
rect 3627 916 4033 924
rect 856 896 913 904
rect 856 886 864 896
rect 2756 904 2764 914
rect 2756 896 2884 904
rect 307 875 333 883
rect 1047 875 1093 883
rect 1187 876 1313 884
rect 1367 876 1433 884
rect 1607 876 1633 884
rect 1887 876 1993 884
rect 2127 876 2193 884
rect 2667 876 2693 884
rect 2876 886 2884 896
rect 2887 875 2933 883
rect 167 856 433 864
rect 447 856 793 864
rect 1087 856 1133 864
rect 1327 856 1493 864
rect 1547 856 1673 864
rect 1687 856 1753 864
rect 2956 864 2964 914
rect 4227 917 4312 925
rect 4347 916 4473 924
rect 4487 916 4593 924
rect 4727 917 4793 925
rect 4867 916 4933 924
rect 5027 916 5053 924
rect 5467 916 5493 924
rect 5507 917 5693 925
rect 5887 917 5933 925
rect 5947 916 6033 924
rect 6147 917 6233 925
rect 6327 917 6453 925
rect 6467 916 6673 924
rect 3187 876 3253 884
rect 3807 876 3953 884
rect 4627 876 4713 884
rect 4787 875 4853 883
rect 4907 875 4953 883
rect 5027 875 5233 883
rect 5427 876 5493 884
rect 5587 875 5613 883
rect 5727 876 5793 884
rect 5907 876 5973 884
rect 5987 875 6053 883
rect 6107 876 6213 884
rect 6367 876 6573 884
rect 2787 856 2964 864
rect 3127 856 3433 864
rect 3547 856 3793 864
rect 4047 856 4193 864
rect 4207 856 4244 864
rect 247 836 353 844
rect 2607 836 2633 844
rect 2987 836 3073 844
rect 3427 836 3493 844
rect 3967 836 4193 844
rect 4236 844 4244 856
rect 5747 856 5813 864
rect 4236 836 4453 844
rect 4467 836 4653 844
rect 4667 836 4693 844
rect 4747 836 5593 844
rect 5607 836 6133 844
rect 6327 836 6533 844
rect 307 816 553 824
rect 727 816 853 824
rect 867 816 993 824
rect 3767 816 3972 824
rect 4007 816 4153 824
rect 4167 816 4253 824
rect 4967 816 5513 824
rect 5527 816 5673 824
rect 2287 796 2533 804
rect 2607 796 3633 804
rect 3647 796 4873 804
rect 4887 796 4913 804
rect 607 776 653 784
rect 1567 776 1913 784
rect 2007 776 2413 784
rect 2427 776 2553 784
rect 2727 776 3133 784
rect 3747 776 3773 784
rect 3827 776 3873 784
rect 3987 776 4153 784
rect 4167 776 4233 784
rect 5347 776 5533 784
rect 5707 776 5793 784
rect 5807 776 5853 784
rect 547 756 593 764
rect 607 756 733 764
rect 947 756 3713 764
rect 4127 756 4273 764
rect 4387 756 4573 764
rect 4587 756 5173 764
rect 5967 756 6213 764
rect 6627 756 6673 764
rect 6687 756 6773 764
rect 507 736 893 744
rect 1747 736 1953 744
rect 2287 736 2313 744
rect 2427 736 2473 744
rect 2547 736 2773 744
rect 2827 736 3073 744
rect 3087 736 3193 744
rect 3207 736 3513 744
rect 3887 736 4033 744
rect 4507 736 5113 744
rect 5847 736 5933 744
rect 5947 736 6533 744
rect 6547 736 6593 744
rect 207 716 253 724
rect 1247 716 1353 724
rect 1420 724 1433 727
rect 1416 716 1433 724
rect 1420 713 1433 716
rect 1447 716 1493 724
rect 2527 716 2693 724
rect 3727 716 3793 724
rect 3807 716 4053 724
rect 4987 716 5033 724
rect 127 696 173 704
rect 267 696 413 704
rect 467 696 532 704
rect 567 696 624 704
rect 616 667 624 696
rect 787 696 813 704
rect 1047 697 1073 705
rect 1147 697 1193 705
rect 1347 697 1393 705
rect 1667 697 1713 705
rect 1847 697 1873 705
rect 1987 697 2013 705
rect 2027 696 2193 704
rect 2207 696 2484 704
rect 756 676 853 684
rect 147 656 233 664
rect 367 655 393 663
rect 616 656 633 667
rect 620 653 633 656
rect 756 666 764 676
rect 2476 684 2484 696
rect 3267 697 3293 705
rect 3387 697 3413 705
rect 3467 697 3493 705
rect 3507 696 3553 704
rect 3607 696 3673 704
rect 2476 676 2773 684
rect 2816 684 2824 694
rect 3927 696 3973 704
rect 4047 696 4124 704
rect 2787 676 2824 684
rect 3227 676 3353 684
rect 847 655 953 663
rect 1107 656 1213 664
rect 1267 656 1373 664
rect 1507 655 1573 663
rect 1587 656 1693 664
rect 1747 656 1973 664
rect 2016 656 2033 664
rect 687 636 913 644
rect 2016 644 2024 656
rect 2047 656 2113 664
rect 2847 656 2933 664
rect 3327 656 3373 664
rect 3527 655 3573 663
rect 3756 664 3764 693
rect 4116 684 4124 696
rect 4247 696 4293 704
rect 4153 684 4167 693
rect 4427 696 4452 704
rect 4487 696 4533 704
rect 4707 697 4793 705
rect 5227 696 5253 704
rect 4876 684 4884 694
rect 5307 696 5353 704
rect 5367 697 5413 705
rect 5667 696 5913 704
rect 4116 676 4144 684
rect 4153 680 4224 684
rect 4836 680 4884 684
rect 4156 676 4224 680
rect 3747 656 3764 664
rect 3807 655 3893 663
rect 3907 656 4013 664
rect 4136 664 4144 676
rect 4216 666 4224 676
rect 4833 676 4884 680
rect 4833 667 4847 676
rect 4136 656 4173 664
rect 4407 656 4493 664
rect 4507 655 4553 663
rect 4687 655 4713 663
rect 4907 655 4953 663
rect 5127 655 5153 663
rect 5247 655 5333 663
rect 5496 664 5504 694
rect 6007 696 6053 704
rect 6187 696 6373 704
rect 6387 696 6433 704
rect 6447 696 6473 704
rect 5347 656 5504 664
rect 5607 655 5633 663
rect 5687 656 5753 664
rect 5767 655 5813 663
rect 6027 656 6073 664
rect 6087 655 6113 663
rect 6347 655 6373 663
rect 6487 655 6593 663
rect 1907 636 2024 644
rect 2047 636 2073 644
rect 2087 636 2233 644
rect 3367 636 3433 644
rect 4367 636 4593 644
rect 4607 636 4753 644
rect 4827 636 4853 644
rect 5427 636 5473 644
rect 287 616 353 624
rect 827 616 1133 624
rect 1227 616 1413 624
rect 1567 616 1653 624
rect 2987 616 3153 624
rect 3267 616 3613 624
rect 3687 616 4253 624
rect 4387 616 4573 624
rect 4756 624 4764 633
rect 4756 616 4973 624
rect 5267 620 5404 624
rect 5267 616 5407 620
rect 5393 607 5407 616
rect 5527 616 5853 624
rect 5867 616 5973 624
rect 6247 616 6553 624
rect 247 596 433 604
rect 1307 596 1533 604
rect 3867 596 3933 604
rect 3987 596 4233 604
rect 4327 596 4353 604
rect 4407 596 4673 604
rect 4727 596 5233 604
rect 6307 596 6393 604
rect 1647 576 1773 584
rect 2787 576 3113 584
rect 4387 576 4793 584
rect 4807 576 5093 584
rect 4027 556 4653 564
rect 5387 556 5433 564
rect 2407 536 2513 544
rect 2527 536 2573 544
rect 2887 536 3033 544
rect 3847 536 3953 544
rect 3967 536 4813 544
rect 147 516 173 524
rect 187 516 353 524
rect 3127 516 3513 524
rect 4167 516 4333 524
rect 5287 516 5413 524
rect 667 496 1233 504
rect 1247 496 1333 504
rect 1347 496 1393 504
rect 1567 496 2613 504
rect 2627 496 2693 504
rect 3047 496 4093 504
rect 987 476 1053 484
rect 1067 476 1193 484
rect 1487 476 1733 484
rect 1807 476 2373 484
rect 2487 476 2633 484
rect 3207 476 3253 484
rect 3507 476 3593 484
rect 3887 476 4453 484
rect 527 456 573 464
rect 827 456 913 464
rect 1127 456 1353 464
rect 1367 456 1373 464
rect 1387 456 2433 464
rect 2476 456 2753 464
rect 667 436 713 444
rect 727 436 833 444
rect 1667 436 2033 444
rect 2047 436 2253 444
rect 2476 444 2484 456
rect 2767 456 2913 464
rect 3087 456 3273 464
rect 3287 456 3393 464
rect 4847 456 5173 464
rect 5927 456 6173 464
rect 6187 456 6313 464
rect 2367 436 2484 444
rect 3867 436 4053 444
rect 4427 436 4713 444
rect 347 416 453 424
rect 647 416 873 424
rect 887 416 1033 424
rect 1047 416 1153 424
rect 1167 416 1313 424
rect 1327 416 1513 424
rect 2507 416 2533 424
rect 2847 416 3073 424
rect 5647 416 5853 424
rect 5867 416 6013 424
rect 607 396 753 404
rect 767 396 813 404
rect 1647 397 1693 405
rect 1827 397 1873 405
rect 2087 396 2153 404
rect 2167 397 2213 405
rect 2387 397 2433 405
rect 2447 396 2573 404
rect 2727 397 2793 405
rect 2807 396 2904 404
rect 116 376 333 384
rect 116 366 124 376
rect 227 355 273 363
rect 367 355 393 363
rect 447 356 512 364
rect 547 356 573 364
rect 587 355 673 363
rect 1167 355 1213 363
rect 1267 356 1292 364
rect 1327 355 1373 363
rect 1427 356 1533 364
rect 1596 364 1604 394
rect 1916 384 1924 394
rect 1916 376 1973 384
rect 1596 356 1713 364
rect 1767 356 1793 364
rect 1947 356 2053 364
rect 2067 356 2233 364
rect 2287 356 2353 364
rect 2896 366 2904 396
rect 2967 397 2993 405
rect 3247 397 3313 405
rect 3467 396 3553 404
rect 3827 397 3913 405
rect 4247 396 4373 404
rect 4507 397 4533 405
rect 4676 396 4713 404
rect 2527 355 2593 363
rect 2707 355 2733 363
rect 3036 364 3044 393
rect 3527 376 3584 384
rect 2947 356 3044 364
rect 3107 356 3313 364
rect 3576 366 3584 376
rect 4007 376 4104 384
rect 3327 356 3433 364
rect 3767 355 3833 363
rect 4027 355 4073 363
rect 4096 364 4104 376
rect 4096 356 4213 364
rect 4367 355 4393 363
rect 2787 336 3093 344
rect 3167 336 3253 344
rect 127 316 313 324
rect 327 316 493 324
rect 507 316 733 324
rect 907 316 1653 324
rect 1767 316 1973 324
rect 1987 316 2393 324
rect 2407 316 2864 324
rect 2107 296 2413 304
rect 2467 296 2833 304
rect 2856 304 2864 316
rect 2887 316 2913 324
rect 2927 316 3053 324
rect 3616 324 3624 352
rect 4676 347 4684 396
rect 5007 397 5213 405
rect 5307 397 5333 405
rect 5527 396 5633 404
rect 5767 397 5813 405
rect 5927 397 5973 405
rect 6147 396 6273 404
rect 6407 397 6433 405
rect 6547 397 6653 405
rect 4756 384 4764 394
rect 4756 376 4833 384
rect 5676 367 5684 394
rect 5007 355 5073 363
rect 5407 356 5613 364
rect 5676 356 5692 367
rect 5680 353 5692 356
rect 5727 356 5953 364
rect 6167 355 6213 363
rect 6227 356 6293 364
rect 6467 356 6553 364
rect 3927 336 4293 344
rect 4307 336 4333 344
rect 5367 336 5433 344
rect 5667 336 5753 344
rect 5767 336 5993 344
rect 6007 336 6393 344
rect 3247 316 3624 324
rect 3687 316 4113 324
rect 4127 316 5133 324
rect 5147 316 5293 324
rect 5707 316 5833 324
rect 5847 316 5913 324
rect 5927 316 6073 324
rect 2856 296 3613 304
rect 5327 296 5633 304
rect 5747 296 5793 304
rect 6387 296 6633 304
rect 787 276 1253 284
rect 1267 276 1393 284
rect 1587 276 1633 284
rect 1647 276 1793 284
rect 2416 284 2424 293
rect 2416 276 2993 284
rect 3327 276 3673 284
rect 3847 276 3873 284
rect 4147 276 4392 284
rect 4427 276 4473 284
rect 5287 276 5333 284
rect 5527 276 5593 284
rect 5967 276 6113 284
rect 6127 276 6233 284
rect 167 256 973 264
rect 987 256 1173 264
rect 1847 256 2024 264
rect 2016 247 2024 256
rect 2087 256 3572 264
rect 3607 256 3853 264
rect 4127 256 4433 264
rect 4447 256 4493 264
rect 5207 256 5393 264
rect 5407 256 5493 264
rect 5507 256 5693 264
rect 5707 256 6493 264
rect 227 236 652 244
rect 687 236 824 244
rect 587 216 633 224
rect 816 224 824 236
rect 927 236 1893 244
rect 2027 236 2213 244
rect 2227 236 3933 244
rect 4247 236 4604 244
rect 4596 227 4604 236
rect 4727 236 4773 244
rect 5787 236 5813 244
rect 6007 236 6093 244
rect 6247 236 6593 244
rect 816 216 904 224
rect 427 196 533 204
rect 896 204 904 216
rect 1016 216 1313 224
rect 1016 204 1024 216
rect 1327 216 1473 224
rect 1687 216 1713 224
rect 2067 216 2133 224
rect 2347 216 2453 224
rect 3067 216 3233 224
rect 3656 216 4093 224
rect 3656 207 3664 216
rect 4407 216 4433 224
rect 4447 216 4553 224
rect 4607 216 4833 224
rect 4847 216 4893 224
rect 5007 216 5213 224
rect 5387 216 5513 224
rect 5567 216 6213 224
rect 896 196 1024 204
rect 1527 196 1733 204
rect 1747 196 1813 204
rect 1827 196 2313 204
rect 2507 196 2553 204
rect 3587 196 3653 204
rect 3767 196 3873 204
rect 3887 196 3993 204
rect 4087 196 4133 204
rect 4327 196 4353 204
rect 4367 196 4924 204
rect 4916 188 4924 196
rect 387 176 493 184
rect 647 177 713 185
rect 767 176 873 184
rect 887 176 1033 184
rect 1087 176 1344 184
rect 1336 164 1344 176
rect 1367 176 1413 184
rect 1456 176 1633 184
rect 1456 164 1464 176
rect 1647 176 1913 184
rect 1987 176 2073 184
rect 2096 176 2113 184
rect 1336 156 1464 164
rect 327 135 353 143
rect 667 135 693 143
rect 747 135 813 143
rect 987 135 1053 143
rect 1267 135 1293 143
rect 1427 135 1653 143
rect 1747 135 1813 143
rect 1867 135 1893 143
rect 1907 136 1953 144
rect 2096 144 2104 176
rect 2367 176 2433 184
rect 2647 176 2673 184
rect 3107 177 3133 185
rect 3307 176 3353 184
rect 3407 176 3553 184
rect 3556 164 3564 174
rect 3647 176 3713 184
rect 3736 176 4033 184
rect 3736 164 3744 176
rect 4100 184 4113 187
rect 3556 156 3744 164
rect 4096 173 4113 184
rect 4167 176 4193 184
rect 4467 176 4524 184
rect 4096 146 4104 173
rect 4516 164 4524 176
rect 4547 176 4613 184
rect 4927 177 4953 185
rect 5487 176 5633 184
rect 5647 176 5913 184
rect 6267 176 6433 184
rect 6447 176 6613 184
rect 6627 177 6733 185
rect 4733 164 4747 173
rect 4147 156 4424 164
rect 4516 160 4747 164
rect 4516 156 4744 160
rect 4416 146 4424 156
rect 4656 146 4664 156
rect 2007 136 2104 144
rect 2307 135 2393 143
rect 2667 135 3033 143
rect 3427 136 3573 144
rect 3667 135 3693 143
rect 3747 136 3833 144
rect 3847 135 3893 143
rect 4227 136 4373 144
rect 4387 140 4404 144
rect 4387 136 4407 140
rect 507 116 613 124
rect 976 124 984 132
rect 4393 127 4407 136
rect 4427 135 4473 143
rect 4707 136 4813 144
rect 4907 135 5013 143
rect 5167 136 5273 144
rect 5327 135 5372 143
rect 5407 135 5453 143
rect 5507 136 5553 144
rect 5567 135 5613 143
rect 5787 136 5813 144
rect 5947 135 5993 143
rect 6007 136 6032 144
rect 6067 136 6233 144
rect 6347 135 6413 143
rect 6427 136 6633 144
rect 867 116 984 124
rect 1207 116 1333 124
rect 1347 116 1373 124
rect 2027 116 2133 124
rect 3087 116 3293 124
rect 3587 116 3633 124
rect 4756 116 4973 124
rect 247 96 393 104
rect 747 96 893 104
rect 907 96 1013 104
rect 1927 96 1993 104
rect 2136 104 2144 113
rect 2136 96 2333 104
rect 2447 96 3933 104
rect 3947 96 4053 104
rect 4756 104 4764 116
rect 4627 96 4764 104
rect 4787 96 5993 104
rect 6047 96 6093 104
rect 107 76 593 84
rect 607 76 633 84
rect 1667 76 1973 84
rect 2907 76 3213 84
rect 3387 76 3533 84
rect 3547 76 4313 84
rect 3147 36 4153 44
rect 5227 36 5893 44
rect 5907 36 6453 44
rect 6467 36 6593 44
rect 1947 16 2053 24
rect 2447 16 2533 24
rect 4467 16 4573 24
use NOR2X1  _922_
timestamp 0
transform -1 0 1050 0 -1 3390
box -6 -8 66 268
use INVX2  _923_
timestamp 0
transform 1 0 1250 0 -1 3390
box -6 -8 46 268
use INVX1  _924_
timestamp 0
transform -1 0 2730 0 1 3390
box -6 -8 46 268
use NAND2X1  _925_
timestamp 0
transform 1 0 2550 0 1 3390
box -6 -8 66 268
use OAI21X1  _926_
timestamp 0
transform -1 0 2650 0 -1 3390
box -6 -8 86 268
use INVX2  _927_
timestamp 0
transform -1 0 1170 0 -1 3390
box -6 -8 46 268
use NOR2X1  _928_
timestamp 0
transform -1 0 2050 0 -1 2870
box -6 -8 66 268
use AOI22X1  _929_
timestamp 0
transform 1 0 2990 0 -1 2870
box -6 -8 106 268
use OAI21X1  _930_
timestamp 0
transform 1 0 2590 0 1 2870
box -6 -8 86 268
use INVX1  _931_
timestamp 0
transform -1 0 3710 0 -1 3390
box -6 -8 46 268
use NAND2X1  _932_
timestamp 0
transform 1 0 3030 0 -1 3390
box -6 -8 66 268
use OAI21X1  _933_
timestamp 0
transform 1 0 2870 0 -1 3390
box -6 -8 86 268
use AOI22X1  _934_
timestamp 0
transform 1 0 2930 0 1 2870
box -6 -8 106 268
use OAI21X1  _935_
timestamp 0
transform 1 0 2750 0 1 2870
box -6 -8 86 268
use INVX1  _936_
timestamp 0
transform -1 0 3550 0 1 3390
box -6 -8 46 268
use NAND2X1  _937_
timestamp 0
transform 1 0 2390 0 1 3390
box -6 -8 66 268
use OAI21X1  _938_
timestamp 0
transform 1 0 2170 0 -1 3390
box -6 -8 86 268
use AOI22X1  _939_
timestamp 0
transform 1 0 2410 0 1 2870
box -6 -8 106 268
use OAI21X1  _940_
timestamp 0
transform 1 0 2070 0 1 2870
box -6 -8 86 268
use INVX1  _941_
timestamp 0
transform 1 0 1470 0 -1 3910
box -6 -8 46 268
use NAND2X1  _942_
timestamp 0
transform -1 0 1750 0 1 3390
box -6 -8 66 268
use OAI21X1  _943_
timestamp 0
transform 1 0 1530 0 1 3390
box -6 -8 86 268
use AOI22X1  _944_
timestamp 0
transform -1 0 2330 0 1 2870
box -6 -8 106 268
use OAI21X1  _945_
timestamp 0
transform 1 0 1530 0 -1 3390
box -6 -8 86 268
use INVX1  _946_
timestamp 0
transform -1 0 4550 0 -1 1830
box -6 -8 46 268
use NAND2X1  _947_
timestamp 0
transform -1 0 1030 0 -1 1830
box -6 -8 66 268
use OAI21X1  _948_
timestamp 0
transform 1 0 650 0 -1 1830
box -6 -8 86 268
use INVX1  _949_
timestamp 0
transform 1 0 3790 0 1 2350
box -6 -8 46 268
use NAND2X1  _950_
timestamp 0
transform 1 0 2210 0 -1 1310
box -6 -8 66 268
use OAI21X1  _951_
timestamp 0
transform -1 0 2430 0 -1 1310
box -6 -8 86 268
use INVX2  _952_
timestamp 0
transform 1 0 3910 0 -1 4430
box -6 -8 46 268
use NAND2X1  _953_
timestamp 0
transform 1 0 550 0 1 2870
box -6 -8 66 268
use OAI21X1  _954_
timestamp 0
transform -1 0 770 0 1 2870
box -6 -8 86 268
use INVX2  _955_
timestamp 0
transform 1 0 2750 0 -1 4950
box -6 -8 46 268
use NAND2X1  _956_
timestamp 0
transform -1 0 410 0 1 3390
box -6 -8 66 268
use OAI21X1  _957_
timestamp 0
transform -1 0 570 0 1 3390
box -6 -8 86 268
use NAND2X1  _958_
timestamp 0
transform 1 0 1130 0 1 1830
box -6 -8 66 268
use OAI21X1  _959_
timestamp 0
transform -1 0 1810 0 1 1830
box -6 -8 86 268
use NAND2X1  _960_
timestamp 0
transform 1 0 2670 0 -1 1830
box -6 -8 66 268
use OAI21X1  _961_
timestamp 0
transform -1 0 2910 0 -1 1830
box -6 -8 86 268
use NAND2X1  _962_
timestamp 0
transform -1 0 3050 0 -1 1830
box -6 -8 66 268
use OAI21X1  _963_
timestamp 0
transform -1 0 3090 0 -1 2350
box -6 -8 86 268
use NAND2X1  _964_
timestamp 0
transform 1 0 1330 0 -1 2870
box -6 -8 66 268
use OAI21X1  _965_
timestamp 0
transform -1 0 1450 0 -1 3390
box -6 -8 86 268
use INVX1  _966_
timestamp 0
transform -1 0 3070 0 1 2350
box -6 -8 46 268
use NAND2X1  _967_
timestamp 0
transform 1 0 2730 0 -1 2350
box -6 -8 66 268
use OAI21X1  _968_
timestamp 0
transform -1 0 2950 0 1 2350
box -6 -8 86 268
use INVX1  _969_
timestamp 0
transform -1 0 3470 0 1 2870
box -6 -8 46 268
use NAND2X1  _970_
timestamp 0
transform -1 0 3190 0 1 2870
box -6 -8 66 268
use OAI21X1  _971_
timestamp 0
transform -1 0 3350 0 1 2870
box -6 -8 86 268
use INVX1  _972_
timestamp 0
transform -1 0 3110 0 1 1830
box -6 -8 46 268
use NAND2X1  _973_
timestamp 0
transform -1 0 2590 0 -1 1830
box -6 -8 66 268
use OAI21X1  _974_
timestamp 0
transform -1 0 2990 0 1 1830
box -6 -8 86 268
use INVX1  _975_
timestamp 0
transform -1 0 2650 0 -1 2870
box -6 -8 46 268
use NAND2X1  _976_
timestamp 0
transform 1 0 2270 0 1 2350
box -6 -8 66 268
use OAI21X1  _977_
timestamp 0
transform -1 0 2490 0 1 2350
box -6 -8 86 268
use INVX1  _978_
timestamp 0
transform -1 0 3790 0 -1 2870
box -6 -8 46 268
use NAND2X1  _979_
timestamp 0
transform 1 0 3330 0 -1 2350
box -6 -8 66 268
use OAI21X1  _980_
timestamp 0
transform -1 0 3670 0 -1 2870
box -6 -8 86 268
use INVX1  _981_
timestamp 0
transform -1 0 3390 0 1 1830
box -6 -8 46 268
use NAND2X1  _982_
timestamp 0
transform -1 0 2990 0 1 1310
box -6 -8 66 268
use OAI21X1  _983_
timestamp 0
transform -1 0 3270 0 1 1830
box -6 -8 86 268
use INVX8  _984_
timestamp 0
transform -1 0 3570 0 -1 3390
box -6 -8 106 268
use INVX1  _985_
timestamp 0
transform 1 0 4170 0 -1 2350
box -6 -8 46 268
use NAND2X1  _986_
timestamp 0
transform 1 0 4110 0 -1 2870
box -6 -8 66 268
use OAI21X1  _987_
timestamp 0
transform -1 0 4330 0 -1 2870
box -6 -8 86 268
use INVX1  _988_
timestamp 0
transform 1 0 3730 0 1 1830
box -6 -8 46 268
use NAND2X1  _989_
timestamp 0
transform 1 0 2570 0 1 2350
box -6 -8 66 268
use OAI21X1  _990_
timestamp 0
transform -1 0 2790 0 1 2350
box -6 -8 86 268
use NAND2X1  _991_
timestamp 0
transform 1 0 2850 0 -1 3910
box -6 -8 66 268
use OAI21X1  _992_
timestamp 0
transform 1 0 2810 0 1 3390
box -6 -8 86 268
use NAND2X1  _993_
timestamp 0
transform 1 0 3990 0 1 3390
box -6 -8 66 268
use OAI21X1  _994_
timestamp 0
transform -1 0 4130 0 -1 3390
box -6 -8 86 268
use NAND2X1  _995_
timestamp 0
transform 1 0 3370 0 1 3390
box -6 -8 66 268
use OAI21X1  _996_
timestamp 0
transform 1 0 3210 0 1 3390
box -6 -8 86 268
use NAND2X1  _997_
timestamp 0
transform 1 0 1770 0 -1 3910
box -6 -8 66 268
use OAI21X1  _998_
timestamp 0
transform 1 0 1590 0 -1 3910
box -6 -8 86 268
use INVX1  _999_
timestamp 0
transform 1 0 2310 0 -1 3910
box -6 -8 46 268
use NAND2X1  _1000_
timestamp 0
transform -1 0 3210 0 1 3910
box -6 -8 66 268
use OAI21X1  _1001_
timestamp 0
transform 1 0 2430 0 -1 3910
box -6 -8 86 268
use INVX1  _1002_
timestamp 0
transform -1 0 2650 0 1 4430
box -6 -8 46 268
use NAND2X1  _1003_
timestamp 0
transform 1 0 2990 0 1 3910
box -6 -8 66 268
use OAI21X1  _1004_
timestamp 0
transform 1 0 2810 0 1 3910
box -6 -8 86 268
use INVX1  _1005_
timestamp 0
transform -1 0 2030 0 1 3390
box -6 -8 46 268
use NAND2X1  _1006_
timestamp 0
transform 1 0 1930 0 -1 3910
box -6 -8 66 268
use OAI21X1  _1007_
timestamp 0
transform 1 0 1830 0 1 3390
box -6 -8 86 268
use INVX1  _1008_
timestamp 0
transform 1 0 1570 0 1 3910
box -6 -8 46 268
use NAND2X1  _1009_
timestamp 0
transform 1 0 1170 0 -1 3910
box -6 -8 66 268
use OAI21X1  _1010_
timestamp 0
transform -1 0 1390 0 -1 3910
box -6 -8 86 268
use NAND3X1  _1011_
timestamp 0
transform 1 0 1070 0 -1 2350
box -6 -8 86 268
use INVX1  _1012_
timestamp 0
transform 1 0 2390 0 1 1310
box -6 -8 46 268
use INVX1  _1013_
timestamp 0
transform -1 0 3510 0 -1 2350
box -6 -8 46 268
use INVX1  _1014_
timestamp 0
transform 1 0 950 0 -1 2350
box -6 -8 46 268
use OAI21X1  _1015_
timestamp 0
transform -1 0 1930 0 -1 2350
box -6 -8 86 268
use NAND2X1  _1016_
timestamp 0
transform 1 0 2010 0 -1 2350
box -6 -8 66 268
use NAND2X1  _1017_
timestamp 0
transform 1 0 2570 0 -1 2350
box -6 -8 66 268
use OAI21X1  _1018_
timestamp 0
transform 1 0 2170 0 -1 2350
box -6 -8 86 268
use AOI21X1  _1019_
timestamp 0
transform -1 0 870 0 1 1830
box -6 -8 86 268
use NAND3X1  _1020_
timestamp 0
transform 1 0 950 0 1 1830
box -6 -8 86 268
use INVX1  _1021_
timestamp 0
transform 1 0 1270 0 -1 1830
box -6 -8 46 268
use NAND2X1  _1022_
timestamp 0
transform -1 0 1550 0 1 1310
box -6 -8 66 268
use OAI21X1  _1023_
timestamp 0
transform 1 0 1390 0 -1 1830
box -6 -8 86 268
use INVX1  _1024_
timestamp 0
transform 1 0 1290 0 1 1830
box -6 -8 46 268
use INVX1  _1025_
timestamp 0
transform -1 0 1590 0 -1 1830
box -6 -8 46 268
use NAND3X1  _1026_
timestamp 0
transform 1 0 1410 0 1 1830
box -6 -8 86 268
use NAND2X1  _1027_
timestamp 0
transform 1 0 1590 0 1 1830
box -6 -8 66 268
use OR2X2  _1028_
timestamp 0
transform -1 0 1610 0 -1 2350
box -6 -8 86 268
use NAND2X1  _1029_
timestamp 0
transform -1 0 1750 0 -1 2350
box -6 -8 66 268
use NAND2X1  _1030_
timestamp 0
transform -1 0 1650 0 1 2350
box -6 -8 66 268
use NAND2X1  _1031_
timestamp 0
transform 1 0 1910 0 1 2870
box -6 -8 66 268
use OAI21X1  _1032_
timestamp 0
transform 1 0 1750 0 1 2870
box -6 -8 86 268
use NAND2X1  _1033_
timestamp 0
transform 1 0 2370 0 -1 1830
box -6 -8 66 268
use INVX1  _1034_
timestamp 0
transform 1 0 1670 0 -1 1830
box -6 -8 46 268
use INVX4  _1035_
timestamp 0
transform 1 0 3910 0 1 2350
box -6 -8 66 268
use OAI21X1  _1036_
timestamp 0
transform -1 0 1410 0 1 1310
box -6 -8 86 268
use INVX1  _1037_
timestamp 0
transform 1 0 1150 0 -1 1310
box -6 -8 46 268
use INVX1  _1038_
timestamp 0
transform -1 0 4670 0 -1 1830
box -6 -8 46 268
use INVX1  _1039_
timestamp 0
transform -1 0 1670 0 -1 1310
box -6 -8 46 268
use AOI21X1  _1040_
timestamp 0
transform 1 0 710 0 1 1310
box -6 -8 86 268
use NAND3X1  _1041_
timestamp 0
transform 1 0 550 0 -1 1310
box -6 -8 86 268
use INVX1  _1042_
timestamp 0
transform 1 0 850 0 1 790
box -6 -8 46 268
use NOR2X1  _1043_
timestamp 0
transform -1 0 770 0 -1 1310
box -6 -8 66 268
use OAI21X1  _1044_
timestamp 0
transform -1 0 1530 0 -1 1310
box -6 -8 86 268
use NAND2X1  _1045_
timestamp 0
transform 1 0 1170 0 1 1310
box -6 -8 66 268
use INVX1  _1046_
timestamp 0
transform 1 0 1030 0 1 1310
box -6 -8 46 268
use OAI21X1  _1047_
timestamp 0
transform 1 0 850 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1048_
timestamp 0
transform 1 0 1290 0 -1 1310
box -6 -8 86 268
use NAND2X1  _1049_
timestamp 0
transform -1 0 1070 0 -1 1310
box -6 -8 66 268
use OAI21X1  _1050_
timestamp 0
transform 1 0 1130 0 1 790
box -6 -8 86 268
use NAND3X1  _1051_
timestamp 0
transform 1 0 1470 0 1 790
box -6 -8 86 268
use NAND2X1  _1052_
timestamp 0
transform -1 0 1810 0 -1 1310
box -6 -8 66 268
use OAI21X1  _1053_
timestamp 0
transform -1 0 2050 0 1 1310
box -6 -8 86 268
use NAND2X1  _1054_
timestamp 0
transform 1 0 2390 0 1 790
box -6 -8 66 268
use INVX1  _1055_
timestamp 0
transform -1 0 2010 0 1 790
box -6 -8 46 268
use NAND3X1  _1056_
timestamp 0
transform -1 0 1710 0 1 790
box -6 -8 86 268
use AOI21X1  _1057_
timestamp 0
transform -1 0 1890 0 1 1310
box -6 -8 86 268
use NAND3X1  _1058_
timestamp 0
transform 1 0 1630 0 1 1310
box -6 -8 86 268
use NAND2X1  _1059_
timestamp 0
transform -1 0 1850 0 -1 1830
box -6 -8 66 268
use OAI21X1  _1060_
timestamp 0
transform 1 0 1950 0 -1 1830
box -6 -8 86 268
use NAND2X1  _1061_
timestamp 0
transform -1 0 2350 0 1 1830
box -6 -8 66 268
use AOI21X1  _1062_
timestamp 0
transform 1 0 1290 0 1 790
box -6 -8 86 268
use OAI21X1  _1063_
timestamp 0
transform -1 0 1890 0 1 790
box -6 -8 86 268
use NAND2X1  _1064_
timestamp 0
transform -1 0 3670 0 1 790
box -6 -8 66 268
use NOR2X1  _1065_
timestamp 0
transform 1 0 2550 0 -1 790
box -6 -8 66 268
use AOI22X1  _1066_
timestamp 0
transform -1 0 2650 0 1 790
box -6 -8 106 268
use NOR2X1  _1067_
timestamp 0
transform 1 0 2410 0 -1 790
box -6 -8 66 268
use OAI21X1  _1068_
timestamp 0
transform -1 0 1050 0 1 790
box -6 -8 86 268
use NAND2X1  _1069_
timestamp 0
transform -1 0 310 0 -1 1310
box -6 -8 66 268
use NAND3X1  _1070_
timestamp 0
transform -1 0 470 0 1 790
box -6 -8 86 268
use INVX1  _1071_
timestamp 0
transform 1 0 270 0 1 270
box -6 -8 46 268
use AOI21X1  _1072_
timestamp 0
transform -1 0 190 0 1 790
box -6 -8 86 268
use OAI21X1  _1073_
timestamp 0
transform 1 0 390 0 1 270
box -6 -8 86 268
use INVX1  _1074_
timestamp 0
transform -1 0 310 0 1 790
box -6 -8 46 268
use INVX1  _1075_
timestamp 0
transform 1 0 110 0 -1 790
box -6 -8 46 268
use NAND3X1  _1076_
timestamp 0
transform 1 0 390 0 -1 790
box -6 -8 86 268
use NAND3X1  _1077_
timestamp 0
transform -1 0 630 0 -1 790
box -6 -8 86 268
use INVX1  _1078_
timestamp 0
transform 1 0 1070 0 -1 790
box -6 -8 46 268
use AOI21X1  _1079_
timestamp 0
transform 1 0 710 0 -1 790
box -6 -8 86 268
use OAI21X1  _1080_
timestamp 0
transform 1 0 1190 0 -1 790
box -6 -8 86 268
use INVX1  _1081_
timestamp 0
transform -1 0 1090 0 1 270
box -6 -8 46 268
use INVX1  _1082_
timestamp 0
transform 1 0 710 0 1 790
box -6 -8 46 268
use AOI21X1  _1083_
timestamp 0
transform 1 0 230 0 -1 790
box -6 -8 86 268
use INVX1  _1084_
timestamp 0
transform 1 0 250 0 1 1310
box -6 -8 46 268
use NAND3X1  _1085_
timestamp 0
transform 1 0 370 0 1 1310
box -6 -8 86 268
use INVX2  _1086_
timestamp 0
transform -1 0 4990 0 1 1830
box -6 -8 46 268
use OAI21X1  _1087_
timestamp 0
transform -1 0 630 0 1 1310
box -6 -8 86 268
use AOI21X1  _1088_
timestamp 0
transform -1 0 470 0 -1 1310
box -6 -8 86 268
use OAI21X1  _1089_
timestamp 0
transform 1 0 550 0 1 790
box -6 -8 86 268
use NAND3X1  _1090_
timestamp 0
transform 1 0 1190 0 1 270
box -6 -8 86 268
use NAND2X1  _1091_
timestamp 0
transform 1 0 1530 0 -1 790
box -6 -8 66 268
use NOR2X1  _1092_
timestamp 0
transform 1 0 1870 0 -1 790
box -6 -8 66 268
use AOI22X1  _1093_
timestamp 0
transform -1 0 1790 0 -1 790
box -6 -8 106 268
use OAI21X1  _1094_
timestamp 0
transform 1 0 2010 0 -1 790
box -6 -8 86 268
use NOR3X1  _1095_
timestamp 0
transform 1 0 2170 0 -1 790
box -6 -8 166 268
use INVX1  _1096_
timestamp 0
transform -1 0 2290 0 1 790
box -6 -8 46 268
use NAND2X1  _1097_
timestamp 0
transform 1 0 2090 0 1 790
box -6 -8 66 268
use OAI21X1  _1098_
timestamp 0
transform 1 0 2130 0 1 1830
box -6 -8 86 268
use NAND2X1  _1099_
timestamp 0
transform -1 0 2910 0 -1 1310
box -6 -8 66 268
use INVX1  _1100_
timestamp 0
transform 1 0 2690 0 -1 790
box -6 -8 46 268
use OAI21X1  _1101_
timestamp 0
transform -1 0 950 0 1 270
box -6 -8 86 268
use OAI21X1  _1102_
timestamp 0
transform 1 0 110 0 1 270
box -6 -8 86 268
use INVX1  _1103_
timestamp 0
transform 1 0 1170 0 -1 270
box -6 -8 46 268
use AOI21X1  _1104_
timestamp 0
transform -1 0 950 0 1 1310
box -6 -8 86 268
use INVX1  _1105_
timestamp 0
transform 1 0 570 0 1 270
box -6 -8 46 268
use NAND3X1  _1106_
timestamp 0
transform -1 0 890 0 -1 1830
box -6 -8 86 268
use NAND2X1  _1107_
timestamp 0
transform -1 0 150 0 -1 1310
box -6 -8 66 268
use NAND3X1  _1108_
timestamp 0
transform 1 0 710 0 1 270
box -6 -8 86 268
use INVX1  _1109_
timestamp 0
transform 1 0 210 0 -1 270
box -6 -8 46 268
use INVX1  _1110_
timestamp 0
transform -1 0 130 0 -1 270
box -6 -8 46 268
use OAI21X1  _1111_
timestamp 0
transform 1 0 530 0 -1 270
box -6 -8 86 268
use NAND3X1  _1112_
timestamp 0
transform 1 0 1450 0 -1 270
box -6 -8 86 268
use NAND3X1  _1113_
timestamp 0
transform 1 0 690 0 -1 270
box -6 -8 86 268
use OAI21X1  _1114_
timestamp 0
transform -1 0 430 0 -1 270
box -6 -8 86 268
use NAND3X1  _1115_
timestamp 0
transform 1 0 850 0 -1 270
box -6 -8 86 268
use NAND2X1  _1116_
timestamp 0
transform 1 0 3930 0 1 1310
box -6 -8 66 268
use INVX1  _1117_
timestamp 0
transform -1 0 4970 0 1 790
box -6 -8 46 268
use AND2X2  _1118_
timestamp 0
transform 1 0 4410 0 1 790
box -6 -8 86 268
use AND2X2  _1119_
timestamp 0
transform 1 0 4410 0 -1 1310
box -6 -8 86 268
use NAND2X1  _1120_
timestamp 0
transform 1 0 4590 0 1 790
box -6 -8 66 268
use INVX2  _1121_
timestamp 0
transform -1 0 4490 0 -1 2350
box -6 -8 46 268
use OAI21X1  _1122_
timestamp 0
transform 1 0 4690 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1123_
timestamp 0
transform 1 0 4750 0 1 790
box -6 -8 86 268
use OAI21X1  _1124_
timestamp 0
transform 1 0 3710 0 -1 1310
box -6 -8 86 268
use INVX2  _1125_
timestamp 0
transform 1 0 3870 0 1 3390
box -6 -8 46 268
use OAI21X1  _1126_
timestamp 0
transform 1 0 4050 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1127_
timestamp 0
transform -1 0 3950 0 -1 1310
box -6 -8 86 268
use AND2X2  _1128_
timestamp 0
transform -1 0 3810 0 1 270
box -6 -8 86 268
use NAND3X1  _1129_
timestamp 0
transform 1 0 1870 0 1 270
box -6 -8 86 268
use AOI21X1  _1130_
timestamp 0
transform 1 0 1010 0 -1 270
box -6 -8 86 268
use AOI21X1  _1131_
timestamp 0
transform 1 0 1290 0 -1 270
box -6 -8 86 268
use NAND2X1  _1132_
timestamp 0
transform -1 0 3970 0 1 270
box -6 -8 66 268
use OAI21X1  _1133_
timestamp 0
transform 1 0 2110 0 -1 270
box -6 -8 86 268
use AOI21X1  _1134_
timestamp 0
transform 1 0 2210 0 1 270
box -6 -8 86 268
use NAND3X1  _1135_
timestamp 0
transform 1 0 1350 0 1 270
box -6 -8 86 268
use NAND3X1  _1136_
timestamp 0
transform -1 0 1870 0 -1 270
box -6 -8 86 268
use OAI21X1  _1137_
timestamp 0
transform 1 0 1630 0 -1 270
box -6 -8 86 268
use AOI22X1  _1138_
timestamp 0
transform 1 0 1510 0 1 270
box -6 -8 106 268
use OAI21X1  _1139_
timestamp 0
transform 1 0 2730 0 1 270
box -6 -8 86 268
use AOI21X1  _1140_
timestamp 0
transform 1 0 1370 0 -1 790
box -6 -8 86 268
use NAND3X1  _1141_
timestamp 0
transform 1 0 1690 0 1 270
box -6 -8 86 268
use NAND3X1  _1142_
timestamp 0
transform 1 0 2030 0 1 270
box -6 -8 86 268
use NAND3X1  _1143_
timestamp 0
transform 1 0 2390 0 1 270
box -6 -8 86 268
use NAND3X1  _1144_
timestamp 0
transform -1 0 3130 0 1 270
box -6 -8 86 268
use INVX1  _1145_
timestamp 0
transform 1 0 2810 0 -1 790
box -6 -8 46 268
use NAND2X1  _1146_
timestamp 0
transform 1 0 3230 0 1 270
box -6 -8 66 268
use NAND2X1  _1147_
timestamp 0
transform 1 0 2930 0 -1 790
box -6 -8 66 268
use AOI21X1  _1148_
timestamp 0
transform 1 0 2910 0 1 790
box -6 -8 86 268
use NAND3X1  _1149_
timestamp 0
transform 1 0 2750 0 1 790
box -6 -8 86 268
use NAND2X1  _1150_
timestamp 0
transform 1 0 3230 0 1 790
box -6 -8 66 268
use OAI21X1  _1151_
timestamp 0
transform 1 0 3070 0 1 790
box -6 -8 86 268
use NAND2X1  _1152_
timestamp 0
transform 1 0 2530 0 -1 1310
box -6 -8 66 268
use INVX1  _1153_
timestamp 0
transform -1 0 2930 0 -1 270
box -6 -8 46 268
use OAI21X1  _1154_
timestamp 0
transform 1 0 2890 0 1 270
box -6 -8 86 268
use INVX1  _1155_
timestamp 0
transform 1 0 4750 0 -1 2870
box -6 -8 46 268
use NOR2X1  _1156_
timestamp 0
transform 1 0 4670 0 1 2350
box -6 -8 66 268
use INVX1  _1157_
timestamp 0
transform -1 0 5090 0 1 270
box -6 -8 46 268
use INVX1  _1158_
timestamp 0
transform -1 0 5590 0 1 790
box -6 -8 46 268
use OAI21X1  _1159_
timestamp 0
transform -1 0 4930 0 -1 790
box -6 -8 86 268
use XOR2X1  _1160_
timestamp 0
transform 1 0 4850 0 1 270
box -6 -8 126 268
use AOI21X1  _1161_
timestamp 0
transform 1 0 2290 0 -1 270
box -6 -8 86 268
use NAND2X1  _1162_
timestamp 0
transform -1 0 4130 0 1 1310
box -6 -8 66 268
use AND2X2  _1163_
timestamp 0
transform -1 0 5090 0 1 1310
box -6 -8 86 268
use OAI21X1  _1164_
timestamp 0
transform 1 0 4570 0 1 1310
box -6 -8 86 268
use AND2X2  _1165_
timestamp 0
transform -1 0 4950 0 -1 1830
box -6 -8 86 268
use OAI21X1  _1166_
timestamp 0
transform 1 0 4210 0 1 1310
box -6 -8 86 268
use NAND3X1  _1167_
timestamp 0
transform -1 0 4470 0 1 1310
box -6 -8 86 268
use INVX1  _1168_
timestamp 0
transform 1 0 4570 0 -1 1310
box -6 -8 46 268
use NAND2X1  _1169_
timestamp 0
transform -1 0 4930 0 1 1310
box -6 -8 66 268
use OAI22X1  _1170_
timestamp 0
transform 1 0 4230 0 -1 1310
box -6 -8 106 268
use NAND3X1  _1171_
timestamp 0
transform 1 0 4850 0 -1 1310
box -6 -8 86 268
use NAND2X1  _1172_
timestamp 0
transform 1 0 5050 0 1 790
box -6 -8 66 268
use OAI21X1  _1173_
timestamp 0
transform 1 0 890 0 -1 790
box -6 -8 86 268
use INVX1  _1174_
timestamp 0
transform 1 0 3710 0 -1 790
box -6 -8 46 268
use NAND2X1  _1175_
timestamp 0
transform 1 0 3310 0 1 1310
box -6 -8 66 268
use NAND3X1  _1176_
timestamp 0
transform 1 0 3390 0 -1 1830
box -6 -8 86 268
use INVX1  _1177_
timestamp 0
transform -1 0 3490 0 1 1310
box -6 -8 46 268
use AOI21X1  _1178_
timestamp 0
transform -1 0 4090 0 -1 1830
box -6 -8 86 268
use OAI21X1  _1179_
timestamp 0
transform 1 0 3590 0 1 1310
box -6 -8 86 268
use INVX1  _1180_
timestamp 0
transform 1 0 3310 0 -1 1310
box -6 -8 46 268
use INVX1  _1181_
timestamp 0
transform 1 0 3590 0 -1 1310
box -6 -8 46 268
use NAND3X1  _1182_
timestamp 0
transform 1 0 3770 0 1 790
box -6 -8 86 268
use NAND3X1  _1183_
timestamp 0
transform 1 0 4170 0 -1 790
box -6 -8 86 268
use AOI21X1  _1184_
timestamp 0
transform 1 0 3930 0 1 790
box -6 -8 86 268
use INVX1  _1185_
timestamp 0
transform 1 0 3570 0 -1 1830
box -6 -8 46 268
use NAND3X1  _1186_
timestamp 0
transform 1 0 3690 0 -1 1830
box -6 -8 86 268
use OAI21X1  _1187_
timestamp 0
transform 1 0 3850 0 -1 1830
box -6 -8 86 268
use AOI21X1  _1188_
timestamp 0
transform 1 0 3770 0 1 1310
box -6 -8 86 268
use OAI21X1  _1189_
timestamp 0
transform -1 0 4170 0 1 790
box -6 -8 86 268
use NAND3X1  _1190_
timestamp 0
transform 1 0 4370 0 1 270
box -6 -8 86 268
use AND2X2  _1191_
timestamp 0
transform -1 0 5290 0 1 790
box -6 -8 86 268
use NAND3X1  _1192_
timestamp 0
transform 1 0 4010 0 -1 790
box -6 -8 86 268
use OAI21X1  _1193_
timestamp 0
transform 1 0 4250 0 1 790
box -6 -8 86 268
use NAND3X1  _1194_
timestamp 0
transform -1 0 4610 0 -1 790
box -6 -8 86 268
use NAND3X1  _1195_
timestamp 0
transform -1 0 4110 0 -1 270
box -6 -8 86 268
use OAI21X1  _1196_
timestamp 0
transform -1 0 2030 0 -1 270
box -6 -8 86 268
use AOI21X1  _1197_
timestamp 0
transform 1 0 4350 0 -1 790
box -6 -8 86 268
use AOI21X1  _1198_
timestamp 0
transform -1 0 4290 0 1 270
box -6 -8 86 268
use OAI21X1  _1199_
timestamp 0
transform -1 0 3770 0 -1 270
box -6 -8 86 268
use NAND3X1  _1200_
timestamp 0
transform 1 0 3530 0 -1 270
box -6 -8 86 268
use INVX1  _1201_
timestamp 0
transform 1 0 4350 0 -1 270
box -6 -8 46 268
use NAND3X1  _1202_
timestamp 0
transform 1 0 4530 0 1 270
box -6 -8 86 268
use OAI21X1  _1203_
timestamp 0
transform 1 0 3870 0 -1 270
box -6 -8 86 268
use NAND3X1  _1204_
timestamp 0
transform -1 0 4770 0 1 270
box -6 -8 86 268
use NAND3X1  _1205_
timestamp 0
transform 1 0 4050 0 1 270
box -6 -8 86 268
use AOI21X1  _1206_
timestamp 0
transform 1 0 2570 0 1 270
box -6 -8 86 268
use AOI21X1  _1207_
timestamp 0
transform -1 0 4270 0 -1 270
box -6 -8 86 268
use AOI21X1  _1208_
timestamp 0
transform -1 0 3430 0 -1 270
box -6 -8 86 268
use OAI21X1  _1209_
timestamp 0
transform -1 0 3110 0 -1 270
box -6 -8 86 268
use NAND3X1  _1210_
timestamp 0
transform -1 0 3270 0 -1 270
box -6 -8 86 268
use INVX1  _1211_
timestamp 0
transform 1 0 3290 0 -1 790
box -6 -8 46 268
use AND2X2  _1212_
timestamp 0
transform 1 0 3390 0 1 270
box -6 -8 86 268
use AOI22X1  _1213_
timestamp 0
transform 1 0 3550 0 1 270
box -6 -8 106 268
use NOR2X1  _1214_
timestamp 0
transform -1 0 3470 0 -1 790
box -6 -8 66 268
use XOR2X1  _1215_
timestamp 0
transform -1 0 3210 0 -1 790
box -6 -8 126 268
use OAI21X1  _1216_
timestamp 0
transform -1 0 2750 0 -1 1310
box -6 -8 86 268
use OAI21X1  _1217_
timestamp 0
transform 1 0 3550 0 -1 790
box -6 -8 86 268
use INVX1  _1218_
timestamp 0
transform 1 0 5130 0 -1 270
box -6 -8 46 268
use NAND2X1  _1219_
timestamp 0
transform -1 0 5230 0 1 270
box -6 -8 66 268
use INVX1  _1220_
timestamp 0
transform -1 0 4850 0 -1 270
box -6 -8 46 268
use AOI21X1  _1221_
timestamp 0
transform 1 0 4650 0 -1 270
box -6 -8 86 268
use AOI22X1  _1222_
timestamp 0
transform 1 0 4550 0 -1 2870
box -6 -8 106 268
use AND2X2  _1223_
timestamp 0
transform 1 0 5050 0 -1 2870
box -6 -8 86 268
use NAND2X1  _1224_
timestamp 0
transform -1 0 5230 0 1 2350
box -6 -8 66 268
use INVX1  _1225_
timestamp 0
transform 1 0 6150 0 -1 2350
box -6 -8 46 268
use NOR2X1  _1226_
timestamp 0
transform 1 0 6010 0 -1 2350
box -6 -8 66 268
use NAND2X1  _1227_
timestamp 0
transform -1 0 5450 0 1 790
box -6 -8 66 268
use OAI21X1  _1228_
timestamp 0
transform 1 0 5670 0 1 790
box -6 -8 86 268
use XNOR2X1  _1229_
timestamp 0
transform -1 0 6470 0 1 790
box -6 -8 126 268
use INVX1  _1230_
timestamp 0
transform 1 0 5030 0 -1 790
box -6 -8 46 268
use AOI21X1  _1231_
timestamp 0
transform 1 0 5150 0 -1 790
box -6 -8 86 268
use NAND2X1  _1232_
timestamp 0
transform 1 0 4890 0 -1 2350
box -6 -8 66 268
use NAND2X1  _1233_
timestamp 0
transform -1 0 5270 0 1 1830
box -6 -8 66 268
use NOR2X1  _1234_
timestamp 0
transform 1 0 5670 0 1 1830
box -6 -8 66 268
use AND2X2  _1235_
timestamp 0
transform -1 0 5590 0 1 1830
box -6 -8 86 268
use OAI21X1  _1236_
timestamp 0
transform -1 0 5590 0 -1 2350
box -6 -8 86 268
use INVX1  _1237_
timestamp 0
transform 1 0 5030 0 -1 2350
box -6 -8 46 268
use AND2X2  _1238_
timestamp 0
transform 1 0 4570 0 -1 2350
box -6 -8 86 268
use NAND2X1  _1239_
timestamp 0
transform -1 0 4810 0 -1 2350
box -6 -8 66 268
use OAI21X1  _1240_
timestamp 0
transform 1 0 5350 0 1 1830
box -6 -8 86 268
use NAND3X1  _1241_
timestamp 0
transform 1 0 5330 0 -1 2350
box -6 -8 86 268
use NAND2X1  _1242_
timestamp 0
transform 1 0 5830 0 1 1830
box -6 -8 66 268
use OAI21X1  _1243_
timestamp 0
transform -1 0 3510 0 -1 1310
box -6 -8 86 268
use INVX1  _1244_
timestamp 0
transform 1 0 5650 0 1 1310
box -6 -8 46 268
use NAND2X1  _1245_
timestamp 0
transform 1 0 4190 0 -1 1830
box -6 -8 66 268
use NAND3X1  _1246_
timestamp 0
transform 1 0 4510 0 1 2350
box -6 -8 86 268
use INVX1  _1247_
timestamp 0
transform -1 0 5070 0 -1 1830
box -6 -8 46 268
use AOI21X1  _1248_
timestamp 0
transform 1 0 4350 0 1 2350
box -6 -8 86 268
use OAI21X1  _1249_
timestamp 0
transform 1 0 5150 0 -1 1830
box -6 -8 86 268
use INVX1  _1250_
timestamp 0
transform 1 0 5450 0 -1 1830
box -6 -8 46 268
use INVX1  _1251_
timestamp 0
transform 1 0 5330 0 -1 1830
box -6 -8 46 268
use NAND3X1  _1252_
timestamp 0
transform 1 0 5750 0 -1 1830
box -6 -8 86 268
use NAND3X1  _1253_
timestamp 0
transform -1 0 5850 0 1 1310
box -6 -8 86 268
use AOI21X1  _1254_
timestamp 0
transform -1 0 5670 0 -1 1830
box -6 -8 86 268
use INVX1  _1255_
timestamp 0
transform -1 0 4090 0 1 2350
box -6 -8 46 268
use NAND3X1  _1256_
timestamp 0
transform 1 0 4170 0 1 2350
box -6 -8 86 268
use OAI21X1  _1257_
timestamp 0
transform 1 0 3750 0 -1 2350
box -6 -8 86 268
use AOI21X1  _1258_
timestamp 0
transform 1 0 4290 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1259_
timestamp 0
transform -1 0 5390 0 1 1310
box -6 -8 86 268
use NAND3X1  _1260_
timestamp 0
transform 1 0 6030 0 1 790
box -6 -8 86 268
use AND2X2  _1261_
timestamp 0
transform 1 0 5970 0 1 1830
box -6 -8 86 268
use NAND3X1  _1262_
timestamp 0
transform 1 0 5910 0 -1 1830
box -6 -8 86 268
use OAI21X1  _1263_
timestamp 0
transform 1 0 5490 0 1 1310
box -6 -8 86 268
use NAND3X1  _1264_
timestamp 0
transform 1 0 5650 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1265_
timestamp 0
transform -1 0 6030 0 -1 790
box -6 -8 86 268
use AOI21X1  _1266_
timestamp 0
transform 1 0 3850 0 -1 790
box -6 -8 86 268
use OAI21X1  _1267_
timestamp 0
transform 1 0 4690 0 -1 790
box -6 -8 86 268
use AOI21X1  _1268_
timestamp 0
transform 1 0 5490 0 -1 1310
box -6 -8 86 268
use AOI21X1  _1269_
timestamp 0
transform -1 0 5930 0 1 790
box -6 -8 86 268
use OAI21X1  _1270_
timestamp 0
transform -1 0 5710 0 -1 790
box -6 -8 86 268
use NAND3X1  _1271_
timestamp 0
transform 1 0 6270 0 1 270
box -6 -8 86 268
use XOR2X1  _1272_
timestamp 0
transform -1 0 6690 0 1 790
box -6 -8 126 268
use NAND3X1  _1273_
timestamp 0
transform 1 0 6110 0 -1 790
box -6 -8 86 268
use OAI21X1  _1274_
timestamp 0
transform 1 0 5790 0 -1 790
box -6 -8 86 268
use NAND3X1  _1275_
timestamp 0
transform -1 0 6730 0 -1 6510
box -6 -8 86 268
use NAND3X1  _1276_
timestamp 0
transform -1 0 6290 0 -1 270
box -6 -8 86 268
use AOI21X1  _1277_
timestamp 0
transform 1 0 4470 0 -1 270
box -6 -8 86 268
use OAI21X1  _1278_
timestamp 0
transform 1 0 4950 0 -1 270
box -6 -8 86 268
use AOI21X1  _1279_
timestamp 0
transform -1 0 6670 0 1 270
box -6 -8 86 268
use AOI21X1  _1280_
timestamp 0
transform -1 0 6190 0 1 270
box -6 -8 86 268
use OAI21X1  _1281_
timestamp 0
transform -1 0 5970 0 -1 270
box -6 -8 86 268
use NAND3X1  _1282_
timestamp 0
transform -1 0 5670 0 -1 270
box -6 -8 86 268
use INVX1  _1283_
timestamp 0
transform 1 0 5490 0 1 270
box -6 -8 46 268
use NAND3X1  _1284_
timestamp 0
transform -1 0 6470 0 -1 270
box -6 -8 86 268
use OAI21X1  _1285_
timestamp 0
transform -1 0 6130 0 -1 270
box -6 -8 86 268
use NAND3X1  _1286_
timestamp 0
transform -1 0 6030 0 1 270
box -6 -8 86 268
use NAND3X1  _1287_
timestamp 0
transform 1 0 5270 0 -1 270
box -6 -8 86 268
use AOI21X1  _1288_
timestamp 0
transform -1 0 5690 0 1 270
box -6 -8 86 268
use AOI21X1  _1289_
timestamp 0
transform -1 0 5510 0 -1 270
box -6 -8 86 268
use OAI21X1  _1290_
timestamp 0
transform -1 0 5410 0 1 270
box -6 -8 86 268
use AOI21X1  _1291_
timestamp 0
transform -1 0 5390 0 -1 790
box -6 -8 86 268
use NAND3X1  _1292_
timestamp 0
transform 1 0 5470 0 -1 790
box -6 -8 86 268
use NAND2X1  _1293_
timestamp 0
transform 1 0 4350 0 -1 1830
box -6 -8 66 268
use OAI22X1  _1294_
timestamp 0
transform 1 0 4270 0 1 1830
box -6 -8 106 268
use INVX1  _1295_
timestamp 0
transform -1 0 4790 0 1 1310
box -6 -8 46 268
use INVX1  _1296_
timestamp 0
transform -1 0 4790 0 -1 1830
box -6 -8 46 268
use INVX1  _1297_
timestamp 0
transform 1 0 5750 0 -1 270
box -6 -8 46 268
use AOI21X1  _1298_
timestamp 0
transform -1 0 5870 0 1 270
box -6 -8 86 268
use NAND2X1  _1299_
timestamp 0
transform 1 0 5970 0 -1 1310
box -6 -8 66 268
use INVX1  _1300_
timestamp 0
transform 1 0 6430 0 -1 790
box -6 -8 46 268
use AOI21X1  _1301_
timestamp 0
transform -1 0 6650 0 -1 790
box -6 -8 86 268
use NAND2X1  _1302_
timestamp 0
transform -1 0 4470 0 -1 2870
box -6 -8 66 268
use INVX1  _1303_
timestamp 0
transform 1 0 5510 0 -1 2870
box -6 -8 46 268
use AND2X2  _1304_
timestamp 0
transform -1 0 4970 0 -1 2870
box -6 -8 86 268
use NAND2X1  _1305_
timestamp 0
transform 1 0 5210 0 -1 2870
box -6 -8 66 268
use NAND2X1  _1306_
timestamp 0
transform 1 0 5130 0 1 2870
box -6 -8 66 268
use OAI21X1  _1307_
timestamp 0
transform 1 0 5430 0 1 2870
box -6 -8 86 268
use AOI21X1  _1308_
timestamp 0
transform 1 0 5810 0 -1 2870
box -6 -8 86 268
use INVX1  _1309_
timestamp 0
transform -1 0 4250 0 -1 3390
box -6 -8 46 268
use OAI21X1  _1310_
timestamp 0
transform 1 0 4830 0 1 2350
box -6 -8 86 268
use OAI21X1  _1311_
timestamp 0
transform -1 0 5430 0 -1 2870
box -6 -8 86 268
use AOI21X1  _1312_
timestamp 0
transform 1 0 5470 0 1 2350
box -6 -8 86 268
use OAI21X1  _1313_
timestamp 0
transform -1 0 5250 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1314_
timestamp 0
transform -1 0 6030 0 1 2350
box -6 -8 86 268
use NAND3X1  _1315_
timestamp 0
transform 1 0 5310 0 1 2350
box -6 -8 86 268
use NAND3X1  _1316_
timestamp 0
transform -1 0 5730 0 -1 2870
box -6 -8 86 268
use AOI21X1  _1317_
timestamp 0
transform 1 0 5670 0 -1 2350
box -6 -8 86 268
use NAND3X1  _1318_
timestamp 0
transform 1 0 5790 0 1 2350
box -6 -8 86 268
use NAND3X1  _1319_
timestamp 0
transform 1 0 5850 0 -1 2350
box -6 -8 86 268
use NAND3X1  _1320_
timestamp 0
transform 1 0 5630 0 1 2350
box -6 -8 86 268
use OAI21X1  _1321_
timestamp 0
transform 1 0 6110 0 1 2350
box -6 -8 86 268
use NAND3X1  _1322_
timestamp 0
transform 1 0 6290 0 1 2350
box -6 -8 86 268
use NAND2X1  _1323_
timestamp 0
transform 1 0 6270 0 -1 2350
box -6 -8 66 268
use INVX1  _1324_
timestamp 0
transform -1 0 6530 0 1 1830
box -6 -8 46 268
use AOI21X1  _1325_
timestamp 0
transform 1 0 6330 0 1 1830
box -6 -8 86 268
use NAND2X1  _1326_
timestamp 0
transform 1 0 4990 0 1 2870
box -6 -8 66 268
use NAND2X1  _1327_
timestamp 0
transform 1 0 4470 0 -1 3390
box -6 -8 66 268
use NAND3X1  _1328_
timestamp 0
transform 1 0 4210 0 1 2870
box -6 -8 86 268
use NAND2X1  _1329_
timestamp 0
transform -1 0 4430 0 1 2870
box -6 -8 66 268
use NAND2X1  _1330_
timestamp 0
transform 1 0 4510 0 1 2870
box -6 -8 66 268
use NAND3X1  _1331_
timestamp 0
transform 1 0 4670 0 1 2870
box -6 -8 86 268
use INVX1  _1332_
timestamp 0
transform 1 0 5130 0 -1 3390
box -6 -8 46 268
use AND2X2  _1333_
timestamp 0
transform 1 0 4490 0 -1 4950
box -6 -8 86 268
use NAND2X1  _1334_
timestamp 0
transform 1 0 4990 0 -1 3390
box -6 -8 66 268
use OAI21X1  _1335_
timestamp 0
transform 1 0 4030 0 1 2870
box -6 -8 86 268
use NAND3X1  _1336_
timestamp 0
transform 1 0 5410 0 -1 3390
box -6 -8 86 268
use NAND2X1  _1337_
timestamp 0
transform 1 0 5590 0 -1 3390
box -6 -8 66 268
use OAI21X1  _1338_
timestamp 0
transform 1 0 4990 0 1 2350
box -6 -8 86 268
use INVX1  _1339_
timestamp 0
transform -1 0 6090 0 -1 3910
box -6 -8 46 268
use NAND2X1  _1340_
timestamp 0
transform -1 0 4770 0 1 3910
box -6 -8 66 268
use INVX1  _1341_
timestamp 0
transform 1 0 3470 0 -1 3910
box -6 -8 46 268
use NAND3X1  _1342_
timestamp 0
transform 1 0 3590 0 -1 3910
box -6 -8 86 268
use NAND2X1  _1343_
timestamp 0
transform -1 0 3970 0 -1 3910
box -6 -8 66 268
use NAND2X1  _1344_
timestamp 0
transform -1 0 4350 0 -1 3910
box -6 -8 66 268
use NAND3X1  _1345_
timestamp 0
transform 1 0 4610 0 -1 3910
box -6 -8 86 268
use INVX1  _1346_
timestamp 0
transform 1 0 5330 0 1 3910
box -6 -8 46 268
use NAND3X1  _1347_
timestamp 0
transform 1 0 4370 0 1 3910
box -6 -8 86 268
use NAND2X1  _1348_
timestamp 0
transform 1 0 3750 0 -1 3910
box -6 -8 66 268
use NAND3X1  _1349_
timestamp 0
transform 1 0 5470 0 1 3910
box -6 -8 86 268
use NAND3X1  _1350_
timestamp 0
transform -1 0 6150 0 1 3390
box -6 -8 86 268
use AOI21X1  _1351_
timestamp 0
transform 1 0 5630 0 1 3910
box -6 -8 86 268
use AOI21X1  _1352_
timestamp 0
transform 1 0 4450 0 -1 3910
box -6 -8 86 268
use OAI21X1  _1353_
timestamp 0
transform 1 0 5570 0 -1 3910
box -6 -8 86 268
use NAND3X1  _1354_
timestamp 0
transform 1 0 6090 0 1 2870
box -6 -8 86 268
use AND2X2  _1355_
timestamp 0
transform 1 0 5750 0 -1 3390
box -6 -8 86 268
use NAND3X1  _1356_
timestamp 0
transform 1 0 6230 0 -1 3390
box -6 -8 86 268
use OAI21X1  _1357_
timestamp 0
transform 1 0 5730 0 -1 3910
box -6 -8 86 268
use NAND3X1  _1358_
timestamp 0
transform 1 0 6570 0 -1 3390
box -6 -8 86 268
use NAND3X1  _1359_
timestamp 0
transform -1 0 6390 0 -1 2870
box -6 -8 86 268
use AOI21X1  _1360_
timestamp 0
transform 1 0 6070 0 -1 1830
box -6 -8 86 268
use OAI21X1  _1361_
timestamp 0
transform 1 0 6150 0 1 1830
box -6 -8 86 268
use AOI21X1  _1362_
timestamp 0
transform -1 0 6470 0 -1 3390
box -6 -8 86 268
use AOI21X1  _1363_
timestamp 0
transform 1 0 5930 0 1 2870
box -6 -8 86 268
use OAI21X1  _1364_
timestamp 0
transform 1 0 5990 0 -1 2870
box -6 -8 86 268
use NAND3X1  _1365_
timestamp 0
transform -1 0 6530 0 1 2350
box -6 -8 86 268
use AND2X2  _1366_
timestamp 0
transform 1 0 6570 0 -1 2350
box -6 -8 86 268
use NAND3X1  _1367_
timestamp 0
transform 1 0 6270 0 1 2870
box -6 -8 86 268
use OAI21X1  _1368_
timestamp 0
transform 1 0 6150 0 -1 2870
box -6 -8 86 268
use NAND3X1  _1369_
timestamp 0
transform 1 0 6610 0 1 1830
box -6 -8 86 268
use NAND3X1  _1370_
timestamp 0
transform -1 0 6390 0 1 1310
box -6 -8 86 268
use AOI21X1  _1371_
timestamp 0
transform 1 0 6190 0 1 790
box -6 -8 86 268
use OAI21X1  _1372_
timestamp 0
transform 1 0 6270 0 -1 790
box -6 -8 86 268
use AOI21X1  _1373_
timestamp 0
transform 1 0 6670 0 1 5990
box -6 -8 86 268
use AOI21X1  _1374_
timestamp 0
transform -1 0 6490 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1375_
timestamp 0
transform -1 0 6310 0 -1 1830
box -6 -8 86 268
use AOI21X1  _1376_
timestamp 0
transform -1 0 6030 0 1 1310
box -6 -8 86 268
use INVX1  _1377_
timestamp 0
transform 1 0 6590 0 -1 1310
box -6 -8 46 268
use NAND3X1  _1378_
timestamp 0
transform -1 0 6550 0 1 1310
box -6 -8 86 268
use OAI21X1  _1379_
timestamp 0
transform -1 0 6490 0 -1 1830
box -6 -8 86 268
use AOI21X1  _1380_
timestamp 0
transform -1 0 6350 0 -1 1310
box -6 -8 86 268
use OAI21X1  _1381_
timestamp 0
transform -1 0 5890 0 -1 1310
box -6 -8 86 268
use AOI21X1  _1382_
timestamp 0
transform -1 0 6650 0 -1 270
box -6 -8 86 268
use OAI21X1  _1383_
timestamp 0
transform -1 0 6510 0 1 270
box -6 -8 86 268
use NAND3X1  _1384_
timestamp 0
transform -1 0 6510 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1385_
timestamp 0
transform -1 0 6210 0 1 1310
box -6 -8 86 268
use NAND3X1  _1386_
timestamp 0
transform -1 0 6190 0 -1 1310
box -6 -8 86 268
use NAND2X1  _1387_
timestamp 0
transform 1 0 5350 0 -1 1310
box -6 -8 66 268
use OAI21X1  _1388_
timestamp 0
transform 1 0 4790 0 1 1830
box -6 -8 86 268
use NOR2X1  _1389_
timestamp 0
transform -1 0 4690 0 1 1830
box -6 -8 66 268
use INVX1  _1390_
timestamp 0
transform -1 0 5110 0 1 1830
box -6 -8 46 268
use AOI21X1  _1391_
timestamp 0
transform 1 0 4470 0 1 1830
box -6 -8 86 268
use AOI22X1  _1392_
timestamp 0
transform 1 0 4090 0 1 1830
box -6 -8 106 268
use NAND2X1  _1393_
timestamp 0
transform 1 0 3930 0 1 3910
box -6 -8 66 268
use INVX1  _1394_
timestamp 0
transform -1 0 5230 0 1 1310
box -6 -8 46 268
use AND2X2  _1395_
timestamp 0
transform -1 0 5270 0 -1 1310
box -6 -8 86 268
use OAI22X1  _1396_
timestamp 0
transform -1 0 5110 0 -1 1310
box -6 -8 106 268
use AOI21X1  _1397_
timestamp 0
transform -1 0 6730 0 1 1310
box -6 -8 86 268
use OAI21X1  _1398_
timestamp 0
transform 1 0 6670 0 1 3390
box -6 -8 86 268
use NAND2X1  _1399_
timestamp 0
transform -1 0 6670 0 1 2350
box -6 -8 66 268
use INVX1  _1400_
timestamp 0
transform -1 0 6590 0 1 3390
box -6 -8 46 268
use INVX1  _1401_
timestamp 0
transform -1 0 6510 0 -1 2870
box -6 -8 46 268
use AOI21X1  _1402_
timestamp 0
transform -1 0 6670 0 -1 2870
box -6 -8 86 268
use AND2X2  _1403_
timestamp 0
transform -1 0 5850 0 1 2870
box -6 -8 86 268
use NAND2X1  _1404_
timestamp 0
transform -1 0 4190 0 1 3390
box -6 -8 66 268
use INVX1  _1405_
timestamp 0
transform 1 0 4970 0 1 3390
box -6 -8 46 268
use AND2X2  _1406_
timestamp 0
transform -1 0 4890 0 -1 3390
box -6 -8 86 268
use AND2X2  _1407_
timestamp 0
transform 1 0 4410 0 -1 4430
box -6 -8 86 268
use NAND2X1  _1408_
timestamp 0
transform -1 0 4830 0 -1 3910
box -6 -8 66 268
use NAND2X1  _1409_
timestamp 0
transform -1 0 4790 0 -1 4430
box -6 -8 66 268
use OAI21X1  _1410_
timestamp 0
transform -1 0 4930 0 1 3910
box -6 -8 86 268
use AOI21X1  _1411_
timestamp 0
transform -1 0 4990 0 -1 3910
box -6 -8 86 268
use OAI21X1  _1412_
timestamp 0
transform 1 0 4470 0 1 3390
box -6 -8 86 268
use OAI21X1  _1413_
timestamp 0
transform -1 0 4910 0 1 2870
box -6 -8 86 268
use AOI21X1  _1414_
timestamp 0
transform 1 0 4810 0 1 3390
box -6 -8 86 268
use AND2X2  _1415_
timestamp 0
transform 1 0 4630 0 -1 3390
box -6 -8 86 268
use OAI21X1  _1416_
timestamp 0
transform 1 0 5250 0 -1 3390
box -6 -8 86 268
use OAI21X1  _1417_
timestamp 0
transform 1 0 5270 0 1 3390
box -6 -8 86 268
use NAND3X1  _1418_
timestamp 0
transform 1 0 4650 0 1 3390
box -6 -8 86 268
use NAND3X1  _1419_
timestamp 0
transform 1 0 5070 0 -1 3910
box -6 -8 86 268
use NOR2X1  _1420_
timestamp 0
transform 1 0 4330 0 -1 3390
box -6 -8 66 268
use AOI21X1  _1421_
timestamp 0
transform 1 0 4290 0 1 3390
box -6 -8 86 268
use NAND3X1  _1422_
timestamp 0
transform 1 0 5430 0 1 3390
box -6 -8 86 268
use NAND3X1  _1423_
timestamp 0
transform 1 0 5750 0 1 3390
box -6 -8 86 268
use INVX1  _1424_
timestamp 0
transform 1 0 5290 0 1 2870
box -6 -8 46 268
use OAI21X1  _1425_
timestamp 0
transform 1 0 5590 0 1 2870
box -6 -8 86 268
use NAND3X1  _1426_
timestamp 0
transform 1 0 5590 0 1 3390
box -6 -8 86 268
use OAI21X1  _1427_
timestamp 0
transform 1 0 5110 0 1 3390
box -6 -8 86 268
use NAND3X1  _1428_
timestamp 0
transform -1 0 5990 0 1 3390
box -6 -8 86 268
use NAND2X1  _1429_
timestamp 0
transform 1 0 5790 0 1 3910
box -6 -8 66 268
use INVX1  _1430_
timestamp 0
transform 1 0 6250 0 1 3390
box -6 -8 46 268
use AOI21X1  _1431_
timestamp 0
transform -1 0 6450 0 1 3390
box -6 -8 86 268
use NAND2X1  _1432_
timestamp 0
transform 1 0 4930 0 -1 5470
box -6 -8 66 268
use NAND2X1  _1433_
timestamp 0
transform -1 0 4410 0 -1 4950
box -6 -8 66 268
use NAND3X1  _1434_
timestamp 0
transform 1 0 4750 0 1 4950
box -6 -8 86 268
use NAND2X1  _1435_
timestamp 0
transform -1 0 4710 0 -1 4950
box -6 -8 66 268
use NAND3X1  _1436_
timestamp 0
transform 1 0 4810 0 -1 4950
box -6 -8 86 268
use NAND3X1  _1437_
timestamp 0
transform 1 0 5090 0 1 4950
box -6 -8 86 268
use INVX1  _1438_
timestamp 0
transform 1 0 5250 0 -1 5470
box -6 -8 46 268
use AND2X2  _1439_
timestamp 0
transform 1 0 3190 0 1 4950
box -6 -8 86 268
use NAND2X1  _1440_
timestamp 0
transform -1 0 5030 0 -1 4950
box -6 -8 66 268
use OAI21X1  _1441_
timestamp 0
transform 1 0 4170 0 -1 4950
box -6 -8 86 268
use NAND3X1  _1442_
timestamp 0
transform 1 0 5430 0 1 4950
box -6 -8 86 268
use NAND2X1  _1443_
timestamp 0
transform 1 0 5590 0 1 4950
box -6 -8 66 268
use AOI21X1  _1444_
timestamp 0
transform 1 0 3730 0 -1 4430
box -6 -8 86 268
use NAND3X1  _1445_
timestamp 0
transform 1 0 3230 0 -1 4430
box -6 -8 86 268
use INVX1  _1446_
timestamp 0
transform -1 0 4030 0 -1 5470
box -6 -8 46 268
use NOR2X1  _1447_
timestamp 0
transform -1 0 4630 0 -1 4430
box -6 -8 66 268
use NAND3X1  _1448_
timestamp 0
transform 1 0 5030 0 -1 4430
box -6 -8 86 268
use AOI21X1  _1449_
timestamp 0
transform 1 0 4530 0 1 3910
box -6 -8 86 268
use OAI21X1  _1450_
timestamp 0
transform 1 0 5010 0 1 3910
box -6 -8 86 268
use OAI21X1  _1451_
timestamp 0
transform 1 0 4730 0 1 4430
box -6 -8 86 268
use NAND3X1  _1452_
timestamp 0
transform 1 0 5370 0 1 4430
box -6 -8 86 268
use AND2X2  _1453_
timestamp 0
transform -1 0 5810 0 1 4950
box -6 -8 86 268
use INVX1  _1454_
timestamp 0
transform 1 0 4230 0 1 4430
box -6 -8 46 268
use NAND2X1  _1455_
timestamp 0
transform 1 0 4070 0 1 4430
box -6 -8 66 268
use NOR2X1  _1456_
timestamp 0
transform -1 0 5490 0 -1 4950
box -6 -8 66 268
use INVX1  _1457_
timestamp 0
transform 1 0 5530 0 1 4430
box -6 -8 46 268
use OAI21X1  _1458_
timestamp 0
transform 1 0 5570 0 -1 4950
box -6 -8 86 268
use NAND3X1  _1459_
timestamp 0
transform 1 0 5690 0 -1 4430
box -6 -8 86 268
use AOI21X1  _1460_
timestamp 0
transform 1 0 5910 0 -1 3390
box -6 -8 86 268
use OAI21X1  _1461_
timestamp 0
transform 1 0 6070 0 -1 3390
box -6 -8 86 268
use NAND2X1  _1462_
timestamp 0
transform -1 0 5190 0 -1 4950
box -6 -8 66 268
use NAND3X1  _1463_
timestamp 0
transform 1 0 5350 0 -1 4430
box -6 -8 86 268
use AOI21X1  _1464_
timestamp 0
transform 1 0 5910 0 -1 4950
box -6 -8 86 268
use AOI21X1  _1465_
timestamp 0
transform 1 0 5210 0 1 4430
box -6 -8 86 268
use OAI21X1  _1466_
timestamp 0
transform 1 0 5810 0 1 4430
box -6 -8 86 268
use NAND3X1  _1467_
timestamp 0
transform 1 0 5930 0 1 3910
box -6 -8 86 268
use AND2X2  _1468_
timestamp 0
transform -1 0 6190 0 1 3910
box -6 -8 86 268
use NAND3X1  _1469_
timestamp 0
transform 1 0 5510 0 -1 4430
box -6 -8 86 268
use OAI21X1  _1470_
timestamp 0
transform 1 0 5970 0 1 4430
box -6 -8 86 268
use NAND3X1  _1471_
timestamp 0
transform -1 0 6110 0 -1 4430
box -6 -8 86 268
use NAND3X1  _1472_
timestamp 0
transform 1 0 6170 0 -1 3910
box -6 -8 86 268
use AOI21X1  _1473_
timestamp 0
transform 1 0 6430 0 1 2870
box -6 -8 86 268
use OAI21X1  _1474_
timestamp 0
transform -1 0 6690 0 1 2870
box -6 -8 86 268
use AOI21X1  _1475_
timestamp 0
transform 1 0 6190 0 -1 4430
box -6 -8 86 268
use AOI21X1  _1476_
timestamp 0
transform 1 0 5850 0 -1 4430
box -6 -8 86 268
use OAI21X1  _1477_
timestamp 0
transform 1 0 6450 0 1 3910
box -6 -8 86 268
use NAND3X1  _1478_
timestamp 0
transform -1 0 6590 0 -1 3910
box -6 -8 86 268
use NAND3X1  _1479_
timestamp 0
transform 1 0 6270 0 1 3910
box -6 -8 86 268
use OAI21X1  _1480_
timestamp 0
transform -1 0 6450 0 -1 4430
box -6 -8 86 268
use NAND3X1  _1481_
timestamp 0
transform 1 0 6610 0 1 3910
box -6 -8 86 268
use NAND3X1  _1482_
timestamp 0
transform 1 0 6670 0 -1 3910
box -6 -8 86 268
use INVX1  _1483_
timestamp 0
transform -1 0 6730 0 1 5470
box -6 -8 46 268
use AOI21X1  _1484_
timestamp 0
transform 1 0 6570 0 -1 1830
box -6 -8 86 268
use AOI21X1  _1485_
timestamp 0
transform -1 0 6770 0 -1 4430
box -6 -8 86 268
use AOI21X1  _1486_
timestamp 0
transform -1 0 6430 0 -1 3910
box -6 -8 86 268
use OAI21X1  _1487_
timestamp 0
transform -1 0 6610 0 -1 4430
box -6 -8 86 268
use NAND2X1  _1488_
timestamp 0
transform -1 0 4930 0 -1 4430
box -6 -8 66 268
use XOR2X1  _1489_
timestamp 0
transform 1 0 4050 0 -1 4430
box -6 -8 126 268
use OAI21X1  _1490_
timestamp 0
transform 1 0 4070 0 1 3910
box -6 -8 86 268
use INVX1  _1491_
timestamp 0
transform -1 0 5110 0 1 4430
box -6 -8 46 268
use AOI21X1  _1492_
timestamp 0
transform 1 0 4910 0 1 4430
box -6 -8 86 268
use INVX1  _1493_
timestamp 0
transform 1 0 6430 0 1 4430
box -6 -8 46 268
use AOI21X1  _1494_
timestamp 0
transform 1 0 6550 0 1 4430
box -6 -8 86 268
use NAND2X1  _1495_
timestamp 0
transform -1 0 5970 0 -1 3910
box -6 -8 66 268
use INVX1  _1496_
timestamp 0
transform 1 0 6330 0 -1 5470
box -6 -8 46 268
use INVX1  _1497_
timestamp 0
transform -1 0 6170 0 1 4430
box -6 -8 46 268
use AOI21X1  _1498_
timestamp 0
transform 1 0 6270 0 1 4430
box -6 -8 86 268
use AND2X2  _1499_
timestamp 0
transform 1 0 5230 0 -1 3910
box -6 -8 86 268
use NAND2X1  _1500_
timestamp 0
transform -1 0 4670 0 -1 5470
box -6 -8 66 268
use NAND2X1  _1501_
timestamp 0
transform 1 0 4150 0 1 5470
box -6 -8 66 268
use NOR2X1  _1502_
timestamp 0
transform 1 0 4870 0 1 5470
box -6 -8 66 268
use AOI22X1  _1503_
timestamp 0
transform -1 0 4850 0 -1 5470
box -6 -8 106 268
use NOR3X1  _1504_
timestamp 0
transform 1 0 5190 0 1 5470
box -6 -8 166 268
use INVX1  _1505_
timestamp 0
transform 1 0 4890 0 -1 5990
box -6 -8 46 268
use AND2X2  _1506_
timestamp 0
transform -1 0 4630 0 -1 5990
box -6 -8 86 268
use NAND2X1  _1507_
timestamp 0
transform 1 0 4590 0 1 5470
box -6 -8 66 268
use INVX1  _1508_
timestamp 0
transform -1 0 5090 0 1 5990
box -6 -8 46 268
use AOI21X1  _1509_
timestamp 0
transform 1 0 5190 0 -1 5990
box -6 -8 86 268
use AND2X2  _1510_
timestamp 0
transform 1 0 4930 0 1 4950
box -6 -8 86 268
use OAI21X1  _1511_
timestamp 0
transform 1 0 5250 0 1 4950
box -6 -8 86 268
use OAI21X1  _1512_
timestamp 0
transform -1 0 5450 0 -1 5470
box -6 -8 86 268
use NAND3X1  _1513_
timestamp 0
transform 1 0 5030 0 -1 5990
box -6 -8 86 268
use OAI21X1  _1514_
timestamp 0
transform 1 0 5010 0 1 5470
box -6 -8 86 268
use AOI22X1  _1515_
timestamp 0
transform 1 0 5070 0 -1 5470
box -6 -8 106 268
use NAND3X1  _1516_
timestamp 0
transform 1 0 5610 0 1 5470
box -6 -8 86 268
use NAND3X1  _1517_
timestamp 0
transform 1 0 5530 0 -1 5470
box -6 -8 86 268
use NAND2X1  _1518_
timestamp 0
transform 1 0 5170 0 1 3910
box -6 -8 66 268
use OAI21X1  _1519_
timestamp 0
transform 1 0 5410 0 -1 3910
box -6 -8 86 268
use NAND3X1  _1520_
timestamp 0
transform 1 0 5350 0 -1 5990
box -6 -8 86 268
use OAI21X1  _1521_
timestamp 0
transform 1 0 5430 0 1 5470
box -6 -8 86 268
use NAND3X1  _1522_
timestamp 0
transform 1 0 5530 0 -1 5990
box -6 -8 86 268
use NAND2X1  _1523_
timestamp 0
transform 1 0 5670 0 1 5990
box -6 -8 66 268
use AOI21X1  _1524_
timestamp 0
transform -1 0 5270 0 -1 4430
box -6 -8 86 268
use AOI21X1  _1525_
timestamp 0
transform -1 0 5990 0 1 4950
box -6 -8 86 268
use NAND2X1  _1526_
timestamp 0
transform 1 0 3690 0 -1 4950
box -6 -8 66 268
use AND2X2  _1527_
timestamp 0
transform 1 0 3190 0 -1 4950
box -6 -8 86 268
use OAI21X1  _1528_
timestamp 0
transform -1 0 4090 0 -1 4950
box -6 -8 86 268
use OAI21X1  _1529_
timestamp 0
transform 1 0 3530 0 -1 4950
box -6 -8 86 268
use NAND3X1  _1530_
timestamp 0
transform 1 0 3830 0 -1 4950
box -6 -8 86 268
use INVX1  _1531_
timestamp 0
transform 1 0 4630 0 1 4950
box -6 -8 46 268
use NAND2X1  _1532_
timestamp 0
transform -1 0 3690 0 1 4950
box -6 -8 66 268
use OAI22X1  _1533_
timestamp 0
transform -1 0 3990 0 1 4430
box -6 -8 106 268
use NAND3X1  _1534_
timestamp 0
transform -1 0 4530 0 1 4950
box -6 -8 86 268
use NAND2X1  _1535_
timestamp 0
transform -1 0 4530 0 -1 5470
box -6 -8 66 268
use XNOR2X1  _1536_
timestamp 0
transform 1 0 4110 0 -1 5470
box -6 -8 126 268
use INVX1  _1537_
timestamp 0
transform 1 0 4310 0 1 5470
box -6 -8 46 268
use NAND2X1  _1538_
timestamp 0
transform 1 0 4430 0 1 5470
box -6 -8 66 268
use NAND3X1  _1539_
timestamp 0
transform 1 0 4310 0 -1 5470
box -6 -8 86 268
use NAND2X1  _1540_
timestamp 0
transform 1 0 5710 0 -1 5470
box -6 -8 66 268
use NOR2X1  _1541_
timestamp 0
transform -1 0 5910 0 -1 5990
box -6 -8 66 268
use NOR2X1  _1542_
timestamp 0
transform -1 0 5330 0 -1 4950
box -6 -8 66 268
use OAI21X1  _1543_
timestamp 0
transform 1 0 5750 0 -1 4950
box -6 -8 86 268
use AOI21X1  _1544_
timestamp 0
transform -1 0 5850 0 1 5470
box -6 -8 86 268
use OAI21X1  _1545_
timestamp 0
transform -1 0 5770 0 -1 5990
box -6 -8 86 268
use AND2X2  _1546_
timestamp 0
transform 1 0 6150 0 1 5990
box -6 -8 86 268
use NAND3X1  _1547_
timestamp 0
transform 1 0 5930 0 1 5470
box -6 -8 86 268
use NAND2X1  _1548_
timestamp 0
transform -1 0 6050 0 -1 5990
box -6 -8 66 268
use NAND3X1  _1549_
timestamp 0
transform 1 0 6330 0 1 5990
box -6 -8 86 268
use NAND3X1  _1550_
timestamp 0
transform -1 0 6390 0 -1 5990
box -6 -8 86 268
use AOI21X1  _1551_
timestamp 0
transform 1 0 5650 0 1 4430
box -6 -8 86 268
use OAI21X1  _1552_
timestamp 0
transform 1 0 6090 0 -1 4950
box -6 -8 86 268
use AOI22X1  _1553_
timestamp 0
transform 1 0 6130 0 -1 5990
box -6 -8 106 268
use NAND3X1  _1554_
timestamp 0
transform 1 0 5850 0 -1 5470
box -6 -8 86 268
use OAI21X1  _1555_
timestamp 0
transform -1 0 6170 0 1 4950
box -6 -8 86 268
use AOI21X1  _1556_
timestamp 0
transform 1 0 6010 0 -1 5470
box -6 -8 86 268
use OAI21X1  _1557_
timestamp 0
transform -1 0 6250 0 -1 5470
box -6 -8 86 268
use AOI21X1  _1558_
timestamp 0
transform 1 0 6450 0 1 4950
box -6 -8 86 268
use NAND3X1  _1559_
timestamp 0
transform 1 0 6630 0 -1 5990
box -6 -8 86 268
use OAI21X1  _1560_
timestamp 0
transform 1 0 6090 0 1 5470
box -6 -8 86 268
use AOI21X1  _1561_
timestamp 0
transform -1 0 6710 0 -1 5470
box -6 -8 86 268
use OAI21X1  _1562_
timestamp 0
transform -1 0 6690 0 1 4950
box -6 -8 86 268
use AOI21X1  _1563_
timestamp 0
transform -1 0 6530 0 -1 5470
box -6 -8 86 268
use AOI21X1  _1564_
timestamp 0
transform 1 0 6270 0 1 4950
box -6 -8 86 268
use OAI22X1  _1565_
timestamp 0
transform 1 0 6410 0 -1 4950
box -6 -8 106 268
use NAND2X1  _1566_
timestamp 0
transform -1 0 6650 0 -1 4950
box -6 -8 66 268
use XNOR2X1  _1567_
timestamp 0
transform -1 0 4630 0 1 4430
box -6 -8 126 268
use NAND2X1  _1568_
timestamp 0
transform 1 0 4230 0 1 3910
box -6 -8 66 268
use OAI21X1  _1569_
timestamp 0
transform -1 0 4330 0 -1 4430
box -6 -8 86 268
use NAND2X1  _1570_
timestamp 0
transform -1 0 3850 0 1 3910
box -6 -8 66 268
use OAI21X1  _1571_
timestamp 0
transform 1 0 6250 0 -1 4950
box -6 -8 86 268
use NOR2X1  _1572_
timestamp 0
transform -1 0 4410 0 1 4430
box -6 -8 66 268
use AOI21X1  _1573_
timestamp 0
transform -1 0 3810 0 1 4430
box -6 -8 86 268
use AOI21X1  _1574_
timestamp 0
transform 1 0 6470 0 -1 5990
box -6 -8 86 268
use OAI21X1  _1575_
timestamp 0
transform 1 0 6490 0 1 5990
box -6 -8 86 268
use NAND2X1  _1576_
timestamp 0
transform 1 0 5530 0 1 5990
box -6 -8 66 268
use INVX1  _1577_
timestamp 0
transform -1 0 5550 0 -1 6510
box -6 -8 46 268
use AOI21X1  _1578_
timestamp 0
transform -1 0 6050 0 1 5990
box -6 -8 86 268
use OAI21X1  _1579_
timestamp 0
transform -1 0 4810 0 -1 5990
box -6 -8 86 268
use INVX1  _1580_
timestamp 0
transform 1 0 4430 0 -1 5990
box -6 -8 46 268
use NAND2X1  _1581_
timestamp 0
transform -1 0 3110 0 -1 5470
box -6 -8 66 268
use AOI22X1  _1582_
timestamp 0
transform -1 0 2970 0 -1 5990
box -6 -8 106 268
use NAND2X1  _1583_
timestamp 0
transform -1 0 2970 0 1 5470
box -6 -8 66 268
use NOR2X1  _1584_
timestamp 0
transform -1 0 3110 0 1 5470
box -6 -8 66 268
use NOR3X1  _1585_
timestamp 0
transform 1 0 3230 0 -1 5990
box -6 -8 166 268
use INVX1  _1586_
timestamp 0
transform 1 0 2730 0 1 5990
box -6 -8 46 268
use INVX1  _1587_
timestamp 0
transform 1 0 2850 0 1 5990
box -6 -8 46 268
use INVX1  _1588_
timestamp 0
transform -1 0 2070 0 1 5470
box -6 -8 46 268
use NAND2X1  _1589_
timestamp 0
transform -1 0 2770 0 -1 5990
box -6 -8 66 268
use AOI21X1  _1590_
timestamp 0
transform 1 0 2970 0 1 5990
box -6 -8 86 268
use NOR2X1  _1591_
timestamp 0
transform 1 0 3950 0 1 4950
box -6 -8 66 268
use OAI21X1  _1592_
timestamp 0
transform -1 0 3850 0 1 4950
box -6 -8 86 268
use OAI21X1  _1593_
timestamp 0
transform -1 0 3870 0 -1 5990
box -6 -8 86 268
use NAND3X1  _1594_
timestamp 0
transform 1 0 3150 0 1 5990
box -6 -8 86 268
use OAI21X1  _1595_
timestamp 0
transform 1 0 3050 0 -1 5990
box -6 -8 86 268
use AND2X2  _1596_
timestamp 0
transform -1 0 4170 0 1 4950
box -6 -8 86 268
use AOI21X1  _1597_
timestamp 0
transform -1 0 4350 0 1 4950
box -6 -8 86 268
use NAND3X1  _1598_
timestamp 0
transform 1 0 4110 0 -1 5990
box -6 -8 86 268
use NAND3X1  _1599_
timestamp 0
transform -1 0 4350 0 -1 5990
box -6 -8 86 268
use NAND3X1  _1600_
timestamp 0
transform 1 0 3630 0 -1 5990
box -6 -8 86 268
use OAI21X1  _1601_
timestamp 0
transform 1 0 3950 0 -1 5990
box -6 -8 86 268
use NAND3X1  _1602_
timestamp 0
transform -1 0 4010 0 1 5990
box -6 -8 86 268
use NAND2X1  _1603_
timestamp 0
transform 1 0 4870 0 -1 6510
box -6 -8 66 268
use INVX1  _1604_
timestamp 0
transform 1 0 3710 0 -1 5470
box -6 -8 46 268
use OAI21X1  _1605_
timestamp 0
transform 1 0 3550 0 -1 5470
box -6 -8 86 268
use INVX1  _1606_
timestamp 0
transform 1 0 1450 0 1 5470
box -6 -8 46 268
use AND2X2  _1607_
timestamp 0
transform -1 0 3470 0 -1 5470
box -6 -8 86 268
use AND2X2  _1608_
timestamp 0
transform -1 0 2830 0 1 5470
box -6 -8 86 268
use AOI22X1  _1609_
timestamp 0
transform 1 0 3210 0 -1 5470
box -6 -8 106 268
use OAI21X1  _1610_
timestamp 0
transform -1 0 2510 0 1 5470
box -6 -8 86 268
use AOI21X1  _1611_
timestamp 0
transform -1 0 2670 0 1 5470
box -6 -8 86 268
use NAND2X1  _1612_
timestamp 0
transform 1 0 1590 0 1 5470
box -6 -8 66 268
use AND2X2  _1613_
timestamp 0
transform 1 0 3330 0 1 5470
box -6 -8 86 268
use NAND2X1  _1614_
timestamp 0
transform 1 0 3470 0 -1 5990
box -6 -8 66 268
use NAND2X1  _1615_
timestamp 0
transform 1 0 3850 0 -1 5470
box -6 -8 66 268
use NAND2X1  _1616_
timestamp 0
transform 1 0 3190 0 1 5470
box -6 -8 66 268
use NAND3X1  _1617_
timestamp 0
transform -1 0 3730 0 1 5470
box -6 -8 86 268
use NAND2X1  _1618_
timestamp 0
transform 1 0 4270 0 -1 6510
box -6 -8 66 268
use NAND2X1  _1619_
timestamp 0
transform -1 0 4770 0 -1 6510
box -6 -8 66 268
use NAND3X1  _1620_
timestamp 0
transform 1 0 3830 0 1 5470
box -6 -8 86 268
use NAND2X1  _1621_
timestamp 0
transform 1 0 3490 0 1 5470
box -6 -8 66 268
use NAND2X1  _1622_
timestamp 0
transform 1 0 3990 0 1 5470
box -6 -8 66 268
use NAND3X1  _1623_
timestamp 0
transform 1 0 5030 0 -1 6510
box -6 -8 86 268
use NAND3X1  _1624_
timestamp 0
transform 1 0 5970 0 -1 6510
box -6 -8 86 268
use OAI21X1  _1625_
timestamp 0
transform 1 0 5810 0 1 5990
box -6 -8 86 268
use AOI21X1  _1626_
timestamp 0
transform 1 0 4270 0 1 5990
box -6 -8 86 268
use NOR2X1  _1627_
timestamp 0
transform -1 0 4630 0 -1 6510
box -6 -8 66 268
use OAI21X1  _1628_
timestamp 0
transform 1 0 4890 0 1 5990
box -6 -8 86 268
use NAND3X1  _1629_
timestamp 0
transform 1 0 6310 0 -1 6510
box -6 -8 86 268
use NAND3X1  _1630_
timestamp 0
transform -1 0 5890 0 -1 6510
box -6 -8 86 268
use OAI21X1  _1631_
timestamp 0
transform 1 0 4730 0 1 5990
box -6 -8 86 268
use NAND3X1  _1632_
timestamp 0
transform 1 0 5650 0 -1 6510
box -6 -8 86 268
use NAND3X1  _1633_
timestamp 0
transform 1 0 6470 0 -1 6510
box -6 -8 86 268
use NOR3X1  _1634_
timestamp 0
transform 1 0 6250 0 1 5470
box -6 -8 166 268
use AOI21X1  _1635_
timestamp 0
transform -1 0 6590 0 1 5470
box -6 -8 86 268
use AOI21X1  _1636_
timestamp 0
transform 1 0 5170 0 1 5990
box -6 -8 86 268
use AOI21X1  _1637_
timestamp 0
transform -1 0 6210 0 -1 6510
box -6 -8 86 268
use OAI21X1  _1638_
timestamp 0
transform 1 0 5350 0 1 5990
box -6 -8 86 268
use NAND2X1  _1639_
timestamp 0
transform 1 0 4730 0 1 5470
box -6 -8 66 268
use AND2X2  _1640_
timestamp 0
transform 1 0 3570 0 -1 4430
box -6 -8 86 268
use OAI21X1  _1641_
timestamp 0
transform 1 0 3410 0 -1 4430
box -6 -8 86 268
use OAI21X1  _1642_
timestamp 0
transform 1 0 3610 0 1 3910
box -6 -8 86 268
use INVX1  _1643_
timestamp 0
transform 1 0 2270 0 1 3910
box -6 -8 46 268
use OAI21X1  _1644_
timestamp 0
transform -1 0 3310 0 1 4430
box -6 -8 86 268
use AOI21X1  _1645_
timestamp 0
transform -1 0 5430 0 -1 6510
box -6 -8 86 268
use OAI21X1  _1646_
timestamp 0
transform -1 0 5270 0 -1 6510
box -6 -8 86 268
use NAND2X1  _1647_
timestamp 0
transform 1 0 3790 0 1 5990
box -6 -8 66 268
use INVX1  _1648_
timestamp 0
transform -1 0 3850 0 -1 6510
box -6 -8 46 268
use AND2X2  _1649_
timestamp 0
transform -1 0 4170 0 1 5990
box -6 -8 86 268
use INVX1  _1650_
timestamp 0
transform -1 0 3530 0 1 5990
box -6 -8 46 268
use AOI21X1  _1651_
timestamp 0
transform -1 0 3690 0 1 5990
box -6 -8 86 268
use OAI21X1  _1652_
timestamp 0
transform -1 0 2650 0 1 5990
box -6 -8 86 268
use NAND2X1  _1653_
timestamp 0
transform 1 0 2570 0 -1 5990
box -6 -8 66 268
use INVX1  _1654_
timestamp 0
transform -1 0 2470 0 -1 5990
box -6 -8 46 268
use AOI22X1  _1655_
timestamp 0
transform -1 0 2330 0 -1 5470
box -6 -8 106 268
use INVX1  _1656_
timestamp 0
transform 1 0 1750 0 1 5470
box -6 -8 46 268
use AND2X2  _1657_
timestamp 0
transform -1 0 2190 0 -1 4950
box -6 -8 86 268
use NAND2X1  _1658_
timestamp 0
transform 1 0 1870 0 1 5470
box -6 -8 66 268
use NAND3X1  _1659_
timestamp 0
transform -1 0 2170 0 -1 5990
box -6 -8 86 268
use NAND2X1  _1660_
timestamp 0
transform -1 0 2350 0 1 5470
box -6 -8 66 268
use NOR2X1  _1661_
timestamp 0
transform 1 0 2150 0 1 5470
box -6 -8 66 268
use OAI21X1  _1662_
timestamp 0
transform 1 0 2270 0 -1 5990
box -6 -8 86 268
use NAND3X1  _1663_
timestamp 0
transform -1 0 2050 0 1 5990
box -6 -8 86 268
use INVX1  _1664_
timestamp 0
transform -1 0 1710 0 1 5990
box -6 -8 46 268
use NOR3X1  _1665_
timestamp 0
transform -1 0 1670 0 -1 5990
box -6 -8 166 268
use AOI21X1  _1666_
timestamp 0
transform -1 0 1990 0 -1 5990
box -6 -8 86 268
use OAI21X1  _1667_
timestamp 0
transform 1 0 1510 0 1 5990
box -6 -8 86 268
use AOI21X1  _1668_
timestamp 0
transform 1 0 2070 0 -1 6510
box -6 -8 86 268
use INVX1  _1669_
timestamp 0
transform 1 0 2390 0 -1 6510
box -6 -8 46 268
use OAI21X1  _1670_
timestamp 0
transform 1 0 1350 0 1 5990
box -6 -8 86 268
use NAND3X1  _1671_
timestamp 0
transform -1 0 1890 0 1 5990
box -6 -8 86 268
use AOI21X1  _1672_
timestamp 0
transform 1 0 1890 0 -1 6510
box -6 -8 86 268
use INVX1  _1673_
timestamp 0
transform -1 0 130 0 -1 5470
box -6 -8 46 268
use XOR2X1  _1674_
timestamp 0
transform -1 0 230 0 1 5470
box -6 -8 126 268
use OR2X2  _1675_
timestamp 0
transform 1 0 90 0 -1 6510
box -6 -8 86 268
use NAND2X1  _1676_
timestamp 0
transform 1 0 250 0 -1 6510
box -6 -8 66 268
use NAND2X1  _1677_
timestamp 0
transform 1 0 410 0 -1 6510
box -6 -8 66 268
use OAI21X1  _1678_
timestamp 0
transform 1 0 2230 0 -1 6510
box -6 -8 86 268
use NAND3X1  _1679_
timestamp 0
transform -1 0 1810 0 -1 6510
box -6 -8 86 268
use NAND3X1  _1680_
timestamp 0
transform -1 0 1650 0 -1 6510
box -6 -8 86 268
use INVX1  _1681_
timestamp 0
transform 1 0 1270 0 -1 6510
box -6 -8 46 268
use NAND3X1  _1682_
timestamp 0
transform -1 0 1470 0 -1 6510
box -6 -8 86 268
use NAND3X1  _1683_
timestamp 0
transform 1 0 2670 0 -1 6510
box -6 -8 86 268
use NAND2X1  _1684_
timestamp 0
transform -1 0 2570 0 -1 6510
box -6 -8 66 268
use OAI21X1  _1685_
timestamp 0
transform -1 0 3390 0 1 5990
box -6 -8 86 268
use NAND3X1  _1686_
timestamp 0
transform 1 0 3950 0 -1 6510
box -6 -8 86 268
use OAI21X1  _1687_
timestamp 0
transform -1 0 4490 0 -1 6510
box -6 -8 86 268
use NAND3X1  _1688_
timestamp 0
transform 1 0 2830 0 -1 6510
box -6 -8 86 268
use NAND2X1  _1689_
timestamp 0
transform -1 0 3070 0 -1 6510
box -6 -8 66 268
use NAND3X1  _1690_
timestamp 0
transform -1 0 3230 0 -1 6510
box -6 -8 86 268
use NAND3X1  _1691_
timestamp 0
transform -1 0 4190 0 -1 6510
box -6 -8 86 268
use INVX1  _1692_
timestamp 0
transform -1 0 4650 0 1 5990
box -6 -8 46 268
use AOI21X1  _1693_
timestamp 0
transform -1 0 4510 0 1 5990
box -6 -8 86 268
use AOI21X1  _1694_
timestamp 0
transform 1 0 3310 0 -1 6510
box -6 -8 86 268
use AOI21X1  _1695_
timestamp 0
transform -1 0 3730 0 -1 6510
box -6 -8 86 268
use OAI21X1  _1696_
timestamp 0
transform 1 0 3470 0 -1 6510
box -6 -8 86 268
use NAND2X1  _1697_
timestamp 0
transform -1 0 3550 0 1 4950
box -6 -8 66 268
use AND2X2  _1698_
timestamp 0
transform -1 0 2990 0 1 4430
box -6 -8 86 268
use NOR2X1  _1699_
timestamp 0
transform 1 0 3070 0 1 4430
box -6 -8 66 268
use OAI21X1  _1700_
timestamp 0
transform -1 0 2990 0 -1 4430
box -6 -8 86 268
use OAI21X1  _1701_
timestamp 0
transform 1 0 2650 0 1 3910
box -6 -8 86 268
use NAND2X1  _1702_
timestamp 0
transform 1 0 3070 0 -1 4430
box -6 -8 66 268
use NOR2X1  _1703_
timestamp 0
transform 1 0 3390 0 1 4430
box -6 -8 66 268
use NAND3X1  _1704_
timestamp 0
transform -1 0 3630 0 1 4430
box -6 -8 86 268
use NAND2X1  _1705_
timestamp 0
transform -1 0 3410 0 1 4950
box -6 -8 66 268
use AOI22X1  _1706_
timestamp 0
transform 1 0 3350 0 -1 4950
box -6 -8 106 268
use NAND2X1  _1707_
timestamp 0
transform -1 0 3110 0 -1 4950
box -6 -8 66 268
use OAI21X1  _1708_
timestamp 0
transform -1 0 2490 0 1 5990
box -6 -8 86 268
use NAND2X1  _1709_
timestamp 0
transform 1 0 1130 0 -1 6510
box -6 -8 66 268
use OAI21X1  _1710_
timestamp 0
transform 1 0 110 0 1 5990
box -6 -8 86 268
use OAI21X1  _1711_
timestamp 0
transform 1 0 1750 0 -1 5990
box -6 -8 86 268
use NAND2X1  _1712_
timestamp 0
transform 1 0 2390 0 1 4950
box -6 -8 66 268
use AOI21X1  _1713_
timestamp 0
transform -1 0 2310 0 1 4950
box -6 -8 86 268
use NAND2X1  _1714_
timestamp 0
transform -1 0 2330 0 -1 4950
box -6 -8 66 268
use NAND2X1  _1715_
timestamp 0
transform 1 0 2070 0 1 4950
box -6 -8 66 268
use NOR2X1  _1716_
timestamp 0
transform 1 0 1970 0 -1 4950
box -6 -8 66 268
use NOR2X1  _1717_
timestamp 0
transform 1 0 1730 0 1 4950
box -6 -8 66 268
use XNOR2X1  _1718_
timestamp 0
transform 1 0 1810 0 -1 5470
box -6 -8 126 268
use NOR2X1  _1719_
timestamp 0
transform -1 0 1250 0 -1 5990
box -6 -8 66 268
use OAI21X1  _1720_
timestamp 0
transform -1 0 1410 0 -1 5990
box -6 -8 86 268
use INVX1  _1721_
timestamp 0
transform -1 0 810 0 1 5470
box -6 -8 46 268
use INVX1  _1722_
timestamp 0
transform 1 0 270 0 1 4950
box -6 -8 46 268
use NAND2X1  _1723_
timestamp 0
transform 1 0 310 0 1 5470
box -6 -8 66 268
use NAND2X1  _1724_
timestamp 0
transform 1 0 270 0 -1 5990
box -6 -8 66 268
use OR2X2  _1725_
timestamp 0
transform -1 0 190 0 -1 5990
box -6 -8 86 268
use NAND2X1  _1726_
timestamp 0
transform 1 0 410 0 -1 5990
box -6 -8 66 268
use OAI21X1  _1727_
timestamp 0
transform -1 0 630 0 -1 5990
box -6 -8 86 268
use OR2X2  _1728_
timestamp 0
transform -1 0 1090 0 -1 5990
box -6 -8 86 268
use INVX1  _1729_
timestamp 0
transform 1 0 710 0 -1 5990
box -6 -8 46 268
use NAND3X1  _1730_
timestamp 0
transform -1 0 910 0 -1 5990
box -6 -8 86 268
use NAND3X1  _1731_
timestamp 0
transform 1 0 290 0 1 5990
box -6 -8 86 268
use NAND2X1  _1732_
timestamp 0
transform 1 0 450 0 1 5990
box -6 -8 66 268
use NAND3X1  _1733_
timestamp 0
transform 1 0 550 0 -1 6510
box -6 -8 86 268
use NAND3X1  _1734_
timestamp 0
transform 1 0 730 0 1 5990
box -6 -8 86 268
use INVX1  _1735_
timestamp 0
transform -1 0 1050 0 -1 6510
box -6 -8 46 268
use INVX1  _1736_
timestamp 0
transform -1 0 630 0 1 5990
box -6 -8 46 268
use INVX1  _1737_
timestamp 0
transform 1 0 730 0 -1 6510
box -6 -8 46 268
use OAI21X1  _1738_
timestamp 0
transform 1 0 850 0 -1 6510
box -6 -8 86 268
use NAND3X1  _1739_
timestamp 0
transform 1 0 1190 0 1 5990
box -6 -8 86 268
use INVX1  _1740_
timestamp 0
transform -1 0 2330 0 1 5990
box -6 -8 46 268
use NAND2X1  _1741_
timestamp 0
transform -1 0 1110 0 1 5990
box -6 -8 66 268
use NAND2X1  _1742_
timestamp 0
transform -1 0 2190 0 1 5990
box -6 -8 66 268
use AND2X2  _1743_
timestamp 0
transform 1 0 2890 0 -1 5470
box -6 -8 86 268
use XNOR2X1  _1744_
timestamp 0
transform -1 0 3090 0 1 4950
box -6 -8 126 268
use OAI21X1  _1745_
timestamp 0
transform 1 0 2730 0 1 4430
box -6 -8 86 268
use INVX1  _1746_
timestamp 0
transform -1 0 2630 0 -1 5470
box -6 -8 46 268
use AND2X2  _1747_
timestamp 0
transform -1 0 2890 0 1 4950
box -6 -8 86 268
use AOI21X1  _1748_
timestamp 0
transform 1 0 890 0 1 5990
box -6 -8 86 268
use OAI22X1  _1749_
timestamp 0
transform -1 0 1990 0 1 4950
box -6 -8 106 268
use INVX1  _1750_
timestamp 0
transform -1 0 2170 0 1 4430
box -6 -8 46 268
use OAI21X1  _1751_
timestamp 0
transform -1 0 2050 0 1 4430
box -6 -8 86 268
use NOR2X1  _1752_
timestamp 0
transform 1 0 1890 0 -1 4430
box -6 -8 66 268
use NAND2X1  _1753_
timestamp 0
transform -1 0 1730 0 1 4430
box -6 -8 66 268
use AND2X2  _1754_
timestamp 0
transform 1 0 1810 0 1 4430
box -6 -8 86 268
use XOR2X1  _1755_
timestamp 0
transform -1 0 1510 0 1 4950
box -6 -8 126 268
use XNOR2X1  _1756_
timestamp 0
transform -1 0 650 0 1 4950
box -6 -8 126 268
use AOI21X1  _1757_
timestamp 0
transform 1 0 450 0 1 5470
box -6 -8 86 268
use INVX1  _1758_
timestamp 0
transform -1 0 510 0 -1 5470
box -6 -8 46 268
use NAND3X1  _1759_
timestamp 0
transform 1 0 610 0 1 5470
box -6 -8 86 268
use NAND3X1  _1760_
timestamp 0
transform 1 0 590 0 -1 5470
box -6 -8 86 268
use INVX1  _1761_
timestamp 0
transform -1 0 1110 0 1 5470
box -6 -8 46 268
use OAI21X1  _1762_
timestamp 0
transform 1 0 890 0 1 5470
box -6 -8 86 268
use NAND2X1  _1763_
timestamp 0
transform -1 0 990 0 -1 5470
box -6 -8 66 268
use XOR2X1  _1764_
timestamp 0
transform 1 0 2030 0 -1 5470
box -6 -8 126 268
use INVX1  _1765_
timestamp 0
transform -1 0 2730 0 1 4950
box -6 -8 46 268
use OAI21X1  _1766_
timestamp 0
transform 1 0 2530 0 1 4950
box -6 -8 86 268
use NOR2X1  _1767_
timestamp 0
transform 1 0 2590 0 -1 4950
box -6 -8 66 268
use AOI21X1  _1768_
timestamp 0
transform -1 0 2490 0 -1 4950
box -6 -8 86 268
use AOI22X1  _1769_
timestamp 0
transform -1 0 2530 0 1 4430
box -6 -8 106 268
use NAND2X1  _1770_
timestamp 0
transform 1 0 2290 0 -1 4430
box -6 -8 66 268
use NAND3X1  _1771_
timestamp 0
transform 1 0 2710 0 -1 5470
box -6 -8 86 268
use AOI21X1  _1772_
timestamp 0
transform -1 0 2950 0 -1 4950
box -6 -8 86 268
use NAND2X1  _1773_
timestamp 0
transform 1 0 2430 0 -1 5470
box -6 -8 66 268
use OAI21X1  _1774_
timestamp 0
transform 1 0 1650 0 -1 5470
box -6 -8 86 268
use NOR2X1  _1775_
timestamp 0
transform 1 0 1590 0 1 4950
box -6 -8 66 268
use AOI21X1  _1776_
timestamp 0
transform 1 0 770 0 -1 5470
box -6 -8 86 268
use NAND2X1  _1777_
timestamp 0
transform -1 0 1290 0 1 4950
box -6 -8 66 268
use OAI21X1  _1778_
timestamp 0
transform -1 0 1790 0 -1 4430
box -6 -8 86 268
use XOR2X1  _1779_
timestamp 0
transform -1 0 1610 0 -1 4430
box -6 -8 126 268
use NAND2X1  _1780_
timestamp 0
transform 1 0 390 0 1 4950
box -6 -8 66 268
use OR2X2  _1781_
timestamp 0
transform 1 0 750 0 1 4950
box -6 -8 86 268
use NAND2X1  _1782_
timestamp 0
transform 1 0 350 0 -1 4950
box -6 -8 66 268
use NAND2X1  _1783_
timestamp 0
transform 1 0 490 0 -1 4950
box -6 -8 66 268
use NAND2X1  _1784_
timestamp 0
transform -1 0 710 0 -1 4950
box -6 -8 66 268
use OAI21X1  _1785_
timestamp 0
transform -1 0 870 0 -1 4950
box -6 -8 86 268
use OR2X2  _1786_
timestamp 0
transform 1 0 1110 0 -1 4950
box -6 -8 86 268
use NAND2X1  _1787_
timestamp 0
transform 1 0 970 0 -1 4950
box -6 -8 66 268
use AND2X2  _1788_
timestamp 0
transform 1 0 1430 0 -1 4950
box -6 -8 86 268
use XOR2X1  _1789_
timestamp 0
transform 1 0 1750 0 -1 4950
box -6 -8 126 268
use OAI21X1  _1790_
timestamp 0
transform -1 0 2350 0 1 4430
box -6 -8 86 268
use OAI21X1  _1791_
timestamp 0
transform -1 0 1670 0 -1 4950
box -6 -8 86 268
use OAI21X1  _1792_
timestamp 0
transform 1 0 1270 0 -1 4950
box -6 -8 86 268
use OAI21X1  _1793_
timestamp 0
transform -1 0 1010 0 1 4950
box -6 -8 86 268
use OAI21X1  _1794_
timestamp 0
transform 1 0 1510 0 1 4430
box -6 -8 86 268
use XOR2X1  _1795_
timestamp 0
transform -1 0 990 0 1 4430
box -6 -8 126 268
use XNOR2X1  _1796_
timestamp 0
transform 1 0 670 0 1 4430
box -6 -8 126 268
use INVX1  _1797_
timestamp 0
transform 1 0 1070 0 1 4430
box -6 -8 46 268
use NAND2X1  _1798_
timestamp 0
transform 1 0 1190 0 1 4430
box -6 -8 66 268
use NAND3X1  _1799_
timestamp 0
transform 1 0 1350 0 1 4430
box -6 -8 86 268
use AND2X2  _1800_
timestamp 0
transform -1 0 1950 0 1 3910
box -6 -8 86 268
use AOI22X1  _1801_
timestamp 0
transform 1 0 1690 0 1 3910
box -6 -8 106 268
use INVX1  _1802_
timestamp 0
transform 1 0 110 0 1 2350
box -6 -8 46 268
use INVX1  _1803_
timestamp 0
transform 1 0 990 0 1 3390
box -6 -8 46 268
use NAND3X1  _1804_
timestamp 0
transform -1 0 1190 0 1 3390
box -6 -8 86 268
use NAND2X1  _1805_
timestamp 0
transform 1 0 230 0 -1 4430
box -6 -8 66 268
use OAI21X1  _1806_
timestamp 0
transform 1 0 330 0 1 3910
box -6 -8 86 268
use INVX1  _1807_
timestamp 0
transform 1 0 230 0 -1 4950
box -6 -8 46 268
use NAND2X1  _1808_
timestamp 0
transform 1 0 510 0 1 4430
box -6 -8 66 268
use OAI21X1  _1809_
timestamp 0
transform 1 0 330 0 1 4430
box -6 -8 86 268
use INVX1  _1810_
timestamp 0
transform 1 0 90 0 -1 4430
box -6 -8 46 268
use NAND2X1  _1811_
timestamp 0
transform -1 0 1170 0 -1 4430
box -6 -8 66 268
use OAI21X1  _1812_
timestamp 0
transform 1 0 930 0 -1 4430
box -6 -8 86 268
use INVX1  _1813_
timestamp 0
transform 1 0 230 0 1 3390
box -6 -8 46 268
use NAND2X1  _1814_
timestamp 0
transform 1 0 910 0 1 3910
box -6 -8 66 268
use OAI21X1  _1815_
timestamp 0
transform 1 0 490 0 1 3910
box -6 -8 86 268
use NOR2X1  _1816_
timestamp 0
transform 1 0 1010 0 -1 3910
box -6 -8 66 268
use NOR2X1  _1817_
timestamp 0
transform -1 0 850 0 -1 4430
box -6 -8 66 268
use AOI21X1  _1818_
timestamp 0
transform 1 0 370 0 -1 4430
box -6 -8 86 268
use NAND2X1  _1819_
timestamp 0
transform -1 0 1150 0 1 4950
box -6 -8 66 268
use OAI21X1  _1820_
timestamp 0
transform -1 0 1330 0 -1 5470
box -6 -8 86 268
use NAND2X1  _1821_
timestamp 0
transform 1 0 90 0 -1 4950
box -6 -8 66 268
use OAI21X1  _1822_
timestamp 0
transform -1 0 1150 0 -1 5470
box -6 -8 86 268
use NAND2X1  _1823_
timestamp 0
transform 1 0 110 0 -1 3910
box -6 -8 66 268
use OAI21X1  _1824_
timestamp 0
transform 1 0 90 0 1 4950
box -6 -8 86 268
use INVX1  _1825_
timestamp 0
transform -1 0 1190 0 1 2870
box -6 -8 46 268
use OAI21X1  _1826_
timestamp 0
transform -1 0 1070 0 -1 2870
box -6 -8 86 268
use OAI21X1  _1827_
timestamp 0
transform 1 0 570 0 -1 2870
box -6 -8 86 268
use OAI21X1  _1828_
timestamp 0
transform 1 0 1810 0 -1 2870
box -6 -8 86 268
use OAI21X1  _1829_
timestamp 0
transform 1 0 1650 0 -1 2870
box -6 -8 86 268
use OAI21X1  _1830_
timestamp 0
transform -1 0 1550 0 -1 2870
box -6 -8 86 268
use OAI21X1  _1831_
timestamp 0
transform 1 0 990 0 1 2870
box -6 -8 86 268
use OAI21X1  _1832_
timestamp 0
transform -1 0 910 0 1 3390
box -6 -8 86 268
use OAI21X1  _1833_
timestamp 0
transform 1 0 650 0 1 3390
box -6 -8 86 268
use NAND2X1  _1834_
timestamp 0
transform -1 0 150 0 -1 2350
box -6 -8 66 268
use OAI21X1  _1835_
timestamp 0
transform -1 0 630 0 -1 2350
box -6 -8 86 268
use NOR2X1  _1836_
timestamp 0
transform 1 0 930 0 1 2350
box -6 -8 66 268
use AOI21X1  _1837_
timestamp 0
transform -1 0 850 0 1 2350
box -6 -8 86 268
use NOR2X1  _1838_
timestamp 0
transform 1 0 490 0 1 1830
box -6 -8 66 268
use AOI21X1  _1839_
timestamp 0
transform -1 0 450 0 -1 2350
box -6 -8 86 268
use NAND2X1  _1840_
timestamp 0
transform -1 0 150 0 1 1830
box -6 -8 66 268
use OAI21X1  _1841_
timestamp 0
transform -1 0 330 0 -1 1830
box -6 -8 86 268
use NAND2X1  _1842_
timestamp 0
transform -1 0 1290 0 -1 2350
box -6 -8 66 268
use OAI21X1  _1843_
timestamp 0
transform -1 0 1450 0 -1 2350
box -6 -8 86 268
use NAND2X1  _1844_
timestamp 0
transform 1 0 1910 0 -1 1310
box -6 -8 66 268
use OAI21X1  _1845_
timestamp 0
transform 1 0 2050 0 -1 1310
box -6 -8 86 268
use NAND2X1  _1846_
timestamp 0
transform -1 0 3050 0 -1 1310
box -6 -8 66 268
use OAI21X1  _1847_
timestamp 0
transform -1 0 3230 0 -1 1310
box -6 -8 86 268
use NAND2X1  _1848_
timestamp 0
transform -1 0 450 0 1 2350
box -6 -8 66 268
use OAI21X1  _1849_
timestamp 0
transform 1 0 230 0 1 2350
box -6 -8 86 268
use DFFPOSX1  _1850_
timestamp 0
transform 1 0 1810 0 1 1830
box -6 -8 246 268
use DFFPOSX1  _1851_
timestamp 0
transform 1 0 3050 0 -1 1830
box -6 -8 246 268
use DFFPOSX1  _1852_
timestamp 0
transform 1 0 3310 0 1 2350
box -6 -8 246 268
use DFFPOSX1  _1853_
timestamp 0
transform 1 0 1190 0 1 3390
box -6 -8 246 268
use DFFPOSX1  _1854_
timestamp 0
transform -1 0 3310 0 1 2350
box -6 -8 246 268
use DFFPOSX1  _1855_
timestamp 0
transform -1 0 3710 0 1 2870
box -6 -8 246 268
use DFFPOSX1  _1856_
timestamp 0
transform 1 0 2590 0 1 1830
box -6 -8 246 268
use DFFPOSX1  _1857_
timestamp 0
transform 1 0 2290 0 -1 2870
box -6 -8 246 268
use DFFPOSX1  _1858_
timestamp 0
transform -1 0 4030 0 -1 2870
box -6 -8 246 268
use DFFPOSX1  _1859_
timestamp 0
transform -1 0 3630 0 1 1830
box -6 -8 246 268
use DFFPOSX1  _1860_
timestamp 0
transform -1 0 3950 0 1 2870
box -6 -8 246 268
use DFFPOSX1  _1861_
timestamp 0
transform 1 0 1930 0 1 2350
box -6 -8 246 268
use DFFPOSX1  _1862_
timestamp 0
transform -1 0 3130 0 1 3390
box -6 -8 246 268
use DFFPOSX1  _1863_
timestamp 0
transform -1 0 3950 0 -1 3390
box -6 -8 246 268
use DFFPOSX1  _1864_
timestamp 0
transform -1 0 3790 0 1 3390
box -6 -8 246 268
use DFFPOSX1  _1865_
timestamp 0
transform -1 0 2190 0 1 3910
box -6 -8 246 268
use DFFPOSX1  _1866_
timestamp 0
transform 1 0 1990 0 -1 3910
box -6 -8 246 268
use DFFPOSX1  _1867_
timestamp 0
transform 1 0 2510 0 -1 3910
box -6 -8 246 268
use DFFPOSX1  _1868_
timestamp 0
transform 1 0 1850 0 -1 3390
box -6 -8 246 268
use DFFPOSX1  _1869_
timestamp 0
transform -1 0 930 0 -1 3910
box -6 -8 246 268
use DFFPOSX1  _1870_
timestamp 0
transform 1 0 2250 0 -1 2350
box -6 -8 246 268
use DFFPOSX1  _1871_
timestamp 0
transform 1 0 1430 0 1 2870
box -6 -8 246 268
use DFFPOSX1  _1872_
timestamp 0
transform 1 0 2030 0 -1 1830
box -6 -8 246 268
use DFFPOSX1  _1873_
timestamp 0
transform -1 0 2590 0 1 1830
box -6 -8 246 268
use DFFPOSX1  _1874_
timestamp 0
transform 1 0 3290 0 1 790
box -6 -8 246 268
use DFFPOSX1  _1875_
timestamp 0
transform 1 0 2590 0 1 1310
box -6 -8 246 268
use DFFPOSX1  _1876_
timestamp 0
transform 1 0 3830 0 -1 2350
box -6 -8 246 268
use DFFPOSX1  _1877_
timestamp 0
transform -1 0 4010 0 1 1830
box -6 -8 246 268
use DFFPOSX1  _1878_
timestamp 0
transform -1 0 3150 0 -1 3910
box -6 -8 246 268
use DFFPOSX1  _1879_
timestamp 0
transform 1 0 3970 0 -1 3910
box -6 -8 246 268
use DFFPOSX1  _1880_
timestamp 0
transform 1 0 3150 0 -1 3910
box -6 -8 246 268
use DFFPOSX1  _1881_
timestamp 0
transform -1 0 2550 0 1 3910
box -6 -8 246 268
use DFFPOSX1  _1882_
timestamp 0
transform 1 0 2590 0 -1 4430
box -6 -8 246 268
use DFFPOSX1  _1883_
timestamp 0
transform 1 0 2350 0 -1 4430
box -6 -8 246 268
use DFFPOSX1  _1884_
timestamp 0
transform -1 0 2190 0 -1 4430
box -6 -8 246 268
use DFFPOSX1  _1885_
timestamp 0
transform 1 0 1250 0 1 3910
box -6 -8 246 268
use DFFPOSX1  _1886_
timestamp 0
transform -1 0 250 0 1 3910
box -6 -8 246 268
use DFFPOSX1  _1887_
timestamp 0
transform -1 0 250 0 1 4430
box -6 -8 246 268
use DFFPOSX1  _1888_
timestamp 0
transform 1 0 1170 0 -1 4430
box -6 -8 246 268
use DFFPOSX1  _1889_
timestamp 0
transform 1 0 570 0 1 3910
box -6 -8 246 268
use DFFPOSX1  _1890_
timestamp 0
transform 1 0 450 0 -1 4430
box -6 -8 246 268
use DFFPOSX1  _1891_
timestamp 0
transform 1 0 1330 0 -1 5470
box -6 -8 246 268
use DFFPOSX1  _1892_
timestamp 0
transform 1 0 1110 0 1 5470
box -6 -8 246 268
use DFFPOSX1  _1893_
timestamp 0
transform -1 0 370 0 -1 5470
box -6 -8 246 268
use DFFPOSX1  _1894_
timestamp 0
transform 1 0 650 0 -1 2870
box -6 -8 246 268
use DFFPOSX1  _1895_
timestamp 0
transform 1 0 2050 0 -1 2870
box -6 -8 246 268
use DFFPOSX1  _1896_
timestamp 0
transform 1 0 1190 0 1 2870
box -6 -8 246 268
use DFFPOSX1  _1897_
timestamp 0
transform 1 0 450 0 -1 3910
box -6 -8 246 268
use DFFPOSX1  _1898_
timestamp 0
transform 1 0 630 0 -1 2350
box -6 -8 246 268
use DFFPOSX1  _1899_
timestamp 0
transform 1 0 450 0 1 2350
box -6 -8 246 268
use DFFPOSX1  _1900_
timestamp 0
transform 1 0 150 0 1 1830
box -6 -8 246 268
use DFFPOSX1  _1901_
timestamp 0
transform 1 0 330 0 -1 1830
box -6 -8 246 268
use DFFPOSX1  _1902_
timestamp 0
transform 1 0 1250 0 1 2350
box -6 -8 246 268
use DFFPOSX1  _1903_
timestamp 0
transform 1 0 2050 0 1 1310
box -6 -8 246 268
use DFFPOSX1  _1904_
timestamp 0
transform -1 0 3230 0 1 1310
box -6 -8 246 268
use DFFPOSX1  _1905_
timestamp 0
transform 1 0 250 0 -1 2870
box -6 -8 246 268
use DFFPOSX1  _1906_
timestamp 0
transform 1 0 10 0 -1 2870
box -6 -8 246 268
use DFFPOSX1  _1907_
timestamp 0
transform 1 0 410 0 -1 3390
box -6 -8 246 268
use DFFPOSX1  _1908_
timestamp 0
transform 1 0 650 0 -1 3390
box -6 -8 246 268
use DFFPOSX1  _1909_
timestamp 0
transform 1 0 1610 0 -1 3390
box -6 -8 246 268
use DFFPOSX1  _1910_
timestamp 0
transform 1 0 2250 0 -1 3390
box -6 -8 246 268
use BUFX2  _1911_
timestamp 0
transform -1 0 2810 0 -1 270
box -6 -8 66 268
use BUFX2  _1912_
timestamp 0
transform -1 0 150 0 -1 1830
box -6 -8 66 268
use BUFX2  _1913_
timestamp 0
transform 1 0 2450 0 -1 270
box -6 -8 66 268
use BUFX2  _1914_
timestamp 0
transform -1 0 170 0 1 2870
box -6 -8 66 268
use BUFX2  _1915_
timestamp 0
transform -1 0 150 0 1 3390
box -6 -8 66 268
use BUFX2  _1916_
timestamp 0
transform -1 0 2650 0 -1 270
box -6 -8 66 268
use BUFX2  _1917_
timestamp 0
transform -1 0 2590 0 1 1310
box -6 -8 66 268
use BUFX2  _1918_
timestamp 0
transform -1 0 310 0 1 2870
box -6 -8 66 268
use BUFX2  _1919_
timestamp 0
transform -1 0 150 0 -1 3390
box -6 -8 66 268
use BUFX2  BUFX2_insert0
timestamp 0
transform 1 0 3170 0 -1 2350
box -6 -8 66 268
use BUFX2  BUFX2_insert1
timestamp 0
transform 1 0 2870 0 -1 2350
box -6 -8 66 268
use BUFX2  BUFX2_insert2
timestamp 0
transform 1 0 3330 0 -1 3390
box -6 -8 66 268
use BUFX2  BUFX2_insert3
timestamp 0
transform 1 0 3310 0 -1 2870
box -6 -8 66 268
use BUFX2  BUFX2_insert4
timestamp 0
transform -1 0 2790 0 -1 3390
box -6 -8 66 268
use BUFX2  BUFX2_insert12
timestamp 0
transform 1 0 3590 0 -1 2350
box -6 -8 66 268
use BUFX2  BUFX2_insert13
timestamp 0
transform 1 0 90 0 1 1310
box -6 -8 66 268
use BUFX2  BUFX2_insert14
timestamp 0
transform 1 0 650 0 1 1830
box -6 -8 66 268
use BUFX2  BUFX2_insert15
timestamp 0
transform 1 0 3630 0 1 2350
box -6 -8 66 268
use BUFX2  BUFX2_insert16
timestamp 0
transform 1 0 850 0 1 2870
box -6 -8 66 268
use BUFX2  BUFX2_insert17
timestamp 0
transform 1 0 1170 0 -1 2870
box -6 -8 66 268
use BUFX2  BUFX2_insert18
timestamp 0
transform -1 0 290 0 -1 2350
box -6 -8 66 268
use BUFX2  BUFX2_insert19
timestamp 0
transform -1 0 1170 0 -1 1830
box -6 -8 66 268
use BUFX2  BUFX2_insert20
timestamp 0
transform -1 0 470 0 1 2870
box -6 -8 66 268
use BUFX2  BUFX2_insert21
timestamp 0
transform 1 0 3450 0 -1 2870
box -6 -8 66 268
use BUFX2  BUFX2_insert22
timestamp 0
transform -1 0 3230 0 -1 2870
box -6 -8 66 268
use BUFX2  BUFX2_insert23
timestamp 0
transform 1 0 3470 0 1 3910
box -6 -8 66 268
use BUFX2  BUFX2_insert24
timestamp 0
transform -1 0 3230 0 -1 3390
box -6 -8 66 268
use BUFX2  BUFX2_insert25
timestamp 0
transform -1 0 3370 0 1 3910
box -6 -8 66 268
use CLKBUF1  CLKBUF1_insert5
timestamp 0
transform -1 0 1250 0 1 3910
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert6
timestamp 0
transform 1 0 2110 0 1 3390
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert7
timestamp 0
transform 1 0 1070 0 1 2350
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert8
timestamp 0
transform -1 0 450 0 -1 3910
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert9
timestamp 0
transform 1 0 230 0 -1 3390
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert10
timestamp 0
transform 1 0 2730 0 -1 2870
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert11
timestamp 0
transform 1 0 1750 0 1 2350
box -6 -8 186 268
use FILL  FILL99450x15750
timestamp 0
transform -1 0 6650 0 -1 1310
box -6 -8 26 268
use FILL  FILL99450x66450
timestamp 0
transform 1 0 6630 0 1 4430
box -6 -8 26 268
use FILL  FILL99750x150
timestamp 0
transform -1 0 6670 0 -1 270
box -6 -8 26 268
use FILL  FILL99750x7950
timestamp 0
transform -1 0 6670 0 -1 790
box -6 -8 26 268
use FILL  FILL99750x15750
timestamp 0
transform -1 0 6670 0 -1 1310
box -6 -8 26 268
use FILL  FILL99750x23550
timestamp 0
transform -1 0 6670 0 -1 1830
box -6 -8 26 268
use FILL  FILL99750x31350
timestamp 0
transform -1 0 6670 0 -1 2350
box -6 -8 26 268
use FILL  FILL99750x46950
timestamp 0
transform -1 0 6670 0 -1 3390
box -6 -8 26 268
use FILL  FILL99750x66450
timestamp 0
transform 1 0 6650 0 1 4430
box -6 -8 26 268
use FILL  FILL99750x70350
timestamp 0
transform -1 0 6670 0 -1 4950
box -6 -8 26 268
use FILL  FILL100050x150
timestamp 0
transform -1 0 6690 0 -1 270
box -6 -8 26 268
use FILL  FILL100050x4050
timestamp 0
transform 1 0 6670 0 1 270
box -6 -8 26 268
use FILL  FILL100050x7950
timestamp 0
transform -1 0 6690 0 -1 790
box -6 -8 26 268
use FILL  FILL100050x15750
timestamp 0
transform -1 0 6690 0 -1 1310
box -6 -8 26 268
use FILL  FILL100050x23550
timestamp 0
transform -1 0 6690 0 -1 1830
box -6 -8 26 268
use FILL  FILL100050x31350
timestamp 0
transform -1 0 6690 0 -1 2350
box -6 -8 26 268
use FILL  FILL100050x35250
timestamp 0
transform 1 0 6670 0 1 2350
box -6 -8 26 268
use FILL  FILL100050x39150
timestamp 0
transform -1 0 6690 0 -1 2870
box -6 -8 26 268
use FILL  FILL100050x46950
timestamp 0
transform -1 0 6690 0 -1 3390
box -6 -8 26 268
use FILL  FILL100050x66450
timestamp 0
transform 1 0 6670 0 1 4430
box -6 -8 26 268
use FILL  FILL100050x70350
timestamp 0
transform -1 0 6690 0 -1 4950
box -6 -8 26 268
use FILL  FILL100350x150
timestamp 0
transform -1 0 6710 0 -1 270
box -6 -8 26 268
use FILL  FILL100350x4050
timestamp 0
transform 1 0 6690 0 1 270
box -6 -8 26 268
use FILL  FILL100350x7950
timestamp 0
transform -1 0 6710 0 -1 790
box -6 -8 26 268
use FILL  FILL100350x11850
timestamp 0
transform 1 0 6690 0 1 790
box -6 -8 26 268
use FILL  FILL100350x15750
timestamp 0
transform -1 0 6710 0 -1 1310
box -6 -8 26 268
use FILL  FILL100350x23550
timestamp 0
transform -1 0 6710 0 -1 1830
box -6 -8 26 268
use FILL  FILL100350x27450
timestamp 0
transform 1 0 6690 0 1 1830
box -6 -8 26 268
use FILL  FILL100350x31350
timestamp 0
transform -1 0 6710 0 -1 2350
box -6 -8 26 268
use FILL  FILL100350x35250
timestamp 0
transform 1 0 6690 0 1 2350
box -6 -8 26 268
use FILL  FILL100350x39150
timestamp 0
transform -1 0 6710 0 -1 2870
box -6 -8 26 268
use FILL  FILL100350x43050
timestamp 0
transform 1 0 6690 0 1 2870
box -6 -8 26 268
use FILL  FILL100350x46950
timestamp 0
transform -1 0 6710 0 -1 3390
box -6 -8 26 268
use FILL  FILL100350x58650
timestamp 0
transform 1 0 6690 0 1 3910
box -6 -8 26 268
use FILL  FILL100350x66450
timestamp 0
transform 1 0 6690 0 1 4430
box -6 -8 26 268
use FILL  FILL100350x70350
timestamp 0
transform -1 0 6710 0 -1 4950
box -6 -8 26 268
use FILL  FILL100350x74250
timestamp 0
transform 1 0 6690 0 1 4950
box -6 -8 26 268
use FILL  FILL100650x150
timestamp 0
transform -1 0 6730 0 -1 270
box -6 -8 26 268
use FILL  FILL100650x4050
timestamp 0
transform 1 0 6710 0 1 270
box -6 -8 26 268
use FILL  FILL100650x7950
timestamp 0
transform -1 0 6730 0 -1 790
box -6 -8 26 268
use FILL  FILL100650x11850
timestamp 0
transform 1 0 6710 0 1 790
box -6 -8 26 268
use FILL  FILL100650x15750
timestamp 0
transform -1 0 6730 0 -1 1310
box -6 -8 26 268
use FILL  FILL100650x23550
timestamp 0
transform -1 0 6730 0 -1 1830
box -6 -8 26 268
use FILL  FILL100650x27450
timestamp 0
transform 1 0 6710 0 1 1830
box -6 -8 26 268
use FILL  FILL100650x31350
timestamp 0
transform -1 0 6730 0 -1 2350
box -6 -8 26 268
use FILL  FILL100650x35250
timestamp 0
transform 1 0 6710 0 1 2350
box -6 -8 26 268
use FILL  FILL100650x39150
timestamp 0
transform -1 0 6730 0 -1 2870
box -6 -8 26 268
use FILL  FILL100650x43050
timestamp 0
transform 1 0 6710 0 1 2870
box -6 -8 26 268
use FILL  FILL100650x46950
timestamp 0
transform -1 0 6730 0 -1 3390
box -6 -8 26 268
use FILL  FILL100650x58650
timestamp 0
transform 1 0 6710 0 1 3910
box -6 -8 26 268
use FILL  FILL100650x66450
timestamp 0
transform 1 0 6710 0 1 4430
box -6 -8 26 268
use FILL  FILL100650x70350
timestamp 0
transform -1 0 6730 0 -1 4950
box -6 -8 26 268
use FILL  FILL100650x74250
timestamp 0
transform 1 0 6710 0 1 4950
box -6 -8 26 268
use FILL  FILL100650x78150
timestamp 0
transform -1 0 6730 0 -1 5470
box -6 -8 26 268
use FILL  FILL100650x85950
timestamp 0
transform -1 0 6730 0 -1 5990
box -6 -8 26 268
use FILL  FILL100950x150
timestamp 0
transform -1 0 6750 0 -1 270
box -6 -8 26 268
use FILL  FILL100950x4050
timestamp 0
transform 1 0 6730 0 1 270
box -6 -8 26 268
use FILL  FILL100950x7950
timestamp 0
transform -1 0 6750 0 -1 790
box -6 -8 26 268
use FILL  FILL100950x11850
timestamp 0
transform 1 0 6730 0 1 790
box -6 -8 26 268
use FILL  FILL100950x15750
timestamp 0
transform -1 0 6750 0 -1 1310
box -6 -8 26 268
use FILL  FILL100950x19650
timestamp 0
transform 1 0 6730 0 1 1310
box -6 -8 26 268
use FILL  FILL100950x23550
timestamp 0
transform -1 0 6750 0 -1 1830
box -6 -8 26 268
use FILL  FILL100950x27450
timestamp 0
transform 1 0 6730 0 1 1830
box -6 -8 26 268
use FILL  FILL100950x31350
timestamp 0
transform -1 0 6750 0 -1 2350
box -6 -8 26 268
use FILL  FILL100950x35250
timestamp 0
transform 1 0 6730 0 1 2350
box -6 -8 26 268
use FILL  FILL100950x39150
timestamp 0
transform -1 0 6750 0 -1 2870
box -6 -8 26 268
use FILL  FILL100950x43050
timestamp 0
transform 1 0 6730 0 1 2870
box -6 -8 26 268
use FILL  FILL100950x46950
timestamp 0
transform -1 0 6750 0 -1 3390
box -6 -8 26 268
use FILL  FILL100950x58650
timestamp 0
transform 1 0 6730 0 1 3910
box -6 -8 26 268
use FILL  FILL100950x66450
timestamp 0
transform 1 0 6730 0 1 4430
box -6 -8 26 268
use FILL  FILL100950x70350
timestamp 0
transform -1 0 6750 0 -1 4950
box -6 -8 26 268
use FILL  FILL100950x74250
timestamp 0
transform 1 0 6730 0 1 4950
box -6 -8 26 268
use FILL  FILL100950x78150
timestamp 0
transform -1 0 6750 0 -1 5470
box -6 -8 26 268
use FILL  FILL100950x82050
timestamp 0
transform 1 0 6730 0 1 5470
box -6 -8 26 268
use FILL  FILL100950x85950
timestamp 0
transform -1 0 6750 0 -1 5990
box -6 -8 26 268
use FILL  FILL100950x93750
timestamp 0
transform -1 0 6750 0 -1 6510
box -6 -8 26 268
use FILL  FILL101250x150
timestamp 0
transform -1 0 6770 0 -1 270
box -6 -8 26 268
use FILL  FILL101250x4050
timestamp 0
transform 1 0 6750 0 1 270
box -6 -8 26 268
use FILL  FILL101250x7950
timestamp 0
transform -1 0 6770 0 -1 790
box -6 -8 26 268
use FILL  FILL101250x11850
timestamp 0
transform 1 0 6750 0 1 790
box -6 -8 26 268
use FILL  FILL101250x15750
timestamp 0
transform -1 0 6770 0 -1 1310
box -6 -8 26 268
use FILL  FILL101250x19650
timestamp 0
transform 1 0 6750 0 1 1310
box -6 -8 26 268
use FILL  FILL101250x23550
timestamp 0
transform -1 0 6770 0 -1 1830
box -6 -8 26 268
use FILL  FILL101250x27450
timestamp 0
transform 1 0 6750 0 1 1830
box -6 -8 26 268
use FILL  FILL101250x31350
timestamp 0
transform -1 0 6770 0 -1 2350
box -6 -8 26 268
use FILL  FILL101250x35250
timestamp 0
transform 1 0 6750 0 1 2350
box -6 -8 26 268
use FILL  FILL101250x39150
timestamp 0
transform -1 0 6770 0 -1 2870
box -6 -8 26 268
use FILL  FILL101250x43050
timestamp 0
transform 1 0 6750 0 1 2870
box -6 -8 26 268
use FILL  FILL101250x46950
timestamp 0
transform -1 0 6770 0 -1 3390
box -6 -8 26 268
use FILL  FILL101250x50850
timestamp 0
transform 1 0 6750 0 1 3390
box -6 -8 26 268
use FILL  FILL101250x54750
timestamp 0
transform -1 0 6770 0 -1 3910
box -6 -8 26 268
use FILL  FILL101250x58650
timestamp 0
transform 1 0 6750 0 1 3910
box -6 -8 26 268
use FILL  FILL101250x66450
timestamp 0
transform 1 0 6750 0 1 4430
box -6 -8 26 268
use FILL  FILL101250x70350
timestamp 0
transform -1 0 6770 0 -1 4950
box -6 -8 26 268
use FILL  FILL101250x74250
timestamp 0
transform 1 0 6750 0 1 4950
box -6 -8 26 268
use FILL  FILL101250x78150
timestamp 0
transform -1 0 6770 0 -1 5470
box -6 -8 26 268
use FILL  FILL101250x82050
timestamp 0
transform 1 0 6750 0 1 5470
box -6 -8 26 268
use FILL  FILL101250x85950
timestamp 0
transform -1 0 6770 0 -1 5990
box -6 -8 26 268
use FILL  FILL101250x89850
timestamp 0
transform 1 0 6750 0 1 5990
box -6 -8 26 268
use FILL  FILL101250x93750
timestamp 0
transform -1 0 6770 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__922_
timestamp 0
transform -1 0 910 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__923_
timestamp 0
transform 1 0 1170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__924_
timestamp 0
transform -1 0 2630 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__925_
timestamp 0
transform 1 0 2450 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__926_
timestamp 0
transform -1 0 2510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__927_
timestamp 0
transform -1 0 1070 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__928_
timestamp 0
transform -1 0 1910 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__929_
timestamp 0
transform 1 0 2910 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__930_
timestamp 0
transform 1 0 2510 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__931_
timestamp 0
transform -1 0 3590 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__932_
timestamp 0
transform 1 0 2950 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__933_
timestamp 0
transform 1 0 2790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__934_
timestamp 0
transform 1 0 2830 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__935_
timestamp 0
transform 1 0 2670 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__936_
timestamp 0
transform -1 0 3450 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__937_
timestamp 0
transform 1 0 2290 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__938_
timestamp 0
transform 1 0 2090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__939_
timestamp 0
transform 1 0 2330 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__940_
timestamp 0
transform 1 0 1970 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__941_
timestamp 0
transform 1 0 1390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__942_
timestamp 0
transform -1 0 1630 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__943_
timestamp 0
transform 1 0 1430 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__944_
timestamp 0
transform -1 0 2170 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__945_
timestamp 0
transform 1 0 1450 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__946_
timestamp 0
transform -1 0 4430 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__947_
timestamp 0
transform -1 0 910 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__948_
timestamp 0
transform 1 0 570 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__949_
timestamp 0
transform 1 0 3690 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__950_
timestamp 0
transform 1 0 2130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__951_
timestamp 0
transform -1 0 2290 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__952_
timestamp 0
transform 1 0 3810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__953_
timestamp 0
transform 1 0 470 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__954_
timestamp 0
transform -1 0 630 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__955_
timestamp 0
transform 1 0 2650 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__956_
timestamp 0
transform -1 0 290 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__957_
timestamp 0
transform -1 0 430 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__958_
timestamp 0
transform 1 0 1030 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__959_
timestamp 0
transform -1 0 1670 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__960_
timestamp 0
transform 1 0 2590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__961_
timestamp 0
transform -1 0 2750 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__962_
timestamp 0
transform -1 0 2930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__963_
timestamp 0
transform -1 0 2950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__964_
timestamp 0
transform 1 0 1230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__965_
timestamp 0
transform -1 0 1310 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__966_
timestamp 0
transform -1 0 2970 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__967_
timestamp 0
transform 1 0 2630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__968_
timestamp 0
transform -1 0 2810 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__969_
timestamp 0
transform -1 0 3370 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__970_
timestamp 0
transform -1 0 3050 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__971_
timestamp 0
transform -1 0 3210 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__972_
timestamp 0
transform -1 0 3010 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__973_
timestamp 0
transform -1 0 2450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__974_
timestamp 0
transform -1 0 2850 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__975_
timestamp 0
transform -1 0 2550 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__976_
timestamp 0
transform 1 0 2170 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__977_
timestamp 0
transform -1 0 2350 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__978_
timestamp 0
transform -1 0 3690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__979_
timestamp 0
transform 1 0 3230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__980_
timestamp 0
transform -1 0 3530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__981_
timestamp 0
transform -1 0 3290 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__982_
timestamp 0
transform -1 0 2850 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__983_
timestamp 0
transform -1 0 3130 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__984_
timestamp 0
transform -1 0 3410 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__985_
timestamp 0
transform 1 0 4070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__986_
timestamp 0
transform 1 0 4030 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__987_
timestamp 0
transform -1 0 4190 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__988_
timestamp 0
transform 1 0 3630 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__989_
timestamp 0
transform 1 0 2490 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__990_
timestamp 0
transform -1 0 2650 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__991_
timestamp 0
transform 1 0 2750 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__992_
timestamp 0
transform 1 0 2730 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__993_
timestamp 0
transform 1 0 3910 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__994_
timestamp 0
transform -1 0 3970 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__995_
timestamp 0
transform 1 0 3290 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__996_
timestamp 0
transform 1 0 3130 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__997_
timestamp 0
transform 1 0 1670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__998_
timestamp 0
transform 1 0 1510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__999_
timestamp 0
transform 1 0 2230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1000_
timestamp 0
transform -1 0 3070 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1001_
timestamp 0
transform 1 0 2350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1002_
timestamp 0
transform -1 0 2550 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1003_
timestamp 0
transform 1 0 2890 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1004_
timestamp 0
transform 1 0 2730 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1005_
timestamp 0
transform -1 0 1930 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1006_
timestamp 0
transform 1 0 1830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1007_
timestamp 0
transform 1 0 1750 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1008_
timestamp 0
transform 1 0 1490 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1009_
timestamp 0
transform 1 0 1070 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1010_
timestamp 0
transform -1 0 1250 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1011_
timestamp 0
transform 1 0 990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1012_
timestamp 0
transform 1 0 2290 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1013_
timestamp 0
transform -1 0 3410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1014_
timestamp 0
transform 1 0 870 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1015_
timestamp 0
transform -1 0 1770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1016_
timestamp 0
transform 1 0 1930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1017_
timestamp 0
transform 1 0 2490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1018_
timestamp 0
transform 1 0 2070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1019_
timestamp 0
transform -1 0 730 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1020_
timestamp 0
transform 1 0 870 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1021_
timestamp 0
transform 1 0 1170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1022_
timestamp 0
transform -1 0 1430 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1023_
timestamp 0
transform 1 0 1310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1024_
timestamp 0
transform 1 0 1190 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1025_
timestamp 0
transform -1 0 1490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1026_
timestamp 0
transform 1 0 1330 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1027_
timestamp 0
transform 1 0 1490 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1028_
timestamp 0
transform -1 0 1470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1029_
timestamp 0
transform -1 0 1630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1030_
timestamp 0
transform -1 0 1510 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1031_
timestamp 0
transform 1 0 1830 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1032_
timestamp 0
transform 1 0 1670 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1033_
timestamp 0
transform 1 0 2270 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1034_
timestamp 0
transform 1 0 1590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1035_
timestamp 0
transform 1 0 3830 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1036_
timestamp 0
transform -1 0 1250 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1037_
timestamp 0
transform 1 0 1070 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1038_
timestamp 0
transform -1 0 4570 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1039_
timestamp 0
transform -1 0 1550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1040_
timestamp 0
transform 1 0 630 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1041_
timestamp 0
transform 1 0 470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1042_
timestamp 0
transform 1 0 750 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1043_
timestamp 0
transform -1 0 650 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1044_
timestamp 0
transform -1 0 1390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1045_
timestamp 0
transform 1 0 1070 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1046_
timestamp 0
transform 1 0 950 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1047_
timestamp 0
transform 1 0 770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1048_
timestamp 0
transform 1 0 1190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1049_
timestamp 0
transform -1 0 950 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1050_
timestamp 0
transform 1 0 1050 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1051_
timestamp 0
transform 1 0 1370 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1052_
timestamp 0
transform -1 0 1690 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1053_
timestamp 0
transform -1 0 1910 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1054_
timestamp 0
transform 1 0 2290 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1055_
timestamp 0
transform -1 0 1910 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1056_
timestamp 0
transform -1 0 1570 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1057_
timestamp 0
transform -1 0 1730 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1058_
timestamp 0
transform 1 0 1550 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1059_
timestamp 0
transform -1 0 1730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1060_
timestamp 0
transform 1 0 1850 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1061_
timestamp 0
transform -1 0 2230 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1062_
timestamp 0
transform 1 0 1210 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1063_
timestamp 0
transform -1 0 1730 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1064_
timestamp 0
transform -1 0 3550 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1065_
timestamp 0
transform 1 0 2470 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1066_
timestamp 0
transform -1 0 2470 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1067_
timestamp 0
transform 1 0 2330 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1068_
timestamp 0
transform -1 0 910 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1069_
timestamp 0
transform -1 0 170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1070_
timestamp 0
transform -1 0 330 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1071_
timestamp 0
transform 1 0 190 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1072_
timestamp 0
transform -1 0 30 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1073_
timestamp 0
transform 1 0 310 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1074_
timestamp 0
transform -1 0 210 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1075_
timestamp 0
transform 1 0 10 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1076_
timestamp 0
transform 1 0 310 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1077_
timestamp 0
transform -1 0 490 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1078_
timestamp 0
transform 1 0 970 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1079_
timestamp 0
transform 1 0 630 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1080_
timestamp 0
transform 1 0 1110 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1081_
timestamp 0
transform -1 0 970 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1082_
timestamp 0
transform 1 0 630 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1083_
timestamp 0
transform 1 0 150 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1084_
timestamp 0
transform 1 0 150 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1085_
timestamp 0
transform 1 0 290 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1086_
timestamp 0
transform -1 0 4890 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1087_
timestamp 0
transform -1 0 470 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1088_
timestamp 0
transform -1 0 330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1089_
timestamp 0
transform 1 0 470 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1090_
timestamp 0
transform 1 0 1090 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1091_
timestamp 0
transform 1 0 1450 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1092_
timestamp 0
transform 1 0 1790 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1093_
timestamp 0
transform -1 0 1610 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1094_
timestamp 0
transform 1 0 1930 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1095_
timestamp 0
transform 1 0 2090 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1096_
timestamp 0
transform -1 0 2170 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1097_
timestamp 0
transform 1 0 2010 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1098_
timestamp 0
transform 1 0 2050 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1099_
timestamp 0
transform -1 0 2770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1100_
timestamp 0
transform 1 0 2610 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1101_
timestamp 0
transform -1 0 810 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1102_
timestamp 0
transform 1 0 10 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1103_
timestamp 0
transform 1 0 1090 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1104_
timestamp 0
transform -1 0 810 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1105_
timestamp 0
transform 1 0 470 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1106_
timestamp 0
transform -1 0 750 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1107_
timestamp 0
transform -1 0 30 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1108_
timestamp 0
transform 1 0 610 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1109_
timestamp 0
transform 1 0 130 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1110_
timestamp 0
transform -1 0 30 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1111_
timestamp 0
transform 1 0 430 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1112_
timestamp 0
transform 1 0 1370 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1113_
timestamp 0
transform 1 0 610 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1114_
timestamp 0
transform -1 0 270 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1115_
timestamp 0
transform 1 0 770 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1116_
timestamp 0
transform 1 0 3850 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1117_
timestamp 0
transform -1 0 4850 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1118_
timestamp 0
transform 1 0 4330 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1119_
timestamp 0
transform 1 0 4330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1120_
timestamp 0
transform 1 0 4490 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1121_
timestamp 0
transform -1 0 4390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1122_
timestamp 0
transform 1 0 4610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1123_
timestamp 0
transform 1 0 4650 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1124_
timestamp 0
transform 1 0 3630 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1125_
timestamp 0
transform 1 0 3790 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1126_
timestamp 0
transform 1 0 3950 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1127_
timestamp 0
transform -1 0 3810 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1128_
timestamp 0
transform -1 0 3670 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1129_
timestamp 0
transform 1 0 1770 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1130_
timestamp 0
transform 1 0 930 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1131_
timestamp 0
transform 1 0 1210 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1132_
timestamp 0
transform -1 0 3830 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1133_
timestamp 0
transform 1 0 2030 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1134_
timestamp 0
transform 1 0 2110 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1135_
timestamp 0
transform 1 0 1270 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1136_
timestamp 0
transform -1 0 1730 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1137_
timestamp 0
transform 1 0 1530 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1138_
timestamp 0
transform 1 0 1430 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1139_
timestamp 0
transform 1 0 2650 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1140_
timestamp 0
transform 1 0 1270 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1141_
timestamp 0
transform 1 0 1610 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1142_
timestamp 0
transform 1 0 1950 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1143_
timestamp 0
transform 1 0 2290 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1144_
timestamp 0
transform -1 0 2990 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1145_
timestamp 0
transform 1 0 2730 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1146_
timestamp 0
transform 1 0 3130 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1147_
timestamp 0
transform 1 0 2850 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1148_
timestamp 0
transform 1 0 2830 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1149_
timestamp 0
transform 1 0 2650 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1150_
timestamp 0
transform 1 0 3150 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1151_
timestamp 0
transform 1 0 2990 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1152_
timestamp 0
transform 1 0 2430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1153_
timestamp 0
transform -1 0 2830 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1154_
timestamp 0
transform 1 0 2810 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1155_
timestamp 0
transform 1 0 4650 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1156_
timestamp 0
transform 1 0 4590 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1157_
timestamp 0
transform -1 0 4990 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1158_
timestamp 0
transform -1 0 5470 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1159_
timestamp 0
transform -1 0 4790 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1160_
timestamp 0
transform 1 0 4770 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1161_
timestamp 0
transform 1 0 2190 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1162_
timestamp 0
transform -1 0 4010 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1163_
timestamp 0
transform -1 0 4950 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1164_
timestamp 0
transform 1 0 4470 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1165_
timestamp 0
transform -1 0 4810 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1166_
timestamp 0
transform 1 0 4130 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1167_
timestamp 0
transform -1 0 4310 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1168_
timestamp 0
transform 1 0 4490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1169_
timestamp 0
transform -1 0 4810 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1170_
timestamp 0
transform 1 0 4130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1171_
timestamp 0
transform 1 0 4770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1172_
timestamp 0
transform 1 0 4970 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1173_
timestamp 0
transform 1 0 790 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1174_
timestamp 0
transform 1 0 3630 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1175_
timestamp 0
transform 1 0 3230 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1176_
timestamp 0
transform 1 0 3290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1177_
timestamp 0
transform -1 0 3390 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1178_
timestamp 0
transform -1 0 3950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1179_
timestamp 0
transform 1 0 3490 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1180_
timestamp 0
transform 1 0 3230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1181_
timestamp 0
transform 1 0 3510 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1182_
timestamp 0
transform 1 0 3670 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1183_
timestamp 0
transform 1 0 4090 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1184_
timestamp 0
transform 1 0 3850 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1185_
timestamp 0
transform 1 0 3470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1186_
timestamp 0
transform 1 0 3610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1187_
timestamp 0
transform 1 0 3770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1188_
timestamp 0
transform 1 0 3670 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1189_
timestamp 0
transform -1 0 4030 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1190_
timestamp 0
transform 1 0 4290 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1191_
timestamp 0
transform -1 0 5130 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1192_
timestamp 0
transform 1 0 3930 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1193_
timestamp 0
transform 1 0 4170 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1194_
timestamp 0
transform -1 0 4450 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1195_
timestamp 0
transform -1 0 3970 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1196_
timestamp 0
transform -1 0 1890 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1197_
timestamp 0
transform 1 0 4250 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1198_
timestamp 0
transform -1 0 4150 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1199_
timestamp 0
transform -1 0 3630 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1200_
timestamp 0
transform 1 0 3430 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1201_
timestamp 0
transform 1 0 4270 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1202_
timestamp 0
transform 1 0 4450 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1203_
timestamp 0
transform 1 0 3770 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1204_
timestamp 0
transform -1 0 4630 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1205_
timestamp 0
transform 1 0 3970 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1206_
timestamp 0
transform 1 0 2470 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1207_
timestamp 0
transform -1 0 4130 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1208_
timestamp 0
transform -1 0 3290 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1209_
timestamp 0
transform -1 0 2950 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1210_
timestamp 0
transform -1 0 3130 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1211_
timestamp 0
transform 1 0 3210 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1212_
timestamp 0
transform 1 0 3290 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1213_
timestamp 0
transform 1 0 3470 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1214_
timestamp 0
transform -1 0 3350 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1215_
timestamp 0
transform -1 0 3010 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1216_
timestamp 0
transform -1 0 2610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1217_
timestamp 0
transform 1 0 3470 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1218_
timestamp 0
transform 1 0 5030 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1219_
timestamp 0
transform -1 0 5110 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1220_
timestamp 0
transform -1 0 4750 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1221_
timestamp 0
transform 1 0 4550 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1222_
timestamp 0
transform 1 0 4470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1223_
timestamp 0
transform 1 0 4970 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1224_
timestamp 0
transform -1 0 5090 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1225_
timestamp 0
transform 1 0 6070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1226_
timestamp 0
transform 1 0 5930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1227_
timestamp 0
transform -1 0 5310 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1228_
timestamp 0
transform 1 0 5590 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1229_
timestamp 0
transform -1 0 6290 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1230_
timestamp 0
transform 1 0 4930 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1231_
timestamp 0
transform 1 0 5070 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1232_
timestamp 0
transform 1 0 4810 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1233_
timestamp 0
transform -1 0 5130 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1234_
timestamp 0
transform 1 0 5590 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1235_
timestamp 0
transform -1 0 5450 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1236_
timestamp 0
transform -1 0 5430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1237_
timestamp 0
transform 1 0 4950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1238_
timestamp 0
transform 1 0 4490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1239_
timestamp 0
transform -1 0 4670 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1240_
timestamp 0
transform 1 0 5270 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1241_
timestamp 0
transform 1 0 5250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1242_
timestamp 0
transform 1 0 5730 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1243_
timestamp 0
transform -1 0 3370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1244_
timestamp 0
transform 1 0 5570 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1245_
timestamp 0
transform 1 0 4090 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1246_
timestamp 0
transform 1 0 4430 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1247_
timestamp 0
transform -1 0 4970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1248_
timestamp 0
transform 1 0 4250 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1249_
timestamp 0
transform 1 0 5070 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1250_
timestamp 0
transform 1 0 5370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1251_
timestamp 0
transform 1 0 5230 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1252_
timestamp 0
transform 1 0 5670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1253_
timestamp 0
transform -1 0 5710 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1254_
timestamp 0
transform -1 0 5510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1255_
timestamp 0
transform -1 0 3990 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1256_
timestamp 0
transform 1 0 4090 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1257_
timestamp 0
transform 1 0 3650 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1258_
timestamp 0
transform 1 0 4210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1259_
timestamp 0
transform -1 0 5250 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1260_
timestamp 0
transform 1 0 5930 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1261_
timestamp 0
transform 1 0 5890 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1262_
timestamp 0
transform 1 0 5830 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1263_
timestamp 0
transform 1 0 5390 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1264_
timestamp 0
transform 1 0 5570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1265_
timestamp 0
transform -1 0 5890 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1266_
timestamp 0
transform 1 0 3750 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1267_
timestamp 0
transform 1 0 4610 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1268_
timestamp 0
transform 1 0 5410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1269_
timestamp 0
transform -1 0 5770 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1270_
timestamp 0
transform -1 0 5570 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1271_
timestamp 0
transform 1 0 6190 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1272_
timestamp 0
transform -1 0 6490 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1273_
timestamp 0
transform 1 0 6030 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1274_
timestamp 0
transform 1 0 5710 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1275_
timestamp 0
transform -1 0 6570 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1276_
timestamp 0
transform -1 0 6150 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1277_
timestamp 0
transform 1 0 4390 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1278_
timestamp 0
transform 1 0 4850 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1279_
timestamp 0
transform -1 0 6530 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1280_
timestamp 0
transform -1 0 6050 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1281_
timestamp 0
transform -1 0 5810 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1282_
timestamp 0
transform -1 0 5530 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1283_
timestamp 0
transform 1 0 5410 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1284_
timestamp 0
transform -1 0 6310 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1285_
timestamp 0
transform -1 0 5990 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1286_
timestamp 0
transform -1 0 5890 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1287_
timestamp 0
transform 1 0 5170 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1288_
timestamp 0
transform -1 0 5550 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1289_
timestamp 0
transform -1 0 5370 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1290_
timestamp 0
transform -1 0 5250 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1291_
timestamp 0
transform -1 0 5250 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1292_
timestamp 0
transform 1 0 5390 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1293_
timestamp 0
transform 1 0 4250 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1294_
timestamp 0
transform 1 0 4190 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1295_
timestamp 0
transform -1 0 4670 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1296_
timestamp 0
transform -1 0 4690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1297_
timestamp 0
transform 1 0 5670 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1298_
timestamp 0
transform -1 0 5710 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1299_
timestamp 0
transform 1 0 5890 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1300_
timestamp 0
transform 1 0 6350 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1301_
timestamp 0
transform -1 0 6490 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1302_
timestamp 0
transform -1 0 4350 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1303_
timestamp 0
transform 1 0 5430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1304_
timestamp 0
transform -1 0 4810 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1305_
timestamp 0
transform 1 0 5130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1306_
timestamp 0
transform 1 0 5050 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1307_
timestamp 0
transform 1 0 5330 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1308_
timestamp 0
transform 1 0 5730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1309_
timestamp 0
transform -1 0 4150 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1310_
timestamp 0
transform 1 0 4730 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1311_
timestamp 0
transform -1 0 5290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1312_
timestamp 0
transform 1 0 5390 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1313_
timestamp 0
transform -1 0 5090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1314_
timestamp 0
transform -1 0 5890 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1315_
timestamp 0
transform 1 0 5230 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1316_
timestamp 0
transform -1 0 5570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1317_
timestamp 0
transform 1 0 5590 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1318_
timestamp 0
transform 1 0 5710 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1319_
timestamp 0
transform 1 0 5750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1320_
timestamp 0
transform 1 0 5550 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1321_
timestamp 0
transform 1 0 6030 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1322_
timestamp 0
transform 1 0 6190 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1323_
timestamp 0
transform 1 0 6190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1324_
timestamp 0
transform -1 0 6430 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1325_
timestamp 0
transform 1 0 6230 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1326_
timestamp 0
transform 1 0 4910 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1327_
timestamp 0
transform 1 0 4390 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1328_
timestamp 0
transform 1 0 4110 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1329_
timestamp 0
transform -1 0 4310 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1330_
timestamp 0
transform 1 0 4430 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1331_
timestamp 0
transform 1 0 4570 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1332_
timestamp 0
transform 1 0 5050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1333_
timestamp 0
transform 1 0 4410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1334_
timestamp 0
transform 1 0 4890 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1335_
timestamp 0
transform 1 0 3950 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1336_
timestamp 0
transform 1 0 5330 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1337_
timestamp 0
transform 1 0 5490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1338_
timestamp 0
transform 1 0 4910 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1339_
timestamp 0
transform -1 0 5990 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1340_
timestamp 0
transform -1 0 4630 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1341_
timestamp 0
transform 1 0 3390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1342_
timestamp 0
transform 1 0 3510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1343_
timestamp 0
transform -1 0 3830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1344_
timestamp 0
transform -1 0 4230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1345_
timestamp 0
transform 1 0 4530 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1346_
timestamp 0
transform 1 0 5230 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1347_
timestamp 0
transform 1 0 4290 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1348_
timestamp 0
transform 1 0 3670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1349_
timestamp 0
transform 1 0 5370 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1350_
timestamp 0
transform -1 0 6010 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1351_
timestamp 0
transform 1 0 5550 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1352_
timestamp 0
transform 1 0 4350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1353_
timestamp 0
transform 1 0 5490 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1354_
timestamp 0
transform 1 0 6010 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1355_
timestamp 0
transform 1 0 5650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1356_
timestamp 0
transform 1 0 6150 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1357_
timestamp 0
transform 1 0 5650 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1358_
timestamp 0
transform 1 0 6470 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1359_
timestamp 0
transform -1 0 6250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1360_
timestamp 0
transform 1 0 5990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1361_
timestamp 0
transform 1 0 6050 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1362_
timestamp 0
transform -1 0 6330 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1363_
timestamp 0
transform 1 0 5850 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1364_
timestamp 0
transform 1 0 5890 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1365_
timestamp 0
transform -1 0 6390 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1366_
timestamp 0
transform 1 0 6490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1367_
timestamp 0
transform 1 0 6170 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1368_
timestamp 0
transform 1 0 6070 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1369_
timestamp 0
transform 1 0 6530 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1370_
timestamp 0
transform -1 0 6230 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1371_
timestamp 0
transform 1 0 6110 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1372_
timestamp 0
transform 1 0 6190 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1373_
timestamp 0
transform 1 0 6570 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1374_
timestamp 0
transform -1 0 6350 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1375_
timestamp 0
transform -1 0 6170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1376_
timestamp 0
transform -1 0 5870 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1377_
timestamp 0
transform 1 0 6510 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1378_
timestamp 0
transform -1 0 6410 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1379_
timestamp 0
transform -1 0 6330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1380_
timestamp 0
transform -1 0 6210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1381_
timestamp 0
transform -1 0 5750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1382_
timestamp 0
transform -1 0 6490 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1383_
timestamp 0
transform -1 0 6370 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1384_
timestamp 0
transform -1 0 6370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1385_
timestamp 0
transform -1 0 6050 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1386_
timestamp 0
transform -1 0 6050 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1387_
timestamp 0
transform 1 0 5270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1388_
timestamp 0
transform 1 0 4690 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1389_
timestamp 0
transform -1 0 4570 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1390_
timestamp 0
transform -1 0 5010 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1391_
timestamp 0
transform 1 0 4370 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1392_
timestamp 0
transform 1 0 4010 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1393_
timestamp 0
transform 1 0 3850 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1394_
timestamp 0
transform -1 0 5110 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1395_
timestamp 0
transform -1 0 5130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1396_
timestamp 0
transform -1 0 4950 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1397_
timestamp 0
transform -1 0 6570 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1398_
timestamp 0
transform 1 0 6590 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1399_
timestamp 0
transform -1 0 6550 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1400_
timestamp 0
transform -1 0 6470 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1401_
timestamp 0
transform -1 0 6410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1402_
timestamp 0
transform -1 0 6530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1403_
timestamp 0
transform -1 0 5690 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1404_
timestamp 0
transform -1 0 4070 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1405_
timestamp 0
transform 1 0 4890 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1406_
timestamp 0
transform -1 0 4730 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1407_
timestamp 0
transform 1 0 4330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1408_
timestamp 0
transform -1 0 4710 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1409_
timestamp 0
transform -1 0 4650 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1410_
timestamp 0
transform -1 0 4790 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1411_
timestamp 0
transform -1 0 4850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1412_
timestamp 0
transform 1 0 4370 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1413_
timestamp 0
transform -1 0 4770 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1414_
timestamp 0
transform 1 0 4730 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1415_
timestamp 0
transform 1 0 4530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1416_
timestamp 0
transform 1 0 5170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1417_
timestamp 0
transform 1 0 5190 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1418_
timestamp 0
transform 1 0 4550 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1419_
timestamp 0
transform 1 0 4990 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1420_
timestamp 0
transform 1 0 4250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1421_
timestamp 0
transform 1 0 4190 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1422_
timestamp 0
transform 1 0 5350 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1423_
timestamp 0
transform 1 0 5670 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1424_
timestamp 0
transform 1 0 5190 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1425_
timestamp 0
transform 1 0 5510 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1426_
timestamp 0
transform 1 0 5510 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1427_
timestamp 0
transform 1 0 5010 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1428_
timestamp 0
transform -1 0 5850 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1429_
timestamp 0
transform 1 0 5710 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1430_
timestamp 0
transform 1 0 6150 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1431_
timestamp 0
transform -1 0 6310 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1432_
timestamp 0
transform 1 0 4850 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1433_
timestamp 0
transform -1 0 4270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1434_
timestamp 0
transform 1 0 4670 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1435_
timestamp 0
transform -1 0 4590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1436_
timestamp 0
transform 1 0 4710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1437_
timestamp 0
transform 1 0 5010 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1438_
timestamp 0
transform 1 0 5170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1439_
timestamp 0
transform 1 0 3090 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1440_
timestamp 0
transform -1 0 4910 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1441_
timestamp 0
transform 1 0 4090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1442_
timestamp 0
transform 1 0 5330 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1443_
timestamp 0
transform 1 0 5510 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1444_
timestamp 0
transform 1 0 3650 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1445_
timestamp 0
transform 1 0 3130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1446_
timestamp 0
transform -1 0 3930 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1447_
timestamp 0
transform -1 0 4510 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1448_
timestamp 0
transform 1 0 4930 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1449_
timestamp 0
transform 1 0 4450 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1450_
timestamp 0
transform 1 0 4930 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1451_
timestamp 0
transform 1 0 4630 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1452_
timestamp 0
transform 1 0 5290 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1453_
timestamp 0
transform -1 0 5670 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1454_
timestamp 0
transform 1 0 4130 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1455_
timestamp 0
transform 1 0 3990 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1456_
timestamp 0
transform -1 0 5350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1457_
timestamp 0
transform 1 0 5450 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1458_
timestamp 0
transform 1 0 5490 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1459_
timestamp 0
transform 1 0 5590 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1460_
timestamp 0
transform 1 0 5830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1461_
timestamp 0
transform 1 0 5990 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1462_
timestamp 0
transform -1 0 5050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1463_
timestamp 0
transform 1 0 5270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1464_
timestamp 0
transform 1 0 5830 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1465_
timestamp 0
transform 1 0 5110 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1466_
timestamp 0
transform 1 0 5730 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1467_
timestamp 0
transform 1 0 5850 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1468_
timestamp 0
transform -1 0 6030 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1469_
timestamp 0
transform 1 0 5430 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1470_
timestamp 0
transform 1 0 5890 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1471_
timestamp 0
transform -1 0 5950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1472_
timestamp 0
transform 1 0 6090 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1473_
timestamp 0
transform 1 0 6350 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1474_
timestamp 0
transform -1 0 6530 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1475_
timestamp 0
transform 1 0 6110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1476_
timestamp 0
transform 1 0 5770 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1477_
timestamp 0
transform 1 0 6350 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1478_
timestamp 0
transform -1 0 6450 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1479_
timestamp 0
transform 1 0 6190 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1480_
timestamp 0
transform -1 0 6290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1481_
timestamp 0
transform 1 0 6530 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1482_
timestamp 0
transform 1 0 6590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1483_
timestamp 0
transform -1 0 6610 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1484_
timestamp 0
transform 1 0 6490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1485_
timestamp 0
transform -1 0 6630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1486_
timestamp 0
transform -1 0 6270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1487_
timestamp 0
transform -1 0 6470 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1488_
timestamp 0
transform -1 0 4810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1489_
timestamp 0
transform 1 0 3950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1490_
timestamp 0
transform 1 0 3990 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1491_
timestamp 0
transform -1 0 5010 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1492_
timestamp 0
transform 1 0 4810 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1493_
timestamp 0
transform 1 0 6350 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1494_
timestamp 0
transform 1 0 6470 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1495_
timestamp 0
transform -1 0 5830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1496_
timestamp 0
transform 1 0 6250 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1497_
timestamp 0
transform -1 0 6070 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1498_
timestamp 0
transform 1 0 6170 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1499_
timestamp 0
transform 1 0 5150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1500_
timestamp 0
transform -1 0 4550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1501_
timestamp 0
transform 1 0 4050 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1502_
timestamp 0
transform 1 0 4790 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1503_
timestamp 0
transform -1 0 4690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1504_
timestamp 0
transform 1 0 5090 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1505_
timestamp 0
transform 1 0 4810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1506_
timestamp 0
transform -1 0 4490 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1507_
timestamp 0
transform 1 0 4490 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1508_
timestamp 0
transform -1 0 4990 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1509_
timestamp 0
transform 1 0 5110 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1510_
timestamp 0
transform 1 0 4830 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1511_
timestamp 0
transform 1 0 5170 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1512_
timestamp 0
transform -1 0 5310 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1513_
timestamp 0
transform 1 0 4930 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1514_
timestamp 0
transform 1 0 4930 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1515_
timestamp 0
transform 1 0 4990 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1516_
timestamp 0
transform 1 0 5510 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1517_
timestamp 0
transform 1 0 5450 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1518_
timestamp 0
transform 1 0 5090 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1519_
timestamp 0
transform 1 0 5310 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1520_
timestamp 0
transform 1 0 5270 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1521_
timestamp 0
transform 1 0 5350 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1522_
timestamp 0
transform 1 0 5430 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1523_
timestamp 0
transform 1 0 5590 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1524_
timestamp 0
transform -1 0 5130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1525_
timestamp 0
transform -1 0 5830 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1526_
timestamp 0
transform 1 0 3610 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1527_
timestamp 0
transform 1 0 3110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1528_
timestamp 0
transform -1 0 3930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1529_
timestamp 0
transform 1 0 3450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1530_
timestamp 0
transform 1 0 3750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1531_
timestamp 0
transform 1 0 4530 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1532_
timestamp 0
transform -1 0 3570 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1533_
timestamp 0
transform -1 0 3830 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1534_
timestamp 0
transform -1 0 4370 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1535_
timestamp 0
transform -1 0 4410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1536_
timestamp 0
transform 1 0 4030 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1537_
timestamp 0
transform 1 0 4210 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1538_
timestamp 0
transform 1 0 4350 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1539_
timestamp 0
transform 1 0 4230 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1540_
timestamp 0
transform 1 0 5610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1541_
timestamp 0
transform -1 0 5790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1542_
timestamp 0
transform -1 0 5210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1543_
timestamp 0
transform 1 0 5650 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1544_
timestamp 0
transform -1 0 5710 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1545_
timestamp 0
transform -1 0 5630 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1546_
timestamp 0
transform 1 0 6050 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1547_
timestamp 0
transform 1 0 5850 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1548_
timestamp 0
transform -1 0 5930 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1549_
timestamp 0
transform 1 0 6230 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1550_
timestamp 0
transform -1 0 6250 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1551_
timestamp 0
transform 1 0 5570 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1552_
timestamp 0
transform 1 0 5990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1553_
timestamp 0
transform 1 0 6050 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1554_
timestamp 0
transform 1 0 5770 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1555_
timestamp 0
transform -1 0 6010 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1556_
timestamp 0
transform 1 0 5930 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1557_
timestamp 0
transform -1 0 6110 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1558_
timestamp 0
transform 1 0 6350 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1559_
timestamp 0
transform 1 0 6550 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1560_
timestamp 0
transform 1 0 6010 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1561_
timestamp 0
transform -1 0 6550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1562_
timestamp 0
transform -1 0 6550 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1563_
timestamp 0
transform -1 0 6390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1564_
timestamp 0
transform 1 0 6170 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1565_
timestamp 0
transform 1 0 6330 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1566_
timestamp 0
transform -1 0 6530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1567_
timestamp 0
transform -1 0 4430 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1568_
timestamp 0
transform 1 0 4150 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1569_
timestamp 0
transform -1 0 4190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1570_
timestamp 0
transform -1 0 3710 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1571_
timestamp 0
transform 1 0 6170 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1572_
timestamp 0
transform -1 0 4290 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1573_
timestamp 0
transform -1 0 3650 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1574_
timestamp 0
transform 1 0 6390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1575_
timestamp 0
transform 1 0 6410 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1576_
timestamp 0
transform 1 0 5430 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1577_
timestamp 0
transform -1 0 5450 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1578_
timestamp 0
transform -1 0 5910 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1579_
timestamp 0
transform -1 0 4650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1580_
timestamp 0
transform 1 0 4350 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1581_
timestamp 0
transform -1 0 2990 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1582_
timestamp 0
transform -1 0 2790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1583_
timestamp 0
transform -1 0 2850 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1584_
timestamp 0
transform -1 0 2990 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1585_
timestamp 0
transform 1 0 3130 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1586_
timestamp 0
transform 1 0 2650 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1587_
timestamp 0
transform 1 0 2770 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1588_
timestamp 0
transform -1 0 1950 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1589_
timestamp 0
transform -1 0 2650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1590_
timestamp 0
transform 1 0 2890 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1591_
timestamp 0
transform 1 0 3850 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1592_
timestamp 0
transform -1 0 3710 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1593_
timestamp 0
transform -1 0 3730 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1594_
timestamp 0
transform 1 0 3050 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1595_
timestamp 0
transform 1 0 2970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1596_
timestamp 0
transform -1 0 4030 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1597_
timestamp 0
transform -1 0 4190 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1598_
timestamp 0
transform 1 0 4030 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1599_
timestamp 0
transform -1 0 4210 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1600_
timestamp 0
transform 1 0 3530 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1601_
timestamp 0
transform 1 0 3870 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1602_
timestamp 0
transform -1 0 3870 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1603_
timestamp 0
transform 1 0 4770 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1604_
timestamp 0
transform 1 0 3630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1605_
timestamp 0
transform 1 0 3470 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1606_
timestamp 0
transform 1 0 1350 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1607_
timestamp 0
transform -1 0 3330 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1608_
timestamp 0
transform -1 0 2690 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1609_
timestamp 0
transform 1 0 3110 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1610_
timestamp 0
transform -1 0 2370 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1611_
timestamp 0
transform -1 0 2530 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1612_
timestamp 0
transform 1 0 1490 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1613_
timestamp 0
transform 1 0 3250 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1614_
timestamp 0
transform 1 0 3390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1615_
timestamp 0
transform 1 0 3750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1616_
timestamp 0
transform 1 0 3110 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1617_
timestamp 0
transform -1 0 3570 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1618_
timestamp 0
transform 1 0 4190 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1619_
timestamp 0
transform -1 0 4650 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1620_
timestamp 0
transform 1 0 3730 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1621_
timestamp 0
transform 1 0 3410 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1622_
timestamp 0
transform 1 0 3910 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1623_
timestamp 0
transform 1 0 4930 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1624_
timestamp 0
transform 1 0 5890 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1625_
timestamp 0
transform 1 0 5730 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1626_
timestamp 0
transform 1 0 4170 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1627_
timestamp 0
transform -1 0 4510 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1628_
timestamp 0
transform 1 0 4810 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1629_
timestamp 0
transform 1 0 6210 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1630_
timestamp 0
transform -1 0 5750 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1631_
timestamp 0
transform 1 0 4650 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1632_
timestamp 0
transform 1 0 5550 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1633_
timestamp 0
transform 1 0 6390 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1634_
timestamp 0
transform 1 0 6170 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1635_
timestamp 0
transform -1 0 6430 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1636_
timestamp 0
transform 1 0 5090 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1637_
timestamp 0
transform -1 0 6070 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1638_
timestamp 0
transform 1 0 5250 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1639_
timestamp 0
transform 1 0 4650 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1640_
timestamp 0
transform 1 0 3490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1641_
timestamp 0
transform 1 0 3310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1642_
timestamp 0
transform 1 0 3530 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1643_
timestamp 0
transform 1 0 2190 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1644_
timestamp 0
transform -1 0 3150 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1645_
timestamp 0
transform -1 0 5290 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1646_
timestamp 0
transform -1 0 5130 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1647_
timestamp 0
transform 1 0 3690 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1648_
timestamp 0
transform -1 0 3750 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1649_
timestamp 0
transform -1 0 4030 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1650_
timestamp 0
transform -1 0 3410 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1651_
timestamp 0
transform -1 0 3550 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1652_
timestamp 0
transform -1 0 2510 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1653_
timestamp 0
transform 1 0 2470 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1654_
timestamp 0
transform -1 0 2370 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1655_
timestamp 0
transform -1 0 2170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1656_
timestamp 0
transform 1 0 1650 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1657_
timestamp 0
transform -1 0 2050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1658_
timestamp 0
transform 1 0 1790 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1659_
timestamp 0
transform -1 0 2010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1660_
timestamp 0
transform -1 0 2230 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1661_
timestamp 0
transform 1 0 2070 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1662_
timestamp 0
transform 1 0 2170 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1663_
timestamp 0
transform -1 0 1910 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1664_
timestamp 0
transform -1 0 1610 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1665_
timestamp 0
transform -1 0 1430 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1666_
timestamp 0
transform -1 0 1850 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1667_
timestamp 0
transform 1 0 1430 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1668_
timestamp 0
transform 1 0 1970 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1669_
timestamp 0
transform 1 0 2310 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1670_
timestamp 0
transform 1 0 1270 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1671_
timestamp 0
transform -1 0 1730 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1672_
timestamp 0
transform 1 0 1810 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1673_
timestamp 0
transform -1 0 30 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1674_
timestamp 0
transform -1 0 30 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1675_
timestamp 0
transform 1 0 10 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1676_
timestamp 0
transform 1 0 170 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1677_
timestamp 0
transform 1 0 310 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1678_
timestamp 0
transform 1 0 2150 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1679_
timestamp 0
transform -1 0 1670 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1680_
timestamp 0
transform -1 0 1490 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1681_
timestamp 0
transform 1 0 1190 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1682_
timestamp 0
transform -1 0 1330 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1683_
timestamp 0
transform 1 0 2570 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1684_
timestamp 0
transform -1 0 2450 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1685_
timestamp 0
transform -1 0 3250 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1686_
timestamp 0
transform 1 0 3850 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1687_
timestamp 0
transform -1 0 4350 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1688_
timestamp 0
transform 1 0 2750 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1689_
timestamp 0
transform -1 0 2930 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1690_
timestamp 0
transform -1 0 3090 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1691_
timestamp 0
transform -1 0 4050 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1692_
timestamp 0
transform -1 0 4530 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1693_
timestamp 0
transform -1 0 4370 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1694_
timestamp 0
transform 1 0 3230 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1695_
timestamp 0
transform -1 0 3570 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1696_
timestamp 0
transform 1 0 3390 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1697_
timestamp 0
transform -1 0 3430 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1698_
timestamp 0
transform -1 0 2830 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1699_
timestamp 0
transform 1 0 2990 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1700_
timestamp 0
transform -1 0 2850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1701_
timestamp 0
transform 1 0 2550 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1702_
timestamp 0
transform 1 0 2990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1703_
timestamp 0
transform 1 0 3310 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1704_
timestamp 0
transform -1 0 3470 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1705_
timestamp 0
transform -1 0 3290 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1706_
timestamp 0
transform 1 0 3270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1707_
timestamp 0
transform -1 0 2970 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1708_
timestamp 0
transform -1 0 2350 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1709_
timestamp 0
transform 1 0 1050 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1710_
timestamp 0
transform 1 0 10 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1711_
timestamp 0
transform 1 0 1670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1712_
timestamp 0
transform 1 0 2310 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1713_
timestamp 0
transform -1 0 2150 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1714_
timestamp 0
transform -1 0 2210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1715_
timestamp 0
transform 1 0 1990 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1716_
timestamp 0
transform 1 0 1870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1717_
timestamp 0
transform 1 0 1650 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1718_
timestamp 0
transform 1 0 1730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1719_
timestamp 0
transform -1 0 1110 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1720_
timestamp 0
transform -1 0 1270 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1721_
timestamp 0
transform -1 0 710 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1722_
timestamp 0
transform 1 0 170 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1723_
timestamp 0
transform 1 0 230 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1724_
timestamp 0
transform 1 0 190 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1725_
timestamp 0
transform -1 0 30 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1726_
timestamp 0
transform 1 0 330 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1727_
timestamp 0
transform -1 0 490 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1728_
timestamp 0
transform -1 0 930 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1729_
timestamp 0
transform 1 0 630 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1730_
timestamp 0
transform -1 0 770 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1731_
timestamp 0
transform 1 0 190 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1732_
timestamp 0
transform 1 0 370 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1733_
timestamp 0
transform 1 0 470 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1734_
timestamp 0
transform 1 0 630 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1735_
timestamp 0
transform -1 0 950 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1736_
timestamp 0
transform -1 0 530 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1737_
timestamp 0
transform 1 0 630 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1738_
timestamp 0
transform 1 0 770 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1739_
timestamp 0
transform 1 0 1110 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1740_
timestamp 0
transform -1 0 2210 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1741_
timestamp 0
transform -1 0 990 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1742_
timestamp 0
transform -1 0 2070 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1743_
timestamp 0
transform 1 0 2790 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1744_
timestamp 0
transform -1 0 2910 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1745_
timestamp 0
transform 1 0 2650 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1746_
timestamp 0
transform -1 0 2510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1747_
timestamp 0
transform -1 0 2750 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1748_
timestamp 0
transform 1 0 810 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1749_
timestamp 0
transform -1 0 1810 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1750_
timestamp 0
transform -1 0 2070 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1751_
timestamp 0
transform -1 0 1910 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1752_
timestamp 0
transform 1 0 1790 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1753_
timestamp 0
transform -1 0 1610 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1754_
timestamp 0
transform 1 0 1730 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1755_
timestamp 0
transform -1 0 1310 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1756_
timestamp 0
transform -1 0 470 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1757_
timestamp 0
transform 1 0 370 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1758_
timestamp 0
transform -1 0 390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1759_
timestamp 0
transform 1 0 530 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1760_
timestamp 0
transform 1 0 510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1761_
timestamp 0
transform -1 0 990 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1762_
timestamp 0
transform 1 0 810 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1763_
timestamp 0
transform -1 0 870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1764_
timestamp 0
transform 1 0 1930 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1765_
timestamp 0
transform -1 0 2630 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1766_
timestamp 0
transform 1 0 2450 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1767_
timestamp 0
transform 1 0 2490 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1768_
timestamp 0
transform -1 0 2350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1769_
timestamp 0
transform -1 0 2370 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1770_
timestamp 0
transform 1 0 2190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1771_
timestamp 0
transform 1 0 2630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1772_
timestamp 0
transform -1 0 2810 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1773_
timestamp 0
transform 1 0 2330 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1774_
timestamp 0
transform 1 0 1570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1775_
timestamp 0
transform 1 0 1510 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1776_
timestamp 0
transform 1 0 670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1777_
timestamp 0
transform -1 0 1170 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1778_
timestamp 0
transform -1 0 1630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1779_
timestamp 0
transform -1 0 1430 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1780_
timestamp 0
transform 1 0 310 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1781_
timestamp 0
transform 1 0 650 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1782_
timestamp 0
transform 1 0 270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1783_
timestamp 0
transform 1 0 410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1784_
timestamp 0
transform -1 0 570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1785_
timestamp 0
transform -1 0 730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1786_
timestamp 0
transform 1 0 1030 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1787_
timestamp 0
transform 1 0 870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1788_
timestamp 0
transform 1 0 1350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1789_
timestamp 0
transform 1 0 1670 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1790_
timestamp 0
transform -1 0 2190 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1791_
timestamp 0
transform -1 0 1530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1792_
timestamp 0
transform 1 0 1190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1793_
timestamp 0
transform -1 0 850 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1794_
timestamp 0
transform 1 0 1430 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1795_
timestamp 0
transform -1 0 810 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1796_
timestamp 0
transform 1 0 570 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1797_
timestamp 0
transform 1 0 990 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1798_
timestamp 0
transform 1 0 1110 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1799_
timestamp 0
transform 1 0 1250 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1800_
timestamp 0
transform -1 0 1810 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1801_
timestamp 0
transform 1 0 1610 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1802_
timestamp 0
transform 1 0 10 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1803_
timestamp 0
transform 1 0 910 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1804_
timestamp 0
transform -1 0 1050 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1805_
timestamp 0
transform 1 0 130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1806_
timestamp 0
transform 1 0 250 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1807_
timestamp 0
transform 1 0 150 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1808_
timestamp 0
transform 1 0 410 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1809_
timestamp 0
transform 1 0 250 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1810_
timestamp 0
transform 1 0 10 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1811_
timestamp 0
transform -1 0 1030 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1812_
timestamp 0
transform 1 0 850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1813_
timestamp 0
transform 1 0 150 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1814_
timestamp 0
transform 1 0 810 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1815_
timestamp 0
transform 1 0 410 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1816_
timestamp 0
transform 1 0 930 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1817_
timestamp 0
transform -1 0 710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1818_
timestamp 0
transform 1 0 290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1819_
timestamp 0
transform -1 0 1030 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1820_
timestamp 0
transform -1 0 1170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1821_
timestamp 0
transform 1 0 10 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1822_
timestamp 0
transform -1 0 1010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1823_
timestamp 0
transform 1 0 10 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1824_
timestamp 0
transform 1 0 10 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1825_
timestamp 0
transform -1 0 1090 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1826_
timestamp 0
transform -1 0 910 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1827_
timestamp 0
transform 1 0 490 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1828_
timestamp 0
transform 1 0 1730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1829_
timestamp 0
transform 1 0 1550 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1830_
timestamp 0
transform -1 0 1410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1831_
timestamp 0
transform 1 0 910 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1832_
timestamp 0
transform -1 0 750 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1833_
timestamp 0
transform 1 0 570 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1834_
timestamp 0
transform -1 0 30 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1835_
timestamp 0
transform -1 0 470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1836_
timestamp 0
transform 1 0 850 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1837_
timestamp 0
transform -1 0 710 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1838_
timestamp 0
transform 1 0 390 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1839_
timestamp 0
transform -1 0 310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1840_
timestamp 0
transform -1 0 30 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1841_
timestamp 0
transform -1 0 170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1842_
timestamp 0
transform -1 0 1170 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1843_
timestamp 0
transform -1 0 1310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1844_
timestamp 0
transform 1 0 1810 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1845_
timestamp 0
transform 1 0 1970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1846_
timestamp 0
transform -1 0 2930 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1847_
timestamp 0
transform -1 0 3070 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1848_
timestamp 0
transform -1 0 330 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1849_
timestamp 0
transform 1 0 150 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1911_
timestamp 0
transform -1 0 2670 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1912_
timestamp 0
transform -1 0 30 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1913_
timestamp 0
transform 1 0 2370 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1914_
timestamp 0
transform -1 0 30 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1915_
timestamp 0
transform -1 0 30 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1916_
timestamp 0
transform -1 0 2530 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1917_
timestamp 0
transform -1 0 2450 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1918_
timestamp 0
transform -1 0 190 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1919_
timestamp 0
transform -1 0 30 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert0
timestamp 0
transform 1 0 3090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert1
timestamp 0
transform 1 0 2790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert2
timestamp 0
transform 1 0 3230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert3
timestamp 0
transform 1 0 3230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert4
timestamp 0
transform -1 0 2670 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert12
timestamp 0
transform 1 0 3510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert13
timestamp 0
transform 1 0 10 0 1 1310
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert14
timestamp 0
transform 1 0 550 0 1 1830
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert15
timestamp 0
transform 1 0 3550 0 1 2350
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert16
timestamp 0
transform 1 0 770 0 1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert17
timestamp 0
transform 1 0 1070 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert18
timestamp 0
transform -1 0 170 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert19
timestamp 0
transform -1 0 1050 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert20
timestamp 0
transform -1 0 330 0 1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert21
timestamp 0
transform 1 0 3370 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert22
timestamp 0
transform -1 0 3110 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert23
timestamp 0
transform 1 0 3370 0 1 3910
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert24
timestamp 0
transform -1 0 3110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert25
timestamp 0
transform -1 0 3230 0 1 3910
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert5
timestamp 0
transform -1 0 990 0 1 3910
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert6
timestamp 0
transform 1 0 2030 0 1 3390
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert7
timestamp 0
transform 1 0 990 0 1 2350
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert8
timestamp 0
transform -1 0 190 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert9
timestamp 0
transform 1 0 150 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert10
timestamp 0
transform 1 0 2650 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert11
timestamp 0
transform 1 0 1650 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__922_
timestamp 0
transform -1 0 930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__923_
timestamp 0
transform 1 0 1190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__924_
timestamp 0
transform -1 0 2650 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__925_
timestamp 0
transform 1 0 2470 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__926_
timestamp 0
transform -1 0 2530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__927_
timestamp 0
transform -1 0 1090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__928_
timestamp 0
transform -1 0 1930 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__929_
timestamp 0
transform 1 0 2930 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__930_
timestamp 0
transform 1 0 2530 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__931_
timestamp 0
transform -1 0 3610 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__932_
timestamp 0
transform 1 0 2970 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__933_
timestamp 0
transform 1 0 2810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__934_
timestamp 0
transform 1 0 2850 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__935_
timestamp 0
transform 1 0 2690 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__936_
timestamp 0
transform -1 0 3470 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__937_
timestamp 0
transform 1 0 2310 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__938_
timestamp 0
transform 1 0 2110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__939_
timestamp 0
transform 1 0 2350 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__940_
timestamp 0
transform 1 0 1990 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__941_
timestamp 0
transform 1 0 1410 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__942_
timestamp 0
transform -1 0 1650 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__943_
timestamp 0
transform 1 0 1450 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__944_
timestamp 0
transform -1 0 2190 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__945_
timestamp 0
transform 1 0 1470 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__946_
timestamp 0
transform -1 0 4450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__947_
timestamp 0
transform -1 0 930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__948_
timestamp 0
transform 1 0 590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__949_
timestamp 0
transform 1 0 3710 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__950_
timestamp 0
transform 1 0 2150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__951_
timestamp 0
transform -1 0 2310 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__952_
timestamp 0
transform 1 0 3830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__953_
timestamp 0
transform 1 0 490 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__954_
timestamp 0
transform -1 0 650 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__955_
timestamp 0
transform 1 0 2670 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__956_
timestamp 0
transform -1 0 310 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__957_
timestamp 0
transform -1 0 450 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__958_
timestamp 0
transform 1 0 1050 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__959_
timestamp 0
transform -1 0 1690 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__960_
timestamp 0
transform 1 0 2610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__961_
timestamp 0
transform -1 0 2770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__962_
timestamp 0
transform -1 0 2950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__963_
timestamp 0
transform -1 0 2970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__964_
timestamp 0
transform 1 0 1250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__965_
timestamp 0
transform -1 0 1330 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__966_
timestamp 0
transform -1 0 2990 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__967_
timestamp 0
transform 1 0 2650 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__968_
timestamp 0
transform -1 0 2830 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__969_
timestamp 0
transform -1 0 3390 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__970_
timestamp 0
transform -1 0 3070 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__971_
timestamp 0
transform -1 0 3230 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__972_
timestamp 0
transform -1 0 3030 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__973_
timestamp 0
transform -1 0 2470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__974_
timestamp 0
transform -1 0 2870 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__975_
timestamp 0
transform -1 0 2570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__976_
timestamp 0
transform 1 0 2190 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__977_
timestamp 0
transform -1 0 2370 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__978_
timestamp 0
transform -1 0 3710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__979_
timestamp 0
transform 1 0 3250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__980_
timestamp 0
transform -1 0 3550 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__981_
timestamp 0
transform -1 0 3310 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__982_
timestamp 0
transform -1 0 2870 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__983_
timestamp 0
transform -1 0 3150 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__984_
timestamp 0
transform -1 0 3430 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__985_
timestamp 0
transform 1 0 4090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__986_
timestamp 0
transform 1 0 4050 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__987_
timestamp 0
transform -1 0 4210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__988_
timestamp 0
transform 1 0 3650 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__989_
timestamp 0
transform 1 0 2510 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__990_
timestamp 0
transform -1 0 2670 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__991_
timestamp 0
transform 1 0 2770 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__992_
timestamp 0
transform 1 0 2750 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__993_
timestamp 0
transform 1 0 3930 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__994_
timestamp 0
transform -1 0 3990 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__995_
timestamp 0
transform 1 0 3310 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__996_
timestamp 0
transform 1 0 3150 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__997_
timestamp 0
transform 1 0 1690 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__998_
timestamp 0
transform 1 0 1530 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__999_
timestamp 0
transform 1 0 2250 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1000_
timestamp 0
transform -1 0 3090 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1001_
timestamp 0
transform 1 0 2370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1002_
timestamp 0
transform -1 0 2570 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1003_
timestamp 0
transform 1 0 2910 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1004_
timestamp 0
transform 1 0 2750 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1005_
timestamp 0
transform -1 0 1950 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1006_
timestamp 0
transform 1 0 1850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1007_
timestamp 0
transform 1 0 1770 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1008_
timestamp 0
transform 1 0 1510 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1009_
timestamp 0
transform 1 0 1090 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1010_
timestamp 0
transform -1 0 1270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1011_
timestamp 0
transform 1 0 1010 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1012_
timestamp 0
transform 1 0 2310 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1013_
timestamp 0
transform -1 0 3430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1014_
timestamp 0
transform 1 0 890 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1015_
timestamp 0
transform -1 0 1790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1016_
timestamp 0
transform 1 0 1950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1017_
timestamp 0
transform 1 0 2510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1018_
timestamp 0
transform 1 0 2090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1019_
timestamp 0
transform -1 0 750 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1020_
timestamp 0
transform 1 0 890 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1021_
timestamp 0
transform 1 0 1190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1022_
timestamp 0
transform -1 0 1450 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1023_
timestamp 0
transform 1 0 1330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1024_
timestamp 0
transform 1 0 1210 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1025_
timestamp 0
transform -1 0 1510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1026_
timestamp 0
transform 1 0 1350 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1027_
timestamp 0
transform 1 0 1510 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1028_
timestamp 0
transform -1 0 1490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1029_
timestamp 0
transform -1 0 1650 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1030_
timestamp 0
transform -1 0 1530 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1031_
timestamp 0
transform 1 0 1850 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1032_
timestamp 0
transform 1 0 1690 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1033_
timestamp 0
transform 1 0 2290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1034_
timestamp 0
transform 1 0 1610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1035_
timestamp 0
transform 1 0 3850 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1036_
timestamp 0
transform -1 0 1270 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1037_
timestamp 0
transform 1 0 1090 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1038_
timestamp 0
transform -1 0 4590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1039_
timestamp 0
transform -1 0 1570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1040_
timestamp 0
transform 1 0 650 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1041_
timestamp 0
transform 1 0 490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1042_
timestamp 0
transform 1 0 770 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1043_
timestamp 0
transform -1 0 670 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1044_
timestamp 0
transform -1 0 1410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1045_
timestamp 0
transform 1 0 1090 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1046_
timestamp 0
transform 1 0 970 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1047_
timestamp 0
transform 1 0 790 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1048_
timestamp 0
transform 1 0 1210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1049_
timestamp 0
transform -1 0 970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1050_
timestamp 0
transform 1 0 1070 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1051_
timestamp 0
transform 1 0 1390 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1052_
timestamp 0
transform -1 0 1710 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1053_
timestamp 0
transform -1 0 1930 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1054_
timestamp 0
transform 1 0 2310 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1055_
timestamp 0
transform -1 0 1930 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1056_
timestamp 0
transform -1 0 1590 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1057_
timestamp 0
transform -1 0 1750 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1058_
timestamp 0
transform 1 0 1570 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1059_
timestamp 0
transform -1 0 1750 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1060_
timestamp 0
transform 1 0 1870 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1061_
timestamp 0
transform -1 0 2250 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1062_
timestamp 0
transform 1 0 1230 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1063_
timestamp 0
transform -1 0 1750 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1064_
timestamp 0
transform -1 0 3570 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1065_
timestamp 0
transform 1 0 2490 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1066_
timestamp 0
transform -1 0 2490 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1067_
timestamp 0
transform 1 0 2350 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1068_
timestamp 0
transform -1 0 930 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1069_
timestamp 0
transform -1 0 190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1070_
timestamp 0
transform -1 0 350 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1071_
timestamp 0
transform 1 0 210 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1072_
timestamp 0
transform -1 0 50 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1073_
timestamp 0
transform 1 0 330 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1074_
timestamp 0
transform -1 0 230 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1075_
timestamp 0
transform 1 0 30 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1076_
timestamp 0
transform 1 0 330 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1077_
timestamp 0
transform -1 0 510 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1078_
timestamp 0
transform 1 0 990 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1079_
timestamp 0
transform 1 0 650 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1080_
timestamp 0
transform 1 0 1130 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1081_
timestamp 0
transform -1 0 990 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1082_
timestamp 0
transform 1 0 650 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1083_
timestamp 0
transform 1 0 170 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1084_
timestamp 0
transform 1 0 170 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1085_
timestamp 0
transform 1 0 310 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1086_
timestamp 0
transform -1 0 4910 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1087_
timestamp 0
transform -1 0 490 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1088_
timestamp 0
transform -1 0 350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1089_
timestamp 0
transform 1 0 490 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1090_
timestamp 0
transform 1 0 1110 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1091_
timestamp 0
transform 1 0 1470 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1092_
timestamp 0
transform 1 0 1810 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1093_
timestamp 0
transform -1 0 1630 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1094_
timestamp 0
transform 1 0 1950 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1095_
timestamp 0
transform 1 0 2110 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1096_
timestamp 0
transform -1 0 2190 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1097_
timestamp 0
transform 1 0 2030 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1098_
timestamp 0
transform 1 0 2070 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1099_
timestamp 0
transform -1 0 2790 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1100_
timestamp 0
transform 1 0 2630 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1101_
timestamp 0
transform -1 0 830 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1102_
timestamp 0
transform 1 0 30 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1103_
timestamp 0
transform 1 0 1110 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1104_
timestamp 0
transform -1 0 830 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1105_
timestamp 0
transform 1 0 490 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1106_
timestamp 0
transform -1 0 770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1107_
timestamp 0
transform -1 0 50 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1108_
timestamp 0
transform 1 0 630 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1109_
timestamp 0
transform 1 0 150 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1110_
timestamp 0
transform -1 0 50 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1111_
timestamp 0
transform 1 0 450 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1112_
timestamp 0
transform 1 0 1390 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1113_
timestamp 0
transform 1 0 630 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1114_
timestamp 0
transform -1 0 290 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1115_
timestamp 0
transform 1 0 790 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1116_
timestamp 0
transform 1 0 3870 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1117_
timestamp 0
transform -1 0 4870 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1118_
timestamp 0
transform 1 0 4350 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1119_
timestamp 0
transform 1 0 4350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1120_
timestamp 0
transform 1 0 4510 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1121_
timestamp 0
transform -1 0 4410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1122_
timestamp 0
transform 1 0 4630 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1123_
timestamp 0
transform 1 0 4670 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1124_
timestamp 0
transform 1 0 3650 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1125_
timestamp 0
transform 1 0 3810 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1126_
timestamp 0
transform 1 0 3970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1127_
timestamp 0
transform -1 0 3830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1128_
timestamp 0
transform -1 0 3690 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1129_
timestamp 0
transform 1 0 1790 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1130_
timestamp 0
transform 1 0 950 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1131_
timestamp 0
transform 1 0 1230 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1132_
timestamp 0
transform -1 0 3850 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1133_
timestamp 0
transform 1 0 2050 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1134_
timestamp 0
transform 1 0 2130 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1135_
timestamp 0
transform 1 0 1290 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1136_
timestamp 0
transform -1 0 1750 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1137_
timestamp 0
transform 1 0 1550 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1138_
timestamp 0
transform 1 0 1450 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1139_
timestamp 0
transform 1 0 2670 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1140_
timestamp 0
transform 1 0 1290 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1141_
timestamp 0
transform 1 0 1630 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1142_
timestamp 0
transform 1 0 1970 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1143_
timestamp 0
transform 1 0 2310 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1144_
timestamp 0
transform -1 0 3010 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1145_
timestamp 0
transform 1 0 2750 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1146_
timestamp 0
transform 1 0 3150 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1147_
timestamp 0
transform 1 0 2870 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1148_
timestamp 0
transform 1 0 2850 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1149_
timestamp 0
transform 1 0 2670 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1150_
timestamp 0
transform 1 0 3170 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1151_
timestamp 0
transform 1 0 3010 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1152_
timestamp 0
transform 1 0 2450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1153_
timestamp 0
transform -1 0 2850 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1154_
timestamp 0
transform 1 0 2830 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1155_
timestamp 0
transform 1 0 4670 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1156_
timestamp 0
transform 1 0 4610 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1157_
timestamp 0
transform -1 0 5010 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1158_
timestamp 0
transform -1 0 5490 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1159_
timestamp 0
transform -1 0 4810 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1160_
timestamp 0
transform 1 0 4790 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1161_
timestamp 0
transform 1 0 2210 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1162_
timestamp 0
transform -1 0 4030 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1163_
timestamp 0
transform -1 0 4970 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1164_
timestamp 0
transform 1 0 4490 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1165_
timestamp 0
transform -1 0 4830 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1166_
timestamp 0
transform 1 0 4150 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1167_
timestamp 0
transform -1 0 4330 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1168_
timestamp 0
transform 1 0 4510 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1169_
timestamp 0
transform -1 0 4830 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1170_
timestamp 0
transform 1 0 4150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1171_
timestamp 0
transform 1 0 4790 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1172_
timestamp 0
transform 1 0 4990 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1173_
timestamp 0
transform 1 0 810 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1174_
timestamp 0
transform 1 0 3650 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1175_
timestamp 0
transform 1 0 3250 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1176_
timestamp 0
transform 1 0 3310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1177_
timestamp 0
transform -1 0 3410 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1178_
timestamp 0
transform -1 0 3970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1179_
timestamp 0
transform 1 0 3510 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1180_
timestamp 0
transform 1 0 3250 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1181_
timestamp 0
transform 1 0 3530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1182_
timestamp 0
transform 1 0 3690 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1183_
timestamp 0
transform 1 0 4110 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1184_
timestamp 0
transform 1 0 3870 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1185_
timestamp 0
transform 1 0 3490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1186_
timestamp 0
transform 1 0 3630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1187_
timestamp 0
transform 1 0 3790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1188_
timestamp 0
transform 1 0 3690 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1189_
timestamp 0
transform -1 0 4050 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1190_
timestamp 0
transform 1 0 4310 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1191_
timestamp 0
transform -1 0 5150 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1192_
timestamp 0
transform 1 0 3950 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1193_
timestamp 0
transform 1 0 4190 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1194_
timestamp 0
transform -1 0 4470 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1195_
timestamp 0
transform -1 0 3990 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1196_
timestamp 0
transform -1 0 1910 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1197_
timestamp 0
transform 1 0 4270 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1198_
timestamp 0
transform -1 0 4170 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1199_
timestamp 0
transform -1 0 3650 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1200_
timestamp 0
transform 1 0 3450 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1201_
timestamp 0
transform 1 0 4290 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1202_
timestamp 0
transform 1 0 4470 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1203_
timestamp 0
transform 1 0 3790 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1204_
timestamp 0
transform -1 0 4650 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1205_
timestamp 0
transform 1 0 3990 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1206_
timestamp 0
transform 1 0 2490 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1207_
timestamp 0
transform -1 0 4150 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1208_
timestamp 0
transform -1 0 3310 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1209_
timestamp 0
transform -1 0 2970 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1210_
timestamp 0
transform -1 0 3150 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1211_
timestamp 0
transform 1 0 3230 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1212_
timestamp 0
transform 1 0 3310 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1213_
timestamp 0
transform 1 0 3490 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1214_
timestamp 0
transform -1 0 3370 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1215_
timestamp 0
transform -1 0 3030 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1216_
timestamp 0
transform -1 0 2630 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1217_
timestamp 0
transform 1 0 3490 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1218_
timestamp 0
transform 1 0 5050 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1219_
timestamp 0
transform -1 0 5130 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1220_
timestamp 0
transform -1 0 4770 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1221_
timestamp 0
transform 1 0 4570 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1222_
timestamp 0
transform 1 0 4490 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1223_
timestamp 0
transform 1 0 4990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1224_
timestamp 0
transform -1 0 5110 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1225_
timestamp 0
transform 1 0 6090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1226_
timestamp 0
transform 1 0 5950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1227_
timestamp 0
transform -1 0 5330 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1228_
timestamp 0
transform 1 0 5610 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1229_
timestamp 0
transform -1 0 6310 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1230_
timestamp 0
transform 1 0 4950 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1231_
timestamp 0
transform 1 0 5090 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1232_
timestamp 0
transform 1 0 4830 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1233_
timestamp 0
transform -1 0 5150 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1234_
timestamp 0
transform 1 0 5610 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1235_
timestamp 0
transform -1 0 5470 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1236_
timestamp 0
transform -1 0 5450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1237_
timestamp 0
transform 1 0 4970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1238_
timestamp 0
transform 1 0 4510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1239_
timestamp 0
transform -1 0 4690 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1240_
timestamp 0
transform 1 0 5290 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1241_
timestamp 0
transform 1 0 5270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1242_
timestamp 0
transform 1 0 5750 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1243_
timestamp 0
transform -1 0 3390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1244_
timestamp 0
transform 1 0 5590 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1245_
timestamp 0
transform 1 0 4110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1246_
timestamp 0
transform 1 0 4450 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1247_
timestamp 0
transform -1 0 4990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1248_
timestamp 0
transform 1 0 4270 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1249_
timestamp 0
transform 1 0 5090 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1250_
timestamp 0
transform 1 0 5390 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1251_
timestamp 0
transform 1 0 5250 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1252_
timestamp 0
transform 1 0 5690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1253_
timestamp 0
transform -1 0 5730 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1254_
timestamp 0
transform -1 0 5530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1255_
timestamp 0
transform -1 0 4010 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1256_
timestamp 0
transform 1 0 4110 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1257_
timestamp 0
transform 1 0 3670 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1258_
timestamp 0
transform 1 0 4230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1259_
timestamp 0
transform -1 0 5270 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1260_
timestamp 0
transform 1 0 5950 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1261_
timestamp 0
transform 1 0 5910 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1262_
timestamp 0
transform 1 0 5850 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1263_
timestamp 0
transform 1 0 5410 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1264_
timestamp 0
transform 1 0 5590 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1265_
timestamp 0
transform -1 0 5910 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1266_
timestamp 0
transform 1 0 3770 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1267_
timestamp 0
transform 1 0 4630 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1268_
timestamp 0
transform 1 0 5430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1269_
timestamp 0
transform -1 0 5790 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1270_
timestamp 0
transform -1 0 5590 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1271_
timestamp 0
transform 1 0 6210 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1272_
timestamp 0
transform -1 0 6510 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1273_
timestamp 0
transform 1 0 6050 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1274_
timestamp 0
transform 1 0 5730 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1275_
timestamp 0
transform -1 0 6590 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1276_
timestamp 0
transform -1 0 6170 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1277_
timestamp 0
transform 1 0 4410 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1278_
timestamp 0
transform 1 0 4870 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1279_
timestamp 0
transform -1 0 6550 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1280_
timestamp 0
transform -1 0 6070 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1281_
timestamp 0
transform -1 0 5830 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1282_
timestamp 0
transform -1 0 5550 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1283_
timestamp 0
transform 1 0 5430 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1284_
timestamp 0
transform -1 0 6330 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1285_
timestamp 0
transform -1 0 6010 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1286_
timestamp 0
transform -1 0 5910 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1287_
timestamp 0
transform 1 0 5190 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1288_
timestamp 0
transform -1 0 5570 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1289_
timestamp 0
transform -1 0 5390 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1290_
timestamp 0
transform -1 0 5270 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1291_
timestamp 0
transform -1 0 5270 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1292_
timestamp 0
transform 1 0 5410 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1293_
timestamp 0
transform 1 0 4270 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1294_
timestamp 0
transform 1 0 4210 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1295_
timestamp 0
transform -1 0 4690 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1296_
timestamp 0
transform -1 0 4710 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1297_
timestamp 0
transform 1 0 5690 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1298_
timestamp 0
transform -1 0 5730 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1299_
timestamp 0
transform 1 0 5910 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1300_
timestamp 0
transform 1 0 6370 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1301_
timestamp 0
transform -1 0 6510 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1302_
timestamp 0
transform -1 0 4370 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1303_
timestamp 0
transform 1 0 5450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1304_
timestamp 0
transform -1 0 4830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1305_
timestamp 0
transform 1 0 5150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1306_
timestamp 0
transform 1 0 5070 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1307_
timestamp 0
transform 1 0 5350 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1308_
timestamp 0
transform 1 0 5750 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1309_
timestamp 0
transform -1 0 4170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1310_
timestamp 0
transform 1 0 4750 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1311_
timestamp 0
transform -1 0 5310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1312_
timestamp 0
transform 1 0 5410 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1313_
timestamp 0
transform -1 0 5110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1314_
timestamp 0
transform -1 0 5910 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1315_
timestamp 0
transform 1 0 5250 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1316_
timestamp 0
transform -1 0 5590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1317_
timestamp 0
transform 1 0 5610 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1318_
timestamp 0
transform 1 0 5730 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1319_
timestamp 0
transform 1 0 5770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1320_
timestamp 0
transform 1 0 5570 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1321_
timestamp 0
transform 1 0 6050 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1322_
timestamp 0
transform 1 0 6210 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1323_
timestamp 0
transform 1 0 6210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1324_
timestamp 0
transform -1 0 6450 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1325_
timestamp 0
transform 1 0 6250 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1326_
timestamp 0
transform 1 0 4930 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1327_
timestamp 0
transform 1 0 4410 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1328_
timestamp 0
transform 1 0 4130 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1329_
timestamp 0
transform -1 0 4330 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1330_
timestamp 0
transform 1 0 4450 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1331_
timestamp 0
transform 1 0 4590 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1332_
timestamp 0
transform 1 0 5070 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1333_
timestamp 0
transform 1 0 4430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1334_
timestamp 0
transform 1 0 4910 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1335_
timestamp 0
transform 1 0 3970 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1336_
timestamp 0
transform 1 0 5350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1337_
timestamp 0
transform 1 0 5510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1338_
timestamp 0
transform 1 0 4930 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1339_
timestamp 0
transform -1 0 6010 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1340_
timestamp 0
transform -1 0 4650 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1341_
timestamp 0
transform 1 0 3410 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1342_
timestamp 0
transform 1 0 3530 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1343_
timestamp 0
transform -1 0 3850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1344_
timestamp 0
transform -1 0 4250 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1345_
timestamp 0
transform 1 0 4550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1346_
timestamp 0
transform 1 0 5250 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1347_
timestamp 0
transform 1 0 4310 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1348_
timestamp 0
transform 1 0 3690 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1349_
timestamp 0
transform 1 0 5390 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1350_
timestamp 0
transform -1 0 6030 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1351_
timestamp 0
transform 1 0 5570 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1352_
timestamp 0
transform 1 0 4370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1353_
timestamp 0
transform 1 0 5510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1354_
timestamp 0
transform 1 0 6030 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1355_
timestamp 0
transform 1 0 5670 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1356_
timestamp 0
transform 1 0 6170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1357_
timestamp 0
transform 1 0 5670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1358_
timestamp 0
transform 1 0 6490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1359_
timestamp 0
transform -1 0 6270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1360_
timestamp 0
transform 1 0 6010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1361_
timestamp 0
transform 1 0 6070 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1362_
timestamp 0
transform -1 0 6350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1363_
timestamp 0
transform 1 0 5870 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1364_
timestamp 0
transform 1 0 5910 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1365_
timestamp 0
transform -1 0 6410 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1366_
timestamp 0
transform 1 0 6510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1367_
timestamp 0
transform 1 0 6190 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1368_
timestamp 0
transform 1 0 6090 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1369_
timestamp 0
transform 1 0 6550 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1370_
timestamp 0
transform -1 0 6250 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1371_
timestamp 0
transform 1 0 6130 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1372_
timestamp 0
transform 1 0 6210 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1373_
timestamp 0
transform 1 0 6590 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1374_
timestamp 0
transform -1 0 6370 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1375_
timestamp 0
transform -1 0 6190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1376_
timestamp 0
transform -1 0 5890 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1377_
timestamp 0
transform 1 0 6530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1378_
timestamp 0
transform -1 0 6430 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1379_
timestamp 0
transform -1 0 6350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1380_
timestamp 0
transform -1 0 6230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1381_
timestamp 0
transform -1 0 5770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1382_
timestamp 0
transform -1 0 6510 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1383_
timestamp 0
transform -1 0 6390 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1384_
timestamp 0
transform -1 0 6390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1385_
timestamp 0
transform -1 0 6070 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1386_
timestamp 0
transform -1 0 6070 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1387_
timestamp 0
transform 1 0 5290 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1388_
timestamp 0
transform 1 0 4710 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1389_
timestamp 0
transform -1 0 4590 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1390_
timestamp 0
transform -1 0 5030 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1391_
timestamp 0
transform 1 0 4390 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1392_
timestamp 0
transform 1 0 4030 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1393_
timestamp 0
transform 1 0 3870 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1394_
timestamp 0
transform -1 0 5130 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1395_
timestamp 0
transform -1 0 5150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1396_
timestamp 0
transform -1 0 4970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1397_
timestamp 0
transform -1 0 6590 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1398_
timestamp 0
transform 1 0 6610 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1399_
timestamp 0
transform -1 0 6570 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1400_
timestamp 0
transform -1 0 6490 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1401_
timestamp 0
transform -1 0 6430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1402_
timestamp 0
transform -1 0 6550 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1403_
timestamp 0
transform -1 0 5710 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1404_
timestamp 0
transform -1 0 4090 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1405_
timestamp 0
transform 1 0 4910 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1406_
timestamp 0
transform -1 0 4750 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1407_
timestamp 0
transform 1 0 4350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1408_
timestamp 0
transform -1 0 4730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1409_
timestamp 0
transform -1 0 4670 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1410_
timestamp 0
transform -1 0 4810 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1411_
timestamp 0
transform -1 0 4870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1412_
timestamp 0
transform 1 0 4390 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1413_
timestamp 0
transform -1 0 4790 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1414_
timestamp 0
transform 1 0 4750 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1415_
timestamp 0
transform 1 0 4550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1416_
timestamp 0
transform 1 0 5190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1417_
timestamp 0
transform 1 0 5210 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1418_
timestamp 0
transform 1 0 4570 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1419_
timestamp 0
transform 1 0 5010 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1420_
timestamp 0
transform 1 0 4270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1421_
timestamp 0
transform 1 0 4210 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1422_
timestamp 0
transform 1 0 5370 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1423_
timestamp 0
transform 1 0 5690 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1424_
timestamp 0
transform 1 0 5210 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1425_
timestamp 0
transform 1 0 5530 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1426_
timestamp 0
transform 1 0 5530 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1427_
timestamp 0
transform 1 0 5030 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1428_
timestamp 0
transform -1 0 5870 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1429_
timestamp 0
transform 1 0 5730 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1430_
timestamp 0
transform 1 0 6170 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1431_
timestamp 0
transform -1 0 6330 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1432_
timestamp 0
transform 1 0 4870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1433_
timestamp 0
transform -1 0 4290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1434_
timestamp 0
transform 1 0 4690 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1435_
timestamp 0
transform -1 0 4610 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1436_
timestamp 0
transform 1 0 4730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1437_
timestamp 0
transform 1 0 5030 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1438_
timestamp 0
transform 1 0 5190 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1439_
timestamp 0
transform 1 0 3110 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1440_
timestamp 0
transform -1 0 4930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1441_
timestamp 0
transform 1 0 4110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1442_
timestamp 0
transform 1 0 5350 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1443_
timestamp 0
transform 1 0 5530 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1444_
timestamp 0
transform 1 0 3670 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1445_
timestamp 0
transform 1 0 3150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1446_
timestamp 0
transform -1 0 3950 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1447_
timestamp 0
transform -1 0 4530 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1448_
timestamp 0
transform 1 0 4950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1449_
timestamp 0
transform 1 0 4470 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1450_
timestamp 0
transform 1 0 4950 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1451_
timestamp 0
transform 1 0 4650 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1452_
timestamp 0
transform 1 0 5310 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1453_
timestamp 0
transform -1 0 5690 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1454_
timestamp 0
transform 1 0 4150 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1455_
timestamp 0
transform 1 0 4010 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1456_
timestamp 0
transform -1 0 5370 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1457_
timestamp 0
transform 1 0 5470 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1458_
timestamp 0
transform 1 0 5510 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1459_
timestamp 0
transform 1 0 5610 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1460_
timestamp 0
transform 1 0 5850 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1461_
timestamp 0
transform 1 0 6010 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1462_
timestamp 0
transform -1 0 5070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1463_
timestamp 0
transform 1 0 5290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1464_
timestamp 0
transform 1 0 5850 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1465_
timestamp 0
transform 1 0 5130 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1466_
timestamp 0
transform 1 0 5750 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1467_
timestamp 0
transform 1 0 5870 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1468_
timestamp 0
transform -1 0 6050 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1469_
timestamp 0
transform 1 0 5450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1470_
timestamp 0
transform 1 0 5910 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1471_
timestamp 0
transform -1 0 5970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1472_
timestamp 0
transform 1 0 6110 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1473_
timestamp 0
transform 1 0 6370 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1474_
timestamp 0
transform -1 0 6550 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1475_
timestamp 0
transform 1 0 6130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1476_
timestamp 0
transform 1 0 5790 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1477_
timestamp 0
transform 1 0 6370 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1478_
timestamp 0
transform -1 0 6470 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1479_
timestamp 0
transform 1 0 6210 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1480_
timestamp 0
transform -1 0 6310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1481_
timestamp 0
transform 1 0 6550 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1482_
timestamp 0
transform 1 0 6610 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1483_
timestamp 0
transform -1 0 6630 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1484_
timestamp 0
transform 1 0 6510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1485_
timestamp 0
transform -1 0 6650 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1486_
timestamp 0
transform -1 0 6290 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1487_
timestamp 0
transform -1 0 6490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1488_
timestamp 0
transform -1 0 4830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1489_
timestamp 0
transform 1 0 3970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1490_
timestamp 0
transform 1 0 4010 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1491_
timestamp 0
transform -1 0 5030 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1492_
timestamp 0
transform 1 0 4830 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1493_
timestamp 0
transform 1 0 6370 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1494_
timestamp 0
transform 1 0 6490 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1495_
timestamp 0
transform -1 0 5850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1496_
timestamp 0
transform 1 0 6270 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1497_
timestamp 0
transform -1 0 6090 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1498_
timestamp 0
transform 1 0 6190 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1499_
timestamp 0
transform 1 0 5170 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1500_
timestamp 0
transform -1 0 4570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1501_
timestamp 0
transform 1 0 4070 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1502_
timestamp 0
transform 1 0 4810 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1503_
timestamp 0
transform -1 0 4710 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1504_
timestamp 0
transform 1 0 5110 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1505_
timestamp 0
transform 1 0 4830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1506_
timestamp 0
transform -1 0 4510 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1507_
timestamp 0
transform 1 0 4510 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1508_
timestamp 0
transform -1 0 5010 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1509_
timestamp 0
transform 1 0 5130 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1510_
timestamp 0
transform 1 0 4850 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1511_
timestamp 0
transform 1 0 5190 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1512_
timestamp 0
transform -1 0 5330 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1513_
timestamp 0
transform 1 0 4950 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1514_
timestamp 0
transform 1 0 4950 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1515_
timestamp 0
transform 1 0 5010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1516_
timestamp 0
transform 1 0 5530 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1517_
timestamp 0
transform 1 0 5470 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1518_
timestamp 0
transform 1 0 5110 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1519_
timestamp 0
transform 1 0 5330 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1520_
timestamp 0
transform 1 0 5290 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1521_
timestamp 0
transform 1 0 5370 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1522_
timestamp 0
transform 1 0 5450 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1523_
timestamp 0
transform 1 0 5610 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1524_
timestamp 0
transform -1 0 5150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1525_
timestamp 0
transform -1 0 5850 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1526_
timestamp 0
transform 1 0 3630 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1527_
timestamp 0
transform 1 0 3130 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1528_
timestamp 0
transform -1 0 3950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1529_
timestamp 0
transform 1 0 3470 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1530_
timestamp 0
transform 1 0 3770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1531_
timestamp 0
transform 1 0 4550 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1532_
timestamp 0
transform -1 0 3590 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1533_
timestamp 0
transform -1 0 3850 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1534_
timestamp 0
transform -1 0 4390 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1535_
timestamp 0
transform -1 0 4430 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1536_
timestamp 0
transform 1 0 4050 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1537_
timestamp 0
transform 1 0 4230 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1538_
timestamp 0
transform 1 0 4370 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1539_
timestamp 0
transform 1 0 4250 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1540_
timestamp 0
transform 1 0 5630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1541_
timestamp 0
transform -1 0 5810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1542_
timestamp 0
transform -1 0 5230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1543_
timestamp 0
transform 1 0 5670 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1544_
timestamp 0
transform -1 0 5730 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1545_
timestamp 0
transform -1 0 5650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1546_
timestamp 0
transform 1 0 6070 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1547_
timestamp 0
transform 1 0 5870 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1548_
timestamp 0
transform -1 0 5950 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1549_
timestamp 0
transform 1 0 6250 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1550_
timestamp 0
transform -1 0 6270 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1551_
timestamp 0
transform 1 0 5590 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1552_
timestamp 0
transform 1 0 6010 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1553_
timestamp 0
transform 1 0 6070 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1554_
timestamp 0
transform 1 0 5790 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1555_
timestamp 0
transform -1 0 6030 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1556_
timestamp 0
transform 1 0 5950 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1557_
timestamp 0
transform -1 0 6130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1558_
timestamp 0
transform 1 0 6370 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1559_
timestamp 0
transform 1 0 6570 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1560_
timestamp 0
transform 1 0 6030 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1561_
timestamp 0
transform -1 0 6570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1562_
timestamp 0
transform -1 0 6570 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1563_
timestamp 0
transform -1 0 6410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1564_
timestamp 0
transform 1 0 6190 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1565_
timestamp 0
transform 1 0 6350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1566_
timestamp 0
transform -1 0 6550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1567_
timestamp 0
transform -1 0 4450 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1568_
timestamp 0
transform 1 0 4170 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1569_
timestamp 0
transform -1 0 4210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1570_
timestamp 0
transform -1 0 3730 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1571_
timestamp 0
transform 1 0 6190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1572_
timestamp 0
transform -1 0 4310 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1573_
timestamp 0
transform -1 0 3670 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1574_
timestamp 0
transform 1 0 6410 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1575_
timestamp 0
transform 1 0 6430 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1576_
timestamp 0
transform 1 0 5450 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1577_
timestamp 0
transform -1 0 5470 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1578_
timestamp 0
transform -1 0 5930 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1579_
timestamp 0
transform -1 0 4670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1580_
timestamp 0
transform 1 0 4370 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1581_
timestamp 0
transform -1 0 3010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1582_
timestamp 0
transform -1 0 2810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1583_
timestamp 0
transform -1 0 2870 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1584_
timestamp 0
transform -1 0 3010 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1585_
timestamp 0
transform 1 0 3150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1586_
timestamp 0
transform 1 0 2670 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1587_
timestamp 0
transform 1 0 2790 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1588_
timestamp 0
transform -1 0 1970 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1589_
timestamp 0
transform -1 0 2670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1590_
timestamp 0
transform 1 0 2910 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1591_
timestamp 0
transform 1 0 3870 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1592_
timestamp 0
transform -1 0 3730 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1593_
timestamp 0
transform -1 0 3750 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1594_
timestamp 0
transform 1 0 3070 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1595_
timestamp 0
transform 1 0 2990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1596_
timestamp 0
transform -1 0 4050 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1597_
timestamp 0
transform -1 0 4210 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1598_
timestamp 0
transform 1 0 4050 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1599_
timestamp 0
transform -1 0 4230 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1600_
timestamp 0
transform 1 0 3550 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1601_
timestamp 0
transform 1 0 3890 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1602_
timestamp 0
transform -1 0 3890 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1603_
timestamp 0
transform 1 0 4790 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1604_
timestamp 0
transform 1 0 3650 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1605_
timestamp 0
transform 1 0 3490 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1606_
timestamp 0
transform 1 0 1370 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1607_
timestamp 0
transform -1 0 3350 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1608_
timestamp 0
transform -1 0 2710 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1609_
timestamp 0
transform 1 0 3130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1610_
timestamp 0
transform -1 0 2390 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1611_
timestamp 0
transform -1 0 2550 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1612_
timestamp 0
transform 1 0 1510 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1613_
timestamp 0
transform 1 0 3270 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1614_
timestamp 0
transform 1 0 3410 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1615_
timestamp 0
transform 1 0 3770 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1616_
timestamp 0
transform 1 0 3130 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1617_
timestamp 0
transform -1 0 3590 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1618_
timestamp 0
transform 1 0 4210 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1619_
timestamp 0
transform -1 0 4670 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1620_
timestamp 0
transform 1 0 3750 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1621_
timestamp 0
transform 1 0 3430 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1622_
timestamp 0
transform 1 0 3930 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1623_
timestamp 0
transform 1 0 4950 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1624_
timestamp 0
transform 1 0 5910 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1625_
timestamp 0
transform 1 0 5750 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1626_
timestamp 0
transform 1 0 4190 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1627_
timestamp 0
transform -1 0 4530 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1628_
timestamp 0
transform 1 0 4830 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1629_
timestamp 0
transform 1 0 6230 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1630_
timestamp 0
transform -1 0 5770 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1631_
timestamp 0
transform 1 0 4670 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1632_
timestamp 0
transform 1 0 5570 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1633_
timestamp 0
transform 1 0 6410 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1634_
timestamp 0
transform 1 0 6190 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1635_
timestamp 0
transform -1 0 6450 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1636_
timestamp 0
transform 1 0 5110 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1637_
timestamp 0
transform -1 0 6090 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1638_
timestamp 0
transform 1 0 5270 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1639_
timestamp 0
transform 1 0 4670 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1640_
timestamp 0
transform 1 0 3510 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1641_
timestamp 0
transform 1 0 3330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1642_
timestamp 0
transform 1 0 3550 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1643_
timestamp 0
transform 1 0 2210 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1644_
timestamp 0
transform -1 0 3170 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1645_
timestamp 0
transform -1 0 5310 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1646_
timestamp 0
transform -1 0 5150 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1647_
timestamp 0
transform 1 0 3710 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1648_
timestamp 0
transform -1 0 3770 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1649_
timestamp 0
transform -1 0 4050 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1650_
timestamp 0
transform -1 0 3430 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1651_
timestamp 0
transform -1 0 3570 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1652_
timestamp 0
transform -1 0 2530 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1653_
timestamp 0
transform 1 0 2490 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1654_
timestamp 0
transform -1 0 2390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1655_
timestamp 0
transform -1 0 2190 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1656_
timestamp 0
transform 1 0 1670 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1657_
timestamp 0
transform -1 0 2070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1658_
timestamp 0
transform 1 0 1810 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1659_
timestamp 0
transform -1 0 2030 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1660_
timestamp 0
transform -1 0 2250 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1661_
timestamp 0
transform 1 0 2090 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1662_
timestamp 0
transform 1 0 2190 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1663_
timestamp 0
transform -1 0 1930 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1664_
timestamp 0
transform -1 0 1630 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1665_
timestamp 0
transform -1 0 1450 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1666_
timestamp 0
transform -1 0 1870 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1667_
timestamp 0
transform 1 0 1450 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1668_
timestamp 0
transform 1 0 1990 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1669_
timestamp 0
transform 1 0 2330 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1670_
timestamp 0
transform 1 0 1290 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1671_
timestamp 0
transform -1 0 1750 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1672_
timestamp 0
transform 1 0 1830 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1673_
timestamp 0
transform -1 0 50 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1674_
timestamp 0
transform -1 0 50 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1675_
timestamp 0
transform 1 0 30 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1676_
timestamp 0
transform 1 0 190 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1677_
timestamp 0
transform 1 0 330 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1678_
timestamp 0
transform 1 0 2170 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1679_
timestamp 0
transform -1 0 1690 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1680_
timestamp 0
transform -1 0 1510 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1681_
timestamp 0
transform 1 0 1210 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1682_
timestamp 0
transform -1 0 1350 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1683_
timestamp 0
transform 1 0 2590 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1684_
timestamp 0
transform -1 0 2470 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1685_
timestamp 0
transform -1 0 3270 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1686_
timestamp 0
transform 1 0 3870 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1687_
timestamp 0
transform -1 0 4370 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1688_
timestamp 0
transform 1 0 2770 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1689_
timestamp 0
transform -1 0 2950 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1690_
timestamp 0
transform -1 0 3110 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1691_
timestamp 0
transform -1 0 4070 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1692_
timestamp 0
transform -1 0 4550 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1693_
timestamp 0
transform -1 0 4390 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1694_
timestamp 0
transform 1 0 3250 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1695_
timestamp 0
transform -1 0 3590 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1696_
timestamp 0
transform 1 0 3410 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1697_
timestamp 0
transform -1 0 3450 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1698_
timestamp 0
transform -1 0 2850 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1699_
timestamp 0
transform 1 0 3010 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1700_
timestamp 0
transform -1 0 2870 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1701_
timestamp 0
transform 1 0 2570 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1702_
timestamp 0
transform 1 0 3010 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1703_
timestamp 0
transform 1 0 3330 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1704_
timestamp 0
transform -1 0 3490 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1705_
timestamp 0
transform -1 0 3310 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1706_
timestamp 0
transform 1 0 3290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1707_
timestamp 0
transform -1 0 2990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1708_
timestamp 0
transform -1 0 2370 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1709_
timestamp 0
transform 1 0 1070 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1710_
timestamp 0
transform 1 0 30 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1711_
timestamp 0
transform 1 0 1690 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1712_
timestamp 0
transform 1 0 2330 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1713_
timestamp 0
transform -1 0 2170 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1714_
timestamp 0
transform -1 0 2230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1715_
timestamp 0
transform 1 0 2010 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1716_
timestamp 0
transform 1 0 1890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1717_
timestamp 0
transform 1 0 1670 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1718_
timestamp 0
transform 1 0 1750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1719_
timestamp 0
transform -1 0 1130 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1720_
timestamp 0
transform -1 0 1290 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1721_
timestamp 0
transform -1 0 730 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1722_
timestamp 0
transform 1 0 190 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1723_
timestamp 0
transform 1 0 250 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1724_
timestamp 0
transform 1 0 210 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1725_
timestamp 0
transform -1 0 50 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1726_
timestamp 0
transform 1 0 350 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1727_
timestamp 0
transform -1 0 510 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1728_
timestamp 0
transform -1 0 950 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1729_
timestamp 0
transform 1 0 650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1730_
timestamp 0
transform -1 0 790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1731_
timestamp 0
transform 1 0 210 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1732_
timestamp 0
transform 1 0 390 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1733_
timestamp 0
transform 1 0 490 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1734_
timestamp 0
transform 1 0 650 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1735_
timestamp 0
transform -1 0 970 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1736_
timestamp 0
transform -1 0 550 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1737_
timestamp 0
transform 1 0 650 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1738_
timestamp 0
transform 1 0 790 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1739_
timestamp 0
transform 1 0 1130 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1740_
timestamp 0
transform -1 0 2230 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1741_
timestamp 0
transform -1 0 1010 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1742_
timestamp 0
transform -1 0 2090 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1743_
timestamp 0
transform 1 0 2810 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1744_
timestamp 0
transform -1 0 2930 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1745_
timestamp 0
transform 1 0 2670 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1746_
timestamp 0
transform -1 0 2530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1747_
timestamp 0
transform -1 0 2770 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1748_
timestamp 0
transform 1 0 830 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1749_
timestamp 0
transform -1 0 1830 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1750_
timestamp 0
transform -1 0 2090 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1751_
timestamp 0
transform -1 0 1930 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1752_
timestamp 0
transform 1 0 1810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1753_
timestamp 0
transform -1 0 1630 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1754_
timestamp 0
transform 1 0 1750 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1755_
timestamp 0
transform -1 0 1330 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1756_
timestamp 0
transform -1 0 490 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1757_
timestamp 0
transform 1 0 390 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1758_
timestamp 0
transform -1 0 410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1759_
timestamp 0
transform 1 0 550 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1760_
timestamp 0
transform 1 0 530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1761_
timestamp 0
transform -1 0 1010 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1762_
timestamp 0
transform 1 0 830 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1763_
timestamp 0
transform -1 0 890 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1764_
timestamp 0
transform 1 0 1950 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1765_
timestamp 0
transform -1 0 2650 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1766_
timestamp 0
transform 1 0 2470 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1767_
timestamp 0
transform 1 0 2510 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1768_
timestamp 0
transform -1 0 2370 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1769_
timestamp 0
transform -1 0 2390 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1770_
timestamp 0
transform 1 0 2210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1771_
timestamp 0
transform 1 0 2650 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1772_
timestamp 0
transform -1 0 2830 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1773_
timestamp 0
transform 1 0 2350 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1774_
timestamp 0
transform 1 0 1590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1775_
timestamp 0
transform 1 0 1530 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1776_
timestamp 0
transform 1 0 690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1777_
timestamp 0
transform -1 0 1190 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1778_
timestamp 0
transform -1 0 1650 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1779_
timestamp 0
transform -1 0 1450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1780_
timestamp 0
transform 1 0 330 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1781_
timestamp 0
transform 1 0 670 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1782_
timestamp 0
transform 1 0 290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1783_
timestamp 0
transform 1 0 430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1784_
timestamp 0
transform -1 0 590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1785_
timestamp 0
transform -1 0 750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1786_
timestamp 0
transform 1 0 1050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1787_
timestamp 0
transform 1 0 890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1788_
timestamp 0
transform 1 0 1370 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1789_
timestamp 0
transform 1 0 1690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1790_
timestamp 0
transform -1 0 2210 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1791_
timestamp 0
transform -1 0 1550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1792_
timestamp 0
transform 1 0 1210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1793_
timestamp 0
transform -1 0 870 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1794_
timestamp 0
transform 1 0 1450 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1795_
timestamp 0
transform -1 0 830 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1796_
timestamp 0
transform 1 0 590 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1797_
timestamp 0
transform 1 0 1010 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1798_
timestamp 0
transform 1 0 1130 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1799_
timestamp 0
transform 1 0 1270 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1800_
timestamp 0
transform -1 0 1830 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1801_
timestamp 0
transform 1 0 1630 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1802_
timestamp 0
transform 1 0 30 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1803_
timestamp 0
transform 1 0 930 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1804_
timestamp 0
transform -1 0 1070 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1805_
timestamp 0
transform 1 0 150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1806_
timestamp 0
transform 1 0 270 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1807_
timestamp 0
transform 1 0 170 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1808_
timestamp 0
transform 1 0 430 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1809_
timestamp 0
transform 1 0 270 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1810_
timestamp 0
transform 1 0 30 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1811_
timestamp 0
transform -1 0 1050 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1812_
timestamp 0
transform 1 0 870 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1813_
timestamp 0
transform 1 0 170 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1814_
timestamp 0
transform 1 0 830 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1815_
timestamp 0
transform 1 0 430 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1816_
timestamp 0
transform 1 0 950 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1817_
timestamp 0
transform -1 0 730 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1818_
timestamp 0
transform 1 0 310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1819_
timestamp 0
transform -1 0 1050 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1820_
timestamp 0
transform -1 0 1190 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1821_
timestamp 0
transform 1 0 30 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1822_
timestamp 0
transform -1 0 1030 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1823_
timestamp 0
transform 1 0 30 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1824_
timestamp 0
transform 1 0 30 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1825_
timestamp 0
transform -1 0 1110 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1826_
timestamp 0
transform -1 0 930 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1827_
timestamp 0
transform 1 0 510 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1828_
timestamp 0
transform 1 0 1750 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1829_
timestamp 0
transform 1 0 1570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1830_
timestamp 0
transform -1 0 1430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1831_
timestamp 0
transform 1 0 930 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1832_
timestamp 0
transform -1 0 770 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1833_
timestamp 0
transform 1 0 590 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1834_
timestamp 0
transform -1 0 50 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1835_
timestamp 0
transform -1 0 490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1836_
timestamp 0
transform 1 0 870 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1837_
timestamp 0
transform -1 0 730 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1838_
timestamp 0
transform 1 0 410 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1839_
timestamp 0
transform -1 0 330 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1840_
timestamp 0
transform -1 0 50 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1841_
timestamp 0
transform -1 0 190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1842_
timestamp 0
transform -1 0 1190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1843_
timestamp 0
transform -1 0 1330 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1844_
timestamp 0
transform 1 0 1830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1845_
timestamp 0
transform 1 0 1990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1846_
timestamp 0
transform -1 0 2950 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1847_
timestamp 0
transform -1 0 3090 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1848_
timestamp 0
transform -1 0 350 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1849_
timestamp 0
transform 1 0 170 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1911_
timestamp 0
transform -1 0 2690 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1912_
timestamp 0
transform -1 0 50 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1913_
timestamp 0
transform 1 0 2390 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1914_
timestamp 0
transform -1 0 50 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1915_
timestamp 0
transform -1 0 50 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1916_
timestamp 0
transform -1 0 2550 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1917_
timestamp 0
transform -1 0 2470 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1918_
timestamp 0
transform -1 0 210 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1919_
timestamp 0
transform -1 0 50 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert0
timestamp 0
transform 1 0 3110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert1
timestamp 0
transform 1 0 2810 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert2
timestamp 0
transform 1 0 3250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert3
timestamp 0
transform 1 0 3250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert4
timestamp 0
transform -1 0 2690 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert12
timestamp 0
transform 1 0 3530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert13
timestamp 0
transform 1 0 30 0 1 1310
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert14
timestamp 0
transform 1 0 570 0 1 1830
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert15
timestamp 0
transform 1 0 3570 0 1 2350
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert16
timestamp 0
transform 1 0 790 0 1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert17
timestamp 0
transform 1 0 1090 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert18
timestamp 0
transform -1 0 190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert19
timestamp 0
transform -1 0 1070 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert20
timestamp 0
transform -1 0 350 0 1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert21
timestamp 0
transform 1 0 3390 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert22
timestamp 0
transform -1 0 3130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert23
timestamp 0
transform 1 0 3390 0 1 3910
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert24
timestamp 0
transform -1 0 3130 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert25
timestamp 0
transform -1 0 3250 0 1 3910
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert5
timestamp 0
transform -1 0 1010 0 1 3910
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert6
timestamp 0
transform 1 0 2050 0 1 3390
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert7
timestamp 0
transform 1 0 1010 0 1 2350
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert8
timestamp 0
transform -1 0 210 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert9
timestamp 0
transform 1 0 170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert10
timestamp 0
transform 1 0 2670 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert11
timestamp 0
transform 1 0 1670 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__922_
timestamp 0
transform -1 0 950 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__923_
timestamp 0
transform 1 0 1210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__924_
timestamp 0
transform -1 0 2670 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__925_
timestamp 0
transform 1 0 2490 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__926_
timestamp 0
transform -1 0 2550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__927_
timestamp 0
transform -1 0 1110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__928_
timestamp 0
transform -1 0 1950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__929_
timestamp 0
transform 1 0 2950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__930_
timestamp 0
transform 1 0 2550 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__931_
timestamp 0
transform -1 0 3630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__932_
timestamp 0
transform 1 0 2990 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__933_
timestamp 0
transform 1 0 2830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__934_
timestamp 0
transform 1 0 2870 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__935_
timestamp 0
transform 1 0 2710 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__936_
timestamp 0
transform -1 0 3490 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__937_
timestamp 0
transform 1 0 2330 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__938_
timestamp 0
transform 1 0 2130 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__939_
timestamp 0
transform 1 0 2370 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__940_
timestamp 0
transform 1 0 2010 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__941_
timestamp 0
transform 1 0 1430 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__942_
timestamp 0
transform -1 0 1670 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__943_
timestamp 0
transform 1 0 1470 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__944_
timestamp 0
transform -1 0 2210 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__945_
timestamp 0
transform 1 0 1490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__946_
timestamp 0
transform -1 0 4470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__947_
timestamp 0
transform -1 0 950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__948_
timestamp 0
transform 1 0 610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__949_
timestamp 0
transform 1 0 3730 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__950_
timestamp 0
transform 1 0 2170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__951_
timestamp 0
transform -1 0 2330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__952_
timestamp 0
transform 1 0 3850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__953_
timestamp 0
transform 1 0 510 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__954_
timestamp 0
transform -1 0 670 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__955_
timestamp 0
transform 1 0 2690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__956_
timestamp 0
transform -1 0 330 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__957_
timestamp 0
transform -1 0 470 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__958_
timestamp 0
transform 1 0 1070 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__959_
timestamp 0
transform -1 0 1710 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__960_
timestamp 0
transform 1 0 2630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__961_
timestamp 0
transform -1 0 2790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__962_
timestamp 0
transform -1 0 2970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__963_
timestamp 0
transform -1 0 2990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__964_
timestamp 0
transform 1 0 1270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__965_
timestamp 0
transform -1 0 1350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__966_
timestamp 0
transform -1 0 3010 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__967_
timestamp 0
transform 1 0 2670 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__968_
timestamp 0
transform -1 0 2850 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__969_
timestamp 0
transform -1 0 3410 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__970_
timestamp 0
transform -1 0 3090 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__971_
timestamp 0
transform -1 0 3250 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__972_
timestamp 0
transform -1 0 3050 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__973_
timestamp 0
transform -1 0 2490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__974_
timestamp 0
transform -1 0 2890 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__975_
timestamp 0
transform -1 0 2590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__976_
timestamp 0
transform 1 0 2210 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__977_
timestamp 0
transform -1 0 2390 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__978_
timestamp 0
transform -1 0 3730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__979_
timestamp 0
transform 1 0 3270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__980_
timestamp 0
transform -1 0 3570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__981_
timestamp 0
transform -1 0 3330 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__982_
timestamp 0
transform -1 0 2890 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__983_
timestamp 0
transform -1 0 3170 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__984_
timestamp 0
transform -1 0 3450 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__985_
timestamp 0
transform 1 0 4110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__986_
timestamp 0
transform 1 0 4070 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__987_
timestamp 0
transform -1 0 4230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__988_
timestamp 0
transform 1 0 3670 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__989_
timestamp 0
transform 1 0 2530 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__990_
timestamp 0
transform -1 0 2690 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__991_
timestamp 0
transform 1 0 2790 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__992_
timestamp 0
transform 1 0 2770 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__993_
timestamp 0
transform 1 0 3950 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__994_
timestamp 0
transform -1 0 4010 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__995_
timestamp 0
transform 1 0 3330 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__996_
timestamp 0
transform 1 0 3170 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__997_
timestamp 0
transform 1 0 1710 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__998_
timestamp 0
transform 1 0 1550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__999_
timestamp 0
transform 1 0 2270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1000_
timestamp 0
transform -1 0 3110 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1001_
timestamp 0
transform 1 0 2390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1002_
timestamp 0
transform -1 0 2590 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1003_
timestamp 0
transform 1 0 2930 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1004_
timestamp 0
transform 1 0 2770 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1005_
timestamp 0
transform -1 0 1970 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1006_
timestamp 0
transform 1 0 1870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1007_
timestamp 0
transform 1 0 1790 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1008_
timestamp 0
transform 1 0 1530 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1009_
timestamp 0
transform 1 0 1110 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1010_
timestamp 0
transform -1 0 1290 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1011_
timestamp 0
transform 1 0 1030 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1012_
timestamp 0
transform 1 0 2330 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1013_
timestamp 0
transform -1 0 3450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1014_
timestamp 0
transform 1 0 910 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1015_
timestamp 0
transform -1 0 1810 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1016_
timestamp 0
transform 1 0 1970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1017_
timestamp 0
transform 1 0 2530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1018_
timestamp 0
transform 1 0 2110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1019_
timestamp 0
transform -1 0 770 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1020_
timestamp 0
transform 1 0 910 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1021_
timestamp 0
transform 1 0 1210 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1022_
timestamp 0
transform -1 0 1470 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1023_
timestamp 0
transform 1 0 1350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1024_
timestamp 0
transform 1 0 1230 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1025_
timestamp 0
transform -1 0 1530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1026_
timestamp 0
transform 1 0 1370 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1027_
timestamp 0
transform 1 0 1530 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1028_
timestamp 0
transform -1 0 1510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1029_
timestamp 0
transform -1 0 1670 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1030_
timestamp 0
transform -1 0 1550 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1031_
timestamp 0
transform 1 0 1870 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1032_
timestamp 0
transform 1 0 1710 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1033_
timestamp 0
transform 1 0 2310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1034_
timestamp 0
transform 1 0 1630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1035_
timestamp 0
transform 1 0 3870 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1036_
timestamp 0
transform -1 0 1290 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1037_
timestamp 0
transform 1 0 1110 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1038_
timestamp 0
transform -1 0 4610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1039_
timestamp 0
transform -1 0 1590 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1040_
timestamp 0
transform 1 0 670 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1041_
timestamp 0
transform 1 0 510 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1042_
timestamp 0
transform 1 0 790 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1043_
timestamp 0
transform -1 0 690 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1044_
timestamp 0
transform -1 0 1430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1045_
timestamp 0
transform 1 0 1110 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1046_
timestamp 0
transform 1 0 990 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1047_
timestamp 0
transform 1 0 810 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1048_
timestamp 0
transform 1 0 1230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1049_
timestamp 0
transform -1 0 990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1050_
timestamp 0
transform 1 0 1090 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1051_
timestamp 0
transform 1 0 1410 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1052_
timestamp 0
transform -1 0 1730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1053_
timestamp 0
transform -1 0 1950 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1054_
timestamp 0
transform 1 0 2330 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1055_
timestamp 0
transform -1 0 1950 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1056_
timestamp 0
transform -1 0 1610 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1057_
timestamp 0
transform -1 0 1770 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1058_
timestamp 0
transform 1 0 1590 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1059_
timestamp 0
transform -1 0 1770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1060_
timestamp 0
transform 1 0 1890 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1061_
timestamp 0
transform -1 0 2270 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1062_
timestamp 0
transform 1 0 1250 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1063_
timestamp 0
transform -1 0 1770 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1064_
timestamp 0
transform -1 0 3590 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1065_
timestamp 0
transform 1 0 2510 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1066_
timestamp 0
transform -1 0 2510 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1067_
timestamp 0
transform 1 0 2370 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1068_
timestamp 0
transform -1 0 950 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1069_
timestamp 0
transform -1 0 210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1070_
timestamp 0
transform -1 0 370 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1071_
timestamp 0
transform 1 0 230 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1072_
timestamp 0
transform -1 0 70 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1073_
timestamp 0
transform 1 0 350 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1074_
timestamp 0
transform -1 0 250 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1075_
timestamp 0
transform 1 0 50 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1076_
timestamp 0
transform 1 0 350 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1077_
timestamp 0
transform -1 0 530 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1078_
timestamp 0
transform 1 0 1010 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1079_
timestamp 0
transform 1 0 670 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1080_
timestamp 0
transform 1 0 1150 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1081_
timestamp 0
transform -1 0 1010 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1082_
timestamp 0
transform 1 0 670 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1083_
timestamp 0
transform 1 0 190 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1084_
timestamp 0
transform 1 0 190 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1085_
timestamp 0
transform 1 0 330 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1086_
timestamp 0
transform -1 0 4930 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1087_
timestamp 0
transform -1 0 510 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1088_
timestamp 0
transform -1 0 370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1089_
timestamp 0
transform 1 0 510 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1090_
timestamp 0
transform 1 0 1130 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1091_
timestamp 0
transform 1 0 1490 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1092_
timestamp 0
transform 1 0 1830 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1093_
timestamp 0
transform -1 0 1650 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1094_
timestamp 0
transform 1 0 1970 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1095_
timestamp 0
transform 1 0 2130 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1096_
timestamp 0
transform -1 0 2210 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1097_
timestamp 0
transform 1 0 2050 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1098_
timestamp 0
transform 1 0 2090 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1099_
timestamp 0
transform -1 0 2810 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1100_
timestamp 0
transform 1 0 2650 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1101_
timestamp 0
transform -1 0 850 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1102_
timestamp 0
transform 1 0 50 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1103_
timestamp 0
transform 1 0 1130 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1104_
timestamp 0
transform -1 0 850 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1105_
timestamp 0
transform 1 0 510 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1106_
timestamp 0
transform -1 0 790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1107_
timestamp 0
transform -1 0 70 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1108_
timestamp 0
transform 1 0 650 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1109_
timestamp 0
transform 1 0 170 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1110_
timestamp 0
transform -1 0 70 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1111_
timestamp 0
transform 1 0 470 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1112_
timestamp 0
transform 1 0 1410 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1113_
timestamp 0
transform 1 0 650 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1114_
timestamp 0
transform -1 0 310 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1115_
timestamp 0
transform 1 0 810 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1116_
timestamp 0
transform 1 0 3890 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1117_
timestamp 0
transform -1 0 4890 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1118_
timestamp 0
transform 1 0 4370 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1119_
timestamp 0
transform 1 0 4370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1120_
timestamp 0
transform 1 0 4530 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1121_
timestamp 0
transform -1 0 4430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1122_
timestamp 0
transform 1 0 4650 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1123_
timestamp 0
transform 1 0 4690 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1124_
timestamp 0
transform 1 0 3670 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1125_
timestamp 0
transform 1 0 3830 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1126_
timestamp 0
transform 1 0 3990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1127_
timestamp 0
transform -1 0 3850 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1128_
timestamp 0
transform -1 0 3710 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1129_
timestamp 0
transform 1 0 1810 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1130_
timestamp 0
transform 1 0 970 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1131_
timestamp 0
transform 1 0 1250 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1132_
timestamp 0
transform -1 0 3870 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1133_
timestamp 0
transform 1 0 2070 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1134_
timestamp 0
transform 1 0 2150 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1135_
timestamp 0
transform 1 0 1310 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1136_
timestamp 0
transform -1 0 1770 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1137_
timestamp 0
transform 1 0 1570 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1138_
timestamp 0
transform 1 0 1470 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1139_
timestamp 0
transform 1 0 2690 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1140_
timestamp 0
transform 1 0 1310 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1141_
timestamp 0
transform 1 0 1650 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1142_
timestamp 0
transform 1 0 1990 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1143_
timestamp 0
transform 1 0 2330 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1144_
timestamp 0
transform -1 0 3030 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1145_
timestamp 0
transform 1 0 2770 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1146_
timestamp 0
transform 1 0 3170 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1147_
timestamp 0
transform 1 0 2890 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1148_
timestamp 0
transform 1 0 2870 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1149_
timestamp 0
transform 1 0 2690 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1150_
timestamp 0
transform 1 0 3190 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1151_
timestamp 0
transform 1 0 3030 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1152_
timestamp 0
transform 1 0 2470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1153_
timestamp 0
transform -1 0 2870 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1154_
timestamp 0
transform 1 0 2850 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1155_
timestamp 0
transform 1 0 4690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1156_
timestamp 0
transform 1 0 4630 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1157_
timestamp 0
transform -1 0 5030 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1158_
timestamp 0
transform -1 0 5510 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1159_
timestamp 0
transform -1 0 4830 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1160_
timestamp 0
transform 1 0 4810 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1161_
timestamp 0
transform 1 0 2230 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1162_
timestamp 0
transform -1 0 4050 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1163_
timestamp 0
transform -1 0 4990 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1164_
timestamp 0
transform 1 0 4510 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1165_
timestamp 0
transform -1 0 4850 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1166_
timestamp 0
transform 1 0 4170 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1167_
timestamp 0
transform -1 0 4350 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1168_
timestamp 0
transform 1 0 4530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1169_
timestamp 0
transform -1 0 4850 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1170_
timestamp 0
transform 1 0 4170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1171_
timestamp 0
transform 1 0 4810 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1172_
timestamp 0
transform 1 0 5010 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1173_
timestamp 0
transform 1 0 830 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1174_
timestamp 0
transform 1 0 3670 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1175_
timestamp 0
transform 1 0 3270 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1176_
timestamp 0
transform 1 0 3330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1177_
timestamp 0
transform -1 0 3430 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1178_
timestamp 0
transform -1 0 3990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1179_
timestamp 0
transform 1 0 3530 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1180_
timestamp 0
transform 1 0 3270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1181_
timestamp 0
transform 1 0 3550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1182_
timestamp 0
transform 1 0 3710 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1183_
timestamp 0
transform 1 0 4130 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1184_
timestamp 0
transform 1 0 3890 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1185_
timestamp 0
transform 1 0 3510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1186_
timestamp 0
transform 1 0 3650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1187_
timestamp 0
transform 1 0 3810 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1188_
timestamp 0
transform 1 0 3710 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1189_
timestamp 0
transform -1 0 4070 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1190_
timestamp 0
transform 1 0 4330 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1191_
timestamp 0
transform -1 0 5170 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1192_
timestamp 0
transform 1 0 3970 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1193_
timestamp 0
transform 1 0 4210 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1194_
timestamp 0
transform -1 0 4490 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1195_
timestamp 0
transform -1 0 4010 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1196_
timestamp 0
transform -1 0 1930 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1197_
timestamp 0
transform 1 0 4290 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1198_
timestamp 0
transform -1 0 4190 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1199_
timestamp 0
transform -1 0 3670 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1200_
timestamp 0
transform 1 0 3470 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1201_
timestamp 0
transform 1 0 4310 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1202_
timestamp 0
transform 1 0 4490 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1203_
timestamp 0
transform 1 0 3810 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1204_
timestamp 0
transform -1 0 4670 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1205_
timestamp 0
transform 1 0 4010 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1206_
timestamp 0
transform 1 0 2510 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1207_
timestamp 0
transform -1 0 4170 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1208_
timestamp 0
transform -1 0 3330 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1209_
timestamp 0
transform -1 0 2990 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1210_
timestamp 0
transform -1 0 3170 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1211_
timestamp 0
transform 1 0 3250 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1212_
timestamp 0
transform 1 0 3330 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1213_
timestamp 0
transform 1 0 3510 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1214_
timestamp 0
transform -1 0 3390 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1215_
timestamp 0
transform -1 0 3050 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1216_
timestamp 0
transform -1 0 2650 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1217_
timestamp 0
transform 1 0 3510 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1218_
timestamp 0
transform 1 0 5070 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1219_
timestamp 0
transform -1 0 5150 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1220_
timestamp 0
transform -1 0 4790 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1221_
timestamp 0
transform 1 0 4590 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1222_
timestamp 0
transform 1 0 4510 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1223_
timestamp 0
transform 1 0 5010 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1224_
timestamp 0
transform -1 0 5130 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1225_
timestamp 0
transform 1 0 6110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1226_
timestamp 0
transform 1 0 5970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1227_
timestamp 0
transform -1 0 5350 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1228_
timestamp 0
transform 1 0 5630 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1229_
timestamp 0
transform -1 0 6330 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1230_
timestamp 0
transform 1 0 4970 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1231_
timestamp 0
transform 1 0 5110 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1232_
timestamp 0
transform 1 0 4850 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1233_
timestamp 0
transform -1 0 5170 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1234_
timestamp 0
transform 1 0 5630 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1235_
timestamp 0
transform -1 0 5490 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1236_
timestamp 0
transform -1 0 5470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1237_
timestamp 0
transform 1 0 4990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1238_
timestamp 0
transform 1 0 4530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1239_
timestamp 0
transform -1 0 4710 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1240_
timestamp 0
transform 1 0 5310 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1241_
timestamp 0
transform 1 0 5290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1242_
timestamp 0
transform 1 0 5770 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1243_
timestamp 0
transform -1 0 3410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1244_
timestamp 0
transform 1 0 5610 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1245_
timestamp 0
transform 1 0 4130 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1246_
timestamp 0
transform 1 0 4470 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1247_
timestamp 0
transform -1 0 5010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1248_
timestamp 0
transform 1 0 4290 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1249_
timestamp 0
transform 1 0 5110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1250_
timestamp 0
transform 1 0 5410 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1251_
timestamp 0
transform 1 0 5270 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1252_
timestamp 0
transform 1 0 5710 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1253_
timestamp 0
transform -1 0 5750 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1254_
timestamp 0
transform -1 0 5550 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1255_
timestamp 0
transform -1 0 4030 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1256_
timestamp 0
transform 1 0 4130 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1257_
timestamp 0
transform 1 0 3690 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1258_
timestamp 0
transform 1 0 4250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1259_
timestamp 0
transform -1 0 5290 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1260_
timestamp 0
transform 1 0 5970 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1261_
timestamp 0
transform 1 0 5930 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1262_
timestamp 0
transform 1 0 5870 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1263_
timestamp 0
transform 1 0 5430 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1264_
timestamp 0
transform 1 0 5610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1265_
timestamp 0
transform -1 0 5930 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1266_
timestamp 0
transform 1 0 3790 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1267_
timestamp 0
transform 1 0 4650 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1268_
timestamp 0
transform 1 0 5450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1269_
timestamp 0
transform -1 0 5810 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1270_
timestamp 0
transform -1 0 5610 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1271_
timestamp 0
transform 1 0 6230 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1272_
timestamp 0
transform -1 0 6530 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1273_
timestamp 0
transform 1 0 6070 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1274_
timestamp 0
transform 1 0 5750 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1275_
timestamp 0
transform -1 0 6610 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1276_
timestamp 0
transform -1 0 6190 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1277_
timestamp 0
transform 1 0 4430 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1278_
timestamp 0
transform 1 0 4890 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1279_
timestamp 0
transform -1 0 6570 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1280_
timestamp 0
transform -1 0 6090 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1281_
timestamp 0
transform -1 0 5850 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1282_
timestamp 0
transform -1 0 5570 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1283_
timestamp 0
transform 1 0 5450 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1284_
timestamp 0
transform -1 0 6350 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1285_
timestamp 0
transform -1 0 6030 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1286_
timestamp 0
transform -1 0 5930 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1287_
timestamp 0
transform 1 0 5210 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1288_
timestamp 0
transform -1 0 5590 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1289_
timestamp 0
transform -1 0 5410 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1290_
timestamp 0
transform -1 0 5290 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1291_
timestamp 0
transform -1 0 5290 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1292_
timestamp 0
transform 1 0 5430 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1293_
timestamp 0
transform 1 0 4290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1294_
timestamp 0
transform 1 0 4230 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1295_
timestamp 0
transform -1 0 4710 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1296_
timestamp 0
transform -1 0 4730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1297_
timestamp 0
transform 1 0 5710 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1298_
timestamp 0
transform -1 0 5750 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1299_
timestamp 0
transform 1 0 5930 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1300_
timestamp 0
transform 1 0 6390 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1301_
timestamp 0
transform -1 0 6530 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1302_
timestamp 0
transform -1 0 4390 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1303_
timestamp 0
transform 1 0 5470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1304_
timestamp 0
transform -1 0 4850 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1305_
timestamp 0
transform 1 0 5170 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1306_
timestamp 0
transform 1 0 5090 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1307_
timestamp 0
transform 1 0 5370 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1308_
timestamp 0
transform 1 0 5770 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1309_
timestamp 0
transform -1 0 4190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1310_
timestamp 0
transform 1 0 4770 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1311_
timestamp 0
transform -1 0 5330 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1312_
timestamp 0
transform 1 0 5430 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1313_
timestamp 0
transform -1 0 5130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1314_
timestamp 0
transform -1 0 5930 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1315_
timestamp 0
transform 1 0 5270 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1316_
timestamp 0
transform -1 0 5610 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1317_
timestamp 0
transform 1 0 5630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1318_
timestamp 0
transform 1 0 5750 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1319_
timestamp 0
transform 1 0 5790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1320_
timestamp 0
transform 1 0 5590 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1321_
timestamp 0
transform 1 0 6070 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1322_
timestamp 0
transform 1 0 6230 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1323_
timestamp 0
transform 1 0 6230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1324_
timestamp 0
transform -1 0 6470 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1325_
timestamp 0
transform 1 0 6270 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1326_
timestamp 0
transform 1 0 4950 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1327_
timestamp 0
transform 1 0 4430 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1328_
timestamp 0
transform 1 0 4150 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1329_
timestamp 0
transform -1 0 4350 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1330_
timestamp 0
transform 1 0 4470 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1331_
timestamp 0
transform 1 0 4610 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1332_
timestamp 0
transform 1 0 5090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1333_
timestamp 0
transform 1 0 4450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1334_
timestamp 0
transform 1 0 4930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1335_
timestamp 0
transform 1 0 3990 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1336_
timestamp 0
transform 1 0 5370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1337_
timestamp 0
transform 1 0 5530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1338_
timestamp 0
transform 1 0 4950 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1339_
timestamp 0
transform -1 0 6030 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1340_
timestamp 0
transform -1 0 4670 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1341_
timestamp 0
transform 1 0 3430 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1342_
timestamp 0
transform 1 0 3550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1343_
timestamp 0
transform -1 0 3870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1344_
timestamp 0
transform -1 0 4270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1345_
timestamp 0
transform 1 0 4570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1346_
timestamp 0
transform 1 0 5270 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1347_
timestamp 0
transform 1 0 4330 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1348_
timestamp 0
transform 1 0 3710 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1349_
timestamp 0
transform 1 0 5410 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1350_
timestamp 0
transform -1 0 6050 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1351_
timestamp 0
transform 1 0 5590 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1352_
timestamp 0
transform 1 0 4390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1353_
timestamp 0
transform 1 0 5530 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1354_
timestamp 0
transform 1 0 6050 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1355_
timestamp 0
transform 1 0 5690 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1356_
timestamp 0
transform 1 0 6190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1357_
timestamp 0
transform 1 0 5690 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1358_
timestamp 0
transform 1 0 6510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1359_
timestamp 0
transform -1 0 6290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1360_
timestamp 0
transform 1 0 6030 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1361_
timestamp 0
transform 1 0 6090 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1362_
timestamp 0
transform -1 0 6370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1363_
timestamp 0
transform 1 0 5890 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1364_
timestamp 0
transform 1 0 5930 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1365_
timestamp 0
transform -1 0 6430 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1366_
timestamp 0
transform 1 0 6530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1367_
timestamp 0
transform 1 0 6210 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1368_
timestamp 0
transform 1 0 6110 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1369_
timestamp 0
transform 1 0 6570 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1370_
timestamp 0
transform -1 0 6270 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1371_
timestamp 0
transform 1 0 6150 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1372_
timestamp 0
transform 1 0 6230 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1373_
timestamp 0
transform 1 0 6610 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1374_
timestamp 0
transform -1 0 6390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1375_
timestamp 0
transform -1 0 6210 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1376_
timestamp 0
transform -1 0 5910 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1377_
timestamp 0
transform 1 0 6550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1378_
timestamp 0
transform -1 0 6450 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1379_
timestamp 0
transform -1 0 6370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1380_
timestamp 0
transform -1 0 6250 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1381_
timestamp 0
transform -1 0 5790 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1382_
timestamp 0
transform -1 0 6530 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1383_
timestamp 0
transform -1 0 6410 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1384_
timestamp 0
transform -1 0 6410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1385_
timestamp 0
transform -1 0 6090 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1386_
timestamp 0
transform -1 0 6090 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1387_
timestamp 0
transform 1 0 5310 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1388_
timestamp 0
transform 1 0 4730 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1389_
timestamp 0
transform -1 0 4610 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1390_
timestamp 0
transform -1 0 5050 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1391_
timestamp 0
transform 1 0 4410 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1392_
timestamp 0
transform 1 0 4050 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1393_
timestamp 0
transform 1 0 3890 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1394_
timestamp 0
transform -1 0 5150 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1395_
timestamp 0
transform -1 0 5170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1396_
timestamp 0
transform -1 0 4990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1397_
timestamp 0
transform -1 0 6610 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1398_
timestamp 0
transform 1 0 6630 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1399_
timestamp 0
transform -1 0 6590 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1400_
timestamp 0
transform -1 0 6510 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1401_
timestamp 0
transform -1 0 6450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1402_
timestamp 0
transform -1 0 6570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1403_
timestamp 0
transform -1 0 5730 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1404_
timestamp 0
transform -1 0 4110 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1405_
timestamp 0
transform 1 0 4930 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1406_
timestamp 0
transform -1 0 4770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1407_
timestamp 0
transform 1 0 4370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1408_
timestamp 0
transform -1 0 4750 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1409_
timestamp 0
transform -1 0 4690 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1410_
timestamp 0
transform -1 0 4830 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1411_
timestamp 0
transform -1 0 4890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1412_
timestamp 0
transform 1 0 4410 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1413_
timestamp 0
transform -1 0 4810 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1414_
timestamp 0
transform 1 0 4770 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1415_
timestamp 0
transform 1 0 4570 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1416_
timestamp 0
transform 1 0 5210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1417_
timestamp 0
transform 1 0 5230 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1418_
timestamp 0
transform 1 0 4590 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1419_
timestamp 0
transform 1 0 5030 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1420_
timestamp 0
transform 1 0 4290 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1421_
timestamp 0
transform 1 0 4230 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1422_
timestamp 0
transform 1 0 5390 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1423_
timestamp 0
transform 1 0 5710 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1424_
timestamp 0
transform 1 0 5230 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1425_
timestamp 0
transform 1 0 5550 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1426_
timestamp 0
transform 1 0 5550 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1427_
timestamp 0
transform 1 0 5050 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1428_
timestamp 0
transform -1 0 5890 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1429_
timestamp 0
transform 1 0 5750 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1430_
timestamp 0
transform 1 0 6190 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1431_
timestamp 0
transform -1 0 6350 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1432_
timestamp 0
transform 1 0 4890 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1433_
timestamp 0
transform -1 0 4310 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1434_
timestamp 0
transform 1 0 4710 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1435_
timestamp 0
transform -1 0 4630 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1436_
timestamp 0
transform 1 0 4750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1437_
timestamp 0
transform 1 0 5050 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1438_
timestamp 0
transform 1 0 5210 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1439_
timestamp 0
transform 1 0 3130 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1440_
timestamp 0
transform -1 0 4950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1441_
timestamp 0
transform 1 0 4130 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1442_
timestamp 0
transform 1 0 5370 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1443_
timestamp 0
transform 1 0 5550 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1444_
timestamp 0
transform 1 0 3690 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1445_
timestamp 0
transform 1 0 3170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1446_
timestamp 0
transform -1 0 3970 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1447_
timestamp 0
transform -1 0 4550 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1448_
timestamp 0
transform 1 0 4970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1449_
timestamp 0
transform 1 0 4490 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1450_
timestamp 0
transform 1 0 4970 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1451_
timestamp 0
transform 1 0 4670 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1452_
timestamp 0
transform 1 0 5330 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1453_
timestamp 0
transform -1 0 5710 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1454_
timestamp 0
transform 1 0 4170 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1455_
timestamp 0
transform 1 0 4030 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1456_
timestamp 0
transform -1 0 5390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1457_
timestamp 0
transform 1 0 5490 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1458_
timestamp 0
transform 1 0 5530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1459_
timestamp 0
transform 1 0 5630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1460_
timestamp 0
transform 1 0 5870 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1461_
timestamp 0
transform 1 0 6030 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1462_
timestamp 0
transform -1 0 5090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1463_
timestamp 0
transform 1 0 5310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1464_
timestamp 0
transform 1 0 5870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1465_
timestamp 0
transform 1 0 5150 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1466_
timestamp 0
transform 1 0 5770 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1467_
timestamp 0
transform 1 0 5890 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1468_
timestamp 0
transform -1 0 6070 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1469_
timestamp 0
transform 1 0 5470 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1470_
timestamp 0
transform 1 0 5930 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1471_
timestamp 0
transform -1 0 5990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1472_
timestamp 0
transform 1 0 6130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1473_
timestamp 0
transform 1 0 6390 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1474_
timestamp 0
transform -1 0 6570 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1475_
timestamp 0
transform 1 0 6150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1476_
timestamp 0
transform 1 0 5810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1477_
timestamp 0
transform 1 0 6390 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1478_
timestamp 0
transform -1 0 6490 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1479_
timestamp 0
transform 1 0 6230 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1480_
timestamp 0
transform -1 0 6330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1481_
timestamp 0
transform 1 0 6570 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1482_
timestamp 0
transform 1 0 6630 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1483_
timestamp 0
transform -1 0 6650 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1484_
timestamp 0
transform 1 0 6530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1485_
timestamp 0
transform -1 0 6670 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1486_
timestamp 0
transform -1 0 6310 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1487_
timestamp 0
transform -1 0 6510 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1488_
timestamp 0
transform -1 0 4850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1489_
timestamp 0
transform 1 0 3990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1490_
timestamp 0
transform 1 0 4030 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1491_
timestamp 0
transform -1 0 5050 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1492_
timestamp 0
transform 1 0 4850 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1493_
timestamp 0
transform 1 0 6390 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1494_
timestamp 0
transform 1 0 6510 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1495_
timestamp 0
transform -1 0 5870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1496_
timestamp 0
transform 1 0 6290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1497_
timestamp 0
transform -1 0 6110 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1498_
timestamp 0
transform 1 0 6210 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1499_
timestamp 0
transform 1 0 5190 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1500_
timestamp 0
transform -1 0 4590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1501_
timestamp 0
transform 1 0 4090 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1502_
timestamp 0
transform 1 0 4830 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1503_
timestamp 0
transform -1 0 4730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1504_
timestamp 0
transform 1 0 5130 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1505_
timestamp 0
transform 1 0 4850 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1506_
timestamp 0
transform -1 0 4530 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1507_
timestamp 0
transform 1 0 4530 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1508_
timestamp 0
transform -1 0 5030 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1509_
timestamp 0
transform 1 0 5150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1510_
timestamp 0
transform 1 0 4870 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1511_
timestamp 0
transform 1 0 5210 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1512_
timestamp 0
transform -1 0 5350 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1513_
timestamp 0
transform 1 0 4970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1514_
timestamp 0
transform 1 0 4970 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1515_
timestamp 0
transform 1 0 5030 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1516_
timestamp 0
transform 1 0 5550 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1517_
timestamp 0
transform 1 0 5490 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1518_
timestamp 0
transform 1 0 5130 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1519_
timestamp 0
transform 1 0 5350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1520_
timestamp 0
transform 1 0 5310 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1521_
timestamp 0
transform 1 0 5390 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1522_
timestamp 0
transform 1 0 5470 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1523_
timestamp 0
transform 1 0 5630 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1524_
timestamp 0
transform -1 0 5170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1525_
timestamp 0
transform -1 0 5870 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1526_
timestamp 0
transform 1 0 3650 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1527_
timestamp 0
transform 1 0 3150 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1528_
timestamp 0
transform -1 0 3970 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1529_
timestamp 0
transform 1 0 3490 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1530_
timestamp 0
transform 1 0 3790 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1531_
timestamp 0
transform 1 0 4570 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1532_
timestamp 0
transform -1 0 3610 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1533_
timestamp 0
transform -1 0 3870 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1534_
timestamp 0
transform -1 0 4410 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1535_
timestamp 0
transform -1 0 4450 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1536_
timestamp 0
transform 1 0 4070 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1537_
timestamp 0
transform 1 0 4250 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1538_
timestamp 0
transform 1 0 4390 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1539_
timestamp 0
transform 1 0 4270 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1540_
timestamp 0
transform 1 0 5650 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1541_
timestamp 0
transform -1 0 5830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1542_
timestamp 0
transform -1 0 5250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1543_
timestamp 0
transform 1 0 5690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1544_
timestamp 0
transform -1 0 5750 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1545_
timestamp 0
transform -1 0 5670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1546_
timestamp 0
transform 1 0 6090 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1547_
timestamp 0
transform 1 0 5890 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1548_
timestamp 0
transform -1 0 5970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1549_
timestamp 0
transform 1 0 6270 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1550_
timestamp 0
transform -1 0 6290 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1551_
timestamp 0
transform 1 0 5610 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1552_
timestamp 0
transform 1 0 6030 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1553_
timestamp 0
transform 1 0 6090 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1554_
timestamp 0
transform 1 0 5810 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1555_
timestamp 0
transform -1 0 6050 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1556_
timestamp 0
transform 1 0 5970 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1557_
timestamp 0
transform -1 0 6150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1558_
timestamp 0
transform 1 0 6390 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1559_
timestamp 0
transform 1 0 6590 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1560_
timestamp 0
transform 1 0 6050 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1561_
timestamp 0
transform -1 0 6590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1562_
timestamp 0
transform -1 0 6590 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1563_
timestamp 0
transform -1 0 6430 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1564_
timestamp 0
transform 1 0 6210 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1565_
timestamp 0
transform 1 0 6370 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1566_
timestamp 0
transform -1 0 6570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1567_
timestamp 0
transform -1 0 4470 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1568_
timestamp 0
transform 1 0 4190 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1569_
timestamp 0
transform -1 0 4230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1570_
timestamp 0
transform -1 0 3750 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1571_
timestamp 0
transform 1 0 6210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1572_
timestamp 0
transform -1 0 4330 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1573_
timestamp 0
transform -1 0 3690 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1574_
timestamp 0
transform 1 0 6430 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1575_
timestamp 0
transform 1 0 6450 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1576_
timestamp 0
transform 1 0 5470 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1577_
timestamp 0
transform -1 0 5490 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1578_
timestamp 0
transform -1 0 5950 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1579_
timestamp 0
transform -1 0 4690 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1580_
timestamp 0
transform 1 0 4390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1581_
timestamp 0
transform -1 0 3030 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1582_
timestamp 0
transform -1 0 2830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1583_
timestamp 0
transform -1 0 2890 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1584_
timestamp 0
transform -1 0 3030 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1585_
timestamp 0
transform 1 0 3170 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1586_
timestamp 0
transform 1 0 2690 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1587_
timestamp 0
transform 1 0 2810 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1588_
timestamp 0
transform -1 0 1990 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1589_
timestamp 0
transform -1 0 2690 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1590_
timestamp 0
transform 1 0 2930 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1591_
timestamp 0
transform 1 0 3890 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1592_
timestamp 0
transform -1 0 3750 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1593_
timestamp 0
transform -1 0 3770 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1594_
timestamp 0
transform 1 0 3090 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1595_
timestamp 0
transform 1 0 3010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1596_
timestamp 0
transform -1 0 4070 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1597_
timestamp 0
transform -1 0 4230 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1598_
timestamp 0
transform 1 0 4070 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1599_
timestamp 0
transform -1 0 4250 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1600_
timestamp 0
transform 1 0 3570 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1601_
timestamp 0
transform 1 0 3910 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1602_
timestamp 0
transform -1 0 3910 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1603_
timestamp 0
transform 1 0 4810 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1604_
timestamp 0
transform 1 0 3670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1605_
timestamp 0
transform 1 0 3510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1606_
timestamp 0
transform 1 0 1390 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1607_
timestamp 0
transform -1 0 3370 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1608_
timestamp 0
transform -1 0 2730 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1609_
timestamp 0
transform 1 0 3150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1610_
timestamp 0
transform -1 0 2410 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1611_
timestamp 0
transform -1 0 2570 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1612_
timestamp 0
transform 1 0 1530 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1613_
timestamp 0
transform 1 0 3290 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1614_
timestamp 0
transform 1 0 3430 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1615_
timestamp 0
transform 1 0 3790 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1616_
timestamp 0
transform 1 0 3150 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1617_
timestamp 0
transform -1 0 3610 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1618_
timestamp 0
transform 1 0 4230 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1619_
timestamp 0
transform -1 0 4690 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1620_
timestamp 0
transform 1 0 3770 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1621_
timestamp 0
transform 1 0 3450 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1622_
timestamp 0
transform 1 0 3950 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1623_
timestamp 0
transform 1 0 4970 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1624_
timestamp 0
transform 1 0 5930 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1625_
timestamp 0
transform 1 0 5770 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1626_
timestamp 0
transform 1 0 4210 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1627_
timestamp 0
transform -1 0 4550 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1628_
timestamp 0
transform 1 0 4850 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1629_
timestamp 0
transform 1 0 6250 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1630_
timestamp 0
transform -1 0 5790 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1631_
timestamp 0
transform 1 0 4690 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1632_
timestamp 0
transform 1 0 5590 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1633_
timestamp 0
transform 1 0 6430 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1634_
timestamp 0
transform 1 0 6210 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1635_
timestamp 0
transform -1 0 6470 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1636_
timestamp 0
transform 1 0 5130 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1637_
timestamp 0
transform -1 0 6110 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1638_
timestamp 0
transform 1 0 5290 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1639_
timestamp 0
transform 1 0 4690 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1640_
timestamp 0
transform 1 0 3530 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1641_
timestamp 0
transform 1 0 3350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1642_
timestamp 0
transform 1 0 3570 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1643_
timestamp 0
transform 1 0 2230 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1644_
timestamp 0
transform -1 0 3190 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1645_
timestamp 0
transform -1 0 5330 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1646_
timestamp 0
transform -1 0 5170 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1647_
timestamp 0
transform 1 0 3730 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1648_
timestamp 0
transform -1 0 3790 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1649_
timestamp 0
transform -1 0 4070 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1650_
timestamp 0
transform -1 0 3450 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1651_
timestamp 0
transform -1 0 3590 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1652_
timestamp 0
transform -1 0 2550 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1653_
timestamp 0
transform 1 0 2510 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1654_
timestamp 0
transform -1 0 2410 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1655_
timestamp 0
transform -1 0 2210 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1656_
timestamp 0
transform 1 0 1690 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1657_
timestamp 0
transform -1 0 2090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1658_
timestamp 0
transform 1 0 1830 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1659_
timestamp 0
transform -1 0 2050 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1660_
timestamp 0
transform -1 0 2270 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1661_
timestamp 0
transform 1 0 2110 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1662_
timestamp 0
transform 1 0 2210 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1663_
timestamp 0
transform -1 0 1950 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1664_
timestamp 0
transform -1 0 1650 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1665_
timestamp 0
transform -1 0 1470 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1666_
timestamp 0
transform -1 0 1890 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1667_
timestamp 0
transform 1 0 1470 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1668_
timestamp 0
transform 1 0 2010 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1669_
timestamp 0
transform 1 0 2350 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1670_
timestamp 0
transform 1 0 1310 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1671_
timestamp 0
transform -1 0 1770 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1672_
timestamp 0
transform 1 0 1850 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1673_
timestamp 0
transform -1 0 70 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1674_
timestamp 0
transform -1 0 70 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1675_
timestamp 0
transform 1 0 50 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1676_
timestamp 0
transform 1 0 210 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1677_
timestamp 0
transform 1 0 350 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1678_
timestamp 0
transform 1 0 2190 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1679_
timestamp 0
transform -1 0 1710 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1680_
timestamp 0
transform -1 0 1530 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1681_
timestamp 0
transform 1 0 1230 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1682_
timestamp 0
transform -1 0 1370 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1683_
timestamp 0
transform 1 0 2610 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1684_
timestamp 0
transform -1 0 2490 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1685_
timestamp 0
transform -1 0 3290 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1686_
timestamp 0
transform 1 0 3890 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1687_
timestamp 0
transform -1 0 4390 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1688_
timestamp 0
transform 1 0 2790 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1689_
timestamp 0
transform -1 0 2970 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1690_
timestamp 0
transform -1 0 3130 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1691_
timestamp 0
transform -1 0 4090 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1692_
timestamp 0
transform -1 0 4570 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1693_
timestamp 0
transform -1 0 4410 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1694_
timestamp 0
transform 1 0 3270 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1695_
timestamp 0
transform -1 0 3610 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1696_
timestamp 0
transform 1 0 3430 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1697_
timestamp 0
transform -1 0 3470 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1698_
timestamp 0
transform -1 0 2870 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1699_
timestamp 0
transform 1 0 3030 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1700_
timestamp 0
transform -1 0 2890 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1701_
timestamp 0
transform 1 0 2590 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1702_
timestamp 0
transform 1 0 3030 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1703_
timestamp 0
transform 1 0 3350 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1704_
timestamp 0
transform -1 0 3510 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1705_
timestamp 0
transform -1 0 3330 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1706_
timestamp 0
transform 1 0 3310 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1707_
timestamp 0
transform -1 0 3010 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1708_
timestamp 0
transform -1 0 2390 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1709_
timestamp 0
transform 1 0 1090 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1710_
timestamp 0
transform 1 0 50 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1711_
timestamp 0
transform 1 0 1710 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1712_
timestamp 0
transform 1 0 2350 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1713_
timestamp 0
transform -1 0 2190 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1714_
timestamp 0
transform -1 0 2250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1715_
timestamp 0
transform 1 0 2030 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1716_
timestamp 0
transform 1 0 1910 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1717_
timestamp 0
transform 1 0 1690 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1718_
timestamp 0
transform 1 0 1770 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1719_
timestamp 0
transform -1 0 1150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1720_
timestamp 0
transform -1 0 1310 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1721_
timestamp 0
transform -1 0 750 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1722_
timestamp 0
transform 1 0 210 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1723_
timestamp 0
transform 1 0 270 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1724_
timestamp 0
transform 1 0 230 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1725_
timestamp 0
transform -1 0 70 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1726_
timestamp 0
transform 1 0 370 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1727_
timestamp 0
transform -1 0 530 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1728_
timestamp 0
transform -1 0 970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1729_
timestamp 0
transform 1 0 670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1730_
timestamp 0
transform -1 0 810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1731_
timestamp 0
transform 1 0 230 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1732_
timestamp 0
transform 1 0 410 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1733_
timestamp 0
transform 1 0 510 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1734_
timestamp 0
transform 1 0 670 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1735_
timestamp 0
transform -1 0 990 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1736_
timestamp 0
transform -1 0 570 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1737_
timestamp 0
transform 1 0 670 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1738_
timestamp 0
transform 1 0 810 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1739_
timestamp 0
transform 1 0 1150 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1740_
timestamp 0
transform -1 0 2250 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1741_
timestamp 0
transform -1 0 1030 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1742_
timestamp 0
transform -1 0 2110 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1743_
timestamp 0
transform 1 0 2830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1744_
timestamp 0
transform -1 0 2950 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1745_
timestamp 0
transform 1 0 2690 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1746_
timestamp 0
transform -1 0 2550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1747_
timestamp 0
transform -1 0 2790 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1748_
timestamp 0
transform 1 0 850 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1749_
timestamp 0
transform -1 0 1850 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1750_
timestamp 0
transform -1 0 2110 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1751_
timestamp 0
transform -1 0 1950 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1752_
timestamp 0
transform 1 0 1830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1753_
timestamp 0
transform -1 0 1650 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1754_
timestamp 0
transform 1 0 1770 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1755_
timestamp 0
transform -1 0 1350 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1756_
timestamp 0
transform -1 0 510 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1757_
timestamp 0
transform 1 0 410 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1758_
timestamp 0
transform -1 0 430 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1759_
timestamp 0
transform 1 0 570 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1760_
timestamp 0
transform 1 0 550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1761_
timestamp 0
transform -1 0 1030 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1762_
timestamp 0
transform 1 0 850 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1763_
timestamp 0
transform -1 0 910 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1764_
timestamp 0
transform 1 0 1970 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1765_
timestamp 0
transform -1 0 2670 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1766_
timestamp 0
transform 1 0 2490 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1767_
timestamp 0
transform 1 0 2530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1768_
timestamp 0
transform -1 0 2390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1769_
timestamp 0
transform -1 0 2410 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1770_
timestamp 0
transform 1 0 2230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1771_
timestamp 0
transform 1 0 2670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1772_
timestamp 0
transform -1 0 2850 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1773_
timestamp 0
transform 1 0 2370 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1774_
timestamp 0
transform 1 0 1610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1775_
timestamp 0
transform 1 0 1550 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1776_
timestamp 0
transform 1 0 710 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1777_
timestamp 0
transform -1 0 1210 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1778_
timestamp 0
transform -1 0 1670 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1779_
timestamp 0
transform -1 0 1470 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1780_
timestamp 0
transform 1 0 350 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1781_
timestamp 0
transform 1 0 690 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1782_
timestamp 0
transform 1 0 310 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1783_
timestamp 0
transform 1 0 450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1784_
timestamp 0
transform -1 0 610 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1785_
timestamp 0
transform -1 0 770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1786_
timestamp 0
transform 1 0 1070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1787_
timestamp 0
transform 1 0 910 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1788_
timestamp 0
transform 1 0 1390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1789_
timestamp 0
transform 1 0 1710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1790_
timestamp 0
transform -1 0 2230 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1791_
timestamp 0
transform -1 0 1570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1792_
timestamp 0
transform 1 0 1230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1793_
timestamp 0
transform -1 0 890 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1794_
timestamp 0
transform 1 0 1470 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1795_
timestamp 0
transform -1 0 850 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1796_
timestamp 0
transform 1 0 610 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1797_
timestamp 0
transform 1 0 1030 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1798_
timestamp 0
transform 1 0 1150 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1799_
timestamp 0
transform 1 0 1290 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1800_
timestamp 0
transform -1 0 1850 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1801_
timestamp 0
transform 1 0 1650 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1802_
timestamp 0
transform 1 0 50 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1803_
timestamp 0
transform 1 0 950 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1804_
timestamp 0
transform -1 0 1090 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1805_
timestamp 0
transform 1 0 170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1806_
timestamp 0
transform 1 0 290 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1807_
timestamp 0
transform 1 0 190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1808_
timestamp 0
transform 1 0 450 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1809_
timestamp 0
transform 1 0 290 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1810_
timestamp 0
transform 1 0 50 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1811_
timestamp 0
transform -1 0 1070 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1812_
timestamp 0
transform 1 0 890 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1813_
timestamp 0
transform 1 0 190 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1814_
timestamp 0
transform 1 0 850 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1815_
timestamp 0
transform 1 0 450 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1816_
timestamp 0
transform 1 0 970 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1817_
timestamp 0
transform -1 0 750 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1818_
timestamp 0
transform 1 0 330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1819_
timestamp 0
transform -1 0 1070 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1820_
timestamp 0
transform -1 0 1210 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1821_
timestamp 0
transform 1 0 50 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1822_
timestamp 0
transform -1 0 1050 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1823_
timestamp 0
transform 1 0 50 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1824_
timestamp 0
transform 1 0 50 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1825_
timestamp 0
transform -1 0 1130 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1826_
timestamp 0
transform -1 0 950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1827_
timestamp 0
transform 1 0 530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1828_
timestamp 0
transform 1 0 1770 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1829_
timestamp 0
transform 1 0 1590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1830_
timestamp 0
transform -1 0 1450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1831_
timestamp 0
transform 1 0 950 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1832_
timestamp 0
transform -1 0 790 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1833_
timestamp 0
transform 1 0 610 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1834_
timestamp 0
transform -1 0 70 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1835_
timestamp 0
transform -1 0 510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1836_
timestamp 0
transform 1 0 890 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1837_
timestamp 0
transform -1 0 750 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1838_
timestamp 0
transform 1 0 430 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1839_
timestamp 0
transform -1 0 350 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1840_
timestamp 0
transform -1 0 70 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1841_
timestamp 0
transform -1 0 210 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1842_
timestamp 0
transform -1 0 1210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1843_
timestamp 0
transform -1 0 1350 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1844_
timestamp 0
transform 1 0 1850 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1845_
timestamp 0
transform 1 0 2010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1846_
timestamp 0
transform -1 0 2970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1847_
timestamp 0
transform -1 0 3110 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1848_
timestamp 0
transform -1 0 370 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1849_
timestamp 0
transform 1 0 190 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1911_
timestamp 0
transform -1 0 2710 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1912_
timestamp 0
transform -1 0 70 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1913_
timestamp 0
transform 1 0 2410 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1914_
timestamp 0
transform -1 0 70 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1915_
timestamp 0
transform -1 0 70 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1916_
timestamp 0
transform -1 0 2570 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1917_
timestamp 0
transform -1 0 2490 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1918_
timestamp 0
transform -1 0 230 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1919_
timestamp 0
transform -1 0 70 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert0
timestamp 0
transform 1 0 3130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert1
timestamp 0
transform 1 0 2830 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert2
timestamp 0
transform 1 0 3270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert3
timestamp 0
transform 1 0 3270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert4
timestamp 0
transform -1 0 2710 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert12
timestamp 0
transform 1 0 3550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert13
timestamp 0
transform 1 0 50 0 1 1310
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert14
timestamp 0
transform 1 0 590 0 1 1830
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert15
timestamp 0
transform 1 0 3590 0 1 2350
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert16
timestamp 0
transform 1 0 810 0 1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert17
timestamp 0
transform 1 0 1110 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert18
timestamp 0
transform -1 0 210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert19
timestamp 0
transform -1 0 1090 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert20
timestamp 0
transform -1 0 370 0 1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert21
timestamp 0
transform 1 0 3410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert22
timestamp 0
transform -1 0 3150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert23
timestamp 0
transform 1 0 3410 0 1 3910
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert24
timestamp 0
transform -1 0 3150 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert25
timestamp 0
transform -1 0 3270 0 1 3910
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert5
timestamp 0
transform -1 0 1030 0 1 3910
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert6
timestamp 0
transform 1 0 2070 0 1 3390
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert7
timestamp 0
transform 1 0 1030 0 1 2350
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert8
timestamp 0
transform -1 0 230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert9
timestamp 0
transform 1 0 190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert10
timestamp 0
transform 1 0 2690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert11
timestamp 0
transform 1 0 1690 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__922_
timestamp 0
transform -1 0 970 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__923_
timestamp 0
transform 1 0 1230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__924_
timestamp 0
transform -1 0 2690 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__925_
timestamp 0
transform 1 0 2510 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__926_
timestamp 0
transform -1 0 2570 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__927_
timestamp 0
transform -1 0 1130 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__928_
timestamp 0
transform -1 0 1970 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__929_
timestamp 0
transform 1 0 2970 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__930_
timestamp 0
transform 1 0 2570 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__931_
timestamp 0
transform -1 0 3650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__932_
timestamp 0
transform 1 0 3010 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__933_
timestamp 0
transform 1 0 2850 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__934_
timestamp 0
transform 1 0 2890 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__935_
timestamp 0
transform 1 0 2730 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__936_
timestamp 0
transform -1 0 3510 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__937_
timestamp 0
transform 1 0 2350 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__938_
timestamp 0
transform 1 0 2150 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__939_
timestamp 0
transform 1 0 2390 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__940_
timestamp 0
transform 1 0 2030 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__941_
timestamp 0
transform 1 0 1450 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__942_
timestamp 0
transform -1 0 1690 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__943_
timestamp 0
transform 1 0 1490 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__944_
timestamp 0
transform -1 0 2230 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__945_
timestamp 0
transform 1 0 1510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__946_
timestamp 0
transform -1 0 4490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__947_
timestamp 0
transform -1 0 970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__948_
timestamp 0
transform 1 0 630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__949_
timestamp 0
transform 1 0 3750 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__950_
timestamp 0
transform 1 0 2190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__951_
timestamp 0
transform -1 0 2350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__952_
timestamp 0
transform 1 0 3870 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__953_
timestamp 0
transform 1 0 530 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__954_
timestamp 0
transform -1 0 690 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__955_
timestamp 0
transform 1 0 2710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__956_
timestamp 0
transform -1 0 350 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__957_
timestamp 0
transform -1 0 490 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__958_
timestamp 0
transform 1 0 1090 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__959_
timestamp 0
transform -1 0 1730 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__960_
timestamp 0
transform 1 0 2650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__961_
timestamp 0
transform -1 0 2810 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__962_
timestamp 0
transform -1 0 2990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__963_
timestamp 0
transform -1 0 3010 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__964_
timestamp 0
transform 1 0 1290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__965_
timestamp 0
transform -1 0 1370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__966_
timestamp 0
transform -1 0 3030 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__967_
timestamp 0
transform 1 0 2690 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__968_
timestamp 0
transform -1 0 2870 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__969_
timestamp 0
transform -1 0 3430 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__970_
timestamp 0
transform -1 0 3110 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__971_
timestamp 0
transform -1 0 3270 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__972_
timestamp 0
transform -1 0 3070 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__973_
timestamp 0
transform -1 0 2510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__974_
timestamp 0
transform -1 0 2910 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__975_
timestamp 0
transform -1 0 2610 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__976_
timestamp 0
transform 1 0 2230 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__977_
timestamp 0
transform -1 0 2410 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__978_
timestamp 0
transform -1 0 3750 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__979_
timestamp 0
transform 1 0 3290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__980_
timestamp 0
transform -1 0 3590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__981_
timestamp 0
transform -1 0 3350 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__982_
timestamp 0
transform -1 0 2910 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__983_
timestamp 0
transform -1 0 3190 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__984_
timestamp 0
transform -1 0 3470 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__985_
timestamp 0
transform 1 0 4130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__986_
timestamp 0
transform 1 0 4090 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__987_
timestamp 0
transform -1 0 4250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__988_
timestamp 0
transform 1 0 3690 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__989_
timestamp 0
transform 1 0 2550 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__990_
timestamp 0
transform -1 0 2710 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__991_
timestamp 0
transform 1 0 2810 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__992_
timestamp 0
transform 1 0 2790 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__993_
timestamp 0
transform 1 0 3970 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__994_
timestamp 0
transform -1 0 4030 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__995_
timestamp 0
transform 1 0 3350 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__996_
timestamp 0
transform 1 0 3190 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__997_
timestamp 0
transform 1 0 1730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__998_
timestamp 0
transform 1 0 1570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__999_
timestamp 0
transform 1 0 2290 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1000_
timestamp 0
transform -1 0 3130 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1001_
timestamp 0
transform 1 0 2410 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1002_
timestamp 0
transform -1 0 2610 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1003_
timestamp 0
transform 1 0 2950 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1004_
timestamp 0
transform 1 0 2790 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1005_
timestamp 0
transform -1 0 1990 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1006_
timestamp 0
transform 1 0 1890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1007_
timestamp 0
transform 1 0 1810 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1008_
timestamp 0
transform 1 0 1550 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1009_
timestamp 0
transform 1 0 1130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1010_
timestamp 0
transform -1 0 1310 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1011_
timestamp 0
transform 1 0 1050 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1012_
timestamp 0
transform 1 0 2350 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1013_
timestamp 0
transform -1 0 3470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1014_
timestamp 0
transform 1 0 930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1015_
timestamp 0
transform -1 0 1830 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1016_
timestamp 0
transform 1 0 1990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1017_
timestamp 0
transform 1 0 2550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1018_
timestamp 0
transform 1 0 2130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1019_
timestamp 0
transform -1 0 790 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1020_
timestamp 0
transform 1 0 930 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1021_
timestamp 0
transform 1 0 1230 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1022_
timestamp 0
transform -1 0 1490 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1023_
timestamp 0
transform 1 0 1370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1024_
timestamp 0
transform 1 0 1250 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1025_
timestamp 0
transform -1 0 1550 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1026_
timestamp 0
transform 1 0 1390 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1027_
timestamp 0
transform 1 0 1550 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1028_
timestamp 0
transform -1 0 1530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1029_
timestamp 0
transform -1 0 1690 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1030_
timestamp 0
transform -1 0 1570 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1031_
timestamp 0
transform 1 0 1890 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1032_
timestamp 0
transform 1 0 1730 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1033_
timestamp 0
transform 1 0 2330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1034_
timestamp 0
transform 1 0 1650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1035_
timestamp 0
transform 1 0 3890 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1036_
timestamp 0
transform -1 0 1310 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1037_
timestamp 0
transform 1 0 1130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1038_
timestamp 0
transform -1 0 4630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1039_
timestamp 0
transform -1 0 1610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1040_
timestamp 0
transform 1 0 690 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1041_
timestamp 0
transform 1 0 530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1042_
timestamp 0
transform 1 0 810 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1043_
timestamp 0
transform -1 0 710 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1044_
timestamp 0
transform -1 0 1450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1045_
timestamp 0
transform 1 0 1130 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1046_
timestamp 0
transform 1 0 1010 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1047_
timestamp 0
transform 1 0 830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1048_
timestamp 0
transform 1 0 1250 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1049_
timestamp 0
transform -1 0 1010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1050_
timestamp 0
transform 1 0 1110 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1051_
timestamp 0
transform 1 0 1430 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1052_
timestamp 0
transform -1 0 1750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1053_
timestamp 0
transform -1 0 1970 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1054_
timestamp 0
transform 1 0 2350 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1055_
timestamp 0
transform -1 0 1970 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1056_
timestamp 0
transform -1 0 1630 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1057_
timestamp 0
transform -1 0 1790 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1058_
timestamp 0
transform 1 0 1610 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1059_
timestamp 0
transform -1 0 1790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1060_
timestamp 0
transform 1 0 1910 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1061_
timestamp 0
transform -1 0 2290 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1062_
timestamp 0
transform 1 0 1270 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1063_
timestamp 0
transform -1 0 1790 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1064_
timestamp 0
transform -1 0 3610 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1065_
timestamp 0
transform 1 0 2530 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1066_
timestamp 0
transform -1 0 2530 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1067_
timestamp 0
transform 1 0 2390 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1068_
timestamp 0
transform -1 0 970 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1069_
timestamp 0
transform -1 0 230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1070_
timestamp 0
transform -1 0 390 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1071_
timestamp 0
transform 1 0 250 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1072_
timestamp 0
transform -1 0 90 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1073_
timestamp 0
transform 1 0 370 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1074_
timestamp 0
transform -1 0 270 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1075_
timestamp 0
transform 1 0 70 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1076_
timestamp 0
transform 1 0 370 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1077_
timestamp 0
transform -1 0 550 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1078_
timestamp 0
transform 1 0 1030 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1079_
timestamp 0
transform 1 0 690 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1080_
timestamp 0
transform 1 0 1170 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1081_
timestamp 0
transform -1 0 1030 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1082_
timestamp 0
transform 1 0 690 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1083_
timestamp 0
transform 1 0 210 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1084_
timestamp 0
transform 1 0 210 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1085_
timestamp 0
transform 1 0 350 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1086_
timestamp 0
transform -1 0 4950 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1087_
timestamp 0
transform -1 0 530 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1088_
timestamp 0
transform -1 0 390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1089_
timestamp 0
transform 1 0 530 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1090_
timestamp 0
transform 1 0 1150 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1091_
timestamp 0
transform 1 0 1510 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1092_
timestamp 0
transform 1 0 1850 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1093_
timestamp 0
transform -1 0 1670 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1094_
timestamp 0
transform 1 0 1990 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1095_
timestamp 0
transform 1 0 2150 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1096_
timestamp 0
transform -1 0 2230 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1097_
timestamp 0
transform 1 0 2070 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1098_
timestamp 0
transform 1 0 2110 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1099_
timestamp 0
transform -1 0 2830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1100_
timestamp 0
transform 1 0 2670 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1101_
timestamp 0
transform -1 0 870 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1102_
timestamp 0
transform 1 0 70 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1103_
timestamp 0
transform 1 0 1150 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1104_
timestamp 0
transform -1 0 870 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1105_
timestamp 0
transform 1 0 530 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1106_
timestamp 0
transform -1 0 810 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1107_
timestamp 0
transform -1 0 90 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1108_
timestamp 0
transform 1 0 670 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1109_
timestamp 0
transform 1 0 190 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1110_
timestamp 0
transform -1 0 90 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1111_
timestamp 0
transform 1 0 490 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1112_
timestamp 0
transform 1 0 1430 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1113_
timestamp 0
transform 1 0 670 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1114_
timestamp 0
transform -1 0 330 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1115_
timestamp 0
transform 1 0 830 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1116_
timestamp 0
transform 1 0 3910 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1117_
timestamp 0
transform -1 0 4910 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1118_
timestamp 0
transform 1 0 4390 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1119_
timestamp 0
transform 1 0 4390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1120_
timestamp 0
transform 1 0 4550 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1121_
timestamp 0
transform -1 0 4450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1122_
timestamp 0
transform 1 0 4670 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1123_
timestamp 0
transform 1 0 4710 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1124_
timestamp 0
transform 1 0 3690 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1125_
timestamp 0
transform 1 0 3850 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1126_
timestamp 0
transform 1 0 4010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1127_
timestamp 0
transform -1 0 3870 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1128_
timestamp 0
transform -1 0 3730 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1129_
timestamp 0
transform 1 0 1830 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1130_
timestamp 0
transform 1 0 990 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1131_
timestamp 0
transform 1 0 1270 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1132_
timestamp 0
transform -1 0 3890 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1133_
timestamp 0
transform 1 0 2090 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1134_
timestamp 0
transform 1 0 2170 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1135_
timestamp 0
transform 1 0 1330 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1136_
timestamp 0
transform -1 0 1790 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1137_
timestamp 0
transform 1 0 1590 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1138_
timestamp 0
transform 1 0 1490 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1139_
timestamp 0
transform 1 0 2710 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1140_
timestamp 0
transform 1 0 1330 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1141_
timestamp 0
transform 1 0 1670 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1142_
timestamp 0
transform 1 0 2010 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1143_
timestamp 0
transform 1 0 2350 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1144_
timestamp 0
transform -1 0 3050 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1145_
timestamp 0
transform 1 0 2790 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1146_
timestamp 0
transform 1 0 3190 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1147_
timestamp 0
transform 1 0 2910 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1148_
timestamp 0
transform 1 0 2890 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1149_
timestamp 0
transform 1 0 2710 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1150_
timestamp 0
transform 1 0 3210 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1151_
timestamp 0
transform 1 0 3050 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1152_
timestamp 0
transform 1 0 2490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1153_
timestamp 0
transform -1 0 2890 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1154_
timestamp 0
transform 1 0 2870 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1155_
timestamp 0
transform 1 0 4710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1156_
timestamp 0
transform 1 0 4650 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1157_
timestamp 0
transform -1 0 5050 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1158_
timestamp 0
transform -1 0 5530 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1159_
timestamp 0
transform -1 0 4850 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1160_
timestamp 0
transform 1 0 4830 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1161_
timestamp 0
transform 1 0 2250 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1162_
timestamp 0
transform -1 0 4070 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1163_
timestamp 0
transform -1 0 5010 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1164_
timestamp 0
transform 1 0 4530 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1165_
timestamp 0
transform -1 0 4870 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1166_
timestamp 0
transform 1 0 4190 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1167_
timestamp 0
transform -1 0 4370 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1168_
timestamp 0
transform 1 0 4550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1169_
timestamp 0
transform -1 0 4870 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1170_
timestamp 0
transform 1 0 4190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1171_
timestamp 0
transform 1 0 4830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1172_
timestamp 0
transform 1 0 5030 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1173_
timestamp 0
transform 1 0 850 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1174_
timestamp 0
transform 1 0 3690 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1175_
timestamp 0
transform 1 0 3290 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1176_
timestamp 0
transform 1 0 3350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1177_
timestamp 0
transform -1 0 3450 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1178_
timestamp 0
transform -1 0 4010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1179_
timestamp 0
transform 1 0 3550 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1180_
timestamp 0
transform 1 0 3290 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1181_
timestamp 0
transform 1 0 3570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1182_
timestamp 0
transform 1 0 3730 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1183_
timestamp 0
transform 1 0 4150 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1184_
timestamp 0
transform 1 0 3910 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1185_
timestamp 0
transform 1 0 3530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1186_
timestamp 0
transform 1 0 3670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1187_
timestamp 0
transform 1 0 3830 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1188_
timestamp 0
transform 1 0 3730 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1189_
timestamp 0
transform -1 0 4090 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1190_
timestamp 0
transform 1 0 4350 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1191_
timestamp 0
transform -1 0 5190 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1192_
timestamp 0
transform 1 0 3990 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1193_
timestamp 0
transform 1 0 4230 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1194_
timestamp 0
transform -1 0 4510 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1195_
timestamp 0
transform -1 0 4030 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1196_
timestamp 0
transform -1 0 1950 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1197_
timestamp 0
transform 1 0 4310 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1198_
timestamp 0
transform -1 0 4210 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1199_
timestamp 0
transform -1 0 3690 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1200_
timestamp 0
transform 1 0 3490 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1201_
timestamp 0
transform 1 0 4330 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1202_
timestamp 0
transform 1 0 4510 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1203_
timestamp 0
transform 1 0 3830 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1204_
timestamp 0
transform -1 0 4690 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1205_
timestamp 0
transform 1 0 4030 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1206_
timestamp 0
transform 1 0 2530 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1207_
timestamp 0
transform -1 0 4190 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1208_
timestamp 0
transform -1 0 3350 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1209_
timestamp 0
transform -1 0 3010 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1210_
timestamp 0
transform -1 0 3190 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1211_
timestamp 0
transform 1 0 3270 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1212_
timestamp 0
transform 1 0 3350 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1213_
timestamp 0
transform 1 0 3530 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1214_
timestamp 0
transform -1 0 3410 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1215_
timestamp 0
transform -1 0 3070 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1216_
timestamp 0
transform -1 0 2670 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1217_
timestamp 0
transform 1 0 3530 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1218_
timestamp 0
transform 1 0 5090 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1219_
timestamp 0
transform -1 0 5170 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1220_
timestamp 0
transform -1 0 4810 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1221_
timestamp 0
transform 1 0 4610 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1222_
timestamp 0
transform 1 0 4530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1223_
timestamp 0
transform 1 0 5030 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1224_
timestamp 0
transform -1 0 5150 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1225_
timestamp 0
transform 1 0 6130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1226_
timestamp 0
transform 1 0 5990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1227_
timestamp 0
transform -1 0 5370 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1228_
timestamp 0
transform 1 0 5650 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1229_
timestamp 0
transform -1 0 6350 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1230_
timestamp 0
transform 1 0 4990 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1231_
timestamp 0
transform 1 0 5130 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1232_
timestamp 0
transform 1 0 4870 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1233_
timestamp 0
transform -1 0 5190 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1234_
timestamp 0
transform 1 0 5650 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1235_
timestamp 0
transform -1 0 5510 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1236_
timestamp 0
transform -1 0 5490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1237_
timestamp 0
transform 1 0 5010 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1238_
timestamp 0
transform 1 0 4550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1239_
timestamp 0
transform -1 0 4730 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1240_
timestamp 0
transform 1 0 5330 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1241_
timestamp 0
transform 1 0 5310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1242_
timestamp 0
transform 1 0 5790 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1243_
timestamp 0
transform -1 0 3430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1244_
timestamp 0
transform 1 0 5630 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1245_
timestamp 0
transform 1 0 4150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1246_
timestamp 0
transform 1 0 4490 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1247_
timestamp 0
transform -1 0 5030 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1248_
timestamp 0
transform 1 0 4310 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1249_
timestamp 0
transform 1 0 5130 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1250_
timestamp 0
transform 1 0 5430 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1251_
timestamp 0
transform 1 0 5290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1252_
timestamp 0
transform 1 0 5730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1253_
timestamp 0
transform -1 0 5770 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1254_
timestamp 0
transform -1 0 5570 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1255_
timestamp 0
transform -1 0 4050 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1256_
timestamp 0
transform 1 0 4150 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1257_
timestamp 0
transform 1 0 3710 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1258_
timestamp 0
transform 1 0 4270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1259_
timestamp 0
transform -1 0 5310 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1260_
timestamp 0
transform 1 0 5990 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1261_
timestamp 0
transform 1 0 5950 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1262_
timestamp 0
transform 1 0 5890 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1263_
timestamp 0
transform 1 0 5450 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1264_
timestamp 0
transform 1 0 5630 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1265_
timestamp 0
transform -1 0 5950 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1266_
timestamp 0
transform 1 0 3810 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1267_
timestamp 0
transform 1 0 4670 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1268_
timestamp 0
transform 1 0 5470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1269_
timestamp 0
transform -1 0 5830 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1270_
timestamp 0
transform -1 0 5630 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1271_
timestamp 0
transform 1 0 6250 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1272_
timestamp 0
transform -1 0 6550 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1273_
timestamp 0
transform 1 0 6090 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1274_
timestamp 0
transform 1 0 5770 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1275_
timestamp 0
transform -1 0 6630 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1276_
timestamp 0
transform -1 0 6210 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1277_
timestamp 0
transform 1 0 4450 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1278_
timestamp 0
transform 1 0 4910 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1279_
timestamp 0
transform -1 0 6590 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1280_
timestamp 0
transform -1 0 6110 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1281_
timestamp 0
transform -1 0 5870 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1282_
timestamp 0
transform -1 0 5590 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1283_
timestamp 0
transform 1 0 5470 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1284_
timestamp 0
transform -1 0 6370 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1285_
timestamp 0
transform -1 0 6050 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1286_
timestamp 0
transform -1 0 5950 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1287_
timestamp 0
transform 1 0 5230 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1288_
timestamp 0
transform -1 0 5610 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1289_
timestamp 0
transform -1 0 5430 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1290_
timestamp 0
transform -1 0 5310 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1291_
timestamp 0
transform -1 0 5310 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1292_
timestamp 0
transform 1 0 5450 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1293_
timestamp 0
transform 1 0 4310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1294_
timestamp 0
transform 1 0 4250 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1295_
timestamp 0
transform -1 0 4730 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1296_
timestamp 0
transform -1 0 4750 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1297_
timestamp 0
transform 1 0 5730 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1298_
timestamp 0
transform -1 0 5770 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1299_
timestamp 0
transform 1 0 5950 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1300_
timestamp 0
transform 1 0 6410 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1301_
timestamp 0
transform -1 0 6550 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1302_
timestamp 0
transform -1 0 4410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1303_
timestamp 0
transform 1 0 5490 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1304_
timestamp 0
transform -1 0 4870 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1305_
timestamp 0
transform 1 0 5190 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1306_
timestamp 0
transform 1 0 5110 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1307_
timestamp 0
transform 1 0 5390 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1308_
timestamp 0
transform 1 0 5790 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1309_
timestamp 0
transform -1 0 4210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1310_
timestamp 0
transform 1 0 4790 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1311_
timestamp 0
transform -1 0 5350 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1312_
timestamp 0
transform 1 0 5450 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1313_
timestamp 0
transform -1 0 5150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1314_
timestamp 0
transform -1 0 5950 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1315_
timestamp 0
transform 1 0 5290 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1316_
timestamp 0
transform -1 0 5630 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1317_
timestamp 0
transform 1 0 5650 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1318_
timestamp 0
transform 1 0 5770 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1319_
timestamp 0
transform 1 0 5810 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1320_
timestamp 0
transform 1 0 5610 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1321_
timestamp 0
transform 1 0 6090 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1322_
timestamp 0
transform 1 0 6250 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1323_
timestamp 0
transform 1 0 6250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1324_
timestamp 0
transform -1 0 6490 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1325_
timestamp 0
transform 1 0 6290 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1326_
timestamp 0
transform 1 0 4970 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1327_
timestamp 0
transform 1 0 4450 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1328_
timestamp 0
transform 1 0 4170 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1329_
timestamp 0
transform -1 0 4370 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1330_
timestamp 0
transform 1 0 4490 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1331_
timestamp 0
transform 1 0 4630 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1332_
timestamp 0
transform 1 0 5110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1333_
timestamp 0
transform 1 0 4470 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1334_
timestamp 0
transform 1 0 4950 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1335_
timestamp 0
transform 1 0 4010 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1336_
timestamp 0
transform 1 0 5390 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1337_
timestamp 0
transform 1 0 5550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1338_
timestamp 0
transform 1 0 4970 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1339_
timestamp 0
transform -1 0 6050 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1340_
timestamp 0
transform -1 0 4690 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1341_
timestamp 0
transform 1 0 3450 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1342_
timestamp 0
transform 1 0 3570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1343_
timestamp 0
transform -1 0 3890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1344_
timestamp 0
transform -1 0 4290 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1345_
timestamp 0
transform 1 0 4590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1346_
timestamp 0
transform 1 0 5290 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1347_
timestamp 0
transform 1 0 4350 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1348_
timestamp 0
transform 1 0 3730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1349_
timestamp 0
transform 1 0 5430 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1350_
timestamp 0
transform -1 0 6070 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1351_
timestamp 0
transform 1 0 5610 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1352_
timestamp 0
transform 1 0 4410 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1353_
timestamp 0
transform 1 0 5550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1354_
timestamp 0
transform 1 0 6070 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1355_
timestamp 0
transform 1 0 5710 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1356_
timestamp 0
transform 1 0 6210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1357_
timestamp 0
transform 1 0 5710 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1358_
timestamp 0
transform 1 0 6530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1359_
timestamp 0
transform -1 0 6310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1360_
timestamp 0
transform 1 0 6050 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1361_
timestamp 0
transform 1 0 6110 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1362_
timestamp 0
transform -1 0 6390 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1363_
timestamp 0
transform 1 0 5910 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1364_
timestamp 0
transform 1 0 5950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1365_
timestamp 0
transform -1 0 6450 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1366_
timestamp 0
transform 1 0 6550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1367_
timestamp 0
transform 1 0 6230 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1368_
timestamp 0
transform 1 0 6130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1369_
timestamp 0
transform 1 0 6590 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1370_
timestamp 0
transform -1 0 6290 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1371_
timestamp 0
transform 1 0 6170 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1372_
timestamp 0
transform 1 0 6250 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1373_
timestamp 0
transform 1 0 6630 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1374_
timestamp 0
transform -1 0 6410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1375_
timestamp 0
transform -1 0 6230 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1376_
timestamp 0
transform -1 0 5930 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1377_
timestamp 0
transform 1 0 6570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1378_
timestamp 0
transform -1 0 6470 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1379_
timestamp 0
transform -1 0 6390 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1380_
timestamp 0
transform -1 0 6270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1381_
timestamp 0
transform -1 0 5810 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1382_
timestamp 0
transform -1 0 6550 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1383_
timestamp 0
transform -1 0 6430 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1384_
timestamp 0
transform -1 0 6430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1385_
timestamp 0
transform -1 0 6110 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1386_
timestamp 0
transform -1 0 6110 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1387_
timestamp 0
transform 1 0 5330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1388_
timestamp 0
transform 1 0 4750 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1389_
timestamp 0
transform -1 0 4630 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1390_
timestamp 0
transform -1 0 5070 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1391_
timestamp 0
transform 1 0 4430 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1392_
timestamp 0
transform 1 0 4070 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1393_
timestamp 0
transform 1 0 3910 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1394_
timestamp 0
transform -1 0 5170 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1395_
timestamp 0
transform -1 0 5190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1396_
timestamp 0
transform -1 0 5010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1397_
timestamp 0
transform -1 0 6630 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1398_
timestamp 0
transform 1 0 6650 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1399_
timestamp 0
transform -1 0 6610 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1400_
timestamp 0
transform -1 0 6530 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1401_
timestamp 0
transform -1 0 6470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1402_
timestamp 0
transform -1 0 6590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1403_
timestamp 0
transform -1 0 5750 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1404_
timestamp 0
transform -1 0 4130 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1405_
timestamp 0
transform 1 0 4950 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1406_
timestamp 0
transform -1 0 4790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1407_
timestamp 0
transform 1 0 4390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1408_
timestamp 0
transform -1 0 4770 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1409_
timestamp 0
transform -1 0 4710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1410_
timestamp 0
transform -1 0 4850 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1411_
timestamp 0
transform -1 0 4910 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1412_
timestamp 0
transform 1 0 4430 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1413_
timestamp 0
transform -1 0 4830 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1414_
timestamp 0
transform 1 0 4790 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1415_
timestamp 0
transform 1 0 4590 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1416_
timestamp 0
transform 1 0 5230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1417_
timestamp 0
transform 1 0 5250 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1418_
timestamp 0
transform 1 0 4610 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1419_
timestamp 0
transform 1 0 5050 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1420_
timestamp 0
transform 1 0 4310 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1421_
timestamp 0
transform 1 0 4250 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1422_
timestamp 0
transform 1 0 5410 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1423_
timestamp 0
transform 1 0 5730 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1424_
timestamp 0
transform 1 0 5250 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1425_
timestamp 0
transform 1 0 5570 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1426_
timestamp 0
transform 1 0 5570 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1427_
timestamp 0
transform 1 0 5070 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1428_
timestamp 0
transform -1 0 5910 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1429_
timestamp 0
transform 1 0 5770 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1430_
timestamp 0
transform 1 0 6210 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1431_
timestamp 0
transform -1 0 6370 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1432_
timestamp 0
transform 1 0 4910 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1433_
timestamp 0
transform -1 0 4330 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1434_
timestamp 0
transform 1 0 4730 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1435_
timestamp 0
transform -1 0 4650 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1436_
timestamp 0
transform 1 0 4770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1437_
timestamp 0
transform 1 0 5070 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1438_
timestamp 0
transform 1 0 5230 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1439_
timestamp 0
transform 1 0 3150 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1440_
timestamp 0
transform -1 0 4970 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1441_
timestamp 0
transform 1 0 4150 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1442_
timestamp 0
transform 1 0 5390 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1443_
timestamp 0
transform 1 0 5570 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1444_
timestamp 0
transform 1 0 3710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1445_
timestamp 0
transform 1 0 3190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1446_
timestamp 0
transform -1 0 3990 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1447_
timestamp 0
transform -1 0 4570 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1448_
timestamp 0
transform 1 0 4990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1449_
timestamp 0
transform 1 0 4510 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1450_
timestamp 0
transform 1 0 4990 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1451_
timestamp 0
transform 1 0 4690 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1452_
timestamp 0
transform 1 0 5350 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1453_
timestamp 0
transform -1 0 5730 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1454_
timestamp 0
transform 1 0 4190 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1455_
timestamp 0
transform 1 0 4050 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1456_
timestamp 0
transform -1 0 5410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1457_
timestamp 0
transform 1 0 5510 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1458_
timestamp 0
transform 1 0 5550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1459_
timestamp 0
transform 1 0 5650 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1460_
timestamp 0
transform 1 0 5890 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1461_
timestamp 0
transform 1 0 6050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1462_
timestamp 0
transform -1 0 5110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1463_
timestamp 0
transform 1 0 5330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1464_
timestamp 0
transform 1 0 5890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1465_
timestamp 0
transform 1 0 5170 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1466_
timestamp 0
transform 1 0 5790 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1467_
timestamp 0
transform 1 0 5910 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1468_
timestamp 0
transform -1 0 6090 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1469_
timestamp 0
transform 1 0 5490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1470_
timestamp 0
transform 1 0 5950 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1471_
timestamp 0
transform -1 0 6010 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1472_
timestamp 0
transform 1 0 6150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1473_
timestamp 0
transform 1 0 6410 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1474_
timestamp 0
transform -1 0 6590 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1475_
timestamp 0
transform 1 0 6170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1476_
timestamp 0
transform 1 0 5830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1477_
timestamp 0
transform 1 0 6410 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1478_
timestamp 0
transform -1 0 6510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1479_
timestamp 0
transform 1 0 6250 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1480_
timestamp 0
transform -1 0 6350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1481_
timestamp 0
transform 1 0 6590 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1482_
timestamp 0
transform 1 0 6650 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1483_
timestamp 0
transform -1 0 6670 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1484_
timestamp 0
transform 1 0 6550 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1485_
timestamp 0
transform -1 0 6690 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1486_
timestamp 0
transform -1 0 6330 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1487_
timestamp 0
transform -1 0 6530 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1488_
timestamp 0
transform -1 0 4870 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1489_
timestamp 0
transform 1 0 4010 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1490_
timestamp 0
transform 1 0 4050 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1491_
timestamp 0
transform -1 0 5070 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1492_
timestamp 0
transform 1 0 4870 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1493_
timestamp 0
transform 1 0 6410 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1494_
timestamp 0
transform 1 0 6530 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1495_
timestamp 0
transform -1 0 5890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1496_
timestamp 0
transform 1 0 6310 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1497_
timestamp 0
transform -1 0 6130 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1498_
timestamp 0
transform 1 0 6230 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1499_
timestamp 0
transform 1 0 5210 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1500_
timestamp 0
transform -1 0 4610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1501_
timestamp 0
transform 1 0 4110 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1502_
timestamp 0
transform 1 0 4850 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1503_
timestamp 0
transform -1 0 4750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1504_
timestamp 0
transform 1 0 5150 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1505_
timestamp 0
transform 1 0 4870 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1506_
timestamp 0
transform -1 0 4550 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1507_
timestamp 0
transform 1 0 4550 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1508_
timestamp 0
transform -1 0 5050 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1509_
timestamp 0
transform 1 0 5170 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1510_
timestamp 0
transform 1 0 4890 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1511_
timestamp 0
transform 1 0 5230 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1512_
timestamp 0
transform -1 0 5370 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1513_
timestamp 0
transform 1 0 4990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1514_
timestamp 0
transform 1 0 4990 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1515_
timestamp 0
transform 1 0 5050 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1516_
timestamp 0
transform 1 0 5570 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1517_
timestamp 0
transform 1 0 5510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1518_
timestamp 0
transform 1 0 5150 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1519_
timestamp 0
transform 1 0 5370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1520_
timestamp 0
transform 1 0 5330 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1521_
timestamp 0
transform 1 0 5410 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1522_
timestamp 0
transform 1 0 5490 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1523_
timestamp 0
transform 1 0 5650 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1524_
timestamp 0
transform -1 0 5190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1525_
timestamp 0
transform -1 0 5890 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1526_
timestamp 0
transform 1 0 3670 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1527_
timestamp 0
transform 1 0 3170 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1528_
timestamp 0
transform -1 0 3990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1529_
timestamp 0
transform 1 0 3510 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1530_
timestamp 0
transform 1 0 3810 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1531_
timestamp 0
transform 1 0 4590 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1532_
timestamp 0
transform -1 0 3630 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1533_
timestamp 0
transform -1 0 3890 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1534_
timestamp 0
transform -1 0 4430 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1535_
timestamp 0
transform -1 0 4470 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1536_
timestamp 0
transform 1 0 4090 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1537_
timestamp 0
transform 1 0 4270 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1538_
timestamp 0
transform 1 0 4410 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1539_
timestamp 0
transform 1 0 4290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1540_
timestamp 0
transform 1 0 5670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1541_
timestamp 0
transform -1 0 5850 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1542_
timestamp 0
transform -1 0 5270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1543_
timestamp 0
transform 1 0 5710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1544_
timestamp 0
transform -1 0 5770 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1545_
timestamp 0
transform -1 0 5690 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1546_
timestamp 0
transform 1 0 6110 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1547_
timestamp 0
transform 1 0 5910 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1548_
timestamp 0
transform -1 0 5990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1549_
timestamp 0
transform 1 0 6290 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1550_
timestamp 0
transform -1 0 6310 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1551_
timestamp 0
transform 1 0 5630 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1552_
timestamp 0
transform 1 0 6050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1553_
timestamp 0
transform 1 0 6110 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1554_
timestamp 0
transform 1 0 5830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1555_
timestamp 0
transform -1 0 6070 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1556_
timestamp 0
transform 1 0 5990 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1557_
timestamp 0
transform -1 0 6170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1558_
timestamp 0
transform 1 0 6410 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1559_
timestamp 0
transform 1 0 6610 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1560_
timestamp 0
transform 1 0 6070 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1561_
timestamp 0
transform -1 0 6610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1562_
timestamp 0
transform -1 0 6610 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1563_
timestamp 0
transform -1 0 6450 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1564_
timestamp 0
transform 1 0 6230 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1565_
timestamp 0
transform 1 0 6390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1566_
timestamp 0
transform -1 0 6590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1567_
timestamp 0
transform -1 0 4490 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1568_
timestamp 0
transform 1 0 4210 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1569_
timestamp 0
transform -1 0 4250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1570_
timestamp 0
transform -1 0 3770 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1571_
timestamp 0
transform 1 0 6230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1572_
timestamp 0
transform -1 0 4350 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1573_
timestamp 0
transform -1 0 3710 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1574_
timestamp 0
transform 1 0 6450 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1575_
timestamp 0
transform 1 0 6470 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1576_
timestamp 0
transform 1 0 5490 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1577_
timestamp 0
transform -1 0 5510 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1578_
timestamp 0
transform -1 0 5970 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1579_
timestamp 0
transform -1 0 4710 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1580_
timestamp 0
transform 1 0 4410 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1581_
timestamp 0
transform -1 0 3050 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1582_
timestamp 0
transform -1 0 2850 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1583_
timestamp 0
transform -1 0 2910 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1584_
timestamp 0
transform -1 0 3050 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1585_
timestamp 0
transform 1 0 3190 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1586_
timestamp 0
transform 1 0 2710 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1587_
timestamp 0
transform 1 0 2830 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1588_
timestamp 0
transform -1 0 2010 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1589_
timestamp 0
transform -1 0 2710 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1590_
timestamp 0
transform 1 0 2950 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1591_
timestamp 0
transform 1 0 3910 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1592_
timestamp 0
transform -1 0 3770 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1593_
timestamp 0
transform -1 0 3790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1594_
timestamp 0
transform 1 0 3110 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1595_
timestamp 0
transform 1 0 3030 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1596_
timestamp 0
transform -1 0 4090 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1597_
timestamp 0
transform -1 0 4250 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1598_
timestamp 0
transform 1 0 4090 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1599_
timestamp 0
transform -1 0 4270 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1600_
timestamp 0
transform 1 0 3590 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1601_
timestamp 0
transform 1 0 3930 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1602_
timestamp 0
transform -1 0 3930 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1603_
timestamp 0
transform 1 0 4830 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1604_
timestamp 0
transform 1 0 3690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1605_
timestamp 0
transform 1 0 3530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1606_
timestamp 0
transform 1 0 1410 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1607_
timestamp 0
transform -1 0 3390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1608_
timestamp 0
transform -1 0 2750 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1609_
timestamp 0
transform 1 0 3170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1610_
timestamp 0
transform -1 0 2430 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1611_
timestamp 0
transform -1 0 2590 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1612_
timestamp 0
transform 1 0 1550 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1613_
timestamp 0
transform 1 0 3310 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1614_
timestamp 0
transform 1 0 3450 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1615_
timestamp 0
transform 1 0 3810 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1616_
timestamp 0
transform 1 0 3170 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1617_
timestamp 0
transform -1 0 3630 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1618_
timestamp 0
transform 1 0 4250 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1619_
timestamp 0
transform -1 0 4710 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1620_
timestamp 0
transform 1 0 3790 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1621_
timestamp 0
transform 1 0 3470 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1622_
timestamp 0
transform 1 0 3970 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1623_
timestamp 0
transform 1 0 4990 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1624_
timestamp 0
transform 1 0 5950 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1625_
timestamp 0
transform 1 0 5790 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1626_
timestamp 0
transform 1 0 4230 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1627_
timestamp 0
transform -1 0 4570 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1628_
timestamp 0
transform 1 0 4870 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1629_
timestamp 0
transform 1 0 6270 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1630_
timestamp 0
transform -1 0 5810 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1631_
timestamp 0
transform 1 0 4710 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1632_
timestamp 0
transform 1 0 5610 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1633_
timestamp 0
transform 1 0 6450 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1634_
timestamp 0
transform 1 0 6230 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1635_
timestamp 0
transform -1 0 6490 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1636_
timestamp 0
transform 1 0 5150 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1637_
timestamp 0
transform -1 0 6130 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1638_
timestamp 0
transform 1 0 5310 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1639_
timestamp 0
transform 1 0 4710 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1640_
timestamp 0
transform 1 0 3550 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1641_
timestamp 0
transform 1 0 3370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1642_
timestamp 0
transform 1 0 3590 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1643_
timestamp 0
transform 1 0 2250 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1644_
timestamp 0
transform -1 0 3210 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1645_
timestamp 0
transform -1 0 5350 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1646_
timestamp 0
transform -1 0 5190 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1647_
timestamp 0
transform 1 0 3750 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1648_
timestamp 0
transform -1 0 3810 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1649_
timestamp 0
transform -1 0 4090 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1650_
timestamp 0
transform -1 0 3470 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1651_
timestamp 0
transform -1 0 3610 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1652_
timestamp 0
transform -1 0 2570 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1653_
timestamp 0
transform 1 0 2530 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1654_
timestamp 0
transform -1 0 2430 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1655_
timestamp 0
transform -1 0 2230 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1656_
timestamp 0
transform 1 0 1710 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1657_
timestamp 0
transform -1 0 2110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1658_
timestamp 0
transform 1 0 1850 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1659_
timestamp 0
transform -1 0 2070 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1660_
timestamp 0
transform -1 0 2290 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1661_
timestamp 0
transform 1 0 2130 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1662_
timestamp 0
transform 1 0 2230 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1663_
timestamp 0
transform -1 0 1970 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1664_
timestamp 0
transform -1 0 1670 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1665_
timestamp 0
transform -1 0 1490 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1666_
timestamp 0
transform -1 0 1910 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1667_
timestamp 0
transform 1 0 1490 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1668_
timestamp 0
transform 1 0 2030 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1669_
timestamp 0
transform 1 0 2370 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1670_
timestamp 0
transform 1 0 1330 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1671_
timestamp 0
transform -1 0 1790 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1672_
timestamp 0
transform 1 0 1870 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1673_
timestamp 0
transform -1 0 90 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1674_
timestamp 0
transform -1 0 90 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1675_
timestamp 0
transform 1 0 70 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1676_
timestamp 0
transform 1 0 230 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1677_
timestamp 0
transform 1 0 370 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1678_
timestamp 0
transform 1 0 2210 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1679_
timestamp 0
transform -1 0 1730 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1680_
timestamp 0
transform -1 0 1550 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1681_
timestamp 0
transform 1 0 1250 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1682_
timestamp 0
transform -1 0 1390 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1683_
timestamp 0
transform 1 0 2630 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1684_
timestamp 0
transform -1 0 2510 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1685_
timestamp 0
transform -1 0 3310 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1686_
timestamp 0
transform 1 0 3910 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1687_
timestamp 0
transform -1 0 4410 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1688_
timestamp 0
transform 1 0 2810 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1689_
timestamp 0
transform -1 0 2990 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1690_
timestamp 0
transform -1 0 3150 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1691_
timestamp 0
transform -1 0 4110 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1692_
timestamp 0
transform -1 0 4590 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1693_
timestamp 0
transform -1 0 4430 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1694_
timestamp 0
transform 1 0 3290 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1695_
timestamp 0
transform -1 0 3630 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1696_
timestamp 0
transform 1 0 3450 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1697_
timestamp 0
transform -1 0 3490 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1698_
timestamp 0
transform -1 0 2890 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1699_
timestamp 0
transform 1 0 3050 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1700_
timestamp 0
transform -1 0 2910 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1701_
timestamp 0
transform 1 0 2610 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1702_
timestamp 0
transform 1 0 3050 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1703_
timestamp 0
transform 1 0 3370 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1704_
timestamp 0
transform -1 0 3530 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1705_
timestamp 0
transform -1 0 3350 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1706_
timestamp 0
transform 1 0 3330 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1707_
timestamp 0
transform -1 0 3030 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1708_
timestamp 0
transform -1 0 2410 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1709_
timestamp 0
transform 1 0 1110 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1710_
timestamp 0
transform 1 0 70 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1711_
timestamp 0
transform 1 0 1730 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1712_
timestamp 0
transform 1 0 2370 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1713_
timestamp 0
transform -1 0 2210 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1714_
timestamp 0
transform -1 0 2270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1715_
timestamp 0
transform 1 0 2050 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1716_
timestamp 0
transform 1 0 1930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1717_
timestamp 0
transform 1 0 1710 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1718_
timestamp 0
transform 1 0 1790 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1719_
timestamp 0
transform -1 0 1170 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1720_
timestamp 0
transform -1 0 1330 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1721_
timestamp 0
transform -1 0 770 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1722_
timestamp 0
transform 1 0 230 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1723_
timestamp 0
transform 1 0 290 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1724_
timestamp 0
transform 1 0 250 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1725_
timestamp 0
transform -1 0 90 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1726_
timestamp 0
transform 1 0 390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1727_
timestamp 0
transform -1 0 550 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1728_
timestamp 0
transform -1 0 990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1729_
timestamp 0
transform 1 0 690 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1730_
timestamp 0
transform -1 0 830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1731_
timestamp 0
transform 1 0 250 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1732_
timestamp 0
transform 1 0 430 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1733_
timestamp 0
transform 1 0 530 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1734_
timestamp 0
transform 1 0 690 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1735_
timestamp 0
transform -1 0 1010 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1736_
timestamp 0
transform -1 0 590 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1737_
timestamp 0
transform 1 0 690 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1738_
timestamp 0
transform 1 0 830 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1739_
timestamp 0
transform 1 0 1170 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1740_
timestamp 0
transform -1 0 2270 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1741_
timestamp 0
transform -1 0 1050 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1742_
timestamp 0
transform -1 0 2130 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1743_
timestamp 0
transform 1 0 2850 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1744_
timestamp 0
transform -1 0 2970 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1745_
timestamp 0
transform 1 0 2710 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1746_
timestamp 0
transform -1 0 2570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1747_
timestamp 0
transform -1 0 2810 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1748_
timestamp 0
transform 1 0 870 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1749_
timestamp 0
transform -1 0 1870 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1750_
timestamp 0
transform -1 0 2130 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1751_
timestamp 0
transform -1 0 1970 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1752_
timestamp 0
transform 1 0 1850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1753_
timestamp 0
transform -1 0 1670 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1754_
timestamp 0
transform 1 0 1790 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1755_
timestamp 0
transform -1 0 1370 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1756_
timestamp 0
transform -1 0 530 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1757_
timestamp 0
transform 1 0 430 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1758_
timestamp 0
transform -1 0 450 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1759_
timestamp 0
transform 1 0 590 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1760_
timestamp 0
transform 1 0 570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1761_
timestamp 0
transform -1 0 1050 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1762_
timestamp 0
transform 1 0 870 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1763_
timestamp 0
transform -1 0 930 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1764_
timestamp 0
transform 1 0 1990 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1765_
timestamp 0
transform -1 0 2690 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1766_
timestamp 0
transform 1 0 2510 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1767_
timestamp 0
transform 1 0 2550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1768_
timestamp 0
transform -1 0 2410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1769_
timestamp 0
transform -1 0 2430 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1770_
timestamp 0
transform 1 0 2250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1771_
timestamp 0
transform 1 0 2690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1772_
timestamp 0
transform -1 0 2870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1773_
timestamp 0
transform 1 0 2390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1774_
timestamp 0
transform 1 0 1630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1775_
timestamp 0
transform 1 0 1570 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1776_
timestamp 0
transform 1 0 730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1777_
timestamp 0
transform -1 0 1230 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1778_
timestamp 0
transform -1 0 1690 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1779_
timestamp 0
transform -1 0 1490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1780_
timestamp 0
transform 1 0 370 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1781_
timestamp 0
transform 1 0 710 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1782_
timestamp 0
transform 1 0 330 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1783_
timestamp 0
transform 1 0 470 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1784_
timestamp 0
transform -1 0 630 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1785_
timestamp 0
transform -1 0 790 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1786_
timestamp 0
transform 1 0 1090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1787_
timestamp 0
transform 1 0 930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1788_
timestamp 0
transform 1 0 1410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1789_
timestamp 0
transform 1 0 1730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1790_
timestamp 0
transform -1 0 2250 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1791_
timestamp 0
transform -1 0 1590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1792_
timestamp 0
transform 1 0 1250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1793_
timestamp 0
transform -1 0 910 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1794_
timestamp 0
transform 1 0 1490 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1795_
timestamp 0
transform -1 0 870 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1796_
timestamp 0
transform 1 0 630 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1797_
timestamp 0
transform 1 0 1050 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1798_
timestamp 0
transform 1 0 1170 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1799_
timestamp 0
transform 1 0 1310 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1800_
timestamp 0
transform -1 0 1870 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1801_
timestamp 0
transform 1 0 1670 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1802_
timestamp 0
transform 1 0 70 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1803_
timestamp 0
transform 1 0 970 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1804_
timestamp 0
transform -1 0 1110 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1805_
timestamp 0
transform 1 0 190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1806_
timestamp 0
transform 1 0 310 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1807_
timestamp 0
transform 1 0 210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1808_
timestamp 0
transform 1 0 470 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1809_
timestamp 0
transform 1 0 310 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1810_
timestamp 0
transform 1 0 70 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1811_
timestamp 0
transform -1 0 1090 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1812_
timestamp 0
transform 1 0 910 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1813_
timestamp 0
transform 1 0 210 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1814_
timestamp 0
transform 1 0 870 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1815_
timestamp 0
transform 1 0 470 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1816_
timestamp 0
transform 1 0 990 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1817_
timestamp 0
transform -1 0 770 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1818_
timestamp 0
transform 1 0 350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1819_
timestamp 0
transform -1 0 1090 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1820_
timestamp 0
transform -1 0 1230 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1821_
timestamp 0
transform 1 0 70 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1822_
timestamp 0
transform -1 0 1070 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1823_
timestamp 0
transform 1 0 70 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1824_
timestamp 0
transform 1 0 70 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1825_
timestamp 0
transform -1 0 1150 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1826_
timestamp 0
transform -1 0 970 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1827_
timestamp 0
transform 1 0 550 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1828_
timestamp 0
transform 1 0 1790 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1829_
timestamp 0
transform 1 0 1610 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1830_
timestamp 0
transform -1 0 1470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1831_
timestamp 0
transform 1 0 970 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1832_
timestamp 0
transform -1 0 810 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1833_
timestamp 0
transform 1 0 630 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1834_
timestamp 0
transform -1 0 90 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1835_
timestamp 0
transform -1 0 530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1836_
timestamp 0
transform 1 0 910 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1837_
timestamp 0
transform -1 0 770 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1838_
timestamp 0
transform 1 0 450 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1839_
timestamp 0
transform -1 0 370 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1840_
timestamp 0
transform -1 0 90 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1841_
timestamp 0
transform -1 0 230 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1842_
timestamp 0
transform -1 0 1230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1843_
timestamp 0
transform -1 0 1370 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1844_
timestamp 0
transform 1 0 1870 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1845_
timestamp 0
transform 1 0 2030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1846_
timestamp 0
transform -1 0 2990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1847_
timestamp 0
transform -1 0 3130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1848_
timestamp 0
transform -1 0 390 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1849_
timestamp 0
transform 1 0 210 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1911_
timestamp 0
transform -1 0 2730 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1912_
timestamp 0
transform -1 0 90 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1913_
timestamp 0
transform 1 0 2430 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1914_
timestamp 0
transform -1 0 90 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1915_
timestamp 0
transform -1 0 90 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1916_
timestamp 0
transform -1 0 2590 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1917_
timestamp 0
transform -1 0 2510 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1918_
timestamp 0
transform -1 0 250 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1919_
timestamp 0
transform -1 0 90 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert0
timestamp 0
transform 1 0 3150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert1
timestamp 0
transform 1 0 2850 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert2
timestamp 0
transform 1 0 3290 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert3
timestamp 0
transform 1 0 3290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert4
timestamp 0
transform -1 0 2730 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert12
timestamp 0
transform 1 0 3570 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert13
timestamp 0
transform 1 0 70 0 1 1310
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert14
timestamp 0
transform 1 0 610 0 1 1830
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert15
timestamp 0
transform 1 0 3610 0 1 2350
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert16
timestamp 0
transform 1 0 830 0 1 2870
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert17
timestamp 0
transform 1 0 1130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert18
timestamp 0
transform -1 0 230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert19
timestamp 0
transform -1 0 1110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert20
timestamp 0
transform -1 0 390 0 1 2870
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert21
timestamp 0
transform 1 0 3430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert22
timestamp 0
transform -1 0 3170 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert23
timestamp 0
transform 1 0 3430 0 1 3910
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert24
timestamp 0
transform -1 0 3170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert25
timestamp 0
transform -1 0 3290 0 1 3910
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert5
timestamp 0
transform -1 0 1050 0 1 3910
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert6
timestamp 0
transform 1 0 2090 0 1 3390
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert7
timestamp 0
transform 1 0 1050 0 1 2350
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert8
timestamp 0
transform -1 0 250 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert9
timestamp 0
transform 1 0 210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert10
timestamp 0
transform 1 0 2710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert11
timestamp 0
transform 1 0 1710 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__922_
timestamp 0
transform -1 0 990 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__925_
timestamp 0
transform 1 0 2530 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__928_
timestamp 0
transform -1 0 1990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__931_
timestamp 0
transform -1 0 3670 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__934_
timestamp 0
transform 1 0 2910 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__937_
timestamp 0
transform 1 0 2370 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__940_
timestamp 0
transform 1 0 2050 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__943_
timestamp 0
transform 1 0 1510 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__946_
timestamp 0
transform -1 0 4510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__949_
timestamp 0
transform 1 0 3770 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__952_
timestamp 0
transform 1 0 3890 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__955_
timestamp 0
transform 1 0 2730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__958_
timestamp 0
transform 1 0 1110 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__961_
timestamp 0
transform -1 0 2830 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__964_
timestamp 0
transform 1 0 1310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__967_
timestamp 0
transform 1 0 2710 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__970_
timestamp 0
transform -1 0 3130 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__973_
timestamp 0
transform -1 0 2530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__976_
timestamp 0
transform 1 0 2250 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__979_
timestamp 0
transform 1 0 3310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__982_
timestamp 0
transform -1 0 2930 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__985_
timestamp 0
transform 1 0 4150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__988_
timestamp 0
transform 1 0 3710 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__991_
timestamp 0
transform 1 0 2830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__994_
timestamp 0
transform -1 0 4050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__997_
timestamp 0
transform 1 0 1750 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1000_
timestamp 0
transform -1 0 3150 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1003_
timestamp 0
transform 1 0 2970 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1006_
timestamp 0
transform 1 0 1910 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1009_
timestamp 0
transform 1 0 1150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1012_
timestamp 0
transform 1 0 2370 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1015_
timestamp 0
transform -1 0 1850 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1018_
timestamp 0
transform 1 0 2150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1021_
timestamp 0
transform 1 0 1250 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1024_
timestamp 0
transform 1 0 1270 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1027_
timestamp 0
transform 1 0 1570 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1030_
timestamp 0
transform -1 0 1590 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1033_
timestamp 0
transform 1 0 2350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1036_
timestamp 0
transform -1 0 1330 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1039_
timestamp 0
transform -1 0 1630 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1042_
timestamp 0
transform 1 0 830 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1045_
timestamp 0
transform 1 0 1150 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1048_
timestamp 0
transform 1 0 1270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1051_
timestamp 0
transform 1 0 1450 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1054_
timestamp 0
transform 1 0 2370 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1057_
timestamp 0
transform -1 0 1810 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1060_
timestamp 0
transform 1 0 1930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1063_
timestamp 0
transform -1 0 1810 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1066_
timestamp 0
transform -1 0 2550 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1069_
timestamp 0
transform -1 0 250 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1072_
timestamp 0
transform -1 0 110 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1075_
timestamp 0
transform 1 0 90 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1078_
timestamp 0
transform 1 0 1050 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1081_
timestamp 0
transform -1 0 1050 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1084_
timestamp 0
transform 1 0 230 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1087_
timestamp 0
transform -1 0 550 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1090_
timestamp 0
transform 1 0 1170 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1093_
timestamp 0
transform -1 0 1690 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1096_
timestamp 0
transform -1 0 2250 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1099_
timestamp 0
transform -1 0 2850 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1102_
timestamp 0
transform 1 0 90 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1105_
timestamp 0
transform 1 0 550 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1108_
timestamp 0
transform 1 0 690 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1111_
timestamp 0
transform 1 0 510 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1114_
timestamp 0
transform -1 0 350 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1117_
timestamp 0
transform -1 0 4930 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1120_
timestamp 0
transform 1 0 4570 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1123_
timestamp 0
transform 1 0 4730 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1126_
timestamp 0
transform 1 0 4030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1129_
timestamp 0
transform 1 0 1850 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1132_
timestamp 0
transform -1 0 3910 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1134_
timestamp 0
transform 1 0 2190 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1137_
timestamp 0
transform 1 0 1610 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1140_
timestamp 0
transform 1 0 1350 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1143_
timestamp 0
transform 1 0 2370 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1146_
timestamp 0
transform 1 0 3210 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1149_
timestamp 0
transform 1 0 2730 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1152_
timestamp 0
transform 1 0 2510 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1155_
timestamp 0
transform 1 0 4730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1158_
timestamp 0
transform -1 0 5550 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1161_
timestamp 0
transform 1 0 2270 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1164_
timestamp 0
transform 1 0 4550 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1167_
timestamp 0
transform -1 0 4390 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1170_
timestamp 0
transform 1 0 4210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1173_
timestamp 0
transform 1 0 870 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1176_
timestamp 0
transform 1 0 3370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1179_
timestamp 0
transform 1 0 3570 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1182_
timestamp 0
transform 1 0 3750 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1185_
timestamp 0
transform 1 0 3550 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1188_
timestamp 0
transform 1 0 3750 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1191_
timestamp 0
transform -1 0 5210 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1194_
timestamp 0
transform -1 0 4530 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1197_
timestamp 0
transform 1 0 4330 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1200_
timestamp 0
transform 1 0 3510 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1203_
timestamp 0
transform 1 0 3850 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1206_
timestamp 0
transform 1 0 2550 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1209_
timestamp 0
transform -1 0 3030 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1212_
timestamp 0
transform 1 0 3370 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1215_
timestamp 0
transform -1 0 3090 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1218_
timestamp 0
transform 1 0 5110 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1221_
timestamp 0
transform 1 0 4630 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1224_
timestamp 0
transform -1 0 5170 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1227_
timestamp 0
transform -1 0 5390 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1230_
timestamp 0
transform 1 0 5010 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1233_
timestamp 0
transform -1 0 5210 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1236_
timestamp 0
transform -1 0 5510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1239_
timestamp 0
transform -1 0 4750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1242_
timestamp 0
transform 1 0 5810 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1245_
timestamp 0
transform 1 0 4170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1248_
timestamp 0
transform 1 0 4330 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1251_
timestamp 0
transform 1 0 5310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1254_
timestamp 0
transform -1 0 5590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1257_
timestamp 0
transform 1 0 3730 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1260_
timestamp 0
transform 1 0 6010 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1263_
timestamp 0
transform 1 0 5470 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1266_
timestamp 0
transform 1 0 3830 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1269_
timestamp 0
transform -1 0 5850 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1272_
timestamp 0
transform -1 0 6570 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1275_
timestamp 0
transform -1 0 6650 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1278_
timestamp 0
transform 1 0 4930 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1281_
timestamp 0
transform -1 0 5890 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1284_
timestamp 0
transform -1 0 6390 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1287_
timestamp 0
transform 1 0 5250 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1290_
timestamp 0
transform -1 0 5330 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1293_
timestamp 0
transform 1 0 4330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1295_
timestamp 0
transform -1 0 4750 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1298_
timestamp 0
transform -1 0 5790 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1301_
timestamp 0
transform -1 0 6570 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1304_
timestamp 0
transform -1 0 4890 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1307_
timestamp 0
transform 1 0 5410 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1310_
timestamp 0
transform 1 0 4810 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1313_
timestamp 0
transform -1 0 5170 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1316_
timestamp 0
transform -1 0 5650 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1319_
timestamp 0
transform 1 0 5830 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1322_
timestamp 0
transform 1 0 6270 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1325_
timestamp 0
transform 1 0 6310 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1328_
timestamp 0
transform 1 0 4190 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1331_
timestamp 0
transform 1 0 4650 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1334_
timestamp 0
transform 1 0 4970 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1337_
timestamp 0
transform 1 0 5570 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1340_
timestamp 0
transform -1 0 4710 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1343_
timestamp 0
transform -1 0 3910 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1346_
timestamp 0
transform 1 0 5310 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1349_
timestamp 0
transform 1 0 5450 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1352_
timestamp 0
transform 1 0 4430 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1355_
timestamp 0
transform 1 0 5730 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1358_
timestamp 0
transform 1 0 6550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1361_
timestamp 0
transform 1 0 6130 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1364_
timestamp 0
transform 1 0 5970 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1367_
timestamp 0
transform 1 0 6250 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1370_
timestamp 0
transform -1 0 6310 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1373_
timestamp 0
transform 1 0 6650 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1376_
timestamp 0
transform -1 0 5950 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1379_
timestamp 0
transform -1 0 6410 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1382_
timestamp 0
transform -1 0 6570 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1385_
timestamp 0
transform -1 0 6130 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1388_
timestamp 0
transform 1 0 4770 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1391_
timestamp 0
transform 1 0 4450 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1394_
timestamp 0
transform -1 0 5190 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1397_
timestamp 0
transform -1 0 6650 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1400_
timestamp 0
transform -1 0 6550 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1403_
timestamp 0
transform -1 0 5770 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1406_
timestamp 0
transform -1 0 4810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1409_
timestamp 0
transform -1 0 4730 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1412_
timestamp 0
transform 1 0 4450 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1415_
timestamp 0
transform 1 0 4610 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1418_
timestamp 0
transform 1 0 4630 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1421_
timestamp 0
transform 1 0 4270 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1424_
timestamp 0
transform 1 0 5270 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1427_
timestamp 0
transform 1 0 5090 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1430_
timestamp 0
transform 1 0 6230 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1433_
timestamp 0
transform -1 0 4350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1436_
timestamp 0
transform 1 0 4790 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1439_
timestamp 0
transform 1 0 3170 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1442_
timestamp 0
transform 1 0 5410 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1445_
timestamp 0
transform 1 0 3210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1448_
timestamp 0
transform 1 0 5010 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1451_
timestamp 0
transform 1 0 4710 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1454_
timestamp 0
transform 1 0 4210 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1456_
timestamp 0
transform -1 0 5430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1459_
timestamp 0
transform 1 0 5670 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1462_
timestamp 0
transform -1 0 5130 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1465_
timestamp 0
transform 1 0 5190 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1468_
timestamp 0
transform -1 0 6110 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1471_
timestamp 0
transform -1 0 6030 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1474_
timestamp 0
transform -1 0 6610 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1477_
timestamp 0
transform 1 0 6430 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1480_
timestamp 0
transform -1 0 6370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1483_
timestamp 0
transform -1 0 6690 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1486_
timestamp 0
transform -1 0 6350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1489_
timestamp 0
transform 1 0 4030 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1492_
timestamp 0
transform 1 0 4890 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1495_
timestamp 0
transform -1 0 5910 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1498_
timestamp 0
transform 1 0 6250 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1501_
timestamp 0
transform 1 0 4130 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1504_
timestamp 0
transform 1 0 5170 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1507_
timestamp 0
transform 1 0 4570 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1510_
timestamp 0
transform 1 0 4910 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1513_
timestamp 0
transform 1 0 5010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1516_
timestamp 0
transform 1 0 5590 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1519_
timestamp 0
transform 1 0 5390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1522_
timestamp 0
transform 1 0 5510 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1525_
timestamp 0
transform -1 0 5910 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1528_
timestamp 0
transform -1 0 4010 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1531_
timestamp 0
transform 1 0 4610 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1534_
timestamp 0
transform -1 0 4450 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1537_
timestamp 0
transform 1 0 4290 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1540_
timestamp 0
transform 1 0 5690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1543_
timestamp 0
transform 1 0 5730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1546_
timestamp 0
transform 1 0 6130 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1549_
timestamp 0
transform 1 0 6310 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1552_
timestamp 0
transform 1 0 6070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1555_
timestamp 0
transform -1 0 6090 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1558_
timestamp 0
transform 1 0 6430 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1561_
timestamp 0
transform -1 0 6630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1564_
timestamp 0
transform 1 0 6250 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1567_
timestamp 0
transform -1 0 4510 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1570_
timestamp 0
transform -1 0 3790 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1573_
timestamp 0
transform -1 0 3730 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1576_
timestamp 0
transform 1 0 5510 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1579_
timestamp 0
transform -1 0 4730 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1582_
timestamp 0
transform -1 0 2870 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1585_
timestamp 0
transform 1 0 3210 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1588_
timestamp 0
transform -1 0 2030 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1591_
timestamp 0
transform 1 0 3930 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1594_
timestamp 0
transform 1 0 3130 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1597_
timestamp 0
transform -1 0 4270 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1600_
timestamp 0
transform 1 0 3610 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1603_
timestamp 0
transform 1 0 4850 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1606_
timestamp 0
transform 1 0 1430 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1609_
timestamp 0
transform 1 0 3190 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1612_
timestamp 0
transform 1 0 1570 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1615_
timestamp 0
transform 1 0 3830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1617_
timestamp 0
transform -1 0 3650 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1620_
timestamp 0
transform 1 0 3810 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1623_
timestamp 0
transform 1 0 5010 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1626_
timestamp 0
transform 1 0 4250 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1629_
timestamp 0
transform 1 0 6290 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1632_
timestamp 0
transform 1 0 5630 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1635_
timestamp 0
transform -1 0 6510 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1638_
timestamp 0
transform 1 0 5330 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1641_
timestamp 0
transform 1 0 3390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1644_
timestamp 0
transform -1 0 3230 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1647_
timestamp 0
transform 1 0 3770 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1650_
timestamp 0
transform -1 0 3490 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1653_
timestamp 0
transform 1 0 2550 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1656_
timestamp 0
transform 1 0 1730 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1659_
timestamp 0
transform -1 0 2090 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1662_
timestamp 0
transform 1 0 2250 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1665_
timestamp 0
transform -1 0 1510 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1668_
timestamp 0
transform 1 0 2050 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1671_
timestamp 0
transform -1 0 1810 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1674_
timestamp 0
transform -1 0 110 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1677_
timestamp 0
transform 1 0 390 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1680_
timestamp 0
transform -1 0 1570 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1683_
timestamp 0
transform 1 0 2650 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1686_
timestamp 0
transform 1 0 3930 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1689_
timestamp 0
transform -1 0 3010 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1692_
timestamp 0
transform -1 0 4610 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1695_
timestamp 0
transform -1 0 3650 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1698_
timestamp 0
transform -1 0 2910 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1701_
timestamp 0
transform 1 0 2630 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1704_
timestamp 0
transform -1 0 3550 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1707_
timestamp 0
transform -1 0 3050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1710_
timestamp 0
transform 1 0 90 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1713_
timestamp 0
transform -1 0 2230 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1716_
timestamp 0
transform 1 0 1950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1719_
timestamp 0
transform -1 0 1190 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1722_
timestamp 0
transform 1 0 250 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1725_
timestamp 0
transform -1 0 110 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1728_
timestamp 0
transform -1 0 1010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1731_
timestamp 0
transform 1 0 270 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1734_
timestamp 0
transform 1 0 710 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1737_
timestamp 0
transform 1 0 710 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1740_
timestamp 0
transform -1 0 2290 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1743_
timestamp 0
transform 1 0 2870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1746_
timestamp 0
transform -1 0 2590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1749_
timestamp 0
transform -1 0 1890 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1752_
timestamp 0
transform 1 0 1870 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1755_
timestamp 0
transform -1 0 1390 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1758_
timestamp 0
transform -1 0 470 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1761_
timestamp 0
transform -1 0 1070 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1764_
timestamp 0
transform 1 0 2010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1767_
timestamp 0
transform 1 0 2570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1770_
timestamp 0
transform 1 0 2270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1773_
timestamp 0
transform 1 0 2410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1776_
timestamp 0
transform 1 0 750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1778_
timestamp 0
transform -1 0 1710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1781_
timestamp 0
transform 1 0 730 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1784_
timestamp 0
transform -1 0 650 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1787_
timestamp 0
transform 1 0 950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1790_
timestamp 0
transform -1 0 2270 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1793_
timestamp 0
transform -1 0 930 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1796_
timestamp 0
transform 1 0 650 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1799_
timestamp 0
transform 1 0 1330 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1802_
timestamp 0
transform 1 0 90 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1805_
timestamp 0
transform 1 0 210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1808_
timestamp 0
transform 1 0 490 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1811_
timestamp 0
transform -1 0 1110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1814_
timestamp 0
transform 1 0 890 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1817_
timestamp 0
transform -1 0 790 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1820_
timestamp 0
transform -1 0 1250 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1823_
timestamp 0
transform 1 0 90 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1826_
timestamp 0
transform -1 0 990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1829_
timestamp 0
transform 1 0 1630 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1832_
timestamp 0
transform -1 0 830 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1835_
timestamp 0
transform -1 0 550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1838_
timestamp 0
transform 1 0 470 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1841_
timestamp 0
transform -1 0 250 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1844_
timestamp 0
transform 1 0 1890 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1847_
timestamp 0
transform -1 0 3150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1911_
timestamp 0
transform -1 0 2750 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1914_
timestamp 0
transform -1 0 110 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1917_
timestamp 0
transform -1 0 2530 0 1 1310
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert2
timestamp 0
transform 1 0 3310 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert14
timestamp 0
transform 1 0 630 0 1 1830
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert17
timestamp 0
transform 1 0 1150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert20
timestamp 0
transform -1 0 410 0 1 2870
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert23
timestamp 0
transform 1 0 3450 0 1 3910
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert25
timestamp 0
transform -1 0 3310 0 1 3910
box -6 -8 26 268
use FILL  FILL_4_CLKBUF1_insert5
timestamp 0
transform -1 0 1070 0 1 3910
box -6 -8 26 268
use FILL  FILL_4_CLKBUF1_insert8
timestamp 0
transform -1 0 270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4_CLKBUF1_insert11
timestamp 0
transform 1 0 1730 0 1 2350
box -6 -8 26 268
<< labels >>
flabel metal1 s 6783 2 6843 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -63 2 -3 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal2 s 2657 6557 2663 6563 3 FreeSans 16 90 0 0 Cin[7]
port 2 nsew
flabel metal2 s 2997 6557 3003 6563 3 FreeSans 16 90 0 0 Cin[6]
port 3 nsew
flabel metal2 s 2837 6557 2843 6563 3 FreeSans 16 90 0 0 Cin[5]
port 4 nsew
flabel metal2 s 3297 6557 3303 6563 3 FreeSans 16 90 0 0 Cin[4]
port 5 nsew
flabel metal2 s 4457 -23 4463 -17 7 FreeSans 16 270 0 0 Cin[3]
port 6 nsew
flabel metal2 s 2557 -23 2563 -17 7 FreeSans 16 270 0 0 Cin[2]
port 7 nsew
flabel metal3 s -24 1176 -16 1184 7 FreeSans 16 0 0 0 Cin[1]
port 8 nsew
flabel metal3 s -24 1436 -16 1444 7 FreeSans 16 0 0 0 Cin[0]
port 9 nsew
flabel metal3 s -24 2736 -16 2744 7 FreeSans 16 0 0 0 Rdy
port 10 nsew
flabel metal2 s 2777 -23 2783 -17 7 FreeSans 16 270 0 0 Vld
port 11 nsew
flabel metal3 s -24 2476 -16 2484 7 FreeSans 16 0 0 0 Xin[3]
port 12 nsew
flabel metal2 s 3017 -23 3023 -17 7 FreeSans 16 270 0 0 Xin[2]
port 13 nsew
flabel metal2 s 1937 -23 1943 -17 7 FreeSans 16 270 0 0 Xin[1]
port 14 nsew
flabel metal3 s -24 1956 -16 1964 7 FreeSans 16 0 0 0 Xin[0]
port 15 nsew
flabel metal3 s -24 3516 -16 3524 7 FreeSans 16 0 0 0 Xout[3]
port 16 nsew
flabel metal3 s -24 3036 -16 3044 7 FreeSans 16 0 0 0 Xout[2]
port 17 nsew
flabel metal2 s 2477 -23 2483 -17 7 FreeSans 16 270 0 0 Xout[1]
port 18 nsew
flabel metal3 s -24 1696 -16 1704 7 FreeSans 16 0 0 0 Xout[0]
port 19 nsew
flabel metal3 s -24 1996 -16 2004 7 FreeSans 16 0 0 0 Yin[3]
port 20 nsew
flabel metal3 s -24 4556 -16 4564 7 FreeSans 16 0 0 0 Yin[2]
port 21 nsew
flabel metal3 s -24 4856 -16 4864 7 FreeSans 16 0 0 0 Yin[1]
port 22 nsew
flabel metal3 s -24 2216 -16 2224 7 FreeSans 16 0 0 0 Yin[0]
port 23 nsew
flabel metal3 s -24 3256 -16 3264 7 FreeSans 16 0 0 0 Yout[3]
port 24 nsew
flabel metal3 s -24 2996 -16 3004 7 FreeSans 16 0 0 0 Yout[2]
port 25 nsew
flabel metal2 s 2437 -23 2443 -17 7 FreeSans 16 270 0 0 Yout[1]
port 26 nsew
flabel metal2 s 2617 -23 2623 -17 7 FreeSans 16 270 0 0 Yout[0]
port 27 nsew
flabel metal3 s -24 3296 -16 3304 7 FreeSans 16 0 0 0 clk
port 28 nsew
<< properties >>
string FIXED_BBOX -40 -40 6780 6560
<< end >>

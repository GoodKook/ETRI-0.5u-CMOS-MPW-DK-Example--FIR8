* NGSPICE file created from fir_pe.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL vdd gnd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A Y vdd gnd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B Y vdd gnd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 D CLK Q vdd gnd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A Y vdd gnd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D Y vdd gnd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D Y vdd gnd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A Y vdd gnd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A Y vdd gnd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B Y vdd gnd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A Y vdd gnd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A Y vdd gnd
.ends

.subckt fir_pe gnd vdd Cin[7] Cin[6] Cin[5] Cin[4] Cin[3] Cin[2] Cin[1] Cin[0] Rdy
+ Vld Xin[3] Xin[2] Xin[1] Xin[0] Xout[3] Xout[2] Xout[1] Xout[0] Yin[3] Yin[2] Yin[1]
+ Yin[0] Yout[3] Yout[2] Yout[1] Yout[0] clk
XFILL_1__1670_ vdd gnd FILL
XFILL_3__1537_ vdd gnd FILL
XFILL_3__1606_ vdd gnd FILL
XFILL_0__1759_ vdd gnd FILL
XFILL_3__1468_ vdd gnd FILL
XFILL_0__1828_ vdd gnd FILL
XFILL_2__992_ vdd gnd FILL
XFILL_3__1399_ vdd gnd FILL
XFILL_1__1104_ vdd gnd FILL
XFILL_1__1035_ vdd gnd FILL
XFILL_1__1799_ vdd gnd FILL
XFILL_2__1213_ vdd gnd FILL
XFILL100050x150 vdd gnd FILL
XFILL_2__1144_ vdd gnd FILL
XFILL_2__1075_ vdd gnd FILL
XFILL_0_CLKBUF1_insert6 vdd gnd FILL
XFILL_0__1544_ vdd gnd FILL
XFILL_0__1613_ vdd gnd FILL
XFILL_3__957_ vdd gnd FILL
XFILL_3__1322_ vdd gnd FILL
X_1270_ _1274_/A _1274_/B _1371_/C _1280_/A vdd gnd OAI21X1
XFILL_0__1475_ vdd gnd FILL
XFILL_3__1184_ vdd gnd FILL
XFILL_3__1253_ vdd gnd FILL
X_1606_ _1892_/Q _1822_/A vdd gnd INVX1
XFILL_1__1653_ vdd gnd FILL
X_1537_ _1539_/A _1538_/A vdd gnd INVX1
XFILL_1__1722_ vdd gnd FILL
X_1468_ _1468_/A _1495_/B _1498_/A vdd gnd AND2X2
X_1399_ _1399_/A _1399_/B _1494_/A vdd gnd NAND2X1
XFILL_1__1584_ vdd gnd FILL
XFILL_4__1293_ vdd gnd FILL
XFILL_2__975_ vdd gnd FILL
XFILL_2__1762_ vdd gnd FILL
XFILL_2__1831_ vdd gnd FILL
XFILL_1__1018_ vdd gnd FILL
X_981_ _981_/A _983_/B vdd gnd INVX1
XFILL_4__1629_ vdd gnd FILL
XFILL_2__1693_ vdd gnd FILL
XFILL_0__1260_ vdd gnd FILL
XFILL_0__1191_ vdd gnd FILL
XFILL_2__1127_ vdd gnd FILL
XFILL_2__1058_ vdd gnd FILL
XFILL_1__993_ vdd gnd FILL
X_1322_ _1322_/A _1399_/A _1322_/C _1399_/B vdd gnd NAND3X1
XFILL99750x15750 vdd gnd FILL
X_1253_ _1360_/B _1360_/A _1263_/C _1269_/B vdd gnd NAND3X1
XFILL_0__1527_ vdd gnd FILL
XFILL_3__1305_ vdd gnd FILL
XFILL_3__1236_ vdd gnd FILL
X_1184_ _1184_/A _1243_/C _1184_/C _1193_/A vdd gnd AOI21X1
XFILL_0__1458_ vdd gnd FILL
XFILL_0__1389_ vdd gnd FILL
XFILL_3__1098_ vdd gnd FILL
XFILL_3__1167_ vdd gnd FILL
XFILL_1__1636_ vdd gnd FILL
XFILL_1__1705_ vdd gnd FILL
XFILL101250x85950 vdd gnd FILL
XFILL_1__1498_ vdd gnd FILL
XFILL_1__1567_ vdd gnd FILL
XFILL_2__958_ vdd gnd FILL
XFILL_2__1745_ vdd gnd FILL
XFILL_2__1814_ vdd gnd FILL
X_964_ Xin[3] _965_/B _965_/C vdd gnd NAND2X1
XFILL_2__1676_ vdd gnd FILL
X_1871_ _1871_/D _1910_/CLK _970_/B vdd gnd DFFPOSX1
XFILL_0__1312_ vdd gnd FILL
XFILL_0__1174_ vdd gnd FILL
XFILL_0__1243_ vdd gnd FILL
XFILL_3__1021_ vdd gnd FILL
XFILL_3__1785_ vdd gnd FILL
X_1305_ _1311_/C _1424_/A _1403_/B vdd gnd NAND2X1
XFILL_1__976_ vdd gnd FILL
X_1236_ _1317_/C _1313_/B _1313_/A _1261_/A vdd gnd OAI21X1
XFILL_1__1352_ vdd gnd FILL
XFILL_1__1421_ vdd gnd FILL
XBUFX2_insert0 _1910_/Q _983_/A vdd gnd BUFX2
X_1098_ _1216_/A _1098_/B _1098_/C _1873_/D vdd gnd OAI21X1
XFILL_1__1283_ vdd gnd FILL
XFILL_3__1219_ vdd gnd FILL
X_1167_ _1168_/A _1167_/B _1167_/C _1191_/A vdd gnd NAND3X1
XFILL_1__1619_ vdd gnd FILL
XFILL_2__1530_ vdd gnd FILL
XFILL_2__1461_ vdd gnd FILL
XFILL_4__1328_ vdd gnd FILL
XFILL_2__1392_ vdd gnd FILL
XFILL_0__994_ vdd gnd FILL
XFILL_2__1659_ vdd gnd FILL
XFILL_2__1728_ vdd gnd FILL
XFILL_0__1792_ vdd gnd FILL
XFILL_3__1570_ vdd gnd FILL
X_947_ _951_/A _947_/B _948_/C vdd gnd NAND2X1
X_1021_ _1036_/C _1023_/B vdd gnd INVX1
X_1785_ _1793_/A _1793_/B _1785_/C _1792_/B vdd gnd OAI21X1
XFILL_3__1004_ vdd gnd FILL
X_1854_ _968_/Y _1904_/CLK _966_/A vdd gnd DFFPOSX1
XFILL_0__1226_ vdd gnd FILL
XFILL_0__1157_ vdd gnd FILL
XFILL_3__1768_ vdd gnd FILL
XFILL_3__1837_ vdd gnd FILL
XFILL_0__1088_ vdd gnd FILL
XFILL_3__1699_ vdd gnd FILL
XFILL_1__1404_ vdd gnd FILL
XFILL_1__959_ vdd gnd FILL
X_1219_ _1224_/B _1219_/B _1383_/A vdd gnd NAND2X1
XFILL_1__1335_ vdd gnd FILL
XFILL_1__1266_ vdd gnd FILL
XFILL_3__990_ vdd gnd FILL
XFILL_1__1197_ vdd gnd FILL
XFILL_2__1513_ vdd gnd FILL
XFILL_2__1444_ vdd gnd FILL
XFILL_2__1375_ vdd gnd FILL
XFILL_0__977_ vdd gnd FILL
XFILL_0__1011_ vdd gnd FILL
XFILL_3__1622_ vdd gnd FILL
X_1570_ _995_/B _1702_/B _1642_/C vdd gnd NAND2X1
XFILL_0__1913_ vdd gnd FILL
XFILL_3__1553_ vdd gnd FILL
XFILL_0__1775_ vdd gnd FILL
XFILL_3__1484_ vdd gnd FILL
XFILL_0__1844_ vdd gnd FILL
XFILL_4__955_ vdd gnd FILL
X_1004_ _1801_/A _1769_/B _1004_/C _1867_/D vdd gnd OAI21X1
XFILL_1__1120_ vdd gnd FILL
XFILL_4__1731_ vdd gnd FILL
X_1768_ _1768_/A _1773_/A _1790_/A _1769_/C vdd gnd AOI21X1
X_1906_ Rdy _1908_/CLK _1906_/Q vdd gnd DFFPOSX1
X_1837_ _1848_/A _1837_/B _1837_/C _1899_/D vdd gnd AOI21X1
XFILL_0__1209_ vdd gnd FILL
XFILL_1__1051_ vdd gnd FILL
XFILL_4__1662_ vdd gnd FILL
X_1699_ _1703_/A _1699_/B _1700_/A vdd gnd NOR2X1
XFILL_2__1160_ vdd gnd FILL
XFILL_1__1318_ vdd gnd FILL
XFILL_4__1027_ vdd gnd FILL
XFILL_2__1091_ vdd gnd FILL
XFILL_1__1249_ vdd gnd FILL
XFILL_3__973_ vdd gnd FILL
XFILL_0__1560_ vdd gnd FILL
XFILL_0__1491_ vdd gnd FILL
XFILL_2__1427_ vdd gnd FILL
XFILL_2__1358_ vdd gnd FILL
XFILL_2__1289_ vdd gnd FILL
X_1622_ _1622_/A _1622_/B _1626_/C vdd gnd NAND2X1
X_1553_ _1553_/A _1576_/B _1578_/B _1625_/C _1634_/A vdd gnd AOI22X1
XFILL_3__1605_ vdd gnd FILL
XFILL_2_BUFX2_insert25 vdd gnd FILL
XFILL_2_BUFX2_insert14 vdd gnd FILL
X_1484_ _1484_/A _1484_/B _1484_/C _1487_/C vdd gnd AOI21X1
XFILL_0__1689_ vdd gnd FILL
XFILL_3__1536_ vdd gnd FILL
XFILL_0__1758_ vdd gnd FILL
XFILL_3__1467_ vdd gnd FILL
XFILL_3__1398_ vdd gnd FILL
XFILL_0__1827_ vdd gnd FILL
XFILL_2__991_ vdd gnd FILL
XFILL_1__1103_ vdd gnd FILL
XFILL_1__1034_ vdd gnd FILL
XFILL_4__1576_ vdd gnd FILL
XFILL_1__1798_ vdd gnd FILL
XFILL_1_BUFX2_insert0 vdd gnd FILL
XFILL_2__1212_ vdd gnd FILL
XFILL_2__1143_ vdd gnd FILL
XFILL_0_CLKBUF1_insert7 vdd gnd FILL
XFILL_2__1074_ vdd gnd FILL
XFILL_3__956_ vdd gnd FILL
XFILL_0__1612_ vdd gnd FILL
XFILL_0__1543_ vdd gnd FILL
XFILL_3__1321_ vdd gnd FILL
XFILL_3__1252_ vdd gnd FILL
XFILL_0__1474_ vdd gnd FILL
XFILL_3__1183_ vdd gnd FILL
X_1536_ _1605_/B _1891_/Q _1539_/A vdd gnd XNOR2X1
X_1605_ _1820_/A _1605_/B _1620_/B _1621_/B vdd gnd OAI21X1
XFILL_1__1652_ vdd gnd FILL
XFILL_1__1583_ vdd gnd FILL
XFILL_1__1721_ vdd gnd FILL
X_1467_ _1552_/A _1476_/B _1476_/A _1479_/A vdd gnd NAND3X1
X_1398_ _1398_/A _1398_/B _1483_/A _1482_/C vdd gnd OAI21X1
XFILL_4__1430_ vdd gnd FILL
XFILL_4__1361_ vdd gnd FILL
XFILL_3__1519_ vdd gnd FILL
XFILL_1__1017_ vdd gnd FILL
XFILL_2__974_ vdd gnd FILL
XFILL_2__1692_ vdd gnd FILL
XFILL_2__1761_ vdd gnd FILL
XFILL_1__1919_ vdd gnd FILL
X_980_ _996_/A _980_/B _980_/C _980_/Y vdd gnd OAI21X1
XFILL_2__1830_ vdd gnd FILL
XFILL_0__1190_ vdd gnd FILL
XFILL_2__1126_ vdd gnd FILL
XFILL_2__1057_ vdd gnd FILL
XFILL_1__992_ vdd gnd FILL
XFILL_3__939_ vdd gnd FILL
X_1321_ _1321_/A _1321_/B _1321_/C _1322_/C vdd gnd OAI21X1
X_1252_ _1254_/C _1338_/C _1254_/A _1360_/B vdd gnd NAND3X1
XFILL_0__1526_ vdd gnd FILL
XFILL_0__1457_ vdd gnd FILL
XFILL_3__1304_ vdd gnd FILL
XFILL_3__1235_ vdd gnd FILL
X_1183_ _1266_/B _1266_/A _1193_/C _1198_/B vdd gnd NAND3X1
XFILL_0__1388_ vdd gnd FILL
XFILL_3__1097_ vdd gnd FILL
XFILL_3__1166_ vdd gnd FILL
X_1519_ _1519_/A _1519_/B _1519_/C _1522_/A vdd gnd OAI21X1
XFILL_1__1635_ vdd gnd FILL
XFILL_1__1566_ vdd gnd FILL
XFILL_1__1704_ vdd gnd FILL
XFILL_4__1275_ vdd gnd FILL
XFILL_1__1497_ vdd gnd FILL
XFILL_2__957_ vdd gnd FILL
XFILL_2__1675_ vdd gnd FILL
XFILL_2__1744_ vdd gnd FILL
XFILL_2__1813_ vdd gnd FILL
X_963_ _963_/A _965_/B _963_/C _963_/Y vdd gnd OAI21X1
XFILL_0__1311_ vdd gnd FILL
XFILL_3__1020_ vdd gnd FILL
X_1870_ _1870_/D _1903_/CLK _967_/A vdd gnd DFFPOSX1
XFILL_0__1242_ vdd gnd FILL
XFILL_2__1109_ vdd gnd FILL
XFILL_0__1173_ vdd gnd FILL
XFILL_3__1784_ vdd gnd FILL
XFILL_1__1420_ vdd gnd FILL
X_1304_ _953_/B Cin[5] _1424_/A vdd gnd AND2X2
XFILL_1__975_ vdd gnd FILL
XBUFX2_insert1 _1910_/Q _977_/A vdd gnd BUFX2
X_1235_ _1240_/C _1235_/B _1313_/B vdd gnd AND2X2
X_1166_ _1847_/B _1533_/B _1239_/A _1167_/C vdd gnd OAI21X1
XFILL_0__1509_ vdd gnd FILL
XFILL_1__1351_ vdd gnd FILL
XFILL_1__1282_ vdd gnd FILL
XFILL_3__1218_ vdd gnd FILL
X_1097_ _1097_/A _1097_/B _1098_/B vdd gnd NAND2X1
XFILL_3__1149_ vdd gnd FILL
XFILL_4__1060_ vdd gnd FILL
XFILL_1__1618_ vdd gnd FILL
XFILL_1__1549_ vdd gnd FILL
XFILL_2__1460_ vdd gnd FILL
XFILL_2__1391_ vdd gnd FILL
XFILL_0__993_ vdd gnd FILL
XFILL_2__1727_ vdd gnd FILL
XFILL_2__1658_ vdd gnd FILL
XFILL_0__1791_ vdd gnd FILL
X_1020_ _950_/B _1106_/B _1899_/Q _1036_/C vdd gnd NAND3X1
X_946_ _946_/A _959_/A vdd gnd INVX1
XFILL_2__1589_ vdd gnd FILL
XFILL_3__1003_ vdd gnd FILL
X_1784_ _1793_/A _1784_/B _1785_/C vdd gnd NAND2X1
X_1853_ _965_/Y _1910_/CLK _955_/A vdd gnd DFFPOSX1
XFILL_0__1156_ vdd gnd FILL
XFILL_0__1225_ vdd gnd FILL
XFILL_0__1087_ vdd gnd FILL
XFILL_3__1767_ vdd gnd FILL
XFILL_3__1836_ vdd gnd FILL
XFILL_3__1698_ vdd gnd FILL
XFILL_1__1403_ vdd gnd FILL
XFILL_1__958_ vdd gnd FILL
X_1218_ _1290_/C _1287_/A vdd gnd INVX1
X_1149_ _1153_/A _1149_/B _1149_/C _1217_/B vdd gnd NAND3X1
XFILL_1__1334_ vdd gnd FILL
XFILL_1__1196_ vdd gnd FILL
XFILL_1__1265_ vdd gnd FILL
XFILL_2__1512_ vdd gnd FILL
XFILL_2__1443_ vdd gnd FILL
XFILL_2__1374_ vdd gnd FILL
XFILL_0__1010_ vdd gnd FILL
XFILL_0__976_ vdd gnd FILL
XFILL_3__1621_ vdd gnd FILL
XFILL_3__1552_ vdd gnd FILL
XFILL_0__1843_ vdd gnd FILL
XFILL_0__1912_ vdd gnd FILL
XFILL_3__1483_ vdd gnd FILL
XFILL_0__1774_ vdd gnd FILL
X_1003_ _933_/B _1790_/A _1004_/C vdd gnd NAND2X1
X_929_ _944_/A _966_/A _965_/B _978_/A _930_/C vdd gnd AOI22X1
X_1905_ _1905_/D _1908_/CLK _956_/B vdd gnd DFFPOSX1
XFILL_1__1050_ vdd gnd FILL
X_1767_ _1773_/B _1767_/B _1768_/A vdd gnd NOR2X1
X_1698_ _1699_/B _1703_/A _1700_/B vdd gnd AND2X2
X_1836_ _1848_/A _1899_/Q _1837_/C vdd gnd NOR2X1
XFILL_0__1208_ vdd gnd FILL
XFILL_0__1139_ vdd gnd FILL
XFILL_3__1819_ vdd gnd FILL
XFILL_1__1317_ vdd gnd FILL
XFILL_1__1248_ vdd gnd FILL
XFILL_2__1090_ vdd gnd FILL
XFILL_1__1179_ vdd gnd FILL
XFILL_3__972_ vdd gnd FILL
XFILL_0__1490_ vdd gnd FILL
XFILL_2__1426_ vdd gnd FILL
XFILL_2__1357_ vdd gnd FILL
XFILL_2__1288_ vdd gnd FILL
X_1621_ _1621_/A _1621_/B _1622_/B vdd gnd NAND2X1
X_1552_ _1552_/A _1552_/B _1552_/C _1574_/C vdd gnd OAI21X1
XFILL_2_BUFX2_insert15 vdd gnd FILL
XFILL_0__959_ vdd gnd FILL
X_1483_ _1483_/A _1484_/C vdd gnd INVX1
XFILL_3__1535_ vdd gnd FILL
XFILL_3__1604_ vdd gnd FILL
XFILL_0__1826_ vdd gnd FILL
XFILL_0__1688_ vdd gnd FILL
XFILL_0__1757_ vdd gnd FILL
XFILL_3__1466_ vdd gnd FILL
XFILL_2__990_ vdd gnd FILL
XFILL_3__1397_ vdd gnd FILL
XFILL_4__937_ vdd gnd FILL
XFILL_1__1102_ vdd gnd FILL
XFILL_1__1033_ vdd gnd FILL
XFILL_4__1713_ vdd gnd FILL
X_1819_ Yin[1] _1824_/B _1820_/C vdd gnd NAND2X1
XFILL_4__1644_ vdd gnd FILL
XFILL_1__1797_ vdd gnd FILL
XFILL_1_BUFX2_insert1 vdd gnd FILL
XFILL_4__1009_ vdd gnd FILL
XFILL_2__1142_ vdd gnd FILL
XFILL_2__1073_ vdd gnd FILL
XFILL_2__1211_ vdd gnd FILL
XFILL_0_CLKBUF1_insert8 vdd gnd FILL
XFILL100050x15750 vdd gnd FILL
XFILL_3__955_ vdd gnd FILL
XFILL_0__1611_ vdd gnd FILL
XFILL_0__1542_ vdd gnd FILL
XFILL_2__1409_ vdd gnd FILL
XFILL_0__1473_ vdd gnd FILL
XFILL_3__1320_ vdd gnd FILL
XFILL_3__1182_ vdd gnd FILL
XFILL_3__1251_ vdd gnd FILL
XFILL_1__1720_ vdd gnd FILL
X_1535_ _1539_/B _1539_/C _1538_/B vdd gnd NAND2X1
X_1604_ _1891_/Q _1820_/A vdd gnd INVX1
XFILL_1__1651_ vdd gnd FILL
XFILL_1__1582_ vdd gnd FILL
X_1466_ _1555_/B _1470_/B _1551_/C _1476_/A vdd gnd OAI21X1
XFILL_0__1809_ vdd gnd FILL
XFILL_3__1518_ vdd gnd FILL
X_1397_ _1397_/A _1397_/B _1397_/C _1398_/B vdd gnd AOI21X1
XFILL_3__1449_ vdd gnd FILL
XFILL_2__973_ vdd gnd FILL
XFILL_1__1016_ vdd gnd FILL
XFILL_2__1691_ vdd gnd FILL
XFILL_2__1760_ vdd gnd FILL
XFILL_1__1918_ vdd gnd FILL
XFILL_1__1849_ vdd gnd FILL
XFILL_4__1558_ vdd gnd FILL
XFILL_4__1489_ vdd gnd FILL
XFILL_2__1125_ vdd gnd FILL
XFILL_2__1056_ vdd gnd FILL
XFILL100650x74250 vdd gnd FILL
X_1320_ _1425_/C _1320_/B _1320_/C _1399_/A vdd gnd NAND3X1
XFILL_1__991_ vdd gnd FILL
XFILL_3__938_ vdd gnd FILL
X_1182_ _1184_/C _1243_/C _1184_/A _1266_/B vdd gnd NAND3X1
X_1251_ _1338_/B _1254_/A vdd gnd INVX1
XFILL_0__1525_ vdd gnd FILL
XFILL_0__1456_ vdd gnd FILL
XFILL_3__1303_ vdd gnd FILL
XFILL_3__1234_ vdd gnd FILL
XFILL_3__1165_ vdd gnd FILL
XFILL_3__1096_ vdd gnd FILL
XFILL_0__1387_ vdd gnd FILL
XFILL_1__1703_ vdd gnd FILL
X_1518_ _956_/B Cin[6] _1519_/B vdd gnd NAND2X1
X_1449_ _955_/A _1449_/B _1897_/Q _1450_/B vdd gnd AOI21X1
XFILL_4__1412_ vdd gnd FILL
XFILL_1__1634_ vdd gnd FILL
XFILL_1__1496_ vdd gnd FILL
XFILL_1__1565_ vdd gnd FILL
XFILL_4__1343_ vdd gnd FILL
XFILL_2__956_ vdd gnd FILL
XFILL_2__1812_ vdd gnd FILL
XFILL_2__1674_ vdd gnd FILL
XFILL_2__1743_ vdd gnd FILL
X_962_ Xin[2] _965_/B _963_/C vdd gnd NAND2X1
XFILL100050x39150 vdd gnd FILL
XFILL_0__1310_ vdd gnd FILL
XFILL_0__1241_ vdd gnd FILL
XFILL_2__1108_ vdd gnd FILL
XFILL_0__1172_ vdd gnd FILL
XFILL_2__1039_ vdd gnd FILL
XFILL_3__1783_ vdd gnd FILL
X_1303_ _1315_/A _1316_/B vdd gnd INVX1
XFILL_1__974_ vdd gnd FILL
XFILL_1__1350_ vdd gnd FILL
XBUFX2_insert2 _1910_/Q _992_/A vdd gnd BUFX2
X_1234_ _1240_/C _1235_/B _1317_/C vdd gnd NOR2X1
X_1096_ _1149_/B _1097_/B vdd gnd INVX1
X_1165_ _956_/B Cin[2] _1239_/A vdd gnd AND2X2
XFILL_0__1508_ vdd gnd FILL
XFILL_0__1439_ vdd gnd FILL
XFILL_1__1281_ vdd gnd FILL
XFILL_3__1217_ vdd gnd FILL
XFILL_3__1148_ vdd gnd FILL
XFILL_3__1079_ vdd gnd FILL
XFILL_1__1548_ vdd gnd FILL
XFILL_1__1617_ vdd gnd FILL
XFILL_1__1479_ vdd gnd FILL
XFILL_4__1257_ vdd gnd FILL
XFILL_2__1390_ vdd gnd FILL
XFILL_4__1188_ vdd gnd FILL
XFILL_0__992_ vdd gnd FILL
XFILL_2__939_ vdd gnd FILL
X_945_ _945_/A _945_/B _945_/C _945_/Y vdd gnd OAI21X1
XFILL99750x150 vdd gnd FILL
XFILL_2__1726_ vdd gnd FILL
XFILL_2__1588_ vdd gnd FILL
XFILL_2__1657_ vdd gnd FILL
XFILL_0__1790_ vdd gnd FILL
XFILL_3__1002_ vdd gnd FILL
XFILL_4__970_ vdd gnd FILL
XFILL_0__1224_ vdd gnd FILL
X_1852_ _963_/Y _1904_/CLK _952_/A vdd gnd DFFPOSX1
X_1783_ _1783_/A _1793_/C _1784_/B vdd gnd NAND2X1
XFILL_0__1155_ vdd gnd FILL
XFILL_3__1835_ vdd gnd FILL
XFILL_0__1086_ vdd gnd FILL
XFILL_3__1697_ vdd gnd FILL
XFILL_3__1766_ vdd gnd FILL
XFILL_1__957_ vdd gnd FILL
XFILL_1__1333_ vdd gnd FILL
XFILL_1__1402_ vdd gnd FILL
XFILL_4__1111_ vdd gnd FILL
X_1079_ _1079_/A _1079_/B _1082_/A _1101_/B vdd gnd AOI21X1
X_1217_ _1217_/A _1217_/B _1217_/C _1292_/B vdd gnd OAI21X1
XFILL_4__1042_ vdd gnd FILL
X_1148_ _1149_/C _1153_/A _1149_/B _1151_/A vdd gnd AOI21X1
XFILL_1__1195_ vdd gnd FILL
XFILL_1__1264_ vdd gnd FILL
XFILL_2__1442_ vdd gnd FILL
XFILL_2__1511_ vdd gnd FILL
XFILL_2__1373_ vdd gnd FILL
XFILL_0__975_ vdd gnd FILL
XFILL_2__1709_ vdd gnd FILL
XFILL_3__1620_ vdd gnd FILL
XFILL_0__1773_ vdd gnd FILL
XFILL_3__1551_ vdd gnd FILL
X_928_ _944_/A _928_/B _965_/B vdd gnd NOR2X1
XFILL_0__1842_ vdd gnd FILL
XFILL_0__1911_ vdd gnd FILL
X_1002_ _1883_/Q _1769_/B vdd gnd INVX1
XFILL_3__1482_ vdd gnd FILL
X_1835_ _1848_/A _1835_/B _1835_/C _1898_/D vdd gnd OAI21X1
XFILL_0__1207_ vdd gnd FILL
X_1904_ _1904_/D _1904_/CLK _953_/B vdd gnd DFFPOSX1
XFILL_4__1591_ vdd gnd FILL
X_1697_ _1705_/A _1706_/A _1703_/A vdd gnd NAND2X1
X_1766_ _1773_/B _1767_/B _1766_/C _1769_/D vdd gnd OAI21X1
XFILL_3__1818_ vdd gnd FILL
XFILL_0__1138_ vdd gnd FILL
XFILL_0__1069_ vdd gnd FILL
XFILL_3__1749_ vdd gnd FILL
XFILL_1__1316_ vdd gnd FILL
XFILL_1__1178_ vdd gnd FILL
XFILL_1__1247_ vdd gnd FILL
XFILL_3__971_ vdd gnd FILL
XFILL_2__1356_ vdd gnd FILL
XFILL_2__1425_ vdd gnd FILL
XFILL_0__958_ vdd gnd FILL
XFILL_2__1287_ vdd gnd FILL
X_1620_ _1620_/A _1620_/B _1620_/C _1622_/A vdd gnd NAND3X1
X_1551_ _1551_/A _1551_/B _1551_/C _1552_/B vdd gnd AOI21X1
X_1482_ _1482_/A _1482_/B _1482_/C _1571_/A vdd gnd NAND3X1
XFILL_2_BUFX2_insert16 vdd gnd FILL
XFILL_3__1603_ vdd gnd FILL
XFILL_3__1534_ vdd gnd FILL
XFILL_0__1756_ vdd gnd FILL
XFILL_3__1465_ vdd gnd FILL
XFILL_0__1825_ vdd gnd FILL
XFILL_0__1687_ vdd gnd FILL
XFILL_1__1101_ vdd gnd FILL
XFILL_3__1396_ vdd gnd FILL
X_1818_ _1827_/A _1824_/B _1818_/C _1890_/D vdd gnd AOI21X1
XFILL_1__1032_ vdd gnd FILL
X_1749_ _1749_/A _1751_/C _1749_/C _1749_/D _1777_/A vdd gnd OAI22X1
XFILL_1__1796_ vdd gnd FILL
XFILL_1_BUFX2_insert2 vdd gnd FILL
XFILL_2__1210_ vdd gnd FILL
XFILL_2__1141_ vdd gnd FILL
XFILL_2__1072_ vdd gnd FILL
XFILL100950x46950 vdd gnd FILL
XFILL_0_CLKBUF1_insert9 vdd gnd FILL
XFILL_0__1610_ vdd gnd FILL
XFILL_3__954_ vdd gnd FILL
XFILL_0__1541_ vdd gnd FILL
XFILL_0__1472_ vdd gnd FILL
XFILL_2__1339_ vdd gnd FILL
XFILL_2__1408_ vdd gnd FILL
XFILL_3__1181_ vdd gnd FILL
XFILL_3__1250_ vdd gnd FILL
X_1603_ _1649_/B _1649_/A _1687_/A vdd gnd NAND2X1
X_1534_ _1597_/A _1597_/B _1592_/C _1539_/B vdd gnd NAND3X1
X_1465_ _1465_/A _1465_/B _1543_/A _1555_/B vdd gnd AOI21X1
XFILL_1__1650_ vdd gnd FILL
XFILL_0__1739_ vdd gnd FILL
XFILL_3__1517_ vdd gnd FILL
XFILL_1__1581_ vdd gnd FILL
XFILL_3__1448_ vdd gnd FILL
XFILL_0__1808_ vdd gnd FILL
XFILL_4__1290_ vdd gnd FILL
X_1396_ _1396_/A _1396_/B _1396_/C _1396_/D _1704_/C vdd gnd OAI22X1
XFILL_2__972_ vdd gnd FILL
XFILL_3__1379_ vdd gnd FILL
XFILL_1__1015_ vdd gnd FILL
XFILL_2__1690_ vdd gnd FILL
XFILL_4__1626_ vdd gnd FILL
XFILL_1__1779_ vdd gnd FILL
XFILL_1__1848_ vdd gnd FILL
XFILL_1__1917_ vdd gnd FILL
XFILL100950x58650 vdd gnd FILL
XFILL_2__1055_ vdd gnd FILL
XFILL_2__1124_ vdd gnd FILL
XFILL_1__990_ vdd gnd FILL
XFILL_0__1524_ vdd gnd FILL
XFILL_3__937_ vdd gnd FILL
XFILL_3__1302_ vdd gnd FILL
X_1181_ _1243_/B _1184_/A vdd gnd INVX1
X_1250_ _1338_/A _1254_/C vdd gnd INVX1
XFILL_0__1455_ vdd gnd FILL
XFILL_3__1233_ vdd gnd FILL
XFILL_3__1095_ vdd gnd FILL
XFILL_0__1386_ vdd gnd FILL
XFILL_3__1164_ vdd gnd FILL
XFILL_1__1633_ vdd gnd FILL
X_1517_ _1517_/A _1517_/B _1517_/C _1553_/A vdd gnd NAND3X1
X_1448_ _1524_/A _1524_/B _1542_/B _1465_/A vdd gnd NAND3X1
XFILL_1__1702_ vdd gnd FILL
XFILL_1__1564_ vdd gnd FILL
XFILL_1__1495_ vdd gnd FILL
X_1379_ _1379_/A _1379_/B _1379_/C _1484_/B vdd gnd OAI21X1
XFILL_2__955_ vdd gnd FILL
XFILL_2__1742_ vdd gnd FILL
XFILL_2__1811_ vdd gnd FILL
X_961_ _961_/A _965_/B _961_/C _961_/Y vdd gnd OAI21X1
XFILL_4__1609_ vdd gnd FILL
XFILL_2__1673_ vdd gnd FILL
XFILL_0__1240_ vdd gnd FILL
XFILL_2__1107_ vdd gnd FILL
XFILL_0__1171_ vdd gnd FILL
XFILL_2__1038_ vdd gnd FILL
XFILL_3__1782_ vdd gnd FILL
X_1302_ _947_/B Cin[7] _1315_/A vdd gnd NAND2X1
X_1233_ _946_/A Cin[2] _1235_/B vdd gnd NAND2X1
XFILL_1__973_ vdd gnd FILL
XFILL_0__1507_ vdd gnd FILL
XBUFX2_insert3 _1910_/Q _996_/A vdd gnd BUFX2
XFILL_1__1280_ vdd gnd FILL
X_1095_ _1213_/B _1095_/B _1095_/C _1149_/B vdd gnd NOR3X1
X_1164_ _1849_/B _1533_/D _1169_/A _1167_/B vdd gnd OAI21X1
XFILL_0__1438_ vdd gnd FILL
XFILL_0__1369_ vdd gnd FILL
XFILL_3__1078_ vdd gnd FILL
XFILL_3__1147_ vdd gnd FILL
XFILL_3__1216_ vdd gnd FILL
XFILL_1__1616_ vdd gnd FILL
XFILL_4__1325_ vdd gnd FILL
XFILL_1__1547_ vdd gnd FILL
XFILL_1__1478_ vdd gnd FILL
XFILL_0__991_ vdd gnd FILL
XFILL_2__938_ vdd gnd FILL
XFILL_2__1725_ vdd gnd FILL
X_944_ _944_/A _975_/A _965_/B _989_/A _945_/C vdd gnd AOI22X1
XFILL_2__1587_ vdd gnd FILL
XFILL_2__1656_ vdd gnd FILL
XFILL_3__1001_ vdd gnd FILL
XFILL_0__1223_ vdd gnd FILL
XFILL_0__1154_ vdd gnd FILL
X_1851_ _961_/Y _1904_/CLK _949_/A vdd gnd DFFPOSX1
X_1782_ _1793_/B _1782_/B _1783_/A vdd gnd NAND2X1
XFILL_3__1834_ vdd gnd FILL
XFILL_0__1085_ vdd gnd FILL
XFILL_3__1696_ vdd gnd FILL
XFILL_3__1765_ vdd gnd FILL
XFILL_1__956_ vdd gnd FILL
X_1216_ _1216_/A _1216_/B _1216_/C _1875_/D vdd gnd OAI21X1
XFILL_1__1332_ vdd gnd FILL
XFILL_1__1401_ vdd gnd FILL
X_1078_ _1138_/A _1140_/C vdd gnd INVX1
X_1147_ _1147_/A _1147_/B _1149_/C vdd gnd NAND2X1
XFILL_1__1263_ vdd gnd FILL
XFILL_1__1194_ vdd gnd FILL
XFILL_2__1510_ vdd gnd FILL
XFILL_2__1441_ vdd gnd FILL
XFILL_2__1372_ vdd gnd FILL
XFILL_4__1239_ vdd gnd FILL
XFILL_0__974_ vdd gnd FILL
XFILL_2__1708_ vdd gnd FILL
XFILL_3__1550_ vdd gnd FILL
XFILL_0__1772_ vdd gnd FILL
XFILL_3__1481_ vdd gnd FILL
X_927_ _927_/A _928_/B vdd gnd INVX2
XFILL_0__1841_ vdd gnd FILL
XFILL_2__1639_ vdd gnd FILL
XFILL_4__952_ vdd gnd FILL
X_1001_ _992_/A _999_/Y _1001_/C _1866_/D vdd gnd OAI21X1
XCLKBUF1_insert10 clk _1904_/CLK vdd gnd CLKBUF1
X_1765_ _1773_/A _1766_/C vdd gnd INVX1
X_1834_ _948_/A Yin[0] _1835_/C vdd gnd NAND2X1
XFILL_0__1206_ vdd gnd FILL
XFILL_0__1137_ vdd gnd FILL
X_1903_ _1903_/D _1903_/CLK _950_/B vdd gnd DFFPOSX1
X_1696_ _1696_/A _1696_/B _1696_/C _1706_/A vdd gnd OAI21X1
XFILL_3__1748_ vdd gnd FILL
XFILL_3__1817_ vdd gnd FILL
XFILL_0__1068_ vdd gnd FILL
XFILL_3__1679_ vdd gnd FILL
XFILL_1__939_ vdd gnd FILL
XFILL_1__1315_ vdd gnd FILL
XFILL_1__1246_ vdd gnd FILL
XFILL_4__1024_ vdd gnd FILL
XFILL_3__970_ vdd gnd FILL
XFILL_1__1177_ vdd gnd FILL
XFILL_2__1355_ vdd gnd FILL
XFILL_2__1424_ vdd gnd FILL
XFILL101250x150 vdd gnd FILL
XFILL_0__957_ vdd gnd FILL
XFILL_2__1286_ vdd gnd FILL
XFILL_3__1602_ vdd gnd FILL
X_1550_ _1574_/B _1574_/A _1634_/C _1564_/A vdd gnd NAND3X1
X_1481_ _1494_/A _1493_/A _1494_/B _1482_/A vdd gnd NAND3X1
XFILL_2_BUFX2_insert17 vdd gnd FILL
XFILL_0__1686_ vdd gnd FILL
XFILL_0__1755_ vdd gnd FILL
XFILL_0__1824_ vdd gnd FILL
XFILL_3__1464_ vdd gnd FILL
XFILL_3__1533_ vdd gnd FILL
XFILL99750x23550 vdd gnd FILL
XFILL_1__1100_ vdd gnd FILL
XFILL_3__1395_ vdd gnd FILL
X_1748_ _1748_/A _1748_/B _1748_/C _1774_/A vdd gnd AOI21X1
X_1817_ _1890_/Q _1824_/B _1818_/C vdd gnd NOR2X1
XFILL_1__1031_ vdd gnd FILL
X_1679_ _1679_/A _1679_/B _1679_/C _1682_/A vdd gnd NAND3X1
XFILL_4__1573_ vdd gnd FILL
XFILL_1__1795_ vdd gnd FILL
XFILL_1_BUFX2_insert3 vdd gnd FILL
XFILL_2__1140_ vdd gnd FILL
XFILL101250x93750 vdd gnd FILL
XFILL_2__1071_ vdd gnd FILL
XFILL_1__1229_ vdd gnd FILL
XFILL_3__953_ vdd gnd FILL
XFILL_0__1540_ vdd gnd FILL
XFILL_0__1471_ vdd gnd FILL
XFILL_2__1407_ vdd gnd FILL
XFILL_2__1338_ vdd gnd FILL
XFILL_2__1269_ vdd gnd FILL
XFILL_3__1180_ vdd gnd FILL
X_1602_ _1602_/A _1647_/A _1602_/C _1649_/B vdd gnd NAND3X1
X_1464_ _1543_/C _1525_/B _1525_/A _1470_/B vdd gnd AOI21X1
X_1533_ _963_/A _1533_/B _965_/A _1533_/D _1597_/B vdd gnd OAI22X1
X_1395_ _1395_/A _1395_/B _1396_/B vdd gnd AND2X2
XFILL_0__1669_ vdd gnd FILL
XFILL_0__1738_ vdd gnd FILL
XFILL_1__1580_ vdd gnd FILL
XFILL_3__1516_ vdd gnd FILL
XFILL_0__1807_ vdd gnd FILL
XFILL_3__1447_ vdd gnd FILL
XFILL_3__1378_ vdd gnd FILL
XFILL_2__971_ vdd gnd FILL
XFILL_1__1014_ vdd gnd FILL
XFILL_1__1916_ vdd gnd FILL
XFILL_1__1778_ vdd gnd FILL
XFILL_1__1847_ vdd gnd FILL
XFILL_2__1123_ vdd gnd FILL
XFILL_2__1054_ vdd gnd FILL
XFILL_3__936_ vdd gnd FILL
XFILL_0__1523_ vdd gnd FILL
XFILL_3__1232_ vdd gnd FILL
XFILL_3__1301_ vdd gnd FILL
X_1180_ _1243_/A _1184_/C vdd gnd INVX1
XFILL_0__1454_ vdd gnd FILL
XFILL_3__1094_ vdd gnd FILL
XFILL_3__1163_ vdd gnd FILL
XFILL_0__1385_ vdd gnd FILL
X_1516_ _1520_/A _1521_/C _1520_/B _1517_/B vdd gnd NAND3X1
XFILL_1__1632_ vdd gnd FILL
X_1447_ _1454_/A _1615_/B _1542_/B vdd gnd NOR2X1
XFILL_1__1701_ vdd gnd FILL
X_1378_ _1397_/B _1397_/A _1397_/C _1483_/A vdd gnd NAND3X1
XFILL_1__1563_ vdd gnd FILL
XFILL_1__1494_ vdd gnd FILL
XFILL_4__1272_ vdd gnd FILL
XFILL_2__954_ vdd gnd FILL
XFILL_2__1672_ vdd gnd FILL
XFILL_2__1741_ vdd gnd FILL
XFILL_2__1810_ vdd gnd FILL
X_960_ Xin[1] _965_/B _961_/C vdd gnd NAND2X1
XFILL_0__1170_ vdd gnd FILL
XFILL_2__1106_ vdd gnd FILL
XFILL_3__1781_ vdd gnd FILL
XFILL_2__1037_ vdd gnd FILL
X_1232_ _953_/B Cin[4] _1313_/A vdd gnd NAND2X1
XFILL_1__972_ vdd gnd FILL
X_1301_ _1301_/A _1301_/B _1301_/C _1379_/C vdd gnd AOI21X1
XFILL_0__1506_ vdd gnd FILL
XFILL_0__1437_ vdd gnd FILL
XBUFX2_insert4 _1910_/Q _998_/A vdd gnd BUFX2
X_1094_ _1213_/B _1095_/C _1095_/B _1097_/A vdd gnd OAI21X1
XFILL_3__1215_ vdd gnd FILL
X_1163_ _953_/B Cin[3] _1169_/A vdd gnd AND2X2
XFILL_0__1368_ vdd gnd FILL
XFILL_3__1146_ vdd gnd FILL
XFILL_3__1077_ vdd gnd FILL
XFILL_0__1299_ vdd gnd FILL
XFILL_1__1546_ vdd gnd FILL
XFILL_1__1615_ vdd gnd FILL
XFILL_1__1477_ vdd gnd FILL
XFILL_2__937_ vdd gnd FILL
XFILL_0__990_ vdd gnd FILL
XFILL_2__1724_ vdd gnd FILL
XFILL_2__1655_ vdd gnd FILL
X_943_ _943_/A _943_/B _943_/C _945_/B vdd gnd OAI21X1
XFILL_2__1586_ vdd gnd FILL
X_1781_ _1782_/B _1793_/B _1793_/C vdd gnd OR2X2
XFILL_3__1000_ vdd gnd FILL
XFILL_0__1222_ vdd gnd FILL
X_1850_ _959_/Y _1903_/CLK _946_/A vdd gnd DFFPOSX1
XFILL_0__1153_ vdd gnd FILL
XFILL_0__1084_ vdd gnd FILL
XFILL_3__1764_ vdd gnd FILL
XFILL_3__1833_ vdd gnd FILL
XFILL_3__1695_ vdd gnd FILL
XFILL_1__955_ vdd gnd FILL
XFILL_1__1400_ vdd gnd FILL
X_1146_ _1212_/B _1212_/A _1147_/B vdd gnd NAND2X1
X_1215_ _1215_/A _1217_/B _1216_/B vdd gnd XOR2X1
XFILL_1__1331_ vdd gnd FILL
XFILL_1__1262_ vdd gnd FILL
XFILL_3__1129_ vdd gnd FILL
X_1077_ _1082_/A _1079_/B _1079_/A _1138_/A vdd gnd NAND3X1
XFILL_1__1193_ vdd gnd FILL
XFILL_2__1440_ vdd gnd FILL
XFILL_1__1529_ vdd gnd FILL
XFILL_4__1307_ vdd gnd FILL
XFILL_2__1371_ vdd gnd FILL
XFILL_0__973_ vdd gnd FILL
XFILL_0__1840_ vdd gnd FILL
XFILL_2__1638_ vdd gnd FILL
XFILL_0__1771_ vdd gnd FILL
XFILL_2__1707_ vdd gnd FILL
XFILL_3__1480_ vdd gnd FILL
X_1000_ _992_/A _1882_/Q _1001_/C vdd gnd NAND2X1
X_926_ _943_/A _999_/A _926_/C _930_/B vdd gnd OAI21X1
XFILL_2__1569_ vdd gnd FILL
XCLKBUF1_insert11 clk _1903_/CLK vdd gnd CLKBUF1
X_1902_ _1902_/D _1910_/CLK _947_/B vdd gnd DFFPOSX1
X_1764_ _1774_/B _1774_/A _1773_/A vdd gnd XOR2X1
X_1833_ _1833_/A _1833_/B _1833_/C _1897_/D vdd gnd OAI21X1
XFILL_0__1205_ vdd gnd FILL
XFILL_0__1136_ vdd gnd FILL
XFILL_0__1067_ vdd gnd FILL
X_1695_ _1695_/A _1695_/B _1695_/C _1696_/B vdd gnd AOI21X1
XFILL_3__1747_ vdd gnd FILL
XFILL_3__1816_ vdd gnd FILL
XFILL_3__1678_ vdd gnd FILL
XFILL_1__938_ vdd gnd FILL
X_1129_ _1161_/B _1196_/C _1161_/A _1142_/B vdd gnd NAND3X1
XFILL_1__1314_ vdd gnd FILL
XFILL_1__1176_ vdd gnd FILL
XFILL_1__1245_ vdd gnd FILL
XFILL_4__1787_ vdd gnd FILL
XFILL_2__1423_ vdd gnd FILL
XFILL_2__1354_ vdd gnd FILL
XFILL_2__1285_ vdd gnd FILL
XFILL_0__956_ vdd gnd FILL
XFILL_3__1601_ vdd gnd FILL
XFILL_3__1532_ vdd gnd FILL
X_1480_ _1480_/A _1480_/B _1480_/C _1494_/B vdd gnd OAI21X1
XFILL_0__1823_ vdd gnd FILL
XFILL_2_BUFX2_insert18 vdd gnd FILL
XFILL_0__1685_ vdd gnd FILL
XFILL_3__1463_ vdd gnd FILL
XFILL_0__1754_ vdd gnd FILL
XFILL_3__1394_ vdd gnd FILL
XFILL_4__934_ vdd gnd FILL
XFILL_1__1030_ vdd gnd FILL
X_1678_ _1678_/A _1678_/B _1681_/A _1688_/A vdd gnd OAI21X1
XFILL_4__1710_ vdd gnd FILL
X_1747_ _1747_/A _1747_/B _1767_/B vdd gnd AND2X2
XFILL_4__1641_ vdd gnd FILL
X_1816_ _1816_/A _945_/A _1824_/B vdd gnd NOR2X1
XFILL_0__1119_ vdd gnd FILL
XFILL_1__1794_ vdd gnd FILL
XFILL_1_BUFX2_insert4 vdd gnd FILL
XFILL_4__1006_ vdd gnd FILL
XFILL_1__1159_ vdd gnd FILL
XFILL_2__1070_ vdd gnd FILL
XFILL_1__1228_ vdd gnd FILL
XFILL_3__952_ vdd gnd FILL
XFILL_0__1470_ vdd gnd FILL
XFILL_2__1406_ vdd gnd FILL
XFILL_2__1337_ vdd gnd FILL
XFILL_2__1268_ vdd gnd FILL
X_1601_ _1601_/A _1601_/B _1601_/C _1602_/C vdd gnd OAI21X1
X_1532_ _1611_/A _1596_/B _1592_/C vdd gnd NAND2X1
XFILL_0__939_ vdd gnd FILL
XFILL_2__1199_ vdd gnd FILL
XFILL_3__1515_ vdd gnd FILL
X_1463_ _1524_/A _1524_/B _1524_/C _1525_/B vdd gnd NAND3X1
XFILL_0__1806_ vdd gnd FILL
X_1394_ _1394_/A _1396_/A vdd gnd INVX1
XFILL_0__1668_ vdd gnd FILL
XFILL_0__1737_ vdd gnd FILL
XFILL_0__1599_ vdd gnd FILL
XFILL_3__1446_ vdd gnd FILL
XFILL_2__970_ vdd gnd FILL
XFILL_3__1377_ vdd gnd FILL
XFILL_1__1013_ vdd gnd FILL
XFILL_1__1915_ vdd gnd FILL
XFILL_4__1555_ vdd gnd FILL
XFILL_1__1777_ vdd gnd FILL
XFILL_4__1486_ vdd gnd FILL
XFILL_1__1846_ vdd gnd FILL
XFILL_2__1122_ vdd gnd FILL
XFILL_2__1053_ vdd gnd FILL
XFILL_3__935_ vdd gnd FILL
XFILL_0__1522_ vdd gnd FILL
XFILL_0__1453_ vdd gnd FILL
XFILL_3__1231_ vdd gnd FILL
XFILL_3__1300_ vdd gnd FILL
XFILL_3__1162_ vdd gnd FILL
XFILL_3__1093_ vdd gnd FILL
XFILL_0__1384_ vdd gnd FILL
X_1515_ _1515_/A _1611_/A _1515_/C _1515_/D _1521_/C vdd gnd AOI22X1
XFILL_1__1700_ vdd gnd FILL
XFILL_1__1631_ vdd gnd FILL
X_1446_ _1605_/B _1615_/B vdd gnd INVX1
XFILL_1__1562_ vdd gnd FILL
XFILL_4__1340_ vdd gnd FILL
X_1377_ _1398_/A _1484_/A vdd gnd INVX1
XFILL_1__1493_ vdd gnd FILL
XFILL_3__1429_ vdd gnd FILL
XFILL_2__953_ vdd gnd FILL
XFILL101250x19650 vdd gnd FILL
XFILL_2__1740_ vdd gnd FILL
XFILL_2__1671_ vdd gnd FILL
XFILL_1__1829_ vdd gnd FILL
XFILL_2__1105_ vdd gnd FILL
XFILL_2__1036_ vdd gnd FILL
XFILL_3__1780_ vdd gnd FILL
XFILL_1__971_ vdd gnd FILL
X_1231_ _1231_/A _1231_/B _1231_/C _1274_/C vdd gnd AOI21X1
X_1300_ _1372_/C _1301_/C vdd gnd INVX1
X_1162_ _950_/B Cin[4] _1168_/A vdd gnd NAND2X1
XFILL_0__1505_ vdd gnd FILL
XFILL_0__1436_ vdd gnd FILL
X_1093_ _1093_/A _1093_/B _1093_/C _1093_/D _1213_/B vdd gnd AOI22X1
XFILL_3__1145_ vdd gnd FILL
XFILL_3__1214_ vdd gnd FILL
XFILL_0__1367_ vdd gnd FILL
XFILL_0__1298_ vdd gnd FILL
XFILL_3__1076_ vdd gnd FILL
X_1429_ _1468_/A _1495_/B _1552_/A vdd gnd NAND2X1
XFILL_1_BUFX2_insert20 vdd gnd FILL
XFILL_1__1545_ vdd gnd FILL
XFILL_1__1614_ vdd gnd FILL
XFILL_1__1476_ vdd gnd FILL
XFILL_4__1254_ vdd gnd FILL
XFILL_2__936_ vdd gnd FILL
XFILL_1_CLKBUF1_insert10 vdd gnd FILL
XFILL_4__1185_ vdd gnd FILL
XFILL_2__1585_ vdd gnd FILL
XFILL_2__1654_ vdd gnd FILL
XFILL_2__1723_ vdd gnd FILL
X_942_ _943_/A _998_/B _943_/C vdd gnd NAND2X1
XFILL_0__1221_ vdd gnd FILL
X_1780_ _1887_/Q _1780_/B _1782_/B vdd gnd NAND2X1
XFILL_2__1019_ vdd gnd FILL
XFILL_0__1083_ vdd gnd FILL
XFILL_0__1152_ vdd gnd FILL
XFILL_3__1694_ vdd gnd FILL
XFILL_3__1763_ vdd gnd FILL
XFILL_3__1832_ vdd gnd FILL
XFILL_1__954_ vdd gnd FILL
XFILL_1__1330_ vdd gnd FILL
X_1145_ _1213_/B _1147_/A vdd gnd INVX1
X_1214_ _1217_/A _1214_/B _1215_/A vdd gnd NOR2X1
XFILL_0__1419_ vdd gnd FILL
XFILL_1__1261_ vdd gnd FILL
XFILL_3__1128_ vdd gnd FILL
X_1076_ _1083_/C _1102_/C _1083_/A _1079_/B vdd gnd NAND3X1
XFILL_1__1192_ vdd gnd FILL
XFILL_3__1059_ vdd gnd FILL
XFILL_1__1528_ vdd gnd FILL
XFILL_1__1459_ vdd gnd FILL
XFILL_2__1370_ vdd gnd FILL
XFILL_0__972_ vdd gnd FILL
XFILL_4__1099_ vdd gnd FILL
X_925_ _943_/A _992_/B _926_/C vdd gnd NAND2X1
XFILL100050x23550 vdd gnd FILL
XFILL_2__1637_ vdd gnd FILL
XFILL100650x70350 vdd gnd FILL
XFILL_2__1706_ vdd gnd FILL
XFILL_0__1770_ vdd gnd FILL
XFILL_2__1568_ vdd gnd FILL
XFILL_2__1499_ vdd gnd FILL
X_1832_ _957_/A _928_/B _1897_/Q _1833_/C vdd gnd OAI21X1
XFILL_0__1204_ vdd gnd FILL
X_1901_ _1901_/D _1908_/CLK _1901_/Q vdd gnd DFFPOSX1
X_1694_ _1694_/A _1694_/B _1694_/C _1696_/A vdd gnd AOI21X1
X_1763_ _1763_/A _1763_/B _1774_/B vdd gnd NAND2X1
XFILL_0__1135_ vdd gnd FILL
XFILL_0__1066_ vdd gnd FILL
XFILL_3__1677_ vdd gnd FILL
XFILL_3__1746_ vdd gnd FILL
XFILL_3__1815_ vdd gnd FILL
XFILL_1__937_ vdd gnd FILL
XFILL_1__1313_ vdd gnd FILL
X_1128_ _1132_/B _1159_/C _1161_/A vdd gnd AND2X2
X_1059_ _977_/A _1095_/B _1060_/B vdd gnd NAND2X1
XFILL_1__1175_ vdd gnd FILL
XFILL_1__1244_ vdd gnd FILL
XFILL_2__1422_ vdd gnd FILL
XFILL_2__1353_ vdd gnd FILL
XFILL_2__1284_ vdd gnd FILL
XFILL_0__955_ vdd gnd FILL
XFILL_1_CLKBUF1_insert5 vdd gnd FILL
XFILL100050x35250 vdd gnd FILL
XFILL_3__1600_ vdd gnd FILL
XFILL_0__1822_ vdd gnd FILL
XFILL_3__1531_ vdd gnd FILL
XFILL_0__1753_ vdd gnd FILL
XFILL_2_BUFX2_insert19 vdd gnd FILL
XFILL_0__1684_ vdd gnd FILL
XFILL_3__1462_ vdd gnd FILL
XFILL_3__1393_ vdd gnd FILL
X_1815_ _1833_/A _1815_/B _1815_/C _1889_/D vdd gnd OAI21X1
X_1677_ _1677_/A _1733_/A _1681_/A vdd gnd NAND2X1
X_1746_ _1771_/A _1773_/B vdd gnd INVX1
XFILL_0__1118_ vdd gnd FILL
XFILL_0__1049_ vdd gnd FILL
XFILL_3__1729_ vdd gnd FILL
XFILL_1__1793_ vdd gnd FILL
XFILL_1__1089_ vdd gnd FILL
XFILL_1__1227_ vdd gnd FILL
XFILL_1__1158_ vdd gnd FILL
XFILL_4__1838_ vdd gnd FILL
XFILL_3__951_ vdd gnd FILL
XFILL_2__1405_ vdd gnd FILL
XFILL_2__1336_ vdd gnd FILL
XFILL_0__938_ vdd gnd FILL
XFILL_2__1198_ vdd gnd FILL
XFILL_2__1267_ vdd gnd FILL
X_1600_ _1600_/A _1600_/B _1600_/C _1647_/A vdd gnd NAND3X1
X_1531_ _1592_/A _1597_/A vdd gnd INVX1
X_1462_ _1542_/A _1542_/B _1543_/C vdd gnd NAND2X1
XFILL_0__1736_ vdd gnd FILL
XFILL_3__1514_ vdd gnd FILL
XFILL_3__1445_ vdd gnd FILL
XFILL_0__1805_ vdd gnd FILL
X_1393_ _991_/B _1702_/B _1490_/C vdd gnd NAND2X1
XFILL_0__1667_ vdd gnd FILL
XFILL_0__1598_ vdd gnd FILL
XFILL_3__1376_ vdd gnd FILL
XFILL_1__1012_ vdd gnd FILL
XFILL_4__1623_ vdd gnd FILL
X_1729_ _1729_/A _1730_/B vdd gnd INVX1
XFILL_1__1914_ vdd gnd FILL
XFILL_1__1845_ vdd gnd FILL
XFILL_1__1776_ vdd gnd FILL
XFILL_2__1121_ vdd gnd FILL
XFILL_2__1052_ vdd gnd FILL
XFILL_3__934_ vdd gnd FILL
XFILL_0__1521_ vdd gnd FILL
XFILL_0__1452_ vdd gnd FILL
XFILL_2__1319_ vdd gnd FILL
XFILL_3__1161_ vdd gnd FILL
XFILL_0__1383_ vdd gnd FILL
XFILL_3__1092_ vdd gnd FILL
XFILL_3__1230_ vdd gnd FILL
X_1514_ _1579_/B _1514_/B _1579_/A _1520_/B vdd gnd OAI21X1
X_1445_ _955_/A Cin[1] _1890_/Q _1605_/B vdd gnd NAND3X1
XFILL_1__1630_ vdd gnd FILL
XFILL_0__1719_ vdd gnd FILL
XFILL_1__1561_ vdd gnd FILL
XFILL_1__1492_ vdd gnd FILL
XFILL_3__1428_ vdd gnd FILL
X_1376_ _1385_/C _1385_/B _1398_/A _1381_/B vdd gnd AOI21X1
XFILL_2__952_ vdd gnd FILL
XFILL_3__1359_ vdd gnd FILL
XFILL_2__1670_ vdd gnd FILL
XFILL_4__1537_ vdd gnd FILL
XFILL_4__1606_ vdd gnd FILL
XFILL_1__1828_ vdd gnd FILL
XFILL_1__1759_ vdd gnd FILL
XFILL_4__1468_ vdd gnd FILL
XFILL_2__1035_ vdd gnd FILL
XFILL_2__1104_ vdd gnd FILL
XFILL_1__970_ vdd gnd FILL
XFILL_2__1799_ vdd gnd FILL
X_1161_ _1161_/A _1161_/B _1161_/C _1203_/C vdd gnd AOI21X1
X_1092_ _1092_/A _1092_/B _1095_/C vdd gnd NOR2X1
X_1230_ _1267_/C _1231_/C vdd gnd INVX1
XFILL_0__1504_ vdd gnd FILL
XFILL_0__1435_ vdd gnd FILL
XFILL_0__1366_ vdd gnd FILL
XFILL_3__1213_ vdd gnd FILL
XFILL_3__1144_ vdd gnd FILL
XFILL_3__1075_ vdd gnd FILL
XFILL_0__1297_ vdd gnd FILL
XFILL_1__1613_ vdd gnd FILL
X_1428_ _1428_/A _1495_/A _1428_/C _1495_/B vdd gnd NAND3X1
XFILL_1_BUFX2_insert21 vdd gnd FILL
XFILL_1__1544_ vdd gnd FILL
XFILL_1__1475_ vdd gnd FILL
X_1359_ _1473_/B _1473_/A _1368_/C _1374_/A vdd gnd NAND3X1
XFILL_4__1322_ vdd gnd FILL
XFILL_1_CLKBUF1_insert11 vdd gnd FILL
XFILL_2__935_ vdd gnd FILL
XFILL_2__1722_ vdd gnd FILL
X_941_ _941_/A _998_/B vdd gnd INVX1
XFILL_2__1653_ vdd gnd FILL
XFILL_2__1584_ vdd gnd FILL
XFILL_0__1220_ vdd gnd FILL
XFILL_3__1831_ vdd gnd FILL
XFILL_2__1018_ vdd gnd FILL
XFILL_0__1082_ vdd gnd FILL
XFILL_0__1151_ vdd gnd FILL
XFILL_3__1693_ vdd gnd FILL
XFILL_3__1762_ vdd gnd FILL
XFILL_1__953_ vdd gnd FILL
X_1213_ _1213_/A _1213_/B _1290_/C _1213_/D _1217_/A vdd gnd AOI22X1
X_1144_ _1213_/B _1212_/B _1212_/A _1153_/A vdd gnd NAND3X1
X_1075_ _1102_/B _1083_/A vdd gnd INVX1
XFILL_1__1260_ vdd gnd FILL
XFILL_0__1349_ vdd gnd FILL
XFILL_0__1418_ vdd gnd FILL
XFILL_1__1191_ vdd gnd FILL
XFILL_3__1127_ vdd gnd FILL
XFILL_3__1058_ vdd gnd FILL
XFILL_1__1458_ vdd gnd FILL
XFILL_1__1527_ vdd gnd FILL
XFILL_0__971_ vdd gnd FILL
XFILL_4__1236_ vdd gnd FILL
XFILL_1__1389_ vdd gnd FILL
XFILL_4__1167_ vdd gnd FILL
XFILL_2__1705_ vdd gnd FILL
X_924_ _924_/A _992_/B vdd gnd INVX1
XFILL_2__1636_ vdd gnd FILL
XFILL_2__1498_ vdd gnd FILL
XFILL_2__1567_ vdd gnd FILL
X_1831_ _1839_/B _1833_/B _1831_/C _1896_/D vdd gnd OAI21X1
X_1900_ _1900_/D _1908_/CLK _1900_/Q vdd gnd DFFPOSX1
XFILL_0__1203_ vdd gnd FILL
XFILL_0__1134_ vdd gnd FILL
X_1693_ _1693_/A _1693_/B _1693_/C _1696_/C vdd gnd AOI21X1
X_1762_ _1776_/C _1762_/B _1762_/C _1763_/B vdd gnd OAI21X1
XFILL_3__1814_ vdd gnd FILL
XFILL_0__1065_ vdd gnd FILL
XFILL_3__1676_ vdd gnd FILL
XFILL_3__1745_ vdd gnd FILL
XFILL_1__936_ vdd gnd FILL
XFILL_1__1312_ vdd gnd FILL
XFILL_1__1243_ vdd gnd FILL
X_1127_ _1127_/A _1127_/B _1127_/C _1132_/B vdd gnd NAND3X1
X_1058_ _1058_/A _1093_/A _1058_/C _1095_/B vdd gnd NAND3X1
XFILL_4__1021_ vdd gnd FILL
XFILL_1__1174_ vdd gnd FILL
XFILL_2__1352_ vdd gnd FILL
XFILL_2__1421_ vdd gnd FILL
XFILL_1_CLKBUF1_insert6 vdd gnd FILL
XFILL_0__954_ vdd gnd FILL
XFILL_2__1283_ vdd gnd FILL
XFILL100950x66450 vdd gnd FILL
XFILL_3__1530_ vdd gnd FILL
XFILL_0__1821_ vdd gnd FILL
XFILL_0__1752_ vdd gnd FILL
XFILL_3__1461_ vdd gnd FILL
XFILL_2__1619_ vdd gnd FILL
XFILL_0__1683_ vdd gnd FILL
XFILL_3__1392_ vdd gnd FILL
X_1745_ _1790_/A _1745_/B _1745_/C _1882_/D vdd gnd OAI21X1
X_1814_ _1889_/Q _1815_/B _1815_/C vdd gnd NAND2X1
XFILL_0__1117_ vdd gnd FILL
X_1676_ _1710_/B _1710_/A _1677_/A vdd gnd NAND2X1
XFILL_3__1728_ vdd gnd FILL
XFILL_1__1792_ vdd gnd FILL
XFILL_4__1570_ vdd gnd FILL
XFILL_0__1048_ vdd gnd FILL
XFILL_3__1659_ vdd gnd FILL
XFILL_1__1226_ vdd gnd FILL
XFILL_1__1157_ vdd gnd FILL
XFILL_1__1088_ vdd gnd FILL
XFILL_3__950_ vdd gnd FILL
XFILL_2__1404_ vdd gnd FILL
XFILL_2__1335_ vdd gnd FILL
XFILL100950x78150 vdd gnd FILL
XFILL_0__937_ vdd gnd FILL
XFILL_2__1266_ vdd gnd FILL
XFILL_2__1197_ vdd gnd FILL
X_1530_ _1592_/A _1530_/B _1530_/C _1539_/C vdd gnd NAND3X1
X_1461_ _1461_/A _1461_/B _1461_/C _1551_/C vdd gnd OAI21X1
X_1392_ _990_/A _990_/B _1392_/C _1392_/D _1877_/D vdd gnd AOI22X1
XFILL_0__1735_ vdd gnd FILL
XFILL_3__1513_ vdd gnd FILL
XFILL_0__1666_ vdd gnd FILL
XFILL_3__1444_ vdd gnd FILL
XFILL_0__1804_ vdd gnd FILL
XFILL_0__1597_ vdd gnd FILL
XFILL_3__1375_ vdd gnd FILL
X_1728_ _1728_/A _1728_/B _1730_/C vdd gnd OR2X2
XFILL_1__1011_ vdd gnd FILL
X_1659_ _1666_/B _1666_/C _1711_/C _1671_/C vdd gnd NAND3X1
XFILL_1__1775_ vdd gnd FILL
XFILL_1__1913_ vdd gnd FILL
XFILL_1__1844_ vdd gnd FILL
XFILL_1__1209_ vdd gnd FILL
XFILL_2__1051_ vdd gnd FILL
XFILL_2__1120_ vdd gnd FILL
XFILL_3__933_ vdd gnd FILL
XFILL_0__1520_ vdd gnd FILL
XFILL_0__1451_ vdd gnd FILL
XFILL_2__1318_ vdd gnd FILL
XFILL_3__1160_ vdd gnd FILL
XFILL_0__1382_ vdd gnd FILL
XFILL_3__1091_ vdd gnd FILL
XFILL_2__1249_ vdd gnd FILL
X_1513_ _1513_/A _1513_/B _1579_/C _1520_/A vdd gnd NAND3X1
X_1444_ _955_/A Cin[1] _1890_/Q _1454_/A vdd gnd AOI21X1
X_1375_ _1379_/A _1379_/B _1397_/C _1385_/B vdd gnd OAI21X1
XFILL_0__1649_ vdd gnd FILL
XFILL_1__1560_ vdd gnd FILL
XFILL_0__1718_ vdd gnd FILL
XFILL_1__1491_ vdd gnd FILL
XFILL_3__1427_ vdd gnd FILL
XFILL_3__1358_ vdd gnd FILL
XFILL_3__1289_ vdd gnd FILL
XFILL_2__951_ vdd gnd FILL
XFILL_1__1758_ vdd gnd FILL
XFILL_1__1827_ vdd gnd FILL
XFILL_1__1689_ vdd gnd FILL
XFILL_2__1103_ vdd gnd FILL
XFILL_2__1034_ vdd gnd FILL
XFILL_0__1503_ vdd gnd FILL
XFILL_2__1798_ vdd gnd FILL
X_1160_ _1219_/B _1160_/B _1278_/A vdd gnd XOR2X1
XFILL_3__1212_ vdd gnd FILL
X_1091_ _1093_/D _1093_/C _1092_/B vdd gnd NAND2X1
XFILL_0__1434_ vdd gnd FILL
XFILL_0__1365_ vdd gnd FILL
XFILL_3__1143_ vdd gnd FILL
XFILL_3__1074_ vdd gnd FILL
XFILL_0__1296_ vdd gnd FILL
XFILL_1__1612_ vdd gnd FILL
X_1427_ _1427_/A _1427_/B _1427_/C _1428_/C vdd gnd OAI21X1
X_1358_ _1461_/C _1431_/B _1431_/A _1473_/A vdd gnd NAND3X1
XFILL_1_BUFX2_insert22 vdd gnd FILL
XFILL_1__1543_ vdd gnd FILL
XFILL_1__1474_ vdd gnd FILL
X_1289_ _1289_/A _1289_/B _1383_/A _1290_/B vdd gnd AOI21X1
XFILL_2__934_ vdd gnd FILL
XFILL_2__1652_ vdd gnd FILL
XFILL_2__1721_ vdd gnd FILL
X_940_ _945_/A _940_/B _940_/C _940_/Y vdd gnd OAI21X1
XFILL_2__1583_ vdd gnd FILL
XFILL_4__1519_ vdd gnd FILL
XFILL_0__1150_ vdd gnd FILL
XFILL_3__1761_ vdd gnd FILL
XFILL_3__1830_ vdd gnd FILL
XFILL_2__1017_ vdd gnd FILL
XFILL_0__1081_ vdd gnd FILL
XFILL_3__1692_ vdd gnd FILL
XFILL_1__952_ vdd gnd FILL
XFILL_2__1919_ vdd gnd FILL
X_1212_ _1212_/A _1212_/B _1213_/A vdd gnd AND2X2
XFILL_0__1417_ vdd gnd FILL
XFILL99750x31350 vdd gnd FILL
X_1143_ _1206_/B _1154_/C _1206_/A _1212_/A vdd gnd NAND3X1
X_1074_ _1102_/A _1083_/C vdd gnd INVX1
XFILL99450x66450 vdd gnd FILL
XFILL_0__1348_ vdd gnd FILL
XFILL_1__1190_ vdd gnd FILL
XFILL_0__1279_ vdd gnd FILL
XFILL_3__1126_ vdd gnd FILL
XFILL_3__1057_ vdd gnd FILL
XFILL_1__1526_ vdd gnd FILL
XFILL_4__1304_ vdd gnd FILL
XFILL_1__1457_ vdd gnd FILL
XFILL_0__970_ vdd gnd FILL
XFILL_1__1388_ vdd gnd FILL
XFILL_2__1635_ vdd gnd FILL
XFILL_2__1704_ vdd gnd FILL
X_923_ _923_/A _945_/A vdd gnd INVX2
XFILL_2__1566_ vdd gnd FILL
XFILL_2__1497_ vdd gnd FILL
X_1761_ _1776_/B _1762_/B vdd gnd INVX1
X_1830_ _944_/A _928_/B _1896_/Q _1831_/C vdd gnd OAI21X1
XFILL_0__1202_ vdd gnd FILL
XFILL_0__1133_ vdd gnd FILL
X_1692_ _1692_/A _1693_/C vdd gnd INVX1
XFILL_3__1744_ vdd gnd FILL
XFILL_3__1813_ vdd gnd FILL
XFILL_0__1064_ vdd gnd FILL
XFILL_3__1675_ vdd gnd FILL
XFILL_1__935_ vdd gnd FILL
X_1126_ _1845_/B _1533_/B _1158_/A _1127_/C vdd gnd OAI21X1
XFILL_1__1311_ vdd gnd FILL
XFILL_1__1242_ vdd gnd FILL
XFILL_3__1109_ vdd gnd FILL
XFILL_1__1173_ vdd gnd FILL
X_1057_ _1058_/C _1093_/A _1058_/A _1060_/A vdd gnd AOI21X1
XFILL_4__1784_ vdd gnd FILL
XFILL_1__1509_ vdd gnd FILL
XFILL_2__1351_ vdd gnd FILL
XFILL_2__1420_ vdd gnd FILL
XFILL_2__1282_ vdd gnd FILL
XFILL_4__1218_ vdd gnd FILL
XFILL_0__953_ vdd gnd FILL
XFILL_1_CLKBUF1_insert7 vdd gnd FILL
XFILL_4__1149_ vdd gnd FILL
XFILL_0__1820_ vdd gnd FILL
XFILL_2__1618_ vdd gnd FILL
XFILL_0__1682_ vdd gnd FILL
XFILL_0__1751_ vdd gnd FILL
XFILL_3__1460_ vdd gnd FILL
XFILL_3__1391_ vdd gnd FILL
XFILL_2__1549_ vdd gnd FILL
XFILL_4__931_ vdd gnd FILL
X_1744_ _1747_/A _1747_/B _1745_/B vdd gnd XNOR2X1
X_1813_ Yin[3] _1833_/A vdd gnd INVX1
XFILL_0__1047_ vdd gnd FILL
XFILL_0__1116_ vdd gnd FILL
X_1675_ _1710_/A _1710_/B _1733_/A vdd gnd OR2X2
XFILL_3__1727_ vdd gnd FILL
XFILL_1__1791_ vdd gnd FILL
XFILL_3__1589_ vdd gnd FILL
XFILL_3__1658_ vdd gnd FILL
X_1109_ _1173_/C _1114_/B vdd gnd INVX1
XFILL_4__1003_ vdd gnd FILL
XFILL_1__1156_ vdd gnd FILL
XFILL_1__1225_ vdd gnd FILL
XFILL_1__1087_ vdd gnd FILL
XFILL_4__1767_ vdd gnd FILL
XFILL_4__1698_ vdd gnd FILL
XFILL_2__1334_ vdd gnd FILL
XFILL_2__1403_ vdd gnd FILL
XFILL_2__1265_ vdd gnd FILL
XFILL_0__936_ vdd gnd FILL
XFILL_2__1196_ vdd gnd FILL
XFILL_0__1803_ vdd gnd FILL
X_1460_ _1460_/A _1524_/B _1460_/C _1461_/B vdd gnd AOI21X1
X_1391_ _1391_/A _1391_/B _990_/A _1392_/C vdd gnd AOI21X1
XFILL_0__1734_ vdd gnd FILL
XFILL_0__1665_ vdd gnd FILL
XFILL_3__1512_ vdd gnd FILL
XFILL_3__1443_ vdd gnd FILL
XFILL_0__1596_ vdd gnd FILL
XFILL_3__1374_ vdd gnd FILL
XFILL_1__1010_ vdd gnd FILL
X_1727_ _1727_/A _1776_/A _1729_/A _1732_/B vdd gnd OAI21X1
X_1658_ _1794_/B _1658_/B _1711_/C vdd gnd NAND2X1
XFILL_1__1912_ vdd gnd FILL
X_1589_ _1589_/A _1658_/B _1652_/C vdd gnd NAND2X1
XFILL_4__1483_ vdd gnd FILL
XFILL_1__1774_ vdd gnd FILL
XFILL_4__1552_ vdd gnd FILL
XFILL_1__1843_ vdd gnd FILL
XFILL_1__1208_ vdd gnd FILL
XFILL_1__1139_ vdd gnd FILL
XFILL_2__1050_ vdd gnd FILL
XFILL_3__932_ vdd gnd FILL
XFILL_0__1450_ vdd gnd FILL
XFILL_2__1248_ vdd gnd FILL
XFILL_2__1317_ vdd gnd FILL
XFILL_3__1090_ vdd gnd FILL
XFILL_0__1381_ vdd gnd FILL
X_1512_ _1521_/A _1521_/B _1520_/C _1517_/C vdd gnd OAI21X1
XFILL_2__1179_ vdd gnd FILL
X_1443_ _1453_/B _1453_/A _1543_/A vdd gnd NAND2X1
X_1374_ _1374_/A _1374_/B _1474_/A _1379_/B vdd gnd AOI21X1
XFILL_0__1648_ vdd gnd FILL
XFILL_0__1579_ vdd gnd FILL
XFILL_0__1717_ vdd gnd FILL
XFILL_1__1490_ vdd gnd FILL
XFILL_3__1357_ vdd gnd FILL
XFILL_3__1426_ vdd gnd FILL
XFILL_3__1288_ vdd gnd FILL
XFILL_2__950_ vdd gnd FILL
XFILL_1__1688_ vdd gnd FILL
XFILL_1__1757_ vdd gnd FILL
XFILL_1__1826_ vdd gnd FILL
XFILL_4__1397_ vdd gnd FILL
XFILL_2__1102_ vdd gnd FILL
XFILL_2__1033_ vdd gnd FILL
XFILL_2__1797_ vdd gnd FILL
XFILL_0__1502_ vdd gnd FILL
XFILL_0__1433_ vdd gnd FILL
XFILL_3__1142_ vdd gnd FILL
X_1090_ _1101_/A _1138_/A _1140_/B _1093_/D vdd gnd NAND3X1
XFILL_3__1211_ vdd gnd FILL
XFILL_0__1364_ vdd gnd FILL
XFILL_3__1073_ vdd gnd FILL
XFILL_0__1295_ vdd gnd FILL
XFILL_1__1611_ vdd gnd FILL
XFILL_1__1542_ vdd gnd FILL
XFILL_1_BUFX2_insert23 vdd gnd FILL
X_1357_ _1357_/A _1357_/B _1357_/C _1431_/B vdd gnd OAI21X1
X_1426_ _1519_/C _1426_/B _1426_/C _1495_/A vdd gnd NAND3X1
XFILL_1_BUFX2_insert12 vdd gnd FILL
X_1288_ _1298_/B _1383_/C _1298_/A _1290_/A vdd gnd AOI21X1
XFILL_4__1251_ vdd gnd FILL
XFILL_3__1409_ vdd gnd FILL
XFILL_2__933_ vdd gnd FILL
XFILL_1__1473_ vdd gnd FILL
XFILL_4__1182_ vdd gnd FILL
XFILL_2__1651_ vdd gnd FILL
XFILL_2__1720_ vdd gnd FILL
XFILL_1__1809_ vdd gnd FILL
XFILL_2__1582_ vdd gnd FILL
XFILL_2__1016_ vdd gnd FILL
XFILL_0__1080_ vdd gnd FILL
XFILL_3__1760_ vdd gnd FILL
XFILL_2__1918_ vdd gnd FILL
XFILL_3__1691_ vdd gnd FILL
X_999_ _999_/A _999_/Y vdd gnd INVX1
XFILL_2__1849_ vdd gnd FILL
X_1142_ _1142_/A _1142_/B _1142_/C _1154_/C vdd gnd NAND3X1
X_1211_ _1217_/C _1214_/B vdd gnd INVX1
XFILL_1__951_ vdd gnd FILL
XFILL_3__1125_ vdd gnd FILL
XFILL_0__1416_ vdd gnd FILL
X_1073_ _1102_/B _1073_/B _1102_/A _1079_/A vdd gnd OAI21X1
XFILL_0__1347_ vdd gnd FILL
XFILL_0__1278_ vdd gnd FILL
XFILL_3__1056_ vdd gnd FILL
X_1409_ _956_/B Cin[5] _1502_/A vdd gnd NAND2X1
XFILL_1__1525_ vdd gnd FILL
XFILL_1__1456_ vdd gnd FILL
XFILL_4__1096_ vdd gnd FILL
XFILL_1__1387_ vdd gnd FILL
XFILL_2__1634_ vdd gnd FILL
XFILL_2__1565_ vdd gnd FILL
XFILL_2__1703_ vdd gnd FILL
X_922_ _927_/A _957_/A _923_/A vdd gnd NOR2X1
XFILL_2__1496_ vdd gnd FILL
XFILL_0__1201_ vdd gnd FILL
X_1691_ _1708_/C _1691_/B _1691_/C _1705_/A vdd gnd NAND3X1
X_1760_ _1776_/A _1776_/B _1760_/C _1763_/A vdd gnd NAND3X1
XFILL_0__1132_ vdd gnd FILL
XFILL_0__1063_ vdd gnd FILL
XFILL_3__1674_ vdd gnd FILL
XFILL_3__1743_ vdd gnd FILL
XFILL_3__1812_ vdd gnd FILL
XFILL_1__934_ vdd gnd FILL
X_1125_ Cin[3] _1533_/B vdd gnd INVX2
XFILL_1__1310_ vdd gnd FILL
XFILL_1__1241_ vdd gnd FILL
XFILL_3__1108_ vdd gnd FILL
X_1056_ _1056_/A _1093_/B _1056_/C _1093_/A vdd gnd NAND3X1
XFILL_1__1172_ vdd gnd FILL
X_1889_ _1889_/D _1897_/CLK _1889_/Q vdd gnd DFFPOSX1
XFILL_3__1039_ vdd gnd FILL
XFILL101250x15750 vdd gnd FILL
XFILL_1__1508_ vdd gnd FILL
XFILL_1__1439_ vdd gnd FILL
XFILL_2__1350_ vdd gnd FILL
XFILL_2__1281_ vdd gnd FILL
XFILL_0__952_ vdd gnd FILL
XFILL_1_CLKBUF1_insert8 vdd gnd FILL
XFILL_0__1681_ vdd gnd FILL
XFILL_2__1548_ vdd gnd FILL
XFILL_2__1617_ vdd gnd FILL
XFILL_0__1750_ vdd gnd FILL
XFILL_3__1390_ vdd gnd FILL
XFILL_2__1479_ vdd gnd FILL
X_1674_ _1723_/B _1824_/A _1710_/B vdd gnd XOR2X1
X_1743_ _1771_/C _1771_/A _1747_/B vdd gnd AND2X2
X_1812_ _1839_/B _1815_/B _1812_/C _1888_/D vdd gnd OAI21X1
XFILL_0__1115_ vdd gnd FILL
XFILL_0__1046_ vdd gnd FILL
XFILL_3__1726_ vdd gnd FILL
XFILL_3__1657_ vdd gnd FILL
XFILL_1__1790_ vdd gnd FILL
XFILL_3__1588_ vdd gnd FILL
X_1108_ _1173_/C _1173_/A _1113_/C _1131_/A vdd gnd NAND3X1
X_1039_ Cin[1] _1044_/B vdd gnd INVX1
XFILL_1__1155_ vdd gnd FILL
XFILL_1__1224_ vdd gnd FILL
XFILL101250x27450 vdd gnd FILL
XFILL_1__1086_ vdd gnd FILL
XFILL_4__1835_ vdd gnd FILL
XFILL_2__1402_ vdd gnd FILL
XFILL_2__1333_ vdd gnd FILL
XFILL_2__1195_ vdd gnd FILL
XFILL_2__1264_ vdd gnd FILL
XFILL_0__935_ vdd gnd FILL
XFILL_0__1733_ vdd gnd FILL
XFILL_3__1511_ vdd gnd FILL
XFILL_0__1802_ vdd gnd FILL
X_1390_ _1396_/C _1391_/B vdd gnd INVX1
XFILL_3__1373_ vdd gnd FILL
XFILL_0__1664_ vdd gnd FILL
XFILL_0__1595_ vdd gnd FILL
XFILL_3__1442_ vdd gnd FILL
X_1726_ _1726_/A _1759_/A _1729_/A vdd gnd NAND2X1
XFILL_4__1620_ vdd gnd FILL
X_1588_ _1661_/A _1658_/B vdd gnd INVX1
X_1657_ _952_/A Cin[6] _1794_/B vdd gnd AND2X2
XFILL_0__1029_ vdd gnd FILL
XFILL_1__1842_ vdd gnd FILL
XFILL_1__1911_ vdd gnd FILL
XFILL_3__1709_ vdd gnd FILL
XFILL_1__1773_ vdd gnd FILL
XFILL101250x39150 vdd gnd FILL
XFILL_1__1207_ vdd gnd FILL
XFILL_1__1138_ vdd gnd FILL
XFILL_1__1069_ vdd gnd FILL
XFILL_4__1749_ vdd gnd FILL
XFILL_3__931_ vdd gnd FILL
XFILL_2__1316_ vdd gnd FILL
XFILL_0__1380_ vdd gnd FILL
XFILL_2__1178_ vdd gnd FILL
XFILL_2__1247_ vdd gnd FILL
X_1442_ _1515_/D _1515_/C _1511_/C _1453_/A vdd gnd NAND3X1
X_1511_ _1511_/A _1511_/B _1511_/C _1520_/C vdd gnd OAI21X1
X_1373_ _1402_/B _1474_/C _1402_/A _1379_/A vdd gnd AOI21X1
XFILL_0__1716_ vdd gnd FILL
XFILL_3__1425_ vdd gnd FILL
XFILL_0__1578_ vdd gnd FILL
XFILL_0__1647_ vdd gnd FILL
XFILL_3__1356_ vdd gnd FILL
XFILL_3__1287_ vdd gnd FILL
XFILL_4__1603_ vdd gnd FILL
X_1709_ _1709_/A _1709_/B _1748_/B vdd gnd NAND2X1
XFILL_4__1534_ vdd gnd FILL
XFILL_1__1825_ vdd gnd FILL
XFILL_1__1687_ vdd gnd FILL
XFILL_1__1756_ vdd gnd FILL
XFILL_4__1465_ vdd gnd FILL
XFILL_2__1032_ vdd gnd FILL
XFILL_2__1101_ vdd gnd FILL
XFILL_2__1796_ vdd gnd FILL
XFILL100050x31350 vdd gnd FILL
XFILL_0__1501_ vdd gnd FILL
XFILL_0__1432_ vdd gnd FILL
XFILL_0__1363_ vdd gnd FILL
XFILL_3__1210_ vdd gnd FILL
XFILL_3__1141_ vdd gnd FILL
XFILL_0__1294_ vdd gnd FILL
XFILL_3__1072_ vdd gnd FILL
XFILL_1_BUFX2_insert24 vdd gnd FILL
X_1425_ _1425_/A _1519_/A _1425_/C _1428_/A vdd gnd OAI21X1
XFILL_1_BUFX2_insert13 vdd gnd FILL
XFILL_1__1541_ vdd gnd FILL
XFILL_1__1610_ vdd gnd FILL
XFILL_1__1472_ vdd gnd FILL
XFILL_3__1408_ vdd gnd FILL
X_1356_ _1460_/C _1524_/B _1460_/A _1461_/C vdd gnd NAND3X1
X_1287_ _1287_/A _1287_/B _1287_/C _1395_/B vdd gnd NAND3X1
XFILL_3__1339_ vdd gnd FILL
XFILL_2__932_ vdd gnd FILL
XFILL_2__1650_ vdd gnd FILL
XFILL_2__1581_ vdd gnd FILL
XFILL_1__1808_ vdd gnd FILL
XFILL100050x4050 vdd gnd FILL
XFILL_1__1739_ vdd gnd FILL
XFILL_4__1448_ vdd gnd FILL
XFILL_4__1379_ vdd gnd FILL
XFILL_2__1015_ vdd gnd FILL
XFILL_3__1690_ vdd gnd FILL
XFILL_2__1848_ vdd gnd FILL
XFILL_1__950_ vdd gnd FILL
XFILL_2__1917_ vdd gnd FILL
XFILL_2__1779_ vdd gnd FILL
X_998_ _998_/A _998_/B _998_/C _998_/Y vdd gnd OAI21X1
X_1210_ _1290_/C _1213_/D _1210_/C _1217_/C vdd gnd NAND3X1
X_1141_ _1141_/A _1141_/B _1141_/C _1206_/A vdd gnd NAND3X1
X_1072_ _956_/B _1104_/B _1901_/Q _1102_/B vdd gnd AOI21X1
XFILL_0__1346_ vdd gnd FILL
XFILL_0__1415_ vdd gnd FILL
XFILL_3__1055_ vdd gnd FILL
XFILL_3__1124_ vdd gnd FILL
XFILL_0__1277_ vdd gnd FILL
X_1408_ _1413_/C _1507_/A _1499_/B vdd gnd NAND2X1
XFILL_1__1524_ vdd gnd FILL
XFILL_1__1455_ vdd gnd FILL
X_1339_ _1460_/C _1357_/C vdd gnd INVX1
XFILL_4__1233_ vdd gnd FILL
XFILL_4__1164_ vdd gnd FILL
XFILL_1__1386_ vdd gnd FILL
XFILL_2__1702_ vdd gnd FILL
XFILL_2__1633_ vdd gnd FILL
XFILL_2__1564_ vdd gnd FILL
XFILL_2__1495_ vdd gnd FILL
XFILL_0__1200_ vdd gnd FILL
X_1690_ _1694_/C _1694_/B _1694_/A _1708_/C vdd gnd NAND3X1
XFILL_3__1811_ vdd gnd FILL
XFILL_0__1131_ vdd gnd FILL
XFILL_0__1062_ vdd gnd FILL
XFILL_3__1742_ vdd gnd FILL
XFILL_3__1673_ vdd gnd FILL
XFILL_1__933_ vdd gnd FILL
X_1055_ _1065_/A _1056_/A vdd gnd INVX1
X_1124_ _1847_/B _1533_/D _1124_/C _1127_/B vdd gnd OAI21X1
XFILL_0__1329_ vdd gnd FILL
XFILL_1__1240_ vdd gnd FILL
XFILL_3__1107_ vdd gnd FILL
XFILL_1__1171_ vdd gnd FILL
XFILL_3__1038_ vdd gnd FILL
X_1888_ _1888_/D _1897_/CLK _1888_/Q vdd gnd DFFPOSX1
XFILL_1__1507_ vdd gnd FILL
XFILL_1__1438_ vdd gnd FILL
XFILL_1__1369_ vdd gnd FILL
XFILL_2__1280_ vdd gnd FILL
XFILL_0__951_ vdd gnd FILL
XFILL_1_CLKBUF1_insert9 vdd gnd FILL
XFILL_4__1078_ vdd gnd FILL
XFILL_0__1680_ vdd gnd FILL
XFILL_2__1547_ vdd gnd FILL
XFILL_2__1616_ vdd gnd FILL
XFILL_2__1478_ vdd gnd FILL
X_1811_ _1888_/Q _1815_/B _1812_/C vdd gnd NAND2X1
XFILL_0__1114_ vdd gnd FILL
X_1742_ _1742_/A _1742_/B _1771_/C vdd gnd NAND2X1
X_1673_ _1893_/Q _1824_/A vdd gnd INVX1
XFILL_0__1045_ vdd gnd FILL
XFILL_3__1587_ vdd gnd FILL
XFILL_3__1725_ vdd gnd FILL
XFILL_3__1656_ vdd gnd FILL
XFILL_1__1223_ vdd gnd FILL
X_1107_ _956_/B Cin[1] _1173_/A vdd gnd NAND2X1
X_1038_ _950_/B _1845_/B vdd gnd INVX1
XFILL_1__1154_ vdd gnd FILL
XFILL_1__1085_ vdd gnd FILL
XFILL_2__1332_ vdd gnd FILL
XFILL_2__1401_ vdd gnd FILL
XFILL_0__934_ vdd gnd FILL
XFILL_2__1194_ vdd gnd FILL
XFILL_2__1263_ vdd gnd FILL
XFILL_0__1732_ vdd gnd FILL
XFILL_3__1510_ vdd gnd FILL
XFILL_3__1441_ vdd gnd FILL
XFILL_0__1801_ vdd gnd FILL
XFILL_0__1594_ vdd gnd FILL
XFILL_0__1663_ vdd gnd FILL
XFILL_3__1372_ vdd gnd FILL
X_1725_ _1725_/A _1725_/B _1759_/A vdd gnd OR2X2
X_1587_ _1652_/B _1594_/A vdd gnd INVX1
X_1656_ _1711_/B _1666_/B vdd gnd INVX1
XFILL_1__1772_ vdd gnd FILL
XFILL_0__1028_ vdd gnd FILL
XFILL_1__1841_ vdd gnd FILL
XFILL_3__1708_ vdd gnd FILL
XFILL_3__1639_ vdd gnd FILL
XFILL_1__1206_ vdd gnd FILL
XFILL_4__1817_ vdd gnd FILL
XFILL_1__1137_ vdd gnd FILL
XFILL_1__1068_ vdd gnd FILL
XFILL_3__930_ vdd gnd FILL
XFILL_2__1315_ vdd gnd FILL
XFILL100650x85950 vdd gnd FILL
XFILL_2__1246_ vdd gnd FILL
XFILL_2__1177_ vdd gnd FILL
X_1510_ _1510_/A _1510_/B _1511_/B vdd gnd AND2X2
X_1441_ _963_/A _1533_/D _1510_/A _1515_/C vdd gnd OAI21X1
XFILL_0__1646_ vdd gnd FILL
XFILL_0__1715_ vdd gnd FILL
XFILL_3__1424_ vdd gnd FILL
X_1372_ _1372_/A _1372_/B _1372_/C _1397_/C vdd gnd OAI21X1
XFILL_0__1577_ vdd gnd FILL
XFILL_3__1355_ vdd gnd FILL
XFILL_3__1286_ vdd gnd FILL
X_1708_ _1708_/A _1708_/B _1708_/C _1740_/A vdd gnd OAI21X1
X_1639_ _1705_/B _1639_/B _1703_/B vdd gnd NAND2X1
XFILL_1__1755_ vdd gnd FILL
XFILL_1__1824_ vdd gnd FILL
XFILL_1__1686_ vdd gnd FILL
XFILL_2__1031_ vdd gnd FILL
XFILL_2__1100_ vdd gnd FILL
XFILL_3_BUFX2_insert0 vdd gnd FILL
XFILL100350x15750 vdd gnd FILL
XFILL_0__1500_ vdd gnd FILL
XFILL_2__1795_ vdd gnd FILL
XFILL_0__1431_ vdd gnd FILL
XFILL_0__1362_ vdd gnd FILL
XFILL_3__1071_ vdd gnd FILL
XFILL_3__1140_ vdd gnd FILL
XFILL_2__1229_ vdd gnd FILL
XFILL_0__1293_ vdd gnd FILL
XFILL_1_BUFX2_insert25 vdd gnd FILL
X_1355_ _1355_/A _1355_/B _1431_/A vdd gnd AND2X2
X_1424_ _1424_/A _1519_/A vdd gnd INVX1
XFILL_1_BUFX2_insert14 vdd gnd FILL
XFILL_0__1629_ vdd gnd FILL
XFILL_1__1540_ vdd gnd FILL
XFILL_1__1471_ vdd gnd FILL
XFILL_3__1407_ vdd gnd FILL
XFILL_3__1338_ vdd gnd FILL
X_1286_ _1298_/A _1383_/C _1298_/B _1287_/B vdd gnd NAND3X1
XFILL_2__931_ vdd gnd FILL
XFILL_3__1269_ vdd gnd FILL
XFILL_1__1738_ vdd gnd FILL
XFILL_2__1580_ vdd gnd FILL
XFILL_4__1516_ vdd gnd FILL
XFILL_1__1807_ vdd gnd FILL
XFILL_1__1669_ vdd gnd FILL
XFILL_2__1014_ vdd gnd FILL
XFILL100350x27450 vdd gnd FILL
XFILL100950x74250 vdd gnd FILL
X_997_ _998_/A _997_/B _998_/C vdd gnd NAND2X1
XFILL_2__1916_ vdd gnd FILL
XFILL_2__1847_ vdd gnd FILL
XFILL_2__1778_ vdd gnd FILL
X_1071_ _1102_/C _1073_/B vdd gnd INVX1
X_1140_ _1140_/A _1140_/B _1140_/C _1141_/C vdd gnd AOI21X1
XFILL_0__1345_ vdd gnd FILL
XFILL_0__1414_ vdd gnd FILL
XFILL_0__1276_ vdd gnd FILL
XFILL_3__1054_ vdd gnd FILL
XFILL_3__1123_ vdd gnd FILL
X_1407_ _956_/B Cin[5] _1507_/A vdd gnd AND2X2
X_1338_ _1338_/A _1338_/B _1338_/C _1460_/C vdd gnd OAI21X1
XFILL_4__1301_ vdd gnd FILL
XFILL_1__1523_ vdd gnd FILL
XFILL_1__1454_ vdd gnd FILL
X_1269_ _1269_/A _1269_/B _1361_/A _1274_/A vdd gnd AOI21X1
XFILL_1__1385_ vdd gnd FILL
XFILL_2__1701_ vdd gnd FILL
XFILL_2__1632_ vdd gnd FILL
XFILL_2__1563_ vdd gnd FILL
XFILL_2__1494_ vdd gnd FILL
XFILL100350x39150 vdd gnd FILL
XFILL_0__1130_ vdd gnd FILL
XFILL_3__1741_ vdd gnd FILL
XFILL_3__1810_ vdd gnd FILL
XFILL_0__1061_ vdd gnd FILL
XFILL_3__1672_ vdd gnd FILL
XFILL_1__932_ vdd gnd FILL
X_1054_ _947_/B Cin[2] _1065_/A vdd gnd NAND2X1
X_1123_ _1123_/A _1123_/B _1123_/C _1159_/C vdd gnd NAND3X1
X_1887_ _1887_/D _1897_/CLK _1887_/Q vdd gnd DFFPOSX1
XFILL_0__1328_ vdd gnd FILL
XFILL_3__1037_ vdd gnd FILL
XFILL_1__1170_ vdd gnd FILL
XFILL_0__1259_ vdd gnd FILL
XFILL_3__1106_ vdd gnd FILL
XFILL_4__1781_ vdd gnd FILL
XFILL_1__1506_ vdd gnd FILL
XFILL_1__1437_ vdd gnd FILL
XFILL_1__1368_ vdd gnd FILL
XFILL_4__1146_ vdd gnd FILL
XFILL_4__1215_ vdd gnd FILL
XFILL_0__950_ vdd gnd FILL
XFILL_1__1299_ vdd gnd FILL
XFILL_2__1615_ vdd gnd FILL
XFILL_2__1546_ vdd gnd FILL
XFILL_2__1477_ vdd gnd FILL
X_1741_ _1741_/A _1741_/B _1742_/B vdd gnd NAND2X1
X_1810_ Yin[2] _1839_/B vdd gnd INVX1
XFILL_0__1113_ vdd gnd FILL
X_1672_ _1679_/C _1679_/B _1679_/A _1678_/B vdd gnd AOI21X1
XFILL_3__1724_ vdd gnd FILL
XFILL_0__1044_ vdd gnd FILL
XFILL_3__1586_ vdd gnd FILL
XFILL_3__1655_ vdd gnd FILL
X_1106_ _946_/A _1106_/B _1894_/Q _1173_/C vdd gnd NAND3X1
XFILL_4__1000_ vdd gnd FILL
XFILL_1__1222_ vdd gnd FILL
XFILL_4__988_ vdd gnd FILL
XFILL_1__1153_ vdd gnd FILL
X_1037_ _1062_/C _1048_/A vdd gnd INVX1
XFILL_1__1084_ vdd gnd FILL
XFILL_4__1695_ vdd gnd FILL
XFILL_4__1764_ vdd gnd FILL
XFILL_2__1400_ vdd gnd FILL
XFILL_2__1331_ vdd gnd FILL
XFILL_2__1262_ vdd gnd FILL
XFILL_0__933_ vdd gnd FILL
XFILL_4__1129_ vdd gnd FILL
XFILL_2__1193_ vdd gnd FILL
XFILL_0__1731_ vdd gnd FILL
XFILL_0__1662_ vdd gnd FILL
XFILL_3__1440_ vdd gnd FILL
XFILL_0__1800_ vdd gnd FILL
XFILL_3__1371_ vdd gnd FILL
XFILL_0__1593_ vdd gnd FILL
XFILL_2__1529_ vdd gnd FILL
X_1724_ _1725_/B _1725_/A _1726_/A vdd gnd NAND2X1
XFILL_0__1027_ vdd gnd FILL
X_1586_ _1652_/A _1594_/B vdd gnd INVX1
XFILL_1__1771_ vdd gnd FILL
X_1655_ _949_/A Cin[6] _952_/A Cin[5] _1711_/B vdd gnd AOI22X1
XFILL_3__1707_ vdd gnd FILL
XFILL_4__1480_ vdd gnd FILL
XFILL_1__1840_ vdd gnd FILL
XFILL_3__1638_ vdd gnd FILL
XFILL_3__1569_ vdd gnd FILL
XFILL_1__1205_ vdd gnd FILL
XFILL_1__1136_ vdd gnd FILL
XFILL_1__1067_ vdd gnd FILL
XFILL_2__1314_ vdd gnd FILL
XFILL_2__1245_ vdd gnd FILL
XFILL_2__1176_ vdd gnd FILL
X_1440_ _1515_/A _1611_/A _1511_/C vdd gnd NAND2X1
X_1371_ _1371_/A _1371_/B _1371_/C _1372_/A vdd gnd AOI21X1
XFILL_0__1645_ vdd gnd FILL
XFILL_0__1714_ vdd gnd FILL
XFILL_3__1423_ vdd gnd FILL
XFILL_3__1354_ vdd gnd FILL
XFILL_3__989_ vdd gnd FILL
XFILL_0__1576_ vdd gnd FILL
XFILL_3__1285_ vdd gnd FILL
X_1638_ _1638_/A _1638_/B _1638_/C _1639_/B vdd gnd OAI21X1
X_1707_ _1772_/B _1772_/A _1747_/A vdd gnd NAND2X1
XFILL_1__1685_ vdd gnd FILL
X_1569_ _1702_/B _1569_/B _1569_/C _1879_/D vdd gnd OAI21X1
XFILL_1__1754_ vdd gnd FILL
XFILL_1__1823_ vdd gnd FILL
XFILL_4__1394_ vdd gnd FILL
XFILL_2__1030_ vdd gnd FILL
XFILL_3_BUFX2_insert1 vdd gnd FILL
XFILL_1__1119_ vdd gnd FILL
XFILL_2__1794_ vdd gnd FILL
XFILL_0__1430_ vdd gnd FILL
XFILL_0__1361_ vdd gnd FILL
XFILL_0__1292_ vdd gnd FILL
XFILL_3__1070_ vdd gnd FILL
XFILL_2__1228_ vdd gnd FILL
XFILL_2__1159_ vdd gnd FILL
X_1423_ _1423_/A _1423_/B _1423_/C _1468_/A vdd gnd NAND3X1
X_1354_ _1461_/A _1363_/B _1363_/A _1473_/B vdd gnd NAND3X1
XFILL_1_BUFX2_insert15 vdd gnd FILL
X_1285_ _1285_/A _1285_/B _1285_/C _1298_/B vdd gnd OAI21X1
XFILL_0__1628_ vdd gnd FILL
XFILL_0__1559_ vdd gnd FILL
XFILL_1__1470_ vdd gnd FILL
XFILL_3__1337_ vdd gnd FILL
XFILL_3__1406_ vdd gnd FILL
XFILL_2__930_ vdd gnd FILL
XFILL_3__1199_ vdd gnd FILL
XFILL_3__1268_ vdd gnd FILL
XFILL_1__1668_ vdd gnd FILL
XFILL_1__1737_ vdd gnd FILL
XFILL_1__1806_ vdd gnd FILL
XFILL_1__1599_ vdd gnd FILL
XFILL_2__1013_ vdd gnd FILL
XFILL_2__1777_ vdd gnd FILL
X_996_ _996_/A _996_/B _996_/C _996_/Y vdd gnd OAI21X1
XFILL_2__1915_ vdd gnd FILL
XFILL_2__1846_ vdd gnd FILL
XFILL_0__1413_ vdd gnd FILL
X_1070_ _956_/B _1104_/B _1901_/Q _1102_/C vdd gnd NAND3X1
XFILL_3__1122_ vdd gnd FILL
XFILL_0__1275_ vdd gnd FILL
XFILL_0__1344_ vdd gnd FILL
XFILL_3__1053_ vdd gnd FILL
XFILL_1__1522_ vdd gnd FILL
X_1337_ _1355_/B _1355_/A _1461_/A vdd gnd NAND2X1
X_1406_ _953_/B Cin[6] _1413_/C vdd gnd AND2X2
X_1268_ _1361_/C _1325_/B _1325_/A _1274_/B vdd gnd AOI21X1
XFILL_1__1453_ vdd gnd FILL
X_1199_ _1203_/A _1203_/B _1277_/C _1208_/A vdd gnd OAI21X1
XFILL_4__1093_ vdd gnd FILL
XFILL_1__1384_ vdd gnd FILL
XFILL_2__1631_ vdd gnd FILL
XFILL_2__1700_ vdd gnd FILL
XFILL_2__1562_ vdd gnd FILL
XFILL_2__1493_ vdd gnd FILL
XFILL_0__1060_ vdd gnd FILL
XFILL_3__1740_ vdd gnd FILL
XFILL_3__1671_ vdd gnd FILL
XFILL_1__931_ vdd gnd FILL
XFILL_2__1829_ vdd gnd FILL
X_979_ _983_/A _979_/B _980_/C vdd gnd NAND2X1
X_1122_ _1847_/B _1533_/D _1159_/A _1123_/A vdd gnd OAI21X1
XFILL_3__1105_ vdd gnd FILL
X_1053_ _1843_/B _1533_/D _1053_/C _1058_/C vdd gnd OAI21X1
X_1886_ _1886_/D _1897_/CLK _1886_/Q vdd gnd DFFPOSX1
XFILL_0__1327_ vdd gnd FILL
XFILL_0__1258_ vdd gnd FILL
XFILL_0__1189_ vdd gnd FILL
XFILL_3__1036_ vdd gnd FILL
XFILL_1__1505_ vdd gnd FILL
XFILL_1__1436_ vdd gnd FILL
XFILL_1__1367_ vdd gnd FILL
XFILL_1__1298_ vdd gnd FILL
XFILL_2__1545_ vdd gnd FILL
XFILL_2__1614_ vdd gnd FILL
XFILL_2__1476_ vdd gnd FILL
X_1740_ _1740_/A _1742_/A vdd gnd INVX1
X_1671_ _1671_/A _1671_/B _1671_/C _1679_/B vdd gnd NAND3X1
XFILL_0__1112_ vdd gnd FILL
XFILL_0__1043_ vdd gnd FILL
XFILL_3__1654_ vdd gnd FILL
XFILL_3__1723_ vdd gnd FILL
XFILL_3__1585_ vdd gnd FILL
X_1105_ _1173_/B _1113_/C vdd gnd INVX1
XFILL_1__1221_ vdd gnd FILL
XFILL_1__1152_ vdd gnd FILL
X_1036_ _1036_/A _1036_/B _1036_/C _1062_/C vdd gnd OAI21X1
X_1869_ _1869_/D _1885_/CLK _943_/B vdd gnd DFFPOSX1
XFILL_4__1832_ vdd gnd FILL
XFILL_3__1019_ vdd gnd FILL
XFILL_1__1083_ vdd gnd FILL
XFILL_1__1419_ vdd gnd FILL
XFILL_2__1330_ vdd gnd FILL
XFILL_2__1261_ vdd gnd FILL
XFILL_0__932_ vdd gnd FILL
XFILL100650x4050 vdd gnd FILL
XFILL_2__1192_ vdd gnd FILL
XFILL_0__1730_ vdd gnd FILL
XFILL_0__1661_ vdd gnd FILL
XFILL_0__1592_ vdd gnd FILL
XFILL_2__1528_ vdd gnd FILL
XFILL_3__1370_ vdd gnd FILL
XFILL_2__1459_ vdd gnd FILL
X_1654_ _1711_/A _1666_/C vdd gnd INVX1
X_1723_ _1893_/Q _1723_/B _1725_/A vdd gnd NAND2X1
XFILL99750x46950 vdd gnd FILL
XFILL_0__1026_ vdd gnd FILL
XFILL_3__1637_ vdd gnd FILL
X_1585_ _1652_/A _1652_/B _1595_/B _1601_/A vdd gnd NOR3X1
XFILL_3__1706_ vdd gnd FILL
XFILL_1__1770_ vdd gnd FILL
XFILL_3__1568_ vdd gnd FILL
XFILL_3__1499_ vdd gnd FILL
X_1019_ _950_/B _1106_/B _1899_/Q _1036_/B vdd gnd AOI21X1
XFILL_1__1204_ vdd gnd FILL
XFILL_1__1135_ vdd gnd FILL
XFILL_1__1066_ vdd gnd FILL
XFILL_4__1746_ vdd gnd FILL
XFILL_4__1677_ vdd gnd FILL
XFILL_2__1313_ vdd gnd FILL
XFILL_2__1175_ vdd gnd FILL
XFILL_2__1244_ vdd gnd FILL
XFILL_0__1713_ vdd gnd FILL
XFILL_3__988_ vdd gnd FILL
X_1370_ _1397_/A _1397_/B _1379_/C _1385_/C vdd gnd NAND3X1
XFILL_0__1575_ vdd gnd FILL
XFILL_0__1644_ vdd gnd FILL
XFILL_3__1353_ vdd gnd FILL
XFILL_3__1422_ vdd gnd FILL
XFILL_3__1284_ vdd gnd FILL
X_1637_ _1637_/A _1637_/B _1646_/A _1638_/B vdd gnd AOI21X1
XFILL_4__1600_ vdd gnd FILL
XFILL_1__1822_ vdd gnd FILL
X_1706_ _1706_/A _1706_/B _1706_/C _1706_/D _1772_/A vdd gnd AOI22X1
XFILL_0__1009_ vdd gnd FILL
XFILL_1__1684_ vdd gnd FILL
XFILL_4__1531_ vdd gnd FILL
XFILL_4__1462_ vdd gnd FILL
XFILL_1__1753_ vdd gnd FILL
X_1568_ _993_/B _1702_/B _1569_/C vdd gnd NAND2X1
X_1499_ _1519_/C _1499_/B _1517_/A vdd gnd AND2X2
XFILL101250x11850 vdd gnd FILL
XFILL_3_BUFX2_insert2 vdd gnd FILL
XFILL_1__1118_ vdd gnd FILL
XFILL_1__1049_ vdd gnd FILL
XFILL_2__1793_ vdd gnd FILL
XFILL_0__1360_ vdd gnd FILL
XFILL_0__1291_ vdd gnd FILL
XFILL_2__1227_ vdd gnd FILL
XFILL_2__1158_ vdd gnd FILL
X_1422_ _1519_/C _1426_/B _1427_/C _1423_/B vdd gnd NAND3X1
XFILL_2__1089_ vdd gnd FILL
X_1353_ _1357_/A _1357_/B _1460_/C _1363_/A vdd gnd OAI21X1
XFILL_3__1405_ vdd gnd FILL
XFILL_1_BUFX2_insert16 vdd gnd FILL
X_1284_ _1382_/C _1382_/B _1382_/A _1383_/C vdd gnd NAND3X1
XFILL_0__1627_ vdd gnd FILL
XFILL_0__1558_ vdd gnd FILL
XFILL_0__1489_ vdd gnd FILL
XFILL_3__1336_ vdd gnd FILL
XFILL_3__1267_ vdd gnd FILL
XFILL_3__1198_ vdd gnd FILL
XFILL_1__1805_ vdd gnd FILL
XFILL101250x23550 vdd gnd FILL
XFILL_1__1667_ vdd gnd FILL
XFILL_1__1736_ vdd gnd FILL
XFILL_1__1598_ vdd gnd FILL
XFILL_4__1445_ vdd gnd FILL
XFILL_4__1376_ vdd gnd FILL
XFILL_2__989_ vdd gnd FILL
XFILL_2__1012_ vdd gnd FILL
XFILL_2__1914_ vdd gnd FILL
XFILL_2__1776_ vdd gnd FILL
X_995_ _996_/A _995_/B _996_/C vdd gnd NAND2X1
XFILL_2__1845_ vdd gnd FILL
XFILL_0__1343_ vdd gnd FILL
XFILL_0__1412_ vdd gnd FILL
XFILL_3__1121_ vdd gnd FILL
XFILL_0__1274_ vdd gnd FILL
XFILL_3__1052_ vdd gnd FILL
X_1405_ _1418_/A _1419_/B vdd gnd INVX1
XFILL_1__1521_ vdd gnd FILL
XFILL_1__1452_ vdd gnd FILL
X_1336_ _1421_/A _1421_/B _1416_/C _1355_/A vdd gnd NAND3X1
X_1198_ _1198_/A _1198_/B _1267_/A _1203_/A vdd gnd AOI21X1
XFILL_4__1161_ vdd gnd FILL
X_1267_ _1267_/A _1267_/B _1267_/C _1371_/C vdd gnd OAI21X1
XFILL_4__1230_ vdd gnd FILL
XFILL_3__1319_ vdd gnd FILL
XFILL_1__1383_ vdd gnd FILL
XFILL101250x35250 vdd gnd FILL
XFILL_2__1630_ vdd gnd FILL
XFILL_2__1561_ vdd gnd FILL
XFILL_1__1719_ vdd gnd FILL
XFILL_2__1492_ vdd gnd FILL
XFILL_2_CLKBUF1_insert5 vdd gnd FILL
XFILL_3__1670_ vdd gnd FILL
XFILL_1__930_ vdd gnd FILL
XFILL_2__1759_ vdd gnd FILL
X_978_ _978_/A _980_/B vdd gnd INVX1
XFILL_2__1828_ vdd gnd FILL
X_1121_ _953_/B _1847_/B vdd gnd INVX2
X_1052_ _1093_/B _1056_/C _1053_/C vdd gnd NAND2X1
XFILL_0__1326_ vdd gnd FILL
XFILL_3__1035_ vdd gnd FILL
XFILL_3__1104_ vdd gnd FILL
X_1885_ _1885_/D _1885_/CLK _1885_/Q vdd gnd DFFPOSX1
XFILL_4_BUFX2_insert20 vdd gnd FILL
XFILL_0__1257_ vdd gnd FILL
XFILL_0__1188_ vdd gnd FILL
XFILL_3__1799_ vdd gnd FILL
XFILL_1__1504_ vdd gnd FILL
XFILL_1__1435_ vdd gnd FILL
X_1319_ _1319_/A _1319_/B _1319_/C _1366_/A vdd gnd NAND3X1
XFILL_1__1366_ vdd gnd FILL
XFILL_1__1297_ vdd gnd FILL
XFILL_4__1075_ vdd gnd FILL
XFILL_2__1544_ vdd gnd FILL
XFILL_2__1613_ vdd gnd FILL
XFILL_2__1475_ vdd gnd FILL
X_1670_ _1720_/B _1670_/B _1670_/C _1679_/C vdd gnd OAI21X1
XFILL_0__1111_ vdd gnd FILL
XFILL_0__1042_ vdd gnd FILL
XFILL_3__1653_ vdd gnd FILL
XFILL_3__1584_ vdd gnd FILL
XFILL_3__1722_ vdd gnd FILL
X_1035_ Cin[2] _1533_/D vdd gnd INVX4
X_1104_ _946_/A _1104_/B _1894_/Q _1173_/B vdd gnd AOI21X1
XFILL_0__1309_ vdd gnd FILL
XFILL_3__1018_ vdd gnd FILL
XFILL_1__1220_ vdd gnd FILL
XFILL_1__1082_ vdd gnd FILL
XFILL_1__1151_ vdd gnd FILL
X_1799_ _1799_/A _1799_/B _1799_/C _1800_/A vdd gnd NAND3X1
X_1868_ _1868_/D _1910_/CLK _938_/B vdd gnd DFFPOSX1
XFILL_1__1349_ vdd gnd FILL
XFILL_1__1418_ vdd gnd FILL
XFILL_0__931_ vdd gnd FILL
XFILL_2__1191_ vdd gnd FILL
XFILL_2__1260_ vdd gnd FILL
XFILL_0__1660_ vdd gnd FILL
XFILL_0__1591_ vdd gnd FILL
XFILL_2__1458_ vdd gnd FILL
XFILL_2__1527_ vdd gnd FILL
XFILL_2__1389_ vdd gnd FILL
X_1653_ _946_/A Cin[7] _1711_/A vdd gnd NAND2X1
X_1584_ _1584_/A _1661_/A _1595_/B vdd gnd NOR2X1
X_1722_ _1886_/Q _1725_/B vdd gnd INVX1
XFILL_0__1025_ vdd gnd FILL
XFILL_3__1636_ vdd gnd FILL
XFILL_3__1705_ vdd gnd FILL
XFILL_3__1567_ vdd gnd FILL
XFILL_0__1789_ vdd gnd FILL
XFILL_3__1498_ vdd gnd FILL
X_1018_ _1216_/A _1018_/B _1018_/C _1870_/D vdd gnd OAI21X1
XFILL_1__1203_ vdd gnd FILL
XFILL101250x4050 vdd gnd FILL
XFILL_1__1134_ vdd gnd FILL
XFILL_1__1065_ vdd gnd FILL
XFILL_4__1814_ vdd gnd FILL
XFILL_2__1312_ vdd gnd FILL
XFILL_2__1174_ vdd gnd FILL
XFILL_2__1243_ vdd gnd FILL
XFILL_0__1712_ vdd gnd FILL
XFILL_3__1421_ vdd gnd FILL
XFILL_3__987_ vdd gnd FILL
XFILL_0__1574_ vdd gnd FILL
XFILL_0__1643_ vdd gnd FILL
XFILL_3__1352_ vdd gnd FILL
XFILL_3__1283_ vdd gnd FILL
X_1705_ _1705_/A _1705_/B _1706_/B vdd gnd NAND2X1
X_1636_ _1693_/B _1692_/A _1693_/A _1638_/A vdd gnd AOI21X1
XFILL_1__1821_ vdd gnd FILL
X_1567_ _1567_/A _1572_/A _1569_/B vdd gnd XNOR2X1
XFILL_0__1008_ vdd gnd FILL
XFILL_3__1619_ vdd gnd FILL
XFILL_1__1683_ vdd gnd FILL
X_1498_ _1498_/A _1498_/B _1498_/C _1634_/C vdd gnd AOI21X1
XFILL_1__1752_ vdd gnd FILL
XFILL_3_BUFX2_insert3 vdd gnd FILL
XFILL_1__1117_ vdd gnd FILL
XFILL_1__1048_ vdd gnd FILL
XFILL_4__1659_ vdd gnd FILL
XFILL_4__1728_ vdd gnd FILL
XFILL_2__1792_ vdd gnd FILL
XFILL_2__1226_ vdd gnd FILL
XFILL_0__1290_ vdd gnd FILL
XFILL_2__1157_ vdd gnd FILL
XFILL_2__1088_ vdd gnd FILL
X_1421_ _1421_/A _1421_/B _1421_/C _1427_/C vdd gnd AOI21X1
XFILL_0__1626_ vdd gnd FILL
X_1352_ _1352_/A _1352_/B _1450_/A _1357_/B vdd gnd AOI21X1
XFILL_3__1404_ vdd gnd FILL
XFILL_1_BUFX2_insert17 vdd gnd FILL
X_1283_ _1383_/A _1298_/A vdd gnd INVX1
XFILL_0__1557_ vdd gnd FILL
XFILL_0__1488_ vdd gnd FILL
XFILL_3__1335_ vdd gnd FILL
XFILL_3__1266_ vdd gnd FILL
XFILL_3__1197_ vdd gnd FILL
X_1619_ _1687_/A _1687_/B _1645_/A vdd gnd NAND2X1
XFILL_1__1735_ vdd gnd FILL
XFILL_4__1513_ vdd gnd FILL
XFILL_1__1804_ vdd gnd FILL
XFILL_1__1666_ vdd gnd FILL
XFILL_1__1597_ vdd gnd FILL
XBUFX2_insert20 _1906_/Q _957_/A vdd gnd BUFX2
XFILL_2__1011_ vdd gnd FILL
XFILL_2__988_ vdd gnd FILL
XFILL_2__1913_ vdd gnd FILL
XFILL_2__1844_ vdd gnd FILL
XFILL_2__1775_ vdd gnd FILL
X_994_ _996_/A _994_/B _994_/C _994_/Y vdd gnd OAI21X1
XFILL_0__1411_ vdd gnd FILL
XFILL_0__1342_ vdd gnd FILL
XFILL_0__1273_ vdd gnd FILL
XFILL_3__1051_ vdd gnd FILL
XFILL_3__1120_ vdd gnd FILL
XFILL_2__1209_ vdd gnd FILL
X_1404_ _950_/B Cin[7] _1418_/A vdd gnd NAND2X1
X_1335_ _961_/A _1533_/D _1420_/A _1421_/B vdd gnd OAI21X1
XFILL_1__1520_ vdd gnd FILL
XFILL_0__1609_ vdd gnd FILL
XFILL_1__1451_ vdd gnd FILL
XFILL_3__1318_ vdd gnd FILL
XFILL_1__1382_ vdd gnd FILL
X_1266_ _1266_/A _1266_/B _1266_/C _1267_/B vdd gnd AOI21X1
X_1197_ _1267_/C _1231_/B _1231_/A _1203_/B vdd gnd AOI21X1
XFILL_3__1249_ vdd gnd FILL
XFILL_2__1560_ vdd gnd FILL
XFILL_1__1718_ vdd gnd FILL
XFILL_2__1491_ vdd gnd FILL
XFILL_4__1427_ vdd gnd FILL
XFILL_1__1649_ vdd gnd FILL
XFILL_2_CLKBUF1_insert6 vdd gnd FILL
XFILL_4__1358_ vdd gnd FILL
XCLKBUF1_insert5 clk _1885_/CLK vdd gnd CLKBUF1
XFILL_2__1827_ vdd gnd FILL
X_977_ _977_/A _977_/B _977_/C _977_/Y vdd gnd OAI21X1
XFILL_2__1689_ vdd gnd FILL
XFILL_2__1758_ vdd gnd FILL
X_1051_ _1062_/C _1062_/B _1062_/A _1093_/B vdd gnd NAND3X1
X_1120_ _1124_/C _1158_/A _1123_/C vdd gnd NAND2X1
X_1884_ _1884_/D _1885_/CLK _1884_/Q vdd gnd DFFPOSX1
XFILL_0__1256_ vdd gnd FILL
XFILL_0__1325_ vdd gnd FILL
XFILL_3__1103_ vdd gnd FILL
XFILL_3__1034_ vdd gnd FILL
XFILL_0__1187_ vdd gnd FILL
XFILL_3__1798_ vdd gnd FILL
X_1318_ _1425_/C _1320_/B _1321_/C _1319_/B vdd gnd NAND3X1
XFILL_1__989_ vdd gnd FILL
XFILL_1__1503_ vdd gnd FILL
XFILL_1__1434_ vdd gnd FILL
XFILL_1__1365_ vdd gnd FILL
XFILL_4__1212_ vdd gnd FILL
XFILL_4__1143_ vdd gnd FILL
X_1249_ _1338_/B _1249_/B _1338_/A _1360_/A vdd gnd OAI21X1
XFILL100050x7950 vdd gnd FILL
XFILL_1__1296_ vdd gnd FILL
XFILL_2__1612_ vdd gnd FILL
XFILL_2__1543_ vdd gnd FILL
XFILL_2__1474_ vdd gnd FILL
XFILL100350x11850 vdd gnd FILL
XFILL100050x46950 vdd gnd FILL
XFILL_0__1110_ vdd gnd FILL
XFILL_3__1721_ vdd gnd FILL
XFILL_0__1041_ vdd gnd FILL
XFILL_3__1652_ vdd gnd FILL
XFILL_3__1583_ vdd gnd FILL
XFILL_4_CLKBUF1_insert11 vdd gnd FILL
X_1103_ _1130_/C _1131_/C vdd gnd INVX1
X_1034_ _1034_/A _1058_/A vdd gnd INVX1
X_1867_ _1867_/D _1885_/CLK _933_/B vdd gnd DFFPOSX1
XFILL_0__1308_ vdd gnd FILL
XFILL_0__1239_ vdd gnd FILL
XFILL_4__985_ vdd gnd FILL
XFILL_3__1017_ vdd gnd FILL
XFILL_1__1081_ vdd gnd FILL
XFILL_1__1150_ vdd gnd FILL
XFILL_4__1692_ vdd gnd FILL
XFILL_4__1761_ vdd gnd FILL
X_1798_ _1798_/A _1798_/B _1801_/D vdd gnd NAND2X1
XFILL_3__1919_ vdd gnd FILL
XFILL_1__1348_ vdd gnd FILL
XFILL_1__1417_ vdd gnd FILL
XFILL_0__930_ vdd gnd FILL
XFILL_2__1190_ vdd gnd FILL
XFILL_4__1126_ vdd gnd FILL
XFILL_4__1057_ vdd gnd FILL
XFILL_1__1279_ vdd gnd FILL
XFILL100350x23550 vdd gnd FILL
XFILL_0__1590_ vdd gnd FILL
XFILL100950x70350 vdd gnd FILL
XFILL_2__1526_ vdd gnd FILL
XFILL_2__1457_ vdd gnd FILL
X_1721_ _1762_/C _1776_/A vdd gnd INVX1
XFILL_2__1388_ vdd gnd FILL
X_1652_ _1652_/A _1652_/B _1652_/C _1680_/A vdd gnd OAI21X1
X_1583_ _949_/A Cin[5] _1661_/A vdd gnd NAND2X1
XFILL_3__1704_ vdd gnd FILL
XFILL_0__1024_ vdd gnd FILL
XFILL_3__1635_ vdd gnd FILL
XFILL_3__1566_ vdd gnd FILL
XFILL_0__1788_ vdd gnd FILL
XFILL_3__1497_ vdd gnd FILL
X_1017_ _967_/A _990_/A _1018_/C vdd gnd NAND2X1
XFILL_1__1202_ vdd gnd FILL
X_1919_ _945_/Y Yout[3] vdd gnd BUFX2
XFILL_1__1133_ vdd gnd FILL
XFILL_1__1064_ vdd gnd FILL
XFILL_2__1311_ vdd gnd FILL
XFILL_2__1242_ vdd gnd FILL
XFILL_2__1173_ vdd gnd FILL
XFILL100350x35250 vdd gnd FILL
XFILL_0__1711_ vdd gnd FILL
XFILL100950x82050 vdd gnd FILL
XFILL_3__1351_ vdd gnd FILL
XFILL_0__1642_ vdd gnd FILL
XFILL_3__1420_ vdd gnd FILL
XFILL_3__986_ vdd gnd FILL
XFILL_2__1509_ vdd gnd FILL
XFILL_0__1573_ vdd gnd FILL
XFILL_0_BUFX2_insert0 vdd gnd FILL
XFILL_3__1282_ vdd gnd FILL
X_1704_ _1704_/A _1706_/C _1704_/C _1772_/B vdd gnd NAND3X1
XFILL_0__1007_ vdd gnd FILL
X_1635_ _1635_/A _1635_/B _1635_/C _1638_/C vdd gnd AOI21X1
XFILL_1__1820_ vdd gnd FILL
X_1566_ _1566_/A _1571_/C _1572_/A vdd gnd NAND2X1
X_1497_ _1552_/C _1498_/C vdd gnd INVX1
XFILL_1__1751_ vdd gnd FILL
XFILL_3__1618_ vdd gnd FILL
XFILL_1__1682_ vdd gnd FILL
XFILL_3__1549_ vdd gnd FILL
XFILL_4__1391_ vdd gnd FILL
XFILL_1__1116_ vdd gnd FILL
XFILL_3_BUFX2_insert4 vdd gnd FILL
XFILL_1__1047_ vdd gnd FILL
XFILL_2__1791_ vdd gnd FILL
XFILL_2__1225_ vdd gnd FILL
XFILL_2__1156_ vdd gnd FILL
XFILL_2__1087_ vdd gnd FILL
X_1351_ _1351_/A _1524_/A _1351_/C _1357_/A vdd gnd AOI21X1
X_1420_ _1420_/A _1420_/B _1421_/C vdd gnd NOR2X1
XFILL_1_BUFX2_insert18 vdd gnd FILL
XFILL99750x7950 vdd gnd FILL
XFILL_0__1625_ vdd gnd FILL
XFILL_3__1334_ vdd gnd FILL
XFILL_3__1403_ vdd gnd FILL
XFILL_3__969_ vdd gnd FILL
X_1282_ _1383_/A _1289_/B _1289_/A _1287_/C vdd gnd NAND3X1
XFILL_0__1556_ vdd gnd FILL
XFILL_0__1487_ vdd gnd FILL
XFILL_3__1196_ vdd gnd FILL
XFILL_3__1265_ vdd gnd FILL
X_1618_ _1651_/B _1687_/C _1687_/B vdd gnd NAND2X1
X_1549_ _1625_/C _1578_/B _1578_/A _1574_/B vdd gnd NAND3X1
XFILL_1__1734_ vdd gnd FILL
XFILL_1__1665_ vdd gnd FILL
XFILL_1__1803_ vdd gnd FILL
XFILL_1__1596_ vdd gnd FILL
XFILL_2__1010_ vdd gnd FILL
XFILL_2__987_ vdd gnd FILL
XBUFX2_insert21 _984_/Y _990_/A vdd gnd BUFX2
XFILL_2__1774_ vdd gnd FILL
X_993_ _996_/A _993_/B _994_/C vdd gnd NAND2X1
XFILL_2__1843_ vdd gnd FILL
XFILL_2__1912_ vdd gnd FILL
XFILL_0__1410_ vdd gnd FILL
XFILL_0__1341_ vdd gnd FILL
XFILL_2__1208_ vdd gnd FILL
XFILL_3__1050_ vdd gnd FILL
XFILL_0__1272_ vdd gnd FILL
XFILL_2__1139_ vdd gnd FILL
X_1334_ _1334_/A _1515_/A _1416_/C vdd gnd NAND2X1
X_1403_ _1425_/C _1403_/B _1423_/A vdd gnd AND2X2
X_1265_ _1371_/B _1371_/A _1274_/C _1280_/B vdd gnd NAND3X1
XFILL_0__1608_ vdd gnd FILL
XFILL_0__1539_ vdd gnd FILL
XFILL_1__1450_ vdd gnd FILL
XFILL_3__1317_ vdd gnd FILL
X_1196_ _1196_/A _1196_/B _1196_/C _1277_/C vdd gnd OAI21X1
XFILL_4__1090_ vdd gnd FILL
XFILL_1__1381_ vdd gnd FILL
XFILL_3__1248_ vdd gnd FILL
XFILL_3__1179_ vdd gnd FILL
XFILL_1__1648_ vdd gnd FILL
XFILL_1__1717_ vdd gnd FILL
XFILL_2__1490_ vdd gnd FILL
XFILL_1__1579_ vdd gnd FILL
XFILL_2_CLKBUF1_insert7 vdd gnd FILL
XCLKBUF1_insert6 clk _1880_/CLK vdd gnd CLKBUF1
XFILL_2__1757_ vdd gnd FILL
XFILL_2__1826_ vdd gnd FILL
X_976_ _977_/A _976_/B _977_/C vdd gnd NAND2X1
XFILL_2__1688_ vdd gnd FILL
XFILL_3__1102_ vdd gnd FILL
X_1050_ _1068_/B _1050_/B _1068_/A _1062_/B vdd gnd OAI21X1
X_1883_ _1883_/D _1885_/CLK _1883_/Q vdd gnd DFFPOSX1
XFILL_0__1255_ vdd gnd FILL
XFILL_0__1324_ vdd gnd FILL
XFILL_3__1033_ vdd gnd FILL
XFILL_0__1186_ vdd gnd FILL
XFILL_1__1502_ vdd gnd FILL
XFILL_3__1797_ vdd gnd FILL
X_1248_ _952_/A _1248_/B _1896_/Q _1338_/B vdd gnd AOI21X1
X_1317_ _1317_/A _1317_/B _1317_/C _1321_/C vdd gnd AOI21X1
XFILL_1__988_ vdd gnd FILL
XFILL_1__1433_ vdd gnd FILL
XFILL_1__1364_ vdd gnd FILL
X_1179_ _1243_/B _1179_/B _1243_/A _1266_/A vdd gnd OAI21X1
XFILL_1__1295_ vdd gnd FILL
XFILL_2__1611_ vdd gnd FILL
XFILL_2__1542_ vdd gnd FILL
XFILL_4__1409_ vdd gnd FILL
XFILL_2__1473_ vdd gnd FILL
XFILL_0__1040_ vdd gnd FILL
XFILL_3__1720_ vdd gnd FILL
XFILL_3__1651_ vdd gnd FILL
XFILL_3__1582_ vdd gnd FILL
XFILL_2__1809_ vdd gnd FILL
X_959_ _959_/A _965_/B _959_/C _959_/Y vdd gnd OAI21X1
X_1102_ _1102_/A _1102_/B _1102_/C _1130_/C vdd gnd OAI21X1
X_1033_ _973_/B _1216_/A _1060_/C vdd gnd NAND2X1
X_1797_ _1799_/B _1798_/A vdd gnd INVX1
X_1866_ _1866_/D _1885_/CLK _999_/A vdd gnd DFFPOSX1
XFILL_0__1307_ vdd gnd FILL
XFILL_0__1238_ vdd gnd FILL
XFILL_3__1016_ vdd gnd FILL
XFILL_1__1080_ vdd gnd FILL
XFILL_0__1169_ vdd gnd FILL
XFILL_3__1918_ vdd gnd FILL
XFILL_3__1849_ vdd gnd FILL
XFILL_0_BUFX2_insert20 vdd gnd FILL
XFILL_1__1347_ vdd gnd FILL
XFILL_1__1416_ vdd gnd FILL
XFILL_1__1278_ vdd gnd FILL
XFILL_2__1525_ vdd gnd FILL
XFILL_2__1456_ vdd gnd FILL
XFILL_2__1387_ vdd gnd FILL
X_1651_ _1651_/A _1651_/B _1685_/A _1708_/A vdd gnd AOI21X1
X_1720_ _1720_/A _1720_/B _1728_/A _1762_/C vdd gnd OAI21X1
XFILL_0__989_ vdd gnd FILL
XFILL_0__1023_ vdd gnd FILL
X_1582_ _946_/A Cin[6] _949_/A Cin[5] _1652_/B vdd gnd AOI22X1
XFILL_3__1634_ vdd gnd FILL
XFILL_3__1703_ vdd gnd FILL
XFILL_3__1496_ vdd gnd FILL
XFILL_3__1565_ vdd gnd FILL
XFILL_0__1787_ vdd gnd FILL
XFILL_4__967_ vdd gnd FILL
X_1016_ _1029_/A _1016_/B _1018_/B vdd gnd NAND2X1
XFILL_1__1201_ vdd gnd FILL
XFILL_1__1132_ vdd gnd FILL
XFILL_4__1743_ vdd gnd FILL
X_1918_ _940_/Y Yout[2] vdd gnd BUFX2
X_1849_ _948_/A _1849_/B _1849_/C _1905_/D vdd gnd OAI21X1
XFILL_1__1063_ vdd gnd FILL
XFILL_4__1674_ vdd gnd FILL
XFILL_2__1310_ vdd gnd FILL
XFILL_2__1241_ vdd gnd FILL
XFILL_4__1108_ vdd gnd FILL
XFILL_2__1172_ vdd gnd FILL
XFILL_4__1039_ vdd gnd FILL
XFILL_3__985_ vdd gnd FILL
XFILL_2__1508_ vdd gnd FILL
XFILL_0__1710_ vdd gnd FILL
XFILL_0__1572_ vdd gnd FILL
XFILL_0__1641_ vdd gnd FILL
XFILL_3__1350_ vdd gnd FILL
XFILL_3__1281_ vdd gnd FILL
XFILL_2__1439_ vdd gnd FILL
XFILL_0_BUFX2_insert1 vdd gnd FILL
X_1634_ _1634_/A _1634_/B _1634_/C _1635_/C vdd gnd NOR3X1
X_1703_ _1703_/A _1703_/B _1706_/C vdd gnd NOR2X1
XFILL_0__1006_ vdd gnd FILL
XFILL_1__1681_ vdd gnd FILL
XFILL_3__1617_ vdd gnd FILL
X_1496_ _1635_/A _1575_/A vdd gnd INVX1
X_1565_ _1565_/A _1565_/B _1565_/C _1565_/D _1571_/C vdd gnd OAI22X1
XFILL_1__1750_ vdd gnd FILL
XFILL_3__1548_ vdd gnd FILL
XFILL_3__1479_ vdd gnd FILL
XFILL_0__1839_ vdd gnd FILL
XFILL_1__1115_ vdd gnd FILL
XFILL_1__1046_ vdd gnd FILL
XFILL_2__1790_ vdd gnd FILL
XFILL_4__1588_ vdd gnd FILL
XFILL_2__1155_ vdd gnd FILL
XFILL_2__1224_ vdd gnd FILL
XFILL_2__1086_ vdd gnd FILL
X_1350_ _1460_/A _1524_/B _1357_/C _1363_/B vdd gnd NAND3X1
XFILL_3__968_ vdd gnd FILL
X_1281_ _1285_/A _1285_/B _1382_/C _1289_/B vdd gnd OAI21X1
XFILL_1_BUFX2_insert19 vdd gnd FILL
XFILL_0__1624_ vdd gnd FILL
XFILL_0__1555_ vdd gnd FILL
XFILL_3__1333_ vdd gnd FILL
XFILL_3__1402_ vdd gnd FILL
XFILL_3__1264_ vdd gnd FILL
XFILL_0__1486_ vdd gnd FILL
XFILL_3__1195_ vdd gnd FILL
X_1617_ _1620_/A _1620_/B _1621_/A _1651_/B vdd gnd NAND3X1
XFILL_1__1802_ vdd gnd FILL
XFILL_1__1733_ vdd gnd FILL
XFILL_4__1373_ vdd gnd FILL
XFILL_1__1664_ vdd gnd FILL
X_1548_ _1554_/C _1555_/C _1578_/B vdd gnd NAND2X1
XFILL_4__1442_ vdd gnd FILL
X_1479_ _1479_/A _1479_/B _1479_/C _1493_/A vdd gnd NAND3X1
XFILL_1__1595_ vdd gnd FILL
XFILL_2__986_ vdd gnd FILL
XBUFX2_insert22 _984_/Y _1216_/A vdd gnd BUFX2
XFILL_1__1029_ vdd gnd FILL
XFILL_2__1911_ vdd gnd FILL
XFILL_2__1773_ vdd gnd FILL
X_992_ _992_/A _992_/B _992_/C _992_/Y vdd gnd OAI21X1
XFILL_2__1842_ vdd gnd FILL
XFILL_0__1340_ vdd gnd FILL
XFILL_2__1207_ vdd gnd FILL
XFILL_2__1138_ vdd gnd FILL
XFILL_0__1271_ vdd gnd FILL
X_1402_ _1402_/A _1402_/B _1402_/C _1480_/C vdd gnd AOI21X1
XFILL_2__1069_ vdd gnd FILL
X_1333_ _949_/A Cin[2] _1515_/A vdd gnd AND2X2
X_1264_ _1361_/C _1325_/B _1325_/A _1371_/A vdd gnd NAND3X1
XFILL_0__1538_ vdd gnd FILL
XFILL_0__1607_ vdd gnd FILL
XFILL_0__1469_ vdd gnd FILL
XFILL_3__1316_ vdd gnd FILL
X_1195_ _1277_/B _1277_/A _1203_/C _1208_/B vdd gnd NAND3X1
XFILL_1__1380_ vdd gnd FILL
XFILL_3__1247_ vdd gnd FILL
XFILL_3__1178_ vdd gnd FILL
XFILL_1__1578_ vdd gnd FILL
XFILL_1__1647_ vdd gnd FILL
XFILL_1__1716_ vdd gnd FILL
XFILL_2_CLKBUF1_insert8 vdd gnd FILL
XFILL_2__969_ vdd gnd FILL
XFILL_4__1287_ vdd gnd FILL
XCLKBUF1_insert7 clk _1910_/CLK vdd gnd CLKBUF1
XFILL_2__1687_ vdd gnd FILL
XFILL_2__1756_ vdd gnd FILL
XFILL_2__1825_ vdd gnd FILL
X_975_ _975_/A _977_/B vdd gnd INVX1
XFILL_0__1323_ vdd gnd FILL
XFILL_3__1101_ vdd gnd FILL
X_1882_ _1882_/D _1885_/CLK _1882_/Q vdd gnd DFFPOSX1
XFILL_4_BUFX2_insert23 vdd gnd FILL
XFILL_3__1032_ vdd gnd FILL
XFILL_0__1185_ vdd gnd FILL
XFILL_0__1254_ vdd gnd FILL
XFILL_3__1796_ vdd gnd FILL
XFILL_1__1501_ vdd gnd FILL
XFILL_1__1432_ vdd gnd FILL
X_1316_ _1316_/A _1316_/B _1403_/B _1425_/C vdd gnd NAND3X1
XFILL_1__987_ vdd gnd FILL
X_1178_ _949_/A _1248_/B _1895_/Q _1243_/B vdd gnd AOI21X1
X_1247_ _1338_/C _1249_/B vdd gnd INVX1
XFILL_1__1363_ vdd gnd FILL
XFILL_1__1294_ vdd gnd FILL
XFILL_4__1072_ vdd gnd FILL
XFILL_2__1541_ vdd gnd FILL
XFILL_2__1610_ vdd gnd FILL
XFILL_2__1472_ vdd gnd FILL
XFILL_3__1650_ vdd gnd FILL
XFILL_2__1739_ vdd gnd FILL
XFILL_3__1581_ vdd gnd FILL
XFILL_2__1808_ vdd gnd FILL
X_1032_ _1801_/A _1032_/B _1032_/C _1871_/D vdd gnd OAI21X1
X_958_ Xin[0] _965_/B _959_/C vdd gnd NAND2X1
X_1101_ _1101_/A _1101_/B _1138_/A _1142_/A vdd gnd OAI21X1
XFILL_0__1306_ vdd gnd FILL
XFILL_3__1015_ vdd gnd FILL
XFILL99750x66450 vdd gnd FILL
X_1796_ _1796_/A _1796_/B _1799_/B vdd gnd XNOR2X1
X_1865_ _998_/Y _1885_/CLK _941_/A vdd gnd DFFPOSX1
XFILL_0__1237_ vdd gnd FILL
XFILL_0__1099_ vdd gnd FILL
XFILL_0__1168_ vdd gnd FILL
XFILL_3__1917_ vdd gnd FILL
XFILL_3__1779_ vdd gnd FILL
XFILL_3__1848_ vdd gnd FILL
XFILL_1__1415_ vdd gnd FILL
XFILL_0_BUFX2_insert21 vdd gnd FILL
XFILL_1__1346_ vdd gnd FILL
XFILL_1__1277_ vdd gnd FILL
XFILL_2__1524_ vdd gnd FILL
XFILL_2__1455_ vdd gnd FILL
XFILL_2__1386_ vdd gnd FILL
X_1650_ _1687_/C _1685_/A vdd gnd INVX1
X_1581_ _956_/B Cin[7] _1652_/A vdd gnd NAND2X1
XFILL_0__988_ vdd gnd FILL
XFILL_0__1022_ vdd gnd FILL
XFILL_3__1633_ vdd gnd FILL
XFILL_3__1702_ vdd gnd FILL
XFILL_3__1564_ vdd gnd FILL
XFILL_0__1786_ vdd gnd FILL
XFILL_3__1495_ vdd gnd FILL
X_1015_ _1843_/B _1257_/B _1835_/B _1016_/B vdd gnd OAI21X1
XFILL_1__1200_ vdd gnd FILL
XFILL_1__1131_ vdd gnd FILL
XFILL_1__1062_ vdd gnd FILL
X_1917_ _935_/Y Yout[1] vdd gnd BUFX2
X_1779_ _1779_/A _1888_/Q _1793_/B vdd gnd XOR2X1
XFILL_4__1811_ vdd gnd FILL
X_1848_ _1848_/A Xin[3] _1849_/C vdd gnd NAND2X1
XFILL101250x31350 vdd gnd FILL
XFILL_2__1240_ vdd gnd FILL
XFILL_2__1171_ vdd gnd FILL
XFILL_1__1329_ vdd gnd FILL
XFILL_3__984_ vdd gnd FILL
XFILL_2__1507_ vdd gnd FILL
XFILL_2__1438_ vdd gnd FILL
XFILL_0__1571_ vdd gnd FILL
XFILL_0__1640_ vdd gnd FILL
XFILL_0_BUFX2_insert2 vdd gnd FILL
XFILL_3__1280_ vdd gnd FILL
XFILL_2__1369_ vdd gnd FILL
X_1633_ _1633_/A _1633_/B _1633_/C _1705_/B vdd gnd NAND3X1
X_1564_ _1564_/A _1564_/B _1635_/A _1565_/B vdd gnd AOI21X1
X_1702_ _1882_/Q _1702_/B _1745_/C vdd gnd NAND2X1
XFILL_0__1005_ vdd gnd FILL
XFILL_1__1680_ vdd gnd FILL
XFILL_3__1547_ vdd gnd FILL
XFILL_3__1616_ vdd gnd FILL
X_1495_ _1495_/A _1495_/B _1635_/A vdd gnd NAND2X1
XFILL_0__1838_ vdd gnd FILL
XFILL_0__1769_ vdd gnd FILL
XFILL_3__1478_ vdd gnd FILL
XFILL_4__949_ vdd gnd FILL
XFILL_1__1114_ vdd gnd FILL
XFILL_1__1045_ vdd gnd FILL
XFILL_4__1725_ vdd gnd FILL
XFILL_4__1656_ vdd gnd FILL
XFILL101250x43050 vdd gnd FILL
XFILL100650x7950 vdd gnd FILL
XFILL_2__1223_ vdd gnd FILL
XFILL_2__1154_ vdd gnd FILL
XFILL_2__1085_ vdd gnd FILL
XFILL_3__1401_ vdd gnd FILL
XFILL_3__967_ vdd gnd FILL
X_1280_ _1280_/A _1280_/B _1372_/B _1285_/B vdd gnd AOI21X1
XFILL_0__1623_ vdd gnd FILL
XFILL_0__1554_ vdd gnd FILL
XFILL_0__1485_ vdd gnd FILL
XFILL_3__1332_ vdd gnd FILL
XFILL_3__1194_ vdd gnd FILL
XFILL_3__1263_ vdd gnd FILL
X_1547_ _1554_/A _1620_/B _1547_/C _1625_/C vdd gnd NAND3X1
X_1616_ _1710_/A _1616_/B _1621_/A vdd gnd NAND2X1
XFILL_4__1510_ vdd gnd FILL
XFILL_1__1801_ vdd gnd FILL
XFILL_1__1594_ vdd gnd FILL
XFILL_1__1663_ vdd gnd FILL
XFILL_1__1732_ vdd gnd FILL
X_1478_ _1486_/C _1486_/B _1486_/A _1482_/B vdd gnd NAND3X1
XFILL_2__985_ vdd gnd FILL
XBUFX2_insert23 _984_/Y _1702_/B vdd gnd BUFX2
XBUFX2_insert12 Cin[0] _1248_/B vdd gnd BUFX2
XFILL_1__1028_ vdd gnd FILL
XFILL_2__1841_ vdd gnd FILL
XFILL_2__1772_ vdd gnd FILL
X_991_ _992_/A _991_/B _992_/C vdd gnd NAND2X1
XFILL_2__1206_ vdd gnd FILL
XFILL_2__1137_ vdd gnd FILL
XFILL_0__1270_ vdd gnd FILL
XFILL_2__1068_ vdd gnd FILL
X_1401_ _1474_/C _1402_/C vdd gnd INVX1
XFILL_0__1606_ vdd gnd FILL
X_1332_ _1416_/A _1421_/A vdd gnd INVX1
X_1194_ _1267_/C _1231_/B _1231_/A _1277_/A vdd gnd NAND3X1
X_1263_ _1263_/A _1263_/B _1263_/C _1325_/B vdd gnd OAI21X1
XFILL_0__1537_ vdd gnd FILL
XFILL_0__1468_ vdd gnd FILL
XFILL_3__1315_ vdd gnd FILL
XFILL_3__1246_ vdd gnd FILL
XFILL_3__1177_ vdd gnd FILL
XFILL_0__1399_ vdd gnd FILL
XFILL_1__1715_ vdd gnd FILL
XFILL_1__1577_ vdd gnd FILL
XFILL_1__1646_ vdd gnd FILL
XFILL_4__1355_ vdd gnd FILL
XFILL_4__1424_ vdd gnd FILL
XFILL_2_CLKBUF1_insert9 vdd gnd FILL
XFILL_2__968_ vdd gnd FILL
XFILL_2__1824_ vdd gnd FILL
XCLKBUF1_insert8 clk _1897_/CLK vdd gnd CLKBUF1
XFILL_2__1686_ vdd gnd FILL
XFILL_2__1755_ vdd gnd FILL
X_974_ _977_/A _974_/B _974_/C _974_/Y vdd gnd OAI21X1
XFILL_3__1031_ vdd gnd FILL
XFILL_0__1322_ vdd gnd FILL
XFILL_3__1100_ vdd gnd FILL
X_1881_ _1881_/D _1885_/CLK _997_/B vdd gnd DFFPOSX1
XFILL_0__1184_ vdd gnd FILL
XFILL_0__1253_ vdd gnd FILL
XFILL_3__1795_ vdd gnd FILL
XFILL_1__986_ vdd gnd FILL
X_1315_ _1315_/A _1315_/B _1315_/C _1320_/B vdd gnd NAND3X1
XFILL_1__1500_ vdd gnd FILL
XFILL_1__1431_ vdd gnd FILL
XFILL_1__1362_ vdd gnd FILL
X_1246_ _952_/A _1248_/B _1896_/Q _1338_/C vdd gnd NAND3X1
XFILL_4__1140_ vdd gnd FILL
X_1177_ _1243_/C _1179_/B vdd gnd INVX1
XFILL_3__1229_ vdd gnd FILL
XFILL_1__1293_ vdd gnd FILL
XFILL_2__1540_ vdd gnd FILL
XFILL_2__1471_ vdd gnd FILL
XFILL_1__1629_ vdd gnd FILL
XFILL_4__1269_ vdd gnd FILL
XFILL_3__1580_ vdd gnd FILL
XFILL_2__1807_ vdd gnd FILL
X_957_ _957_/A _965_/A _957_/C _957_/Y vdd gnd OAI21X1
XFILL_2__1669_ vdd gnd FILL
XFILL_2__1738_ vdd gnd FILL
X_1031_ _970_/B _1801_/A _1032_/C vdd gnd NAND2X1
X_1100_ _1206_/B _1154_/A vdd gnd INVX1
XFILL_0__1305_ vdd gnd FILL
XFILL_0__1236_ vdd gnd FILL
XFILL_3__1014_ vdd gnd FILL
XFILL_4__982_ vdd gnd FILL
X_1795_ _1795_/A _1889_/Q _1796_/B vdd gnd XOR2X1
X_1864_ _996_/Y _1880_/CLK _936_/A vdd gnd DFFPOSX1
XFILL_0__1098_ vdd gnd FILL
XFILL_3__1916_ vdd gnd FILL
XFILL_0__1167_ vdd gnd FILL
XFILL_3__1778_ vdd gnd FILL
XFILL_1__969_ vdd gnd FILL
XFILL_0_BUFX2_insert22 vdd gnd FILL
XFILL_3__1847_ vdd gnd FILL
XFILL_1__1345_ vdd gnd FILL
XFILL_1__1414_ vdd gnd FILL
XFILL_4__1054_ vdd gnd FILL
XFILL_4__1123_ vdd gnd FILL
X_1229_ _1299_/B _1299_/A _1372_/B vdd gnd XNOR2X1
XFILL_1__1276_ vdd gnd FILL
XFILL_2__1523_ vdd gnd FILL
XFILL_2__1454_ vdd gnd FILL
XFILL_2__1385_ vdd gnd FILL
X_1580_ _1602_/A _1599_/A vdd gnd INVX1
XFILL_3__1701_ vdd gnd FILL
XFILL_0__987_ vdd gnd FILL
XFILL_0__1021_ vdd gnd FILL
XFILL_3__1632_ vdd gnd FILL
XFILL_3__1563_ vdd gnd FILL
XFILL_0__1785_ vdd gnd FILL
XFILL_3__1494_ vdd gnd FILL
X_1014_ _1898_/Q _1835_/B vdd gnd INVX1
XFILL_1__1061_ vdd gnd FILL
XFILL_0__1219_ vdd gnd FILL
X_1916_ _930_/Y Yout[0] vdd gnd BUFX2
XFILL_1__1130_ vdd gnd FILL
X_1847_ _951_/A _1847_/B _1847_/C _1904_/D vdd gnd OAI21X1
X_1778_ _963_/A _1778_/B _1794_/C _1779_/A vdd gnd OAI21X1
XFILL_1__1328_ vdd gnd FILL
XFILL_2__1170_ vdd gnd FILL
XFILL_1__1259_ vdd gnd FILL
XFILL_3__983_ vdd gnd FILL
XFILL_2__1506_ vdd gnd FILL
XFILL_2__1437_ vdd gnd FILL
XFILL_0__1570_ vdd gnd FILL
XFILL_0_BUFX2_insert3 vdd gnd FILL
X_1701_ _998_/A _1701_/B _1701_/C _1881_/D vdd gnd OAI21X1
XFILL_2__1368_ vdd gnd FILL
XFILL_2__1299_ vdd gnd FILL
X_1632_ _1692_/A _1693_/A _1693_/B _1633_/B vdd gnd NAND3X1
X_1563_ _1635_/B _1575_/C _1575_/A _1565_/A vdd gnd AOI21X1
X_1494_ _1494_/A _1494_/B _1565_/C _1562_/C vdd gnd AOI21X1
XFILL_0__1004_ vdd gnd FILL
XFILL_3__1546_ vdd gnd FILL
XFILL_3__1615_ vdd gnd FILL
XFILL_0__1768_ vdd gnd FILL
XFILL_3__1477_ vdd gnd FILL
XFILL_0__1837_ vdd gnd FILL
XFILL_0__1699_ vdd gnd FILL
XFILL_1__1113_ vdd gnd FILL
XFILL_1__1044_ vdd gnd FILL
XFILL_2__1222_ vdd gnd FILL
XFILL_2__1153_ vdd gnd FILL
XFILL_2__1084_ vdd gnd FILL
XFILL_0__1622_ vdd gnd FILL
XFILL_3__1400_ vdd gnd FILL
XFILL_3__1331_ vdd gnd FILL
XFILL_3__966_ vdd gnd FILL
XFILL_0__1553_ vdd gnd FILL
XFILL_0__1484_ vdd gnd FILL
XFILL_3__1262_ vdd gnd FILL
XFILL_3__1193_ vdd gnd FILL
X_1546_ _1553_/A _1576_/B _1578_/A vdd gnd AND2X2
XFILL_1__1731_ vdd gnd FILL
X_1615_ _1891_/Q _1615_/B _1620_/A vdd gnd NAND2X1
X_1477_ _1480_/B _1480_/A _1479_/C _1486_/B vdd gnd OAI21X1
XFILL_1__1800_ vdd gnd FILL
XFILL101250x7950 vdd gnd FILL
XFILL_1__1593_ vdd gnd FILL
XFILL_1__1662_ vdd gnd FILL
XFILL_3__1529_ vdd gnd FILL
XFILL_2__984_ vdd gnd FILL
XBUFX2_insert24 _984_/Y _1801_/A vdd gnd BUFX2
XBUFX2_insert13 Cin[0] _1104_/B vdd gnd BUFX2
X_990_ _990_/A _990_/B _990_/C _990_/Y vdd gnd OAI21X1
XFILL_1__1027_ vdd gnd FILL
XFILL_2__1840_ vdd gnd FILL
XFILL_4__1638_ vdd gnd FILL
XFILL_2__1771_ vdd gnd FILL
XFILL_4__1707_ vdd gnd FILL
XFILL_2__1205_ vdd gnd FILL
XFILL_2__1136_ vdd gnd FILL
XFILL_2__1067_ vdd gnd FILL
X_1400_ _1494_/A _1486_/C vdd gnd INVX1
X_1331_ _1416_/A _1331_/B _1331_/C _1355_/B vdd gnd NAND3X1
XFILL_0__1605_ vdd gnd FILL
XFILL_3__1314_ vdd gnd FILL
XFILL_3__949_ vdd gnd FILL
X_1262_ _1360_/C _1360_/B _1360_/A _1361_/C vdd gnd NAND3X1
X_1193_ _1193_/A _1193_/B _1193_/C _1231_/B vdd gnd OAI21X1
XFILL_0__1536_ vdd gnd FILL
XFILL_0__1467_ vdd gnd FILL
XFILL_0__1398_ vdd gnd FILL
XFILL_3__1176_ vdd gnd FILL
XFILL_3__1245_ vdd gnd FILL
XFILL_1__1645_ vdd gnd FILL
X_1529_ _965_/A _1533_/D _1611_/A _1530_/C vdd gnd OAI21X1
XFILL_1__1714_ vdd gnd FILL
XFILL_1__1576_ vdd gnd FILL
XFILL_2__967_ vdd gnd FILL
XFILL_2__1754_ vdd gnd FILL
XFILL_2__1823_ vdd gnd FILL
XCLKBUF1_insert9 clk _1908_/CLK vdd gnd CLKBUF1
X_973_ _977_/A _973_/B _974_/C vdd gnd NAND2X1
XFILL_2__1685_ vdd gnd FILL
XFILL100350x31350 vdd gnd FILL
XFILL100050x66450 vdd gnd FILL
X_1880_ _1880_/D _1880_/CLK _995_/B vdd gnd DFFPOSX1
XFILL_0__1321_ vdd gnd FILL
XFILL_3__1030_ vdd gnd FILL
XFILL_4_BUFX2_insert14 vdd gnd FILL
XFILL_0__1252_ vdd gnd FILL
XFILL_4_BUFX2_insert25 vdd gnd FILL
XFILL_0__1183_ vdd gnd FILL
XFILL_2__1119_ vdd gnd FILL
XFILL_3__1794_ vdd gnd FILL
X_1314_ _1321_/A _1321_/B _1320_/C _1319_/C vdd gnd OAI21X1
XFILL_1__985_ vdd gnd FILL
XFILL_0__1519_ vdd gnd FILL
XFILL_1__1430_ vdd gnd FILL
XFILL_1__1361_ vdd gnd FILL
X_1176_ _949_/A _1248_/B _1895_/Q _1243_/C vdd gnd NAND3X1
X_1245_ _949_/A Cin[1] _1338_/A vdd gnd NAND2X1
XFILL_3__1159_ vdd gnd FILL
XFILL_1__1292_ vdd gnd FILL
XFILL_3__1228_ vdd gnd FILL
XFILL_1__1628_ vdd gnd FILL
XFILL_2__1470_ vdd gnd FILL
XFILL_4__1406_ vdd gnd FILL
XFILL_1__1559_ vdd gnd FILL
XFILL_4__1337_ vdd gnd FILL
XFILL_2__1737_ vdd gnd FILL
XFILL_2__1806_ vdd gnd FILL
X_956_ _957_/A _956_/B _957_/C vdd gnd NAND2X1
XFILL100350x43050 vdd gnd FILL
XFILL_2__1668_ vdd gnd FILL
XFILL_2__1599_ vdd gnd FILL
X_1030_ _1030_/A _1034_/A _1032_/B vdd gnd NAND2X1
X_1863_ _994_/Y _1880_/CLK _931_/A vdd gnd DFFPOSX1
XFILL_0__1304_ vdd gnd FILL
XFILL_3__1013_ vdd gnd FILL
XFILL_0__1235_ vdd gnd FILL
XFILL_0__1166_ vdd gnd FILL
X_1794_ _1888_/Q _1794_/B _1794_/C _1795_/A vdd gnd OAI21X1
XFILL_3__1915_ vdd gnd FILL
XFILL_0__1097_ vdd gnd FILL
XFILL_3__1846_ vdd gnd FILL
XFILL_3__1777_ vdd gnd FILL
XFILL_0_BUFX2_insert23 vdd gnd FILL
XFILL_1__968_ vdd gnd FILL
XFILL_0_BUFX2_insert12 vdd gnd FILL
X_1228_ _1228_/A _1240_/C _1228_/C _1299_/A vdd gnd OAI21X1
XFILL_1__1275_ vdd gnd FILL
XFILL_1__1344_ vdd gnd FILL
XFILL_1__1413_ vdd gnd FILL
X_1159_ _1159_/A _1228_/A _1159_/C _1219_/B vdd gnd OAI21X1
XFILL_2__1522_ vdd gnd FILL
XFILL_2__1453_ vdd gnd FILL
XFILL_2__1384_ vdd gnd FILL
XFILL_0__986_ vdd gnd FILL
XFILL_0__1020_ vdd gnd FILL
XFILL_3__1700_ vdd gnd FILL
XFILL_3__1631_ vdd gnd FILL
XFILL_3__1562_ vdd gnd FILL
XFILL_0__1784_ vdd gnd FILL
XFILL_3__1493_ vdd gnd FILL
X_939_ _944_/A _972_/A _965_/B _986_/A _940_/C vdd gnd AOI22X1
XFILL_4__964_ vdd gnd FILL
X_1013_ _1248_/B _1257_/B vdd gnd INVX1
X_1777_ _1777_/A _1777_/B _1793_/A vdd gnd NAND2X1
X_1915_ _957_/Y Xout[3] vdd gnd BUFX2
XFILL_0__1218_ vdd gnd FILL
XFILL_0__1149_ vdd gnd FILL
X_1846_ _951_/A Xin[2] _1847_/C vdd gnd NAND2X1
XFILL_1__1060_ vdd gnd FILL
XFILL_4__1740_ vdd gnd FILL
XFILL_4__1671_ vdd gnd FILL
XFILL_3__1829_ vdd gnd FILL
XFILL_1__1327_ vdd gnd FILL
XFILL_1__1258_ vdd gnd FILL
XFILL_4__1105_ vdd gnd FILL
XFILL_4__1036_ vdd gnd FILL
XFILL_1__1189_ vdd gnd FILL
XFILL_3__982_ vdd gnd FILL
XFILL_2__1505_ vdd gnd FILL
XFILL_2__1436_ vdd gnd FILL
XFILL_0_BUFX2_insert4 vdd gnd FILL
XFILL_2__1367_ vdd gnd FILL
X_1631_ _1685_/B _1631_/B _1631_/C _1693_/B vdd gnd OAI21X1
X_1700_ _1700_/A _1700_/B _992_/A _1701_/C vdd gnd OAI21X1
XFILL_0__1003_ vdd gnd FILL
XFILL_0__969_ vdd gnd FILL
XFILL_2__1298_ vdd gnd FILL
XFILL_3__1614_ vdd gnd FILL
X_1562_ _1562_/A _1562_/B _1562_/C _1566_/A vdd gnd OAI21X1
X_1493_ _1493_/A _1565_/C vdd gnd INVX1
XFILL_3__1545_ vdd gnd FILL
XFILL_0__1767_ vdd gnd FILL
XFILL_3__1476_ vdd gnd FILL
XFILL_0__1698_ vdd gnd FILL
XFILL_0__1836_ vdd gnd FILL
XFILL_1__1112_ vdd gnd FILL
X_1829_ _1837_/B _1833_/B _1829_/C _1895_/D vdd gnd OAI21X1
XFILL_1__1043_ vdd gnd FILL
XFILL_4__1585_ vdd gnd FILL
XFILL_2__1221_ vdd gnd FILL
XFILL_2__1083_ vdd gnd FILL
XFILL_2__1152_ vdd gnd FILL
XFILL_3__965_ vdd gnd FILL
XFILL_0__1621_ vdd gnd FILL
XFILL_0__1552_ vdd gnd FILL
XFILL_3__1330_ vdd gnd FILL
XFILL_0__1483_ vdd gnd FILL
XFILL_2__1419_ vdd gnd FILL
XFILL_3__1261_ vdd gnd FILL
XFILL_3__1192_ vdd gnd FILL
X_1614_ _1620_/C _1621_/B _1687_/C vdd gnd NAND2X1
X_1545_ _1625_/A _1578_/C _1625_/B _1574_/A vdd gnd OAI21X1
XFILL_1__1730_ vdd gnd FILL
XFILL_1__1661_ vdd gnd FILL
X_1476_ _1476_/A _1476_/B _1552_/A _1480_/B vdd gnd AOI21X1
XFILL_4__1370_ vdd gnd FILL
XFILL_1__1592_ vdd gnd FILL
XFILL_0__1819_ vdd gnd FILL
XFILL_3__1528_ vdd gnd FILL
XFILL_3__1459_ vdd gnd FILL
XBUFX2_insert25 _984_/Y _1790_/A vdd gnd BUFX2
XFILL_2__983_ vdd gnd FILL
XBUFX2_insert14 Cin[0] _1106_/B vdd gnd BUFX2
XFILL_2__1770_ vdd gnd FILL
XFILL_1__1026_ vdd gnd FILL
XFILL_2__1204_ vdd gnd FILL
XFILL_2__1135_ vdd gnd FILL
XFILL100950x85950 vdd gnd FILL
XFILL_2__1066_ vdd gnd FILL
X_1330_ _1420_/B _1334_/A _1331_/C vdd gnd NAND2X1
X_1261_ _1261_/A _1261_/B _1325_/A vdd gnd AND2X2
XFILL_3__948_ vdd gnd FILL
XFILL_0__1535_ vdd gnd FILL
XFILL_0__1604_ vdd gnd FILL
XFILL_3__1313_ vdd gnd FILL
X_1192_ _1266_/C _1266_/B _1266_/A _1267_/C vdd gnd NAND3X1
XFILL_3__1244_ vdd gnd FILL
XFILL_0__1466_ vdd gnd FILL
XFILL_3__1175_ vdd gnd FILL
XFILL_0__1397_ vdd gnd FILL
XFILL_1__1713_ vdd gnd FILL
X_1528_ _963_/A _1533_/B _1596_/B _1530_/B vdd gnd OAI21X1
X_1459_ _1551_/B _1551_/A _1470_/C _1476_/B vdd gnd NAND3X1
XFILL_1__1644_ vdd gnd FILL
XFILL_1__1575_ vdd gnd FILL
XFILL_4__1284_ vdd gnd FILL
XFILL_1__1009_ vdd gnd FILL
XFILL_2__966_ vdd gnd FILL
XFILL_2__1822_ vdd gnd FILL
XFILL_2__1753_ vdd gnd FILL
X_972_ _972_/A _974_/B vdd gnd INVX1
XFILL100650x15750 vdd gnd FILL
XFILL_2__1684_ vdd gnd FILL
XFILL_0__1320_ vdd gnd FILL
XFILL_0__1182_ vdd gnd FILL
XFILL_2__1118_ vdd gnd FILL
XFILL_0__1251_ vdd gnd FILL
XFILL_3__1793_ vdd gnd FILL
XFILL_2__1049_ vdd gnd FILL
XFILL_1__984_ vdd gnd FILL
X_1313_ _1313_/A _1313_/B _1313_/C _1320_/C vdd gnd OAI21X1
X_1244_ _1360_/C _1263_/C vdd gnd INVX1
XFILL_0__1518_ vdd gnd FILL
XFILL_1__1360_ vdd gnd FILL
XFILL_1__1291_ vdd gnd FILL
XFILL_3__1227_ vdd gnd FILL
X_1175_ _946_/A Cin[1] _1243_/A vdd gnd NAND2X1
XFILL_0__1449_ vdd gnd FILL
XFILL_3__1089_ vdd gnd FILL
XFILL_3__1158_ vdd gnd FILL
XFILL_1__1627_ vdd gnd FILL
XFILL_1__1558_ vdd gnd FILL
XFILL_1__1489_ vdd gnd FILL
XFILL_2__949_ vdd gnd FILL
XFILL100650x27450 vdd gnd FILL
XFILL_2__1667_ vdd gnd FILL
XFILL_2__1736_ vdd gnd FILL
X_955_ _955_/A _965_/A vdd gnd INVX2
XFILL_2__1805_ vdd gnd FILL
XFILL_2__1598_ vdd gnd FILL
XFILL_0__1303_ vdd gnd FILL
X_1793_ _1793_/A _1793_/B _1793_/C _1796_/A vdd gnd OAI21X1
X_1862_ _992_/Y _1880_/CLK _924_/A vdd gnd DFFPOSX1
XFILL_0__1234_ vdd gnd FILL
XFILL_3__1012_ vdd gnd FILL
XFILL_0__1165_ vdd gnd FILL
XFILL_3__1776_ vdd gnd FILL
XFILL_3__1914_ vdd gnd FILL
XFILL_0__1096_ vdd gnd FILL
XFILL_3__1845_ vdd gnd FILL
XFILL_1__1412_ vdd gnd FILL
XFILL_0_BUFX2_insert24 vdd gnd FILL
XFILL_1__967_ vdd gnd FILL
X_1227_ _956_/B Cin[3] _1240_/C vdd gnd NAND2X1
X_1158_ _1158_/A _1228_/A vdd gnd INVX1
XFILL_0_BUFX2_insert13 vdd gnd FILL
XFILL_1__1343_ vdd gnd FILL
XFILL_1__1274_ vdd gnd FILL
X_1089_ _1089_/A _1089_/B _1089_/C _1140_/B vdd gnd OAI21X1
XFILL_2__1521_ vdd gnd FILL
XFILL_2__1452_ vdd gnd FILL
XFILL_4__1319_ vdd gnd FILL
XFILL_2__1383_ vdd gnd FILL
XFILL100650x39150 vdd gnd FILL
XFILL_0__985_ vdd gnd FILL
XFILL_3__1630_ vdd gnd FILL
XFILL_2__1719_ vdd gnd FILL
XFILL_3__1561_ vdd gnd FILL
XFILL_0__1783_ vdd gnd FILL
XFILL_3__1492_ vdd gnd FILL
X_938_ _943_/A _938_/B _938_/C _940_/B vdd gnd OAI21X1
X_1012_ _947_/B _1843_/B vdd gnd INVX1
X_1914_ _954_/Y Xout[2] vdd gnd BUFX2
X_1776_ _1776_/A _1776_/B _1776_/C _1792_/A vdd gnd AOI21X1
XFILL_0__1079_ vdd gnd FILL
XFILL_0__1217_ vdd gnd FILL
XFILL_0__1148_ vdd gnd FILL
X_1845_ _951_/A _1845_/B _1845_/C _1903_/D vdd gnd OAI21X1
XFILL_3__1759_ vdd gnd FILL
XFILL_3__1828_ vdd gnd FILL
XFILL_1__1326_ vdd gnd FILL
XFILL_1__1257_ vdd gnd FILL
XFILL_1__1188_ vdd gnd FILL
XFILL_3__981_ vdd gnd FILL
XFILL_2__1504_ vdd gnd FILL
XFILL_4__1799_ vdd gnd FILL
XFILL_2__1435_ vdd gnd FILL
XFILL_2__1366_ vdd gnd FILL
XFILL_2__1297_ vdd gnd FILL
X_1630_ _1645_/A _1645_/B _1645_/C _1692_/A vdd gnd NAND3X1
XFILL_0__1002_ vdd gnd FILL
XFILL_0__968_ vdd gnd FILL
XFILL_3__1613_ vdd gnd FILL
X_1561_ _1635_/B _1575_/C _1635_/A _1562_/B vdd gnd AOI21X1
X_1492_ _1704_/C _1492_/B _1492_/C _1567_/A vdd gnd AOI21X1
XFILL_0__1835_ vdd gnd FILL
XFILL_3__1544_ vdd gnd FILL
XFILL_0__1697_ vdd gnd FILL
XFILL_0__1766_ vdd gnd FILL
XFILL_3__1475_ vdd gnd FILL
XFILL_1__1111_ vdd gnd FILL
XFILL_1__1042_ vdd gnd FILL
XFILL_4__946_ vdd gnd FILL
XFILL_4__1653_ vdd gnd FILL
X_1759_ _1759_/A _1759_/B _1759_/C _1776_/B vdd gnd NAND3X1
XFILL_4__1722_ vdd gnd FILL
X_1828_ _944_/A _928_/B _1895_/Q _1829_/C vdd gnd OAI21X1
XFILL_2__1220_ vdd gnd FILL
XFILL_2__1151_ vdd gnd FILL
XFILL_1__1309_ vdd gnd FILL
XFILL_4__1018_ vdd gnd FILL
XFILL_2__1082_ vdd gnd FILL
XFILL_3__964_ vdd gnd FILL
XFILL_0__1620_ vdd gnd FILL
XFILL_0__1551_ vdd gnd FILL
XFILL_0__1482_ vdd gnd FILL
XFILL_2__1418_ vdd gnd FILL
XFILL_3__1260_ vdd gnd FILL
XFILL_2__1349_ vdd gnd FILL
XFILL_3__1191_ vdd gnd FILL
X_1544_ _1554_/A _1620_/B _1547_/C _1625_/A vdd gnd AOI21X1
X_1613_ _1616_/B _1710_/A _1620_/C vdd gnd AND2X2
XFILL_1__1660_ vdd gnd FILL
XFILL_1__1591_ vdd gnd FILL
XFILL_3__1527_ vdd gnd FILL
X_1475_ _1552_/C _1498_/B _1498_/A _1480_/A vdd gnd AOI21X1
XFILL_0__1818_ vdd gnd FILL
XFILL_0__1749_ vdd gnd FILL
XFILL_3__1458_ vdd gnd FILL
XFILL_3__1389_ vdd gnd FILL
XFILL_2__982_ vdd gnd FILL
XBUFX2_insert15 Cin[0] _1449_/B vdd gnd BUFX2
XFILL_1__1025_ vdd gnd FILL
XFILL_1__1789_ vdd gnd FILL
XFILL_4__1498_ vdd gnd FILL
XFILL_4__1567_ vdd gnd FILL
XFILL_3_CLKBUF1_insert5 vdd gnd FILL
XFILL_2__1203_ vdd gnd FILL
XFILL_2__1134_ vdd gnd FILL
XFILL_2__1065_ vdd gnd FILL
X_1191_ _1191_/A _1228_/C _1231_/A vdd gnd AND2X2
X_1260_ _1361_/A _1269_/B _1269_/A _1371_/B vdd gnd NAND3X1
XFILL_3__947_ vdd gnd FILL
XFILL_0__1603_ vdd gnd FILL
XFILL_0__1534_ vdd gnd FILL
XFILL_0__1465_ vdd gnd FILL
XFILL_3__1312_ vdd gnd FILL
XFILL_3__1174_ vdd gnd FILL
XFILL_3__1243_ vdd gnd FILL
XFILL_0__1396_ vdd gnd FILL
X_1527_ _955_/A Cin[2] _1596_/B vdd gnd AND2X2
XFILL_1__1574_ vdd gnd FILL
XFILL_1__1712_ vdd gnd FILL
X_1458_ _1458_/A _1458_/B _1525_/A _1551_/A vdd gnd OAI21X1
XFILL_1__1643_ vdd gnd FILL
XFILL_4__1352_ vdd gnd FILL
XFILL_4__1421_ vdd gnd FILL
X_1389_ _1389_/A _1389_/B _1391_/A vdd gnd NOR2X1
XFILL_2__965_ vdd gnd FILL
XFILL_1__1008_ vdd gnd FILL
XFILL_2__1683_ vdd gnd FILL
XFILL_2__1821_ vdd gnd FILL
XFILL_2__1752_ vdd gnd FILL
X_971_ _996_/A _971_/B _971_/C _971_/Y vdd gnd OAI21X1
XFILL_2__1117_ vdd gnd FILL
XFILL_2__1048_ vdd gnd FILL
XFILL_0__1181_ vdd gnd FILL
XFILL_0__1250_ vdd gnd FILL
XFILL_3__1792_ vdd gnd FILL
X_1312_ _1315_/B _1315_/C _1315_/A _1321_/B vdd gnd AOI21X1
XFILL_1__983_ vdd gnd FILL
X_1174_ _1266_/C _1193_/C vdd gnd INVX1
X_1243_ _1243_/A _1243_/B _1243_/C _1360_/C vdd gnd OAI21X1
XFILL_0__1517_ vdd gnd FILL
XFILL_0__1448_ vdd gnd FILL
XFILL_3__1226_ vdd gnd FILL
XFILL_1__1290_ vdd gnd FILL
XFILL_3__1157_ vdd gnd FILL
XFILL_0__1379_ vdd gnd FILL
XFILL_3__1088_ vdd gnd FILL
XFILL_1__1626_ vdd gnd FILL
XFILL_1__1557_ vdd gnd FILL
XFILL_4__1266_ vdd gnd FILL
XFILL_1__1488_ vdd gnd FILL
XFILL_4__1197_ vdd gnd FILL
XFILL_2__948_ vdd gnd FILL
XFILL_2__1804_ vdd gnd FILL
XFILL_2__1735_ vdd gnd FILL
XFILL_2__1666_ vdd gnd FILL
XFILL_2__1597_ vdd gnd FILL
X_954_ _957_/A _963_/A _954_/C _954_/Y vdd gnd OAI21X1
XFILL_0__1302_ vdd gnd FILL
XFILL_3__1011_ vdd gnd FILL
X_1792_ _1792_/A _1792_/B _1799_/C _1798_/B vdd gnd OAI21X1
XFILL_2_CLKBUF1_insert10 vdd gnd FILL
X_1861_ _990_/Y _1903_/CLK _989_/A vdd gnd DFFPOSX1
XFILL_0__1233_ vdd gnd FILL
XFILL_3__1913_ vdd gnd FILL
XFILL_0__1095_ vdd gnd FILL
XFILL_0__1164_ vdd gnd FILL
XFILL_3__1775_ vdd gnd FILL
XFILL_1__966_ vdd gnd FILL
XFILL_3__1844_ vdd gnd FILL
XFILL_0_BUFX2_insert25 vdd gnd FILL
XFILL_1__1411_ vdd gnd FILL
XFILL_1__1342_ vdd gnd FILL
X_1226_ _1226_/A _1322_/A _1299_/B vdd gnd NOR2X1
XFILL_0_BUFX2_insert14 vdd gnd FILL
X_1157_ _1224_/B _1160_/B vdd gnd INVX1
XFILL_4__1120_ vdd gnd FILL
XFILL_3__1209_ vdd gnd FILL
XFILL_1__1273_ vdd gnd FILL
XFILL_4__1051_ vdd gnd FILL
X_1088_ _1088_/A _1088_/B _1102_/A _1089_/B vdd gnd AOI21X1
XFILL_2__1520_ vdd gnd FILL
XFILL_2__1451_ vdd gnd FILL
XFILL_1__1609_ vdd gnd FILL
XFILL_2__1382_ vdd gnd FILL
XFILL_0__984_ vdd gnd FILL
XFILL_3__1560_ vdd gnd FILL
XFILL_2__1649_ vdd gnd FILL
XFILL_2__1718_ vdd gnd FILL
XFILL_0__1782_ vdd gnd FILL
XFILL_3__1491_ vdd gnd FILL
X_937_ _943_/A _996_/B _938_/C vdd gnd NAND2X1
X_1011_ _947_/B _1106_/B _1898_/Q _1029_/A vdd gnd NAND3X1
X_1913_ _951_/Y Xout[1] vdd gnd BUFX2
XFILL_0__1216_ vdd gnd FILL
X_1775_ _1791_/A _1791_/B _1789_/A vdd gnd NOR2X1
XFILL_0__1078_ vdd gnd FILL
XFILL_0__1147_ vdd gnd FILL
X_1844_ _951_/A Xin[1] _1845_/C vdd gnd NAND2X1
XFILL_3__1689_ vdd gnd FILL
XFILL_3__1758_ vdd gnd FILL
XFILL_3__1827_ vdd gnd FILL
XFILL_1__949_ vdd gnd FILL
XFILL_1__1325_ vdd gnd FILL
X_1209_ _1209_/A _1209_/B _1209_/C _1213_/D vdd gnd OAI21X1
XFILL_1__1256_ vdd gnd FILL
XFILL_1__1187_ vdd gnd FILL
XFILL_3__980_ vdd gnd FILL
XFILL_2__1503_ vdd gnd FILL
XFILL_2__1434_ vdd gnd FILL
XFILL_2__1365_ vdd gnd FILL
XFILL_2__1296_ vdd gnd FILL
X_1560_ _1634_/A _1634_/B _1634_/C _1635_/B vdd gnd OAI21X1
XFILL_0__1001_ vdd gnd FILL
XFILL_0__967_ vdd gnd FILL
XFILL_3__1612_ vdd gnd FILL
XFILL_0__1765_ vdd gnd FILL
XFILL_3__1543_ vdd gnd FILL
X_1491_ _1571_/A _1492_/C vdd gnd INVX1
XFILL_0__1834_ vdd gnd FILL
XFILL_0__1696_ vdd gnd FILL
XFILL_3__1474_ vdd gnd FILL
X_1827_ _1827_/A _1833_/B _1827_/C _1894_/D vdd gnd OAI21X1
XFILL_1__1110_ vdd gnd FILL
XFILL_1__1041_ vdd gnd FILL
X_1689_ _1708_/B _1708_/A _1694_/A vdd gnd NAND2X1
X_1758_ _1776_/C _1760_/C vdd gnd INVX1
XFILL_1__1308_ vdd gnd FILL
XFILL_2__1081_ vdd gnd FILL
XFILL_2__1150_ vdd gnd FILL
XFILL_1__1239_ vdd gnd FILL
XFILL_3__963_ vdd gnd FILL
XFILL_0__1550_ vdd gnd FILL
XFILL_0__1481_ vdd gnd FILL
XFILL_2__1417_ vdd gnd FILL
XFILL_3__1190_ vdd gnd FILL
XFILL_2__1348_ vdd gnd FILL
XFILL_2__1279_ vdd gnd FILL
X_1612_ _1892_/Q _1612_/B _1710_/A vdd gnd NAND2X1
X_1543_ _1543_/A _1543_/B _1543_/C _1547_/C vdd gnd OAI21X1
X_1474_ _1474_/A _1474_/B _1474_/C _1479_/C vdd gnd OAI21X1
XFILL_1__1590_ vdd gnd FILL
XFILL_0__1748_ vdd gnd FILL
XFILL_3__1526_ vdd gnd FILL
XFILL_0__1817_ vdd gnd FILL
XFILL_0__1679_ vdd gnd FILL
XFILL_3__1457_ vdd gnd FILL
XFILL_4__928_ vdd gnd FILL
XFILL_3__1388_ vdd gnd FILL
XFILL_2__981_ vdd gnd FILL
XBUFX2_insert16 _1906_/Q _944_/A vdd gnd BUFX2
XFILL_1__1024_ vdd gnd FILL
XFILL_4__1635_ vdd gnd FILL
XFILL_4__1704_ vdd gnd FILL
XFILL_1__1788_ vdd gnd FILL
XFILL_3_CLKBUF1_insert6 vdd gnd FILL
XFILL_2__1202_ vdd gnd FILL
XFILL_2__1133_ vdd gnd FILL
XFILL_2__1064_ vdd gnd FILL
XFILL_0__1602_ vdd gnd FILL
XFILL_3__1311_ vdd gnd FILL
X_1190_ _1267_/A _1198_/B _1198_/A _1277_/B vdd gnd NAND3X1
XFILL_3__946_ vdd gnd FILL
XFILL_0__1464_ vdd gnd FILL
XFILL_0__1533_ vdd gnd FILL
XFILL_3__1242_ vdd gnd FILL
XFILL_3__1173_ vdd gnd FILL
XFILL_0__1395_ vdd gnd FILL
XFILL_1__1711_ vdd gnd FILL
X_1526_ _949_/A Cin[4] _1592_/A vdd gnd NAND2X1
X_1457_ _1465_/B _1458_/B vdd gnd INVX1
XFILL_3__1509_ vdd gnd FILL
XFILL_1__1573_ vdd gnd FILL
XFILL_1__1642_ vdd gnd FILL
X_1388_ _1389_/A _1389_/B _1396_/C _1392_/D vdd gnd OAI21X1
XFILL101250x46950 vdd gnd FILL
XFILL_2__964_ vdd gnd FILL
XFILL_2__1820_ vdd gnd FILL
XFILL_1__1007_ vdd gnd FILL
X_970_ _996_/A _970_/B _971_/C vdd gnd NAND2X1
XFILL_2__1682_ vdd gnd FILL
XFILL_4__1549_ vdd gnd FILL
XFILL_2__1751_ vdd gnd FILL
XFILL_4_BUFX2_insert17 vdd gnd FILL
XFILL_2__1047_ vdd gnd FILL
XFILL_0__1180_ vdd gnd FILL
XFILL_2__1116_ vdd gnd FILL
XFILL_3__1791_ vdd gnd FILL
X_1311_ _1847_/B _1413_/B _1311_/C _1315_/C vdd gnd OAI21X1
XFILL_1__982_ vdd gnd FILL
XFILL_3__929_ vdd gnd FILL
X_1242_ _1261_/B _1261_/A _1361_/A vdd gnd NAND2X1
X_1173_ _1173_/A _1173_/B _1173_/C _1266_/C vdd gnd OAI21X1
XFILL_0__1516_ vdd gnd FILL
XFILL_0__1447_ vdd gnd FILL
XFILL_3__1156_ vdd gnd FILL
XFILL_3__1225_ vdd gnd FILL
XFILL_3__1087_ vdd gnd FILL
XFILL_0__1378_ vdd gnd FILL
X_1509_ _1579_/C _1513_/B _1513_/A _1521_/A vdd gnd AOI21X1
XFILL_4__1403_ vdd gnd FILL
XFILL_1__1625_ vdd gnd FILL
XFILL_1__1556_ vdd gnd FILL
XFILL_1__1487_ vdd gnd FILL
XFILL101250x58650 vdd gnd FILL
XFILL_4__1334_ vdd gnd FILL
XFILL_2__947_ vdd gnd FILL
XFILL_2__1734_ vdd gnd FILL
XFILL_2__1803_ vdd gnd FILL
X_953_ _957_/A _953_/B _954_/C vdd gnd NAND2X1
XFILL_2__1665_ vdd gnd FILL
XFILL_2__1596_ vdd gnd FILL
XFILL_3__1010_ vdd gnd FILL
X_1860_ _987_/Y _1880_/CLK _986_/A vdd gnd DFFPOSX1
XFILL_0__1232_ vdd gnd FILL
XFILL_0__1301_ vdd gnd FILL
X_1791_ _1791_/A _1791_/B _1791_/C _1799_/C vdd gnd OAI21X1
XFILL_2_CLKBUF1_insert11 vdd gnd FILL
XFILL_3__1843_ vdd gnd FILL
XFILL_0__1094_ vdd gnd FILL
XFILL_0__1163_ vdd gnd FILL
XFILL_3__1912_ vdd gnd FILL
XFILL_3__1774_ vdd gnd FILL
XFILL_1__965_ vdd gnd FILL
XFILL_0_BUFX2_insert15 vdd gnd FILL
XFILL_1__1410_ vdd gnd FILL
XFILL_1__1341_ vdd gnd FILL
X_1156_ _1843_/B _1413_/B _1224_/B vdd gnd NOR2X1
X_1225_ _1319_/A _1322_/A vdd gnd INVX1
X_1087_ _1849_/B _1257_/B _1901_/Q _1088_/A vdd gnd OAI21X1
XFILL_3__1208_ vdd gnd FILL
XFILL_3__1139_ vdd gnd FILL
XFILL_1__1272_ vdd gnd FILL
XFILL_1__1608_ vdd gnd FILL
XFILL_2__1450_ vdd gnd FILL
XFILL_1__1539_ vdd gnd FILL
XFILL_4__1248_ vdd gnd FILL
XFILL_0__983_ vdd gnd FILL
XFILL_2__1381_ vdd gnd FILL
XFILL_4__1179_ vdd gnd FILL
XFILL_2__1717_ vdd gnd FILL
XFILL_0__1781_ vdd gnd FILL
XFILL_3__1490_ vdd gnd FILL
X_936_ _936_/A _996_/B vdd gnd INVX1
XFILL_2__1648_ vdd gnd FILL
XFILL_2__1579_ vdd gnd FILL
X_1010_ _1801_/A _1801_/B _1010_/C _1869_/D vdd gnd OAI21X1
XFILL_4__961_ vdd gnd FILL
X_1843_ _1848_/A _1843_/B _1843_/C _1902_/D vdd gnd OAI21X1
XFILL_0__1215_ vdd gnd FILL
X_1912_ _948_/Y Xout[0] vdd gnd BUFX2
X_1774_ _1774_/A _1774_/B _1774_/C _1791_/A vdd gnd OAI21X1
XFILL_3__1826_ vdd gnd FILL
XFILL_0__1146_ vdd gnd FILL
XFILL_0__1077_ vdd gnd FILL
XFILL_3__1688_ vdd gnd FILL
XFILL_3__1757_ vdd gnd FILL
X_1208_ _1208_/A _1208_/B _1278_/A _1209_/B vdd gnd AOI21X1
XFILL_1__948_ vdd gnd FILL
XFILL_1__1255_ vdd gnd FILL
XFILL_1__1324_ vdd gnd FILL
X_1139_ _1206_/C _1154_/B _1154_/A _1212_/B vdd gnd OAI21X1
XFILL_4__1102_ vdd gnd FILL
XFILL_4__1033_ vdd gnd FILL
XFILL_1__1186_ vdd gnd FILL
XFILL_2__1502_ vdd gnd FILL
XFILL_2__1433_ vdd gnd FILL
XFILL_2__1364_ vdd gnd FILL
XFILL_0__1000_ vdd gnd FILL
XFILL_0__966_ vdd gnd FILL
XFILL_2__1295_ vdd gnd FILL
X_1490_ _1702_/B _1490_/B _1490_/C _1878_/D vdd gnd OAI21X1
XFILL_3__1611_ vdd gnd FILL
XFILL_0__1764_ vdd gnd FILL
XFILL_3__1542_ vdd gnd FILL
XFILL_0__1833_ vdd gnd FILL
XFILL_3__1473_ vdd gnd FILL
XFILL_0__1695_ vdd gnd FILL
X_1826_ _1848_/A _928_/B _1894_/Q _1827_/C vdd gnd OAI21X1
XFILL_0__1129_ vdd gnd FILL
XFILL_1__1040_ vdd gnd FILL
X_1688_ _1688_/A _1733_/B _1688_/C _1694_/B vdd gnd NAND3X1
XFILL_4__1582_ vdd gnd FILL
X_1757_ _1759_/C _1759_/A _1759_/B _1776_/C vdd gnd AOI21X1
XFILL_3__1809_ vdd gnd FILL
XFILL_1__1307_ vdd gnd FILL
XFILL_1__1238_ vdd gnd FILL
XFILL_2__1080_ vdd gnd FILL
XFILL_1__1169_ vdd gnd FILL
XFILL_3__962_ vdd gnd FILL
XFILL_0__1480_ vdd gnd FILL
XFILL_2__1347_ vdd gnd FILL
XFILL_2__1416_ vdd gnd FILL
X_1611_ _1611_/A _1723_/B _1611_/C _1612_/B vdd gnd AOI21X1
XFILL_0__949_ vdd gnd FILL
XFILL_2__1278_ vdd gnd FILL
X_1542_ _1542_/A _1542_/B _1543_/B vdd gnd NOR2X1
X_1473_ _1473_/A _1473_/B _1473_/C _1474_/B vdd gnd AOI21X1
XFILL_0__1678_ vdd gnd FILL
XFILL_3__1525_ vdd gnd FILL
XFILL_0__1747_ vdd gnd FILL
XFILL_3__1456_ vdd gnd FILL
XFILL_0__1816_ vdd gnd FILL
XFILL_2__980_ vdd gnd FILL
XFILL_3__1387_ vdd gnd FILL
X_1809_ _1837_/B _1815_/B _1809_/C _1887_/D vdd gnd OAI21X1
XBUFX2_insert17 _1906_/Q _1848_/A vdd gnd BUFX2
XFILL_1__1023_ vdd gnd FILL
XFILL_1__1787_ vdd gnd FILL
XFILL_3_CLKBUF1_insert7 vdd gnd FILL
XFILL_2__1201_ vdd gnd FILL
XFILL_2__1132_ vdd gnd FILL
XFILL_2__1063_ vdd gnd FILL
XFILL_3__945_ vdd gnd FILL
XFILL_0__1601_ vdd gnd FILL
XFILL_0__1532_ vdd gnd FILL
XFILL_3__1310_ vdd gnd FILL
XFILL_0__1463_ vdd gnd FILL
XFILL_3__1241_ vdd gnd FILL
XFILL_3__1172_ vdd gnd FILL
XFILL_0__1394_ vdd gnd FILL
XFILL_1__1710_ vdd gnd FILL
X_1525_ _1525_/A _1525_/B _1555_/A _1554_/C vdd gnd AOI21X1
X_1456_ _1542_/A _1524_/C _1458_/A vdd gnd NOR2X1
XFILL_1__1641_ vdd gnd FILL
X_1387_ _1395_/A _1394_/A _1396_/C vdd gnd NAND2X1
XFILL_3__1508_ vdd gnd FILL
XFILL_3__1439_ vdd gnd FILL
XFILL_1__1572_ vdd gnd FILL
XFILL_4__1281_ vdd gnd FILL
XFILL_2__963_ vdd gnd FILL
XFILL_2__1750_ vdd gnd FILL
XFILL_1__1006_ vdd gnd FILL
XFILL_2__1681_ vdd gnd FILL
XFILL_4__1617_ vdd gnd FILL
XFILL_1__1839_ vdd gnd FILL
XFILL_2__1115_ vdd gnd FILL
XFILL_2__1046_ vdd gnd FILL
XFILL_3__1790_ vdd gnd FILL
XFILL_3__928_ vdd gnd FILL
X_1310_ _1845_/B _1778_/B _1424_/A _1315_/B vdd gnd OAI21X1
X_1241_ _1317_/B _1317_/A _1313_/C _1261_/B vdd gnd NAND3X1
XFILL_1__981_ vdd gnd FILL
XFILL_0__1515_ vdd gnd FILL
XFILL_3__1224_ vdd gnd FILL
X_1172_ _1228_/C _1191_/A _1267_/A vdd gnd NAND2X1
XFILL_0__1446_ vdd gnd FILL
XFILL_3__1155_ vdd gnd FILL
XFILL_3__1086_ vdd gnd FILL
XFILL_0__1377_ vdd gnd FILL
XFILL_1__1624_ vdd gnd FILL
X_1508_ _1579_/B _1513_/B vdd gnd INVX1
X_1439_ _952_/A Cin[3] _1611_/A vdd gnd AND2X2
XFILL_1__1555_ vdd gnd FILL
XFILL_1__1486_ vdd gnd FILL
XFILL_2__946_ vdd gnd FILL
XFILL_2__1733_ vdd gnd FILL
X_952_ _952_/A _963_/A vdd gnd INVX2
XFILL_2__1802_ vdd gnd FILL
XFILL_2__1664_ vdd gnd FILL
XFILL_2__1595_ vdd gnd FILL
X_1790_ _1790_/A _1790_/B _1790_/C _1884_/D vdd gnd OAI21X1
XFILL_0__1231_ vdd gnd FILL
XFILL_0__1300_ vdd gnd FILL
XFILL_0__1162_ vdd gnd FILL
XFILL_3__1773_ vdd gnd FILL
XFILL_2__1029_ vdd gnd FILL
XFILL_3__1842_ vdd gnd FILL
XFILL_3__1911_ vdd gnd FILL
XFILL_0__1093_ vdd gnd FILL
XFILL_0_BUFX2_insert16 vdd gnd FILL
XFILL_1__964_ vdd gnd FILL
X_1224_ _1311_/C _1224_/B _1319_/A vdd gnd NAND2X1
XFILL_1__1340_ vdd gnd FILL
X_1155_ Cin[5] _1413_/B vdd gnd INVX1
X_1086_ _956_/B _1849_/B vdd gnd INVX2
XFILL_3__1207_ vdd gnd FILL
XFILL_1__1271_ vdd gnd FILL
XFILL_0__1429_ vdd gnd FILL
XFILL_3__1138_ vdd gnd FILL
XFILL_3__1069_ vdd gnd FILL
XFILL_1__1538_ vdd gnd FILL
XFILL_1__1607_ vdd gnd FILL
XFILL_4__1316_ vdd gnd FILL
XFILL_2__1380_ vdd gnd FILL
XFILL_1__1469_ vdd gnd FILL
XFILL_0__982_ vdd gnd FILL
XFILL_2__929_ vdd gnd FILL
XFILL_2__1647_ vdd gnd FILL
XFILL_0__1780_ vdd gnd FILL
XFILL_2__1716_ vdd gnd FILL
X_935_ _945_/A _935_/B _935_/C _935_/Y vdd gnd OAI21X1
XFILL_2__1578_ vdd gnd FILL
X_1773_ _1773_/A _1773_/B _1774_/C vdd gnd NAND2X1
X_1842_ _1848_/A Xin[0] _1843_/C vdd gnd NAND2X1
X_1911_ _983_/A Vld vdd gnd BUFX2
XFILL_0__1145_ vdd gnd FILL
XFILL_0__1214_ vdd gnd FILL
XFILL_3__1756_ vdd gnd FILL
XFILL_3__1825_ vdd gnd FILL
XFILL_0__1076_ vdd gnd FILL
XFILL_3__1687_ vdd gnd FILL
X_1207_ _1221_/B _1278_/C _1221_/A _1209_/A vdd gnd AOI21X1
XFILL_1__947_ vdd gnd FILL
XFILL_1__1323_ vdd gnd FILL
X_1138_ _1138_/A _1138_/B _1141_/B _1141_/A _1206_/C vdd gnd AOI22X1
X_1069_ _953_/B Cin[1] _1102_/A vdd gnd NAND2X1
XFILL_1__1254_ vdd gnd FILL
XFILL_1__1185_ vdd gnd FILL
XFILL_2__1501_ vdd gnd FILL
XFILL_4__1796_ vdd gnd FILL
XFILL_2__1432_ vdd gnd FILL
XFILL_2__1363_ vdd gnd FILL
XFILL_2__1294_ vdd gnd FILL
XFILL100650x11850 vdd gnd FILL
XFILL100350x46950 vdd gnd FILL
XFILL_0__965_ vdd gnd FILL
XFILL100950x93750 vdd gnd FILL
XFILL_3__1610_ vdd gnd FILL
XFILL_0__1694_ vdd gnd FILL
XFILL_3__1541_ vdd gnd FILL
XFILL_0__1763_ vdd gnd FILL
XFILL_3__1472_ vdd gnd FILL
XFILL_0__1832_ vdd gnd FILL
XFILL_4__943_ vdd gnd FILL
X_1756_ _1780_/B _1887_/Q _1759_/B vdd gnd XNOR2X1
X_1825_ _965_/B _1833_/B vdd gnd INVX1
XFILL_3_BUFX2_insert20 vdd gnd FILL
XFILL_0__1128_ vdd gnd FILL
XFILL_0__1059_ vdd gnd FILL
X_1687_ _1687_/A _1687_/B _1687_/C _1688_/C vdd gnd OAI21X1
XFILL_4__1650_ vdd gnd FILL
XFILL_3__1739_ vdd gnd FILL
XFILL_3__1808_ vdd gnd FILL
XFILL_1__1306_ vdd gnd FILL
XFILL_1__1237_ vdd gnd FILL
XFILL_4__1015_ vdd gnd FILL
XFILL_1__1168_ vdd gnd FILL
XFILL_1__1099_ vdd gnd FILL
XFILL_4__1917_ vdd gnd FILL
XFILL_3__961_ vdd gnd FILL
XFILL100650x23550 vdd gnd FILL
XFILL100350x58650 vdd gnd FILL
XFILL_2__1346_ vdd gnd FILL
XFILL_2__1415_ vdd gnd FILL
XFILL_2__1277_ vdd gnd FILL
X_1610_ _1611_/C _1670_/C _1822_/A _1616_/B vdd gnd OAI21X1
XFILL_0__948_ vdd gnd FILL
X_1541_ _1554_/C _1555_/C _1578_/C vdd gnd NOR2X1
XFILL_0__1815_ vdd gnd FILL
X_1472_ _1479_/A _1479_/B _1480_/C _1486_/A vdd gnd NAND3X1
XFILL_0__1677_ vdd gnd FILL
XFILL_0__1746_ vdd gnd FILL
XFILL_3__1524_ vdd gnd FILL
XFILL_3__1455_ vdd gnd FILL
XFILL_3__1386_ vdd gnd FILL
XBUFX2_insert18 _1906_/Q _948_/A vdd gnd BUFX2
XFILL_1__1022_ vdd gnd FILL
X_1739_ _1740_/A _1741_/A _1741_/B _1771_/A vdd gnd NAND3X1
X_1808_ _1887_/Q _1815_/B _1809_/C vdd gnd NAND2X1
XFILL_4__1564_ vdd gnd FILL
XFILL_1__1786_ vdd gnd FILL
XFILL_4__1495_ vdd gnd FILL
XFILL_3_CLKBUF1_insert8 vdd gnd FILL
XFILL_2__1200_ vdd gnd FILL
XFILL_2__1131_ vdd gnd FILL
XFILL_2__1062_ vdd gnd FILL
XFILL_3__944_ vdd gnd FILL
XFILL100650x35250 vdd gnd FILL
XFILL_0__1600_ vdd gnd FILL
XFILL_0__1531_ vdd gnd FILL
XFILL_0__1462_ vdd gnd FILL
XFILL_3__1240_ vdd gnd FILL
XFILL_0__1393_ vdd gnd FILL
XFILL_2__1329_ vdd gnd FILL
XFILL_3__1171_ vdd gnd FILL
X_1524_ _1524_/A _1524_/B _1524_/C _1555_/A vdd gnd AOI21X1
XFILL_3__1507_ vdd gnd FILL
XFILL_1__1571_ vdd gnd FILL
X_1455_ _1605_/B _1455_/B _1524_/C vdd gnd NAND2X1
XFILL_1__1640_ vdd gnd FILL
X_1386_ _1386_/A _1386_/B _1386_/C _1395_/A vdd gnd NAND3X1
XFILL_0__1729_ vdd gnd FILL
XFILL_3__1438_ vdd gnd FILL
XFILL_3__1369_ vdd gnd FILL
XFILL_2__962_ vdd gnd FILL
XFILL_1__1005_ vdd gnd FILL
XFILL_2__1680_ vdd gnd FILL
XFILL_1__1769_ vdd gnd FILL
XFILL_1__1838_ vdd gnd FILL
XFILL_2__1114_ vdd gnd FILL
XFILL_2__1045_ vdd gnd FILL
XFILL_3__927_ vdd gnd FILL
XFILL_1__980_ vdd gnd FILL
X_1240_ _959_/A _1533_/D _1240_/C _1317_/B vdd gnd OAI21X1
X_1171_ _1171_/A _1171_/B _1171_/C _1228_/C vdd gnd NAND3X1
XFILL_0__1514_ vdd gnd FILL
XFILL_0__1445_ vdd gnd FILL
XFILL_3__1223_ vdd gnd FILL
XFILL_3__1154_ vdd gnd FILL
XFILL_3__1085_ vdd gnd FILL
XFILL_0__1376_ vdd gnd FILL
X_1507_ _1507_/A _1589_/A _1579_/C vdd gnd NAND2X1
XFILL_1__1623_ vdd gnd FILL
XFILL_1__1554_ vdd gnd FILL
X_1438_ _1511_/A _1515_/D vdd gnd INVX1
X_1369_ _1474_/C _1402_/A _1402_/B _1397_/B vdd gnd NAND3X1
XFILL_4__1263_ vdd gnd FILL
XFILL_1__1485_ vdd gnd FILL
XFILL_2__945_ vdd gnd FILL
XFILL_4__1194_ vdd gnd FILL
XFILL_2__1663_ vdd gnd FILL
XFILL_2__1732_ vdd gnd FILL
XFILL_2__1801_ vdd gnd FILL
X_951_ _951_/A _961_/A _951_/C _951_/Y vdd gnd OAI21X1
XFILL_2__1594_ vdd gnd FILL
XFILL_2__1028_ vdd gnd FILL
XFILL_0__1161_ vdd gnd FILL
XFILL_0__1092_ vdd gnd FILL
XFILL_0__1230_ vdd gnd FILL
XFILL_3__1772_ vdd gnd FILL
XFILL_3__1841_ vdd gnd FILL
X_1223_ _950_/B Cin[6] _1311_/C vdd gnd AND2X2
XFILL_0_BUFX2_insert17 vdd gnd FILL
XFILL_1__963_ vdd gnd FILL
X_1154_ _1154_/A _1154_/B _1154_/C _1205_/C vdd gnd OAI21X1
XFILL_0__1428_ vdd gnd FILL
XFILL_3__1206_ vdd gnd FILL
XFILL_3__1137_ vdd gnd FILL
XFILL_1__1270_ vdd gnd FILL
X_1085_ _956_/B _1104_/B _1841_/B _1088_/B vdd gnd NAND3X1
XFILL_0__1359_ vdd gnd FILL
XFILL_3__1068_ vdd gnd FILL
XFILL_1__1537_ vdd gnd FILL
XFILL_1__1606_ vdd gnd FILL
XFILL_1__1468_ vdd gnd FILL
XFILL_2__928_ vdd gnd FILL
XFILL_1__1399_ vdd gnd FILL
XFILL_0__981_ vdd gnd FILL
XFILL_2__1646_ vdd gnd FILL
XFILL_2__1715_ vdd gnd FILL
X_934_ _944_/A _969_/A _965_/B _981_/A _935_/C vdd gnd AOI22X1
XFILL_2__1577_ vdd gnd FILL
X_1910_ _1910_/D _1910_/CLK _1910_/Q vdd gnd DFFPOSX1
X_1772_ _1772_/A _1772_/B _1772_/C _1791_/B vdd gnd AOI21X1
XFILL_0__1213_ vdd gnd FILL
XFILL_0__1144_ vdd gnd FILL
XFILL_0__1075_ vdd gnd FILL
X_1841_ _948_/A _1841_/B _1841_/C _1901_/D vdd gnd OAI21X1
XFILL_3__1686_ vdd gnd FILL
XFILL_3__1755_ vdd gnd FILL
XFILL_3__1824_ vdd gnd FILL
XFILL99750x70350 vdd gnd FILL
X_1206_ _1206_/A _1206_/B _1206_/C _1209_/C vdd gnd AOI21X1
X_1137_ _1196_/B _1161_/C _1161_/A _1141_/B vdd gnd OAI21X1
XFILL_1__946_ vdd gnd FILL
XFILL_1__1322_ vdd gnd FILL
X_1068_ _1068_/A _1068_/B _1068_/C _1082_/A vdd gnd OAI21X1
XFILL_1__1184_ vdd gnd FILL
XFILL_1__1253_ vdd gnd FILL
XFILL_2__1500_ vdd gnd FILL
XFILL_2__1431_ vdd gnd FILL
XFILL_2__1362_ vdd gnd FILL
XFILL_2__1293_ vdd gnd FILL
XFILL_0__964_ vdd gnd FILL
XFILL_3__1540_ vdd gnd FILL
XFILL_0__1831_ vdd gnd FILL
XFILL_2__1629_ vdd gnd FILL
XFILL_0__1693_ vdd gnd FILL
XFILL_0__1762_ vdd gnd FILL
XFILL_3__1471_ vdd gnd FILL
X_1686_ _1695_/C _1695_/B _1695_/A _1691_/C vdd gnd NAND3X1
X_1755_ _1777_/B _1777_/A _1780_/B vdd gnd XOR2X1
X_1824_ _1824_/A _1824_/B _1824_/C _1893_/D vdd gnd OAI21X1
XFILL_3_BUFX2_insert21 vdd gnd FILL
XFILL_0__1127_ vdd gnd FILL
XFILL_0__1058_ vdd gnd FILL
XFILL_3__1669_ vdd gnd FILL
XFILL_3__1738_ vdd gnd FILL
XFILL_3__1807_ vdd gnd FILL
XFILL_1__929_ vdd gnd FILL
XFILL_1__1305_ vdd gnd FILL
XFILL_1__1236_ vdd gnd FILL
XFILL_1__1098_ vdd gnd FILL
XFILL_1__1167_ vdd gnd FILL
XFILL_4__1778_ vdd gnd FILL
XFILL_4__1847_ vdd gnd FILL
XFILL_3__960_ vdd gnd FILL
XFILL_2__1414_ vdd gnd FILL
XFILL_2__1345_ vdd gnd FILL
XFILL_2__1276_ vdd gnd FILL
X_1540_ _1620_/B _1554_/A _1555_/C vdd gnd NAND2X1
XFILL_0__947_ vdd gnd FILL
XFILL_3__1523_ vdd gnd FILL
X_1471_ _1552_/C _1498_/B _1498_/A _1479_/B vdd gnd NAND3X1
XFILL_0__1814_ vdd gnd FILL
XFILL_0__1676_ vdd gnd FILL
XFILL_3__1454_ vdd gnd FILL
XFILL_0__1745_ vdd gnd FILL
XFILL_3__1385_ vdd gnd FILL
X_1807_ Yin[1] _1837_/B vdd gnd INVX1
XFILL_4__925_ vdd gnd FILL
XBUFX2_insert19 _1906_/Q _951_/A vdd gnd BUFX2
XFILL_1__1021_ vdd gnd FILL
XFILL_4__1632_ vdd gnd FILL
X_1669_ _1680_/A _1679_/A vdd gnd INVX1
X_1738_ _1748_/C _1738_/B _1738_/C _1741_/B vdd gnd OAI21X1
XFILL_4__1701_ vdd gnd FILL
XFILL_1__1785_ vdd gnd FILL
XFILL_3_CLKBUF1_insert9 vdd gnd FILL
XFILL_2__1061_ vdd gnd FILL
XFILL_2__1130_ vdd gnd FILL
XFILL_1__1219_ vdd gnd FILL
XFILL100950x19650 vdd gnd FILL
XFILL_3__943_ vdd gnd FILL
XFILL_0__1530_ vdd gnd FILL
XFILL_0__1461_ vdd gnd FILL
XFILL_3__1170_ vdd gnd FILL
XFILL_2__1328_ vdd gnd FILL
XFILL_0__1392_ vdd gnd FILL
XFILL_2__1259_ vdd gnd FILL
X_1523_ _1553_/A _1576_/B _1625_/B vdd gnd NAND2X1
X_1454_ _1454_/A _1455_/B vdd gnd INVX1
XFILL_2_BUFX2_insert0 vdd gnd FILL
XFILL_3__1506_ vdd gnd FILL
XFILL_0__1728_ vdd gnd FILL
XFILL_1__1570_ vdd gnd FILL
X_1385_ _1398_/A _1385_/B _1385_/C _1386_/C vdd gnd NAND3X1
XFILL_0__1659_ vdd gnd FILL
XFILL_3__1437_ vdd gnd FILL
XFILL_3__1368_ vdd gnd FILL
XFILL_3__1299_ vdd gnd FILL
XFILL_2__961_ vdd gnd FILL
XFILL_1__1004_ vdd gnd FILL
XFILL_4__1546_ vdd gnd FILL
XFILL_4__1615_ vdd gnd FILL
XFILL_1__1837_ vdd gnd FILL
XFILL_1__1768_ vdd gnd FILL
XFILL_1__1699_ vdd gnd FILL
XFILL_4__1477_ vdd gnd FILL
XFILL_2__1113_ vdd gnd FILL
XFILL_2__1044_ vdd gnd FILL
XFILL_3__926_ vdd gnd FILL
X_1170_ _1847_/B _1533_/B _1849_/B _1533_/D _1171_/B vdd gnd OAI22X1
XFILL_0__1513_ vdd gnd FILL
XFILL_0__1444_ vdd gnd FILL
XFILL_3__1222_ vdd gnd FILL
XFILL_0__1375_ vdd gnd FILL
XFILL_3__1153_ vdd gnd FILL
XFILL_3__1084_ vdd gnd FILL
X_1506_ _946_/A Cin[6] _1589_/A vdd gnd AND2X2
X_1437_ _1511_/A _1437_/B _1437_/C _1453_/B vdd gnd NAND3X1
XFILL_4__1400_ vdd gnd FILL
XFILL_1__1553_ vdd gnd FILL
XFILL_1__1622_ vdd gnd FILL
XFILL_4__1331_ vdd gnd FILL
X_1368_ _1368_/A _1368_/B _1368_/C _1402_/B vdd gnd OAI21X1
XFILL_1__1484_ vdd gnd FILL
X_1299_ _1299_/A _1299_/B _1398_/A vdd gnd NAND2X1
XFILL_2__944_ vdd gnd FILL
XFILL_2__1800_ vdd gnd FILL
X_950_ _951_/A _950_/B _951_/C vdd gnd NAND2X1
XFILL_2__1731_ vdd gnd FILL
XFILL_2__1593_ vdd gnd FILL
XFILL_2__1662_ vdd gnd FILL
XFILL_2__1027_ vdd gnd FILL
XFILL_0__1160_ vdd gnd FILL
XFILL_0__1091_ vdd gnd FILL
XFILL_3__1771_ vdd gnd FILL
XFILL_3__1840_ vdd gnd FILL
XFILL_1__962_ vdd gnd FILL
X_1222_ _947_/B Cin[6] _950_/B Cin[5] _1226_/A vdd gnd AOI22X1
XFILL_0_BUFX2_insert18 vdd gnd FILL
X_1153_ _1153_/A _1210_/C vdd gnd INVX1
X_1084_ _1901_/Q _1841_/B vdd gnd INVX1
XFILL_0__1427_ vdd gnd FILL
XFILL_0__1358_ vdd gnd FILL
XFILL_3__1205_ vdd gnd FILL
XFILL_3__1136_ vdd gnd FILL
XFILL_3__1067_ vdd gnd FILL
XFILL_0__1289_ vdd gnd FILL
XFILL_1__1536_ vdd gnd FILL
XFILL_1__1605_ vdd gnd FILL
XFILL_1__1467_ vdd gnd FILL
XFILL_4__1176_ vdd gnd FILL
XFILL_4__1245_ vdd gnd FILL
XFILL_1__1398_ vdd gnd FILL
XFILL_2__927_ vdd gnd FILL
XFILL_0__980_ vdd gnd FILL
XFILL_2__1714_ vdd gnd FILL
X_933_ _943_/A _933_/B _933_/C _935_/B vdd gnd OAI21X1
XFILL_2__1645_ vdd gnd FILL
XFILL_2__1576_ vdd gnd FILL
X_1840_ _948_/A Yin[3] _1841_/C vdd gnd NAND2X1
XFILL_0__1212_ vdd gnd FILL
X_1771_ _1771_/A _1773_/A _1771_/C _1772_/C vdd gnd NAND3X1
XFILL_3__1823_ vdd gnd FILL
XFILL_0__1143_ vdd gnd FILL
XFILL_0__1074_ vdd gnd FILL
XFILL_3__1685_ vdd gnd FILL
XFILL_3__1754_ vdd gnd FILL
XFILL_1__945_ vdd gnd FILL
XFILL_1__1321_ vdd gnd FILL
XFILL_4__1030_ vdd gnd FILL
X_1205_ _1205_/A _1205_/B _1205_/C _1290_/C vdd gnd NAND3X1
X_1136_ _1196_/C _1196_/A _1161_/B _1141_/A vdd gnd NAND3X1
X_1067_ _1067_/A _1206_/B _1140_/A vdd gnd NOR2X1
XFILL_1__1183_ vdd gnd FILL
XFILL_3__1119_ vdd gnd FILL
XFILL_1__1252_ vdd gnd FILL
XFILL_2__1430_ vdd gnd FILL
XFILL_1__1519_ vdd gnd FILL
XFILL_2__1361_ vdd gnd FILL
XFILL_2__1292_ vdd gnd FILL
XFILL_0__963_ vdd gnd FILL
XFILL_0__1761_ vdd gnd FILL
XFILL_3__1470_ vdd gnd FILL
XFILL_0__1830_ vdd gnd FILL
XFILL_2__1628_ vdd gnd FILL
XFILL_0__1692_ vdd gnd FILL
XFILL_2__1559_ vdd gnd FILL
X_1823_ Yin[3] _1824_/B _1824_/C vdd gnd NAND2X1
X_1685_ _1685_/A _1685_/B _1708_/B _1695_/B vdd gnd OAI21X1
X_1754_ _1754_/A _1754_/B _1777_/B vdd gnd AND2X2
XFILL_3__1806_ vdd gnd FILL
XFILL_3_BUFX2_insert22 vdd gnd FILL
XFILL_0__1126_ vdd gnd FILL
XFILL_0__1057_ vdd gnd FILL
XFILL_3__1668_ vdd gnd FILL
XFILL_3__1737_ vdd gnd FILL
XFILL_3__1599_ vdd gnd FILL
XFILL_1__928_ vdd gnd FILL
XFILL_1__1304_ vdd gnd FILL
XFILL_1__1235_ vdd gnd FILL
X_1119_ _953_/B Cin[2] _1158_/A vdd gnd AND2X2
XFILL101250x54750 vdd gnd FILL
XFILL_1__1097_ vdd gnd FILL
XFILL_1__1166_ vdd gnd FILL
XFILL_2__1344_ vdd gnd FILL
XFILL_2__1413_ vdd gnd FILL
XFILL_2__1275_ vdd gnd FILL
XFILL100950x150 vdd gnd FILL
XFILL_0__946_ vdd gnd FILL
X_1470_ _1555_/B _1470_/B _1470_/C _1498_/B vdd gnd OAI21X1
XFILL_3__1522_ vdd gnd FILL
XFILL_3__1453_ vdd gnd FILL
XFILL_0__1744_ vdd gnd FILL
XFILL_0__1813_ vdd gnd FILL
XFILL_0__1675_ vdd gnd FILL
XFILL_3__1384_ vdd gnd FILL
X_1806_ _1827_/A _1815_/B _1806_/C _1886_/D vdd gnd OAI21X1
XFILL_1__1020_ vdd gnd FILL
XFILL_0__1109_ vdd gnd FILL
X_1668_ _1680_/C _1709_/A _1680_/A _1678_/A vdd gnd AOI21X1
X_1737_ _1748_/A _1738_/B vdd gnd INVX1
X_1599_ _1599_/A _1599_/B _1599_/C _1649_/A vdd gnd NAND3X1
XFILL_1__1784_ vdd gnd FILL
XFILL101250x66450 vdd gnd FILL
XFILL_1__1218_ vdd gnd FILL
XFILL_2__1060_ vdd gnd FILL
XFILL_1__1149_ vdd gnd FILL
XFILL_3__942_ vdd gnd FILL
XFILL_4__1829_ vdd gnd FILL
XFILL_0__1460_ vdd gnd FILL
XFILL_2__1327_ vdd gnd FILL
XFILL_0__1391_ vdd gnd FILL
XFILL_0__929_ vdd gnd FILL
XFILL_2__1258_ vdd gnd FILL
XFILL_2__1189_ vdd gnd FILL
X_1522_ _1522_/A _1576_/A _1522_/C _1576_/B vdd gnd NAND3X1
X_1453_ _1453_/A _1453_/B _1525_/A vdd gnd AND2X2
XFILL_2_BUFX2_insert1 vdd gnd FILL
XFILL_3__1505_ vdd gnd FILL
XFILL_0__1727_ vdd gnd FILL
XFILL_0__1658_ vdd gnd FILL
XFILL_3__1436_ vdd gnd FILL
X_1384_ _1484_/A _1483_/A _1484_/B _1386_/B vdd gnd NAND3X1
XFILL_0__1589_ vdd gnd FILL
XFILL_3__1367_ vdd gnd FILL
XFILL_3__1298_ vdd gnd FILL
XFILL_2__960_ vdd gnd FILL
XFILL_1__1003_ vdd gnd FILL
XFILL_1__1767_ vdd gnd FILL
XFILL_1__1836_ vdd gnd FILL
XFILL101250x78150 vdd gnd FILL
XFILL_1__1698_ vdd gnd FILL
XFILL_2__1112_ vdd gnd FILL
XFILL_2__1043_ vdd gnd FILL
XFILL_3__925_ vdd gnd FILL
XFILL_0__1512_ vdd gnd FILL
XFILL_0__1443_ vdd gnd FILL
XFILL_0__1374_ vdd gnd FILL
XFILL_3__1221_ vdd gnd FILL
XFILL_3__1083_ vdd gnd FILL
XFILL_3__1152_ vdd gnd FILL
X_1505_ _1579_/A _1513_/A vdd gnd INVX1
XFILL_1__1621_ vdd gnd FILL
X_1436_ _949_/A Cin[3] _1510_/B _1437_/C vdd gnd NAND3X1
X_1367_ _1473_/B _1473_/A _1473_/C _1474_/C vdd gnd NAND3X1
XFILL_1__1483_ vdd gnd FILL
XFILL_1__1552_ vdd gnd FILL
XFILL_3__1419_ vdd gnd FILL
X_1298_ _1298_/A _1298_/B _1298_/C _1381_/C vdd gnd AOI21X1
XFILL_2__943_ vdd gnd FILL
XFILL_2__1730_ vdd gnd FILL
XFILL_2__1661_ vdd gnd FILL
XFILL_2__1592_ vdd gnd FILL
XFILL_1__1819_ vdd gnd FILL
XFILL_4__1528_ vdd gnd FILL
XFILL_4__1459_ vdd gnd FILL
XFILL_2__1026_ vdd gnd FILL
XFILL_0__1090_ vdd gnd FILL
XFILL100050x70350 vdd gnd FILL
XFILL_3__1770_ vdd gnd FILL
X_1221_ _1221_/A _1221_/B _1221_/C _1285_/C vdd gnd AOI21X1
XFILL_1__961_ vdd gnd FILL
XFILL_3__1204_ vdd gnd FILL
X_1083_ _1083_/A _1102_/C _1083_/C _1089_/A vdd gnd AOI21X1
X_1152_ _982_/B _1216_/A _1216_/C vdd gnd NAND2X1
XFILL_0_BUFX2_insert19 vdd gnd FILL
XFILL_0__1357_ vdd gnd FILL
XFILL_0__1426_ vdd gnd FILL
XFILL_0__1288_ vdd gnd FILL
XFILL_3__1135_ vdd gnd FILL
XFILL_3__1066_ vdd gnd FILL
XFILL_1__1604_ vdd gnd FILL
X_1419_ _1419_/A _1419_/B _1499_/B _1519_/C vdd gnd NAND3X1
XFILL_4__1313_ vdd gnd FILL
XFILL_1__1535_ vdd gnd FILL
XFILL_1__1466_ vdd gnd FILL
XFILL_1__1397_ vdd gnd FILL
XFILL_2__926_ vdd gnd FILL
XFILL_2__1713_ vdd gnd FILL
X_932_ _943_/A _994_/B _933_/C vdd gnd NAND2X1
XFILL_2__1575_ vdd gnd FILL
XFILL_2__1644_ vdd gnd FILL
X_1770_ _1884_/Q _1790_/A _1790_/C vdd gnd NAND2X1
XFILL_0__1142_ vdd gnd FILL
XFILL_0__1211_ vdd gnd FILL
XFILL_3__1822_ vdd gnd FILL
XFILL_2__1009_ vdd gnd FILL
XFILL_0__1073_ vdd gnd FILL
XFILL_3__1684_ vdd gnd FILL
XFILL_3__1753_ vdd gnd FILL
XFILL_1__944_ vdd gnd FILL
X_1204_ _1278_/C _1221_/A _1221_/B _1205_/B vdd gnd NAND3X1
XFILL_1__1320_ vdd gnd FILL
X_1135_ _1140_/A _1138_/A _1140_/B _1138_/B vdd gnd NAND3X1
X_1066_ _947_/B Cin[3] _950_/B Cin[2] _1067_/A vdd gnd AOI22X1
XFILL_1__1251_ vdd gnd FILL
XFILL_0__1409_ vdd gnd FILL
X_1899_ _1899_/D _1908_/CLK _1899_/Q vdd gnd DFFPOSX1
XFILL_1__1182_ vdd gnd FILL
XFILL_3__1118_ vdd gnd FILL
XFILL_3__1049_ vdd gnd FILL
XFILL_4__1793_ vdd gnd FILL
XFILL_2__1360_ vdd gnd FILL
XFILL_1__1518_ vdd gnd FILL
XFILL_1__1449_ vdd gnd FILL
XFILL_2__1291_ vdd gnd FILL
XFILL_4__1227_ vdd gnd FILL
XFILL_4__1158_ vdd gnd FILL
XFILL_0__962_ vdd gnd FILL
XFILL_2__1627_ vdd gnd FILL
XFILL_0__1691_ vdd gnd FILL
XFILL_0__1760_ vdd gnd FILL
XFILL_2__1558_ vdd gnd FILL
XFILL_2__1489_ vdd gnd FILL
XFILL_4__940_ vdd gnd FILL
X_1822_ _1822_/A _1824_/B _1822_/C _1892_/D vdd gnd OAI21X1
X_1753_ _1794_/B _1794_/C _1754_/A vdd gnd NAND2X1
XFILL_0__1125_ vdd gnd FILL
XFILL_3_BUFX2_insert12 vdd gnd FILL
X_1684_ _1688_/A _1733_/B _1708_/B vdd gnd NAND2X1
XFILL_3__1736_ vdd gnd FILL
XFILL_3__1805_ vdd gnd FILL
XFILL_3_BUFX2_insert23 vdd gnd FILL
XFILL_0__1056_ vdd gnd FILL
XFILL_3__1667_ vdd gnd FILL
XFILL_3__1598_ vdd gnd FILL
XFILL_1__927_ vdd gnd FILL
XFILL_1__1303_ vdd gnd FILL
XFILL_1__1234_ vdd gnd FILL
X_1118_ _950_/B Cin[3] _1124_/C vdd gnd AND2X2
X_1049_ _1049_/A _1049_/B _1062_/A vdd gnd NAND2X1
XFILL_4__1012_ vdd gnd FILL
XFILL_4__1914_ vdd gnd FILL
XFILL_1__1096_ vdd gnd FILL
XFILL_1__1165_ vdd gnd FILL
XFILL_4__1776_ vdd gnd FILL
XFILL_2__1343_ vdd gnd FILL
XFILL_2__1412_ vdd gnd FILL
XFILL_2__1274_ vdd gnd FILL
XFILL_0__945_ vdd gnd FILL
XFILL_3__1521_ vdd gnd FILL
XFILL_0__1674_ vdd gnd FILL
XFILL_0__1743_ vdd gnd FILL
XFILL_3__1452_ vdd gnd FILL
XFILL_0__1812_ vdd gnd FILL
XFILL_3__1383_ vdd gnd FILL
X_1736_ _1736_/A _1748_/C vdd gnd INVX1
X_1805_ _1886_/Q _1815_/B _1806_/C vdd gnd NAND2X1
XFILL_0__1108_ vdd gnd FILL
XFILL_0__1039_ vdd gnd FILL
X_1667_ _1720_/B _1670_/B _1671_/B _1680_/C vdd gnd OAI21X1
X_1598_ _1600_/A _1600_/B _1601_/C _1599_/B vdd gnd NAND3X1
XFILL_3__1719_ vdd gnd FILL
XFILL_4__1561_ vdd gnd FILL
XFILL_1__1783_ vdd gnd FILL
XFILL_4__1492_ vdd gnd FILL
XFILL_1__1217_ vdd gnd FILL
XFILL_1__1148_ vdd gnd FILL
XFILL_3__941_ vdd gnd FILL
XFILL_1__1079_ vdd gnd FILL
XFILL_2__1326_ vdd gnd FILL
XFILL_2__1257_ vdd gnd FILL
XFILL_0__1390_ vdd gnd FILL
XFILL_0__928_ vdd gnd FILL
XFILL_2__1188_ vdd gnd FILL
X_1521_ _1521_/A _1521_/B _1521_/C _1522_/C vdd gnd OAI21X1
X_1452_ _1465_/B _1543_/A _1465_/A _1551_/B vdd gnd NAND3X1
XFILL_2_BUFX2_insert2 vdd gnd FILL
X_1383_ _1383_/A _1383_/B _1383_/C _1386_/A vdd gnd OAI21X1
XFILL_0__1726_ vdd gnd FILL
XFILL_3__1504_ vdd gnd FILL
XFILL_3__1435_ vdd gnd FILL
XFILL_0__1657_ vdd gnd FILL
XFILL_3__1366_ vdd gnd FILL
XFILL_0__1588_ vdd gnd FILL
XFILL_1__1002_ vdd gnd FILL
XFILL_3__1297_ vdd gnd FILL
X_1719_ _1728_/B _1728_/A _1727_/A vdd gnd NOR2X1
XFILL_1__1766_ vdd gnd FILL
XFILL_1__1835_ vdd gnd FILL
XFILL_1__1697_ vdd gnd FILL
XFILL_2__1111_ vdd gnd FILL
XFILL_2__1042_ vdd gnd FILL
XFILL_3__924_ vdd gnd FILL
XFILL_0__1511_ vdd gnd FILL
XFILL_3__1220_ vdd gnd FILL
XFILL_0__1373_ vdd gnd FILL
XFILL_0__1442_ vdd gnd FILL
XFILL_2__1309_ vdd gnd FILL
XFILL_3__1082_ vdd gnd FILL
XFILL_3__1151_ vdd gnd FILL
X_1504_ _1579_/A _1579_/B _1514_/B _1521_/B vdd gnd NOR3X1
XFILL_1__1620_ vdd gnd FILL
X_1435_ _952_/A Cin[2] _1510_/B vdd gnd NAND2X1
XFILL_1__1551_ vdd gnd FILL
X_1366_ _1366_/A _1399_/B _1402_/A vdd gnd AND2X2
XFILL_0__1709_ vdd gnd FILL
XFILL_3__1349_ vdd gnd FILL
XFILL_1__1482_ vdd gnd FILL
XFILL_3__1418_ vdd gnd FILL
XFILL_2__942_ vdd gnd FILL
X_1297_ _1383_/C _1298_/C vdd gnd INVX1
XFILL_4__1191_ vdd gnd FILL
XFILL_4__1260_ vdd gnd FILL
XFILL_2__1660_ vdd gnd FILL
XFILL_2__1591_ vdd gnd FILL
XFILL_1__1749_ vdd gnd FILL
XFILL_1__1818_ vdd gnd FILL
XFILL_2__1025_ vdd gnd FILL
XFILL_2__1789_ vdd gnd FILL
X_1220_ _1278_/C _1221_/C vdd gnd INVX1
X_1151_ _1151_/A _1151_/B _1151_/C _1874_/D vdd gnd OAI21X1
XFILL_1__960_ vdd gnd FILL
XFILL_0__1425_ vdd gnd FILL
XFILL_3__1203_ vdd gnd FILL
X_1082_ _1082_/A _1089_/C vdd gnd INVX1
XFILL_0__1356_ vdd gnd FILL
XFILL_0__1287_ vdd gnd FILL
XFILL_3__1134_ vdd gnd FILL
XFILL_3__1065_ vdd gnd FILL
XFILL_1__1603_ vdd gnd FILL
XFILL_1__1534_ vdd gnd FILL
X_1349_ _1524_/A _1351_/C _1351_/A _1524_/B vdd gnd NAND3X1
X_1418_ _1418_/A _1418_/B _1418_/C _1426_/B vdd gnd NAND3X1
XFILL_1__1465_ vdd gnd FILL
XFILL_2__925_ vdd gnd FILL
XFILL_1__1396_ vdd gnd FILL
XFILL_2__1712_ vdd gnd FILL
XFILL_2__1643_ vdd gnd FILL
X_931_ _931_/A _994_/B vdd gnd INVX1
XFILL_2__1574_ vdd gnd FILL
XFILL100650x31350 vdd gnd FILL
XFILL100350x66450 vdd gnd FILL
XFILL_2__1008_ vdd gnd FILL
XFILL_0__1210_ vdd gnd FILL
XFILL_0__1141_ vdd gnd FILL
XFILL_0__1072_ vdd gnd FILL
XFILL_3__1821_ vdd gnd FILL
XFILL_3__1752_ vdd gnd FILL
XFILL_3__1683_ vdd gnd FILL
XFILL_1__943_ vdd gnd FILL
X_1203_ _1203_/A _1203_/B _1203_/C _1221_/B vdd gnd OAI21X1
X_1134_ _1142_/C _1142_/B _1142_/A _1154_/B vdd gnd AOI21X1
XFILL_0__1408_ vdd gnd FILL
X_1065_ _1065_/A _1159_/A _1206_/B vdd gnd NOR2X1
XFILL_3__1117_ vdd gnd FILL
XFILL_1__1181_ vdd gnd FILL
XFILL_1__1250_ vdd gnd FILL
XFILL_0__1339_ vdd gnd FILL
X_1898_ _1898_/D _1908_/CLK _1898_/Q vdd gnd DFFPOSX1
XFILL_3__1048_ vdd gnd FILL
XFILL_1__1517_ vdd gnd FILL
XFILL_2__1290_ vdd gnd FILL
XFILL_1__1448_ vdd gnd FILL
XFILL_1__1379_ vdd gnd FILL
XFILL_0__961_ vdd gnd FILL
XFILL_0__1690_ vdd gnd FILL
XFILL_2__1626_ vdd gnd FILL
XFILL100650x43050 vdd gnd FILL
XFILL_2__1557_ vdd gnd FILL
XFILL_2__1488_ vdd gnd FILL
X_1683_ _1688_/A _1733_/B _1708_/A _1695_/A vdd gnd NAND3X1
X_1821_ Yin[2] _1824_/B _1822_/C vdd gnd NAND2X1
X_1752_ _965_/A _1752_/B _1794_/C vdd gnd NOR2X1
XFILL_3_BUFX2_insert24 vdd gnd FILL
XFILL_0__1055_ vdd gnd FILL
XFILL_0__1124_ vdd gnd FILL
XFILL_3_BUFX2_insert13 vdd gnd FILL
XFILL_3__1735_ vdd gnd FILL
XFILL_3__1666_ vdd gnd FILL
XFILL_3__1804_ vdd gnd FILL
XFILL_3__1597_ vdd gnd FILL
XFILL_1__926_ vdd gnd FILL
X_1117_ _1127_/A _1123_/B vdd gnd INVX1
XFILL_1__1302_ vdd gnd FILL
XFILL_1__1233_ vdd gnd FILL
X_1048_ _1048_/A _1048_/B _1048_/C _1056_/C vdd gnd NAND3X1
XFILL_1__1164_ vdd gnd FILL
XFILL_1__1095_ vdd gnd FILL
XFILL_4__1844_ vdd gnd FILL
XFILL_4_CLKBUF1_insert5 vdd gnd FILL
XFILL_2__1411_ vdd gnd FILL
XFILL_2__1342_ vdd gnd FILL
XFILL_4__1209_ vdd gnd FILL
XFILL_2__1273_ vdd gnd FILL
XFILL_0__944_ vdd gnd FILL
XFILL_3__1520_ vdd gnd FILL
XFILL_0__1811_ vdd gnd FILL
XFILL_0__1742_ vdd gnd FILL
XFILL_2__1609_ vdd gnd FILL
XFILL_0__1673_ vdd gnd FILL
XFILL_3__1451_ vdd gnd FILL
XFILL_3__1382_ vdd gnd FILL
XFILL_4__922_ vdd gnd FILL
X_1735_ _1748_/B _1738_/C vdd gnd INVX1
X_1666_ _1711_/C _1666_/B _1666_/C _1670_/B vdd gnd AOI21X1
X_1804_ _1910_/D _1816_/A _923_/A _1815_/B vdd gnd NAND3X1
XFILL_0__1107_ vdd gnd FILL
XFILL_0__1038_ vdd gnd FILL
XFILL_3__1649_ vdd gnd FILL
XFILL_3__1718_ vdd gnd FILL
X_1597_ _1597_/A _1597_/B _1597_/C _1601_/C vdd gnd AOI21X1
XFILL_1__1782_ vdd gnd FILL
XFILL_1__1147_ vdd gnd FILL
XFILL_1__1216_ vdd gnd FILL
XFILL_4__1758_ vdd gnd FILL
XFILL_3__940_ vdd gnd FILL
XFILL_1__1078_ vdd gnd FILL
XFILL_4__1689_ vdd gnd FILL
XFILL_2__1256_ vdd gnd FILL
XFILL_2__1325_ vdd gnd FILL
XFILL_2__1187_ vdd gnd FILL
X_1520_ _1520_/A _1520_/B _1520_/C _1576_/A vdd gnd NAND3X1
XFILL_0__927_ vdd gnd FILL
XFILL_3__1503_ vdd gnd FILL
X_1451_ _1454_/A _1615_/B _1542_/A _1465_/B vdd gnd OAI21X1
XFILL_2_BUFX2_insert3 vdd gnd FILL
X_1382_ _1382_/A _1382_/B _1382_/C _1383_/B vdd gnd AOI21X1
XFILL_0__1587_ vdd gnd FILL
XFILL_0__1725_ vdd gnd FILL
XFILL_0__1656_ vdd gnd FILL
XFILL_3__1434_ vdd gnd FILL
XFILL_3__1365_ vdd gnd FILL
XFILL_3__1296_ vdd gnd FILL
XFILL_1__1001_ vdd gnd FILL
X_1649_ _1649_/A _1649_/B _1651_/A vdd gnd AND2X2
XFILL_4__1612_ vdd gnd FILL
X_1718_ _1718_/A _1749_/C _1728_/A vdd gnd XNOR2X1
XFILL_1__1834_ vdd gnd FILL
XFILL_1__1696_ vdd gnd FILL
XFILL_1__1765_ vdd gnd FILL
XFILL_4__1543_ vdd gnd FILL
XFILL_4__1474_ vdd gnd FILL
XFILL_2__1110_ vdd gnd FILL
XFILL_2__1041_ vdd gnd FILL
XFILL_3__923_ vdd gnd FILL
XFILL_0__1510_ vdd gnd FILL
XFILL_0__1441_ vdd gnd FILL
XFILL_3__1150_ vdd gnd FILL
XFILL_2__1308_ vdd gnd FILL
XFILL_2__1239_ vdd gnd FILL
XFILL_3__1081_ vdd gnd FILL
XFILL_0__1372_ vdd gnd FILL
X_1503_ _946_/A Cin[5] _956_/B Cin[6] _1579_/B vdd gnd AOI22X1
XFILL_0__1708_ vdd gnd FILL
XFILL_1__1550_ vdd gnd FILL
X_1434_ _952_/A Cin[2] _1510_/A _1437_/B vdd gnd NAND3X1
X_1365_ _1474_/A _1374_/B _1374_/A _1397_/A vdd gnd NAND3X1
X_1296_ _1396_/D _1389_/B vdd gnd INVX1
XFILL_0__1639_ vdd gnd FILL
XFILL_1__1481_ vdd gnd FILL
XFILL_3__1348_ vdd gnd FILL
XFILL_2__941_ vdd gnd FILL
XFILL_3__1417_ vdd gnd FILL
XFILL_3__1279_ vdd gnd FILL
XFILL_2__1590_ vdd gnd FILL
XFILL_1__1817_ vdd gnd FILL
XFILL_1__1679_ vdd gnd FILL
XFILL_1__1748_ vdd gnd FILL
XFILL_4__1388_ vdd gnd FILL
XFILL_2__1024_ vdd gnd FILL
XFILL_2__1788_ vdd gnd FILL
XFILL_0_CLKBUF1_insert10 vdd gnd FILL
X_1150_ _983_/A _1217_/B _1151_/B vdd gnd NAND2X1
XFILL_0__1355_ vdd gnd FILL
XFILL_0__1424_ vdd gnd FILL
XFILL_3__1202_ vdd gnd FILL
XFILL_3__1133_ vdd gnd FILL
X_1081_ _1140_/A _1101_/A vdd gnd INVX1
XFILL_0__1286_ vdd gnd FILL
XFILL_3__1064_ vdd gnd FILL
X_1417_ _1427_/A _1427_/B _1426_/C _1423_/C vdd gnd OAI21X1
XFILL_1__1602_ vdd gnd FILL
XFILL_1__1464_ vdd gnd FILL
XFILL_1__1533_ vdd gnd FILL
X_1348_ _1348_/A _1348_/B _1351_/A vdd gnd NAND2X1
XFILL_4__1242_ vdd gnd FILL
X_1279_ _1301_/B _1372_/C _1301_/A _1285_/A vdd gnd AOI21X1
XFILL_2__924_ vdd gnd FILL
XFILL_4__1173_ vdd gnd FILL
XFILL_1__1395_ vdd gnd FILL
X_930_ _945_/A _930_/B _930_/C _930_/Y vdd gnd OAI21X1
XFILL_2__1711_ vdd gnd FILL
XFILL_2__1573_ vdd gnd FILL
XFILL_2__1642_ vdd gnd FILL
XFILL100950x15750 vdd gnd FILL
XFILL_2__1007_ vdd gnd FILL
XFILL_0__1071_ vdd gnd FILL
XFILL_0__1140_ vdd gnd FILL
XFILL_3__1682_ vdd gnd FILL
XFILL_3__1820_ vdd gnd FILL
XFILL_3__1751_ vdd gnd FILL
XFILL_1__942_ vdd gnd FILL
X_1202_ _1277_/B _1277_/C _1277_/A _1278_/C vdd gnd NAND3X1
X_1133_ _1196_/B _1161_/C _1196_/A _1142_/C vdd gnd OAI21X1
X_1064_ _950_/B Cin[3] _1159_/A vdd gnd NAND2X1
XFILL_0__1407_ vdd gnd FILL
XFILL_0__1338_ vdd gnd FILL
XFILL_3__1047_ vdd gnd FILL
XFILL_1__1180_ vdd gnd FILL
XFILL_3__1116_ vdd gnd FILL
X_1897_ _1897_/D _1897_/CLK _1897_/Q vdd gnd DFFPOSX1
XFILL_0__1269_ vdd gnd FILL
XFILL_1__1516_ vdd gnd FILL
XFILL_1__1447_ vdd gnd FILL
XFILL_4__1087_ vdd gnd FILL
XFILL_1__1378_ vdd gnd FILL
XFILL_0__960_ vdd gnd FILL
XFILL100950x27450 vdd gnd FILL
XFILL_2__1625_ vdd gnd FILL
XFILL_2__1556_ vdd gnd FILL
X_1820_ _1820_/A _1824_/B _1820_/C _1891_/D vdd gnd OAI21X1
XFILL_2__1487_ vdd gnd FILL
X_1682_ _1682_/A _1709_/B _1682_/C _1733_/B vdd gnd NAND3X1
X_1751_ _963_/A _1752_/B _1751_/C _1754_/B vdd gnd OAI21X1
XFILL_3_BUFX2_insert25 vdd gnd FILL
XFILL_3__1803_ vdd gnd FILL
XFILL_3_BUFX2_insert14 vdd gnd FILL
XFILL_0__1054_ vdd gnd FILL
XFILL_0__1123_ vdd gnd FILL
XFILL_3__1734_ vdd gnd FILL
XFILL_3__1665_ vdd gnd FILL
XFILL_1__925_ vdd gnd FILL
XFILL_3__1596_ vdd gnd FILL
XFILL_1__1301_ vdd gnd FILL
X_1047_ _1068_/B _1050_/B _1049_/A _1048_/B vdd gnd OAI21X1
X_1116_ _947_/B Cin[4] _1127_/A vdd gnd NAND2X1
XFILL_1__1232_ vdd gnd FILL
XFILL_1__1094_ vdd gnd FILL
XFILL_1__1163_ vdd gnd FILL
XFILL_2__1410_ vdd gnd FILL
XFILL_2__1341_ vdd gnd FILL
XFILL_2__1272_ vdd gnd FILL
XFILL_0__943_ vdd gnd FILL
XFILL100950x39150 vdd gnd FILL
XFILL_0__1741_ vdd gnd FILL
XFILL_0__1810_ vdd gnd FILL
XFILL_3__1450_ vdd gnd FILL
XFILL_0__1672_ vdd gnd FILL
XFILL_2__1608_ vdd gnd FILL
XFILL_2__1539_ vdd gnd FILL
XFILL_3__1381_ vdd gnd FILL
X_1803_ _943_/A _1816_/A vdd gnd INVX1
X_1734_ _1748_/B _1736_/A _1748_/A _1741_/A vdd gnd NAND3X1
X_1665_ _1711_/A _1711_/B _1720_/A _1720_/B vdd gnd NOR3X1
X_1596_ _1611_/A _1596_/B _1597_/C vdd gnd AND2X2
XFILL_0__1037_ vdd gnd FILL
XFILL_0__1106_ vdd gnd FILL
XFILL_3__1648_ vdd gnd FILL
XFILL_3__1579_ vdd gnd FILL
XFILL_3__1717_ vdd gnd FILL
XFILL_1__1781_ vdd gnd FILL
XFILL_1__1215_ vdd gnd FILL
XFILL_1__1146_ vdd gnd FILL
XFILL_1__1077_ vdd gnd FILL
XFILL_4__1826_ vdd gnd FILL
XFILL_2__1324_ vdd gnd FILL
XFILL_0__926_ vdd gnd FILL
XFILL_2__1255_ vdd gnd FILL
XFILL_2__1186_ vdd gnd FILL
X_1450_ _1450_/A _1450_/B _1524_/A _1542_/A vdd gnd OAI21X1
XFILL_2_BUFX2_insert4 vdd gnd FILL
XFILL_0__1724_ vdd gnd FILL
XFILL_3__1502_ vdd gnd FILL
XFILL_3__1433_ vdd gnd FILL
XFILL_3__999_ vdd gnd FILL
X_1381_ _1381_/A _1381_/B _1381_/C _1394_/A vdd gnd OAI21X1
XFILL_0__1586_ vdd gnd FILL
XFILL_0__1655_ vdd gnd FILL
XFILL_3__1364_ vdd gnd FILL
XFILL_3__1295_ vdd gnd FILL
XFILL_1__1000_ vdd gnd FILL
X_1648_ _1694_/C _1695_/C vdd gnd INVX1
X_1579_ _1579_/A _1579_/B _1579_/C _1602_/A vdd gnd OAI21X1
X_1717_ _1717_/A _1749_/D _1718_/A vdd gnd NOR2X1
XFILL_1__1833_ vdd gnd FILL
XFILL_1__1695_ vdd gnd FILL
XFILL_1__1764_ vdd gnd FILL
XFILL_2__1040_ vdd gnd FILL
XFILL_1__1129_ vdd gnd FILL
XFILL_3__922_ vdd gnd FILL
XFILL_0__1440_ vdd gnd FILL
XFILL_2__1307_ vdd gnd FILL
XFILL_3__1080_ vdd gnd FILL
XFILL_0__1371_ vdd gnd FILL
XFILL_2__1238_ vdd gnd FILL
XFILL_2__1169_ vdd gnd FILL
X_1502_ _1502_/A _1584_/A _1514_/B vdd gnd NOR2X1
X_1433_ _949_/A Cin[3] _1510_/A vdd gnd NAND2X1
XFILL99450x15750 vdd gnd FILL
XFILL_0__1707_ vdd gnd FILL
XFILL_1__1480_ vdd gnd FILL
XFILL_3__1416_ vdd gnd FILL
X_1364_ _1368_/A _1368_/B _1473_/C _1374_/B vdd gnd OAI21X1
X_1295_ _1395_/B _1389_/A vdd gnd INVX1
XFILL_0__1638_ vdd gnd FILL
XFILL_0__1569_ vdd gnd FILL
XFILL_3__1347_ vdd gnd FILL
XFILL_2__940_ vdd gnd FILL
XFILL_3__1278_ vdd gnd FILL
XFILL_4__1525_ vdd gnd FILL
XFILL_1__1747_ vdd gnd FILL
XFILL_1__1816_ vdd gnd FILL
XFILL101250x50850 vdd gnd FILL
XFILL_1__1678_ vdd gnd FILL
XFILL_4__1456_ vdd gnd FILL
XFILL_2__1023_ vdd gnd FILL
XFILL_2__1787_ vdd gnd FILL
XFILL_0_CLKBUF1_insert11 vdd gnd FILL
X_1080_ _1101_/B _1140_/C _1140_/A _1093_/C vdd gnd OAI21X1
XFILL_0__1423_ vdd gnd FILL
XFILL_0__1354_ vdd gnd FILL
XFILL_3__1201_ vdd gnd FILL
XFILL_3__1132_ vdd gnd FILL
XFILL_3__1063_ vdd gnd FILL
XFILL_0__1285_ vdd gnd FILL
XFILL_1__1601_ vdd gnd FILL
X_1347_ _955_/A _1449_/B _1897_/Q _1524_/A vdd gnd NAND3X1
X_1416_ _1416_/A _1416_/B _1416_/C _1426_/C vdd gnd OAI21X1
XFILL_1__1532_ vdd gnd FILL
XFILL_1__1463_ vdd gnd FILL
XFILL_4__1310_ vdd gnd FILL
X_1278_ _1278_/A _1278_/B _1278_/C _1382_/C vdd gnd OAI21X1
XFILL_1__1394_ vdd gnd FILL
XFILL_2__923_ vdd gnd FILL
XFILL_2__1710_ vdd gnd FILL
XFILL_4__1439_ vdd gnd FILL
XFILL_2__1572_ vdd gnd FILL
XFILL_2__1641_ vdd gnd FILL
XFILL_2__1006_ vdd gnd FILL
XFILL_0__1070_ vdd gnd FILL
XFILL_3__1681_ vdd gnd FILL
XFILL_3__1750_ vdd gnd FILL
XFILL_1__941_ vdd gnd FILL
XFILL_2__1839_ vdd gnd FILL
X_1201_ _1278_/A _1221_/A vdd gnd INVX1
X_989_ _989_/A _990_/A _990_/C vdd gnd NAND2X1
X_1132_ _1159_/C _1132_/B _1196_/A vdd gnd NAND2X1
X_1063_ _1065_/A _1063_/B _1093_/B _1092_/A vdd gnd OAI21X1
XFILL_0__1337_ vdd gnd FILL
XFILL_0__1406_ vdd gnd FILL
XFILL_3__1115_ vdd gnd FILL
XFILL_0__1268_ vdd gnd FILL
XFILL_3__1046_ vdd gnd FILL
XFILL_4__1790_ vdd gnd FILL
X_1896_ _1896_/D _1910_/CLK _1896_/Q vdd gnd DFFPOSX1
XFILL_0__1199_ vdd gnd FILL
XFILL_1__1515_ vdd gnd FILL
XFILL_1__1446_ vdd gnd FILL
XFILL_4__1155_ vdd gnd FILL
XFILL_4__1224_ vdd gnd FILL
XFILL_1__1377_ vdd gnd FILL
XFILL101250x74250 vdd gnd FILL
XFILL_2__1624_ vdd gnd FILL
XFILL_2__1555_ vdd gnd FILL
XFILL_2__1486_ vdd gnd FILL
XFILL100650x150 vdd gnd FILL
X_1750_ Cin[7] _1752_/B vdd gnd INVX1
XFILL_0__1122_ vdd gnd FILL
X_1681_ _1681_/A _1682_/C vdd gnd INVX1
XFILL_3_BUFX2_insert15 vdd gnd FILL
XFILL_3__1802_ vdd gnd FILL
XFILL_0__1053_ vdd gnd FILL
XFILL_3__1733_ vdd gnd FILL
XFILL_3__1664_ vdd gnd FILL
XFILL_3__1595_ vdd gnd FILL
XFILL_1__924_ vdd gnd FILL
X_1115_ _1130_/C _1130_/B _1130_/A _1196_/C vdd gnd NAND3X1
XFILL_1__1231_ vdd gnd FILL
XFILL_1__1300_ vdd gnd FILL
X_1046_ _1068_/A _1049_/A vdd gnd INVX1
X_1879_ _1879_/D _1880_/CLK _993_/B vdd gnd DFFPOSX1
XFILL_4__997_ vdd gnd FILL
XFILL_3__1029_ vdd gnd FILL
XFILL_4__1911_ vdd gnd FILL
XFILL_1__1093_ vdd gnd FILL
XFILL_1__1162_ vdd gnd FILL
XFILL_4__1773_ vdd gnd FILL
XFILL_2__1340_ vdd gnd FILL
XFILL_1__1429_ vdd gnd FILL
XFILL_0__942_ vdd gnd FILL
XFILL_2__1271_ vdd gnd FILL
XFILL_4__1069_ vdd gnd FILL
XFILL_0__1740_ vdd gnd FILL
XFILL_0__1671_ vdd gnd FILL
XFILL_2__1607_ vdd gnd FILL
XFILL_2__1538_ vdd gnd FILL
XFILL_2__1469_ vdd gnd FILL
XFILL_3__1380_ vdd gnd FILL
X_1733_ _1733_/A _1733_/B _1733_/C _1748_/A vdd gnd NAND3X1
X_1802_ Yin[0] _1827_/A vdd gnd INVX1
XFILL_0__1105_ vdd gnd FILL
X_1664_ _1670_/C _1671_/B vdd gnd INVX1
X_1595_ _1652_/B _1595_/B _1652_/A _1600_/B vdd gnd OAI21X1
XFILL_1__1780_ vdd gnd FILL
XFILL_3__1716_ vdd gnd FILL
XFILL_0__1036_ vdd gnd FILL
XFILL_3__1578_ vdd gnd FILL
XFILL_3__1647_ vdd gnd FILL
X_1029_ _1029_/A _1029_/B _1030_/A vdd gnd NAND2X1
XFILL_1__1214_ vdd gnd FILL
XFILL_1__1076_ vdd gnd FILL
XFILL_1__1145_ vdd gnd FILL
XFILL_2__1323_ vdd gnd FILL
XFILL_0__925_ vdd gnd FILL
XFILL_2__1185_ vdd gnd FILL
XFILL_2__1254_ vdd gnd FILL
X_1380_ _1484_/B _1483_/A _1484_/A _1381_/A vdd gnd AOI21X1
XFILL_0__1654_ vdd gnd FILL
XFILL_3__1501_ vdd gnd FILL
XFILL_0__1723_ vdd gnd FILL
XFILL_3__1432_ vdd gnd FILL
XFILL_3__998_ vdd gnd FILL
XFILL_3__1363_ vdd gnd FILL
XFILL_0__1585_ vdd gnd FILL
XFILL_3__1294_ vdd gnd FILL
X_1716_ _1749_/A _1751_/C _1717_/A vdd gnd NOR2X1
X_1578_ _1578_/A _1578_/B _1578_/C _1631_/C vdd gnd AOI21X1
X_1647_ _1647_/A _1649_/B _1694_/C vdd gnd NAND2X1
XFILL_1__1763_ vdd gnd FILL
XFILL_1__1832_ vdd gnd FILL
XFILL_0__1019_ vdd gnd FILL
XFILL_1__1694_ vdd gnd FILL
XFILL_1__1128_ vdd gnd FILL
XFILL_4__1808_ vdd gnd FILL
XFILL100350x4050 vdd gnd FILL
XFILL_1__1059_ vdd gnd FILL
XFILL_2__1306_ vdd gnd FILL
XFILL_2__1237_ vdd gnd FILL
XFILL_0__1370_ vdd gnd FILL
XFILL_2__1099_ vdd gnd FILL
XFILL_2__1168_ vdd gnd FILL
X_1501_ _946_/A Cin[6] _1584_/A vdd gnd NAND2X1
X_1432_ _946_/A Cin[4] _1511_/A vdd gnd NAND2X1
X_1363_ _1363_/A _1363_/B _1461_/A _1368_/A vdd gnd AOI21X1
XFILL_0__1637_ vdd gnd FILL
XFILL_0__1706_ vdd gnd FILL
XFILL_3__1346_ vdd gnd FILL
XFILL_3__1415_ vdd gnd FILL
X_1294_ _983_/A _987_/B _1294_/C _1294_/D _1876_/D vdd gnd OAI22X1
XFILL_0__1568_ vdd gnd FILL
XFILL_0__1499_ vdd gnd FILL
XFILL_3__1277_ vdd gnd FILL
XFILL_1__1746_ vdd gnd FILL
XFILL_1__1815_ vdd gnd FILL
XFILL_1__1677_ vdd gnd FILL
XFILL_2__999_ vdd gnd FILL
XFILL_2__1022_ vdd gnd FILL
XFILL_2__1786_ vdd gnd FILL
XFILL_3__1200_ vdd gnd FILL
XFILL_0__1353_ vdd gnd FILL
XFILL_0__1422_ vdd gnd FILL
XFILL_3__1131_ vdd gnd FILL
XFILL_0__1284_ vdd gnd FILL
XFILL_3__1062_ vdd gnd FILL
XFILL_1__1600_ vdd gnd FILL
XFILL_1__1531_ vdd gnd FILL
X_1346_ _1450_/A _1351_/C vdd gnd INVX1
X_1415_ _1420_/A _1420_/B _1416_/B vdd gnd AND2X2
XFILL_1__1462_ vdd gnd FILL
XFILL_1__1393_ vdd gnd FILL
XFILL_2__922_ vdd gnd FILL
XFILL_3__1329_ vdd gnd FILL
X_1277_ _1277_/A _1277_/B _1277_/C _1278_/B vdd gnd AOI21X1
XFILL_2__1640_ vdd gnd FILL
XFILL_1__1729_ vdd gnd FILL
XFILL_4__1507_ vdd gnd FILL
XFILL_2__1571_ vdd gnd FILL
XFILL_2__1005_ vdd gnd FILL
XFILL_3__1680_ vdd gnd FILL
XFILL_2__1769_ vdd gnd FILL
XFILL_1__940_ vdd gnd FILL
X_988_ _988_/A _990_/B vdd gnd INVX1
XFILL_2__1838_ vdd gnd FILL
X_1200_ _1278_/A _1208_/B _1208_/A _1205_/A vdd gnd NAND3X1
XFILL_0__1405_ vdd gnd FILL
X_1131_ _1131_/A _1131_/B _1131_/C _1161_/C vdd gnd AOI21X1
X_1062_ _1062_/A _1062_/B _1062_/C _1063_/B vdd gnd AOI21X1
XFILL_0__1336_ vdd gnd FILL
X_1895_ _1895_/D _1910_/CLK _1895_/Q vdd gnd DFFPOSX1
XFILL_3__1114_ vdd gnd FILL
XFILL_0__1267_ vdd gnd FILL
XFILL_3__1045_ vdd gnd FILL
XFILL_0__1198_ vdd gnd FILL
XFILL_1__1514_ vdd gnd FILL
X_1329_ _949_/A Cin[2] _1420_/B vdd gnd NAND2X1
XFILL_1__1445_ vdd gnd FILL
XFILL_1__1376_ vdd gnd FILL
XFILL_2__1623_ vdd gnd FILL
XFILL_2__1554_ vdd gnd FILL
XFILL_2__1485_ vdd gnd FILL
XFILL_0__1121_ vdd gnd FILL
XFILL_0__1052_ vdd gnd FILL
X_1680_ _1680_/A _1709_/A _1680_/C _1709_/B vdd gnd NAND3X1
XFILL_3__1732_ vdd gnd FILL
XFILL_3__1801_ vdd gnd FILL
XFILL_3_BUFX2_insert16 vdd gnd FILL
XFILL_3__1594_ vdd gnd FILL
XFILL_3__1663_ vdd gnd FILL
XFILL_1__923_ vdd gnd FILL
X_1114_ _1173_/B _1114_/B _1173_/A _1130_/A vdd gnd OAI21X1
XFILL_1__1161_ vdd gnd FILL
XFILL_1__1230_ vdd gnd FILL
X_1045_ _950_/B Cin[1] _1068_/A vdd gnd NAND2X1
X_1878_ _1878_/D _1880_/CLK _991_/B vdd gnd DFFPOSX1
XFILL_0__1319_ vdd gnd FILL
XFILL_3__1028_ vdd gnd FILL
XFILL_1__1092_ vdd gnd FILL
XFILL_4__1841_ vdd gnd FILL
XFILL_4_CLKBUF1_insert8 vdd gnd FILL
XFILL_4__1206_ vdd gnd FILL
XFILL_2__1270_ vdd gnd FILL
XFILL_0__941_ vdd gnd FILL
XFILL_1__1428_ vdd gnd FILL
XFILL_1__1359_ vdd gnd FILL
XFILL_4__1137_ vdd gnd FILL
XFILL_0__1670_ vdd gnd FILL
XFILL_2__1606_ vdd gnd FILL
XFILL_2__1537_ vdd gnd FILL
XFILL_2__1468_ vdd gnd FILL
XFILL_2__1399_ vdd gnd FILL
X_1663_ _1670_/C _1671_/A _1671_/C _1709_/A vdd gnd NAND3X1
X_1732_ _1759_/C _1732_/B _1733_/C vdd gnd NAND2X1
X_1801_ _1801_/A _1801_/B _1801_/C _1801_/D _1885_/D vdd gnd AOI22X1
XFILL_0__1035_ vdd gnd FILL
XFILL_0__1104_ vdd gnd FILL
X_1594_ _1594_/A _1594_/B _1652_/C _1600_/A vdd gnd NAND3X1
XFILL_3__1715_ vdd gnd FILL
XFILL_3__1577_ vdd gnd FILL
XFILL_3__1646_ vdd gnd FILL
XFILL_0__1799_ vdd gnd FILL
XFILL_4__979_ vdd gnd FILL
X_1028_ _1029_/B _1029_/A _1034_/A vdd gnd OR2X2
XFILL_1__1213_ vdd gnd FILL
XFILL_1__1144_ vdd gnd FILL
XFILL_4__1755_ vdd gnd FILL
XFILL_1__1075_ vdd gnd FILL
XFILL_4__1686_ vdd gnd FILL
XFILL_2__1322_ vdd gnd FILL
XFILL_2__1253_ vdd gnd FILL
XFILL_0__924_ vdd gnd FILL
XFILL_2__1184_ vdd gnd FILL
XFILL_3__1500_ vdd gnd FILL
XFILL_3__997_ vdd gnd FILL
XFILL_0__1653_ vdd gnd FILL
XFILL_0__1584_ vdd gnd FILL
XFILL_0__1722_ vdd gnd FILL
XFILL_3__1431_ vdd gnd FILL
XFILL_3__1362_ vdd gnd FILL
XFILL_3__1293_ vdd gnd FILL
X_1646_ _1646_/A _1646_/B _1692_/A _1691_/B vdd gnd OAI21X1
X_1715_ _955_/A Cin[6] _1751_/C vdd gnd NAND2X1
XFILL_0__1018_ vdd gnd FILL
XFILL_3__1629_ vdd gnd FILL
X_1577_ _1693_/A _1646_/A vdd gnd INVX1
XFILL_1__1693_ vdd gnd FILL
XFILL_1__1762_ vdd gnd FILL
XFILL_4__1540_ vdd gnd FILL
XFILL_4__1471_ vdd gnd FILL
XFILL_1__1831_ vdd gnd FILL
XFILL_1__1127_ vdd gnd FILL
XFILL_1__1058_ vdd gnd FILL
XFILL_2__1305_ vdd gnd FILL
XFILL_2__1236_ vdd gnd FILL
XFILL_2__1167_ vdd gnd FILL
X_1500_ _953_/B Cin[7] _1579_/A vdd gnd NAND2X1
XFILL100350x74250 vdd gnd FILL
XFILL_2__1098_ vdd gnd FILL
X_1431_ _1431_/A _1431_/B _1431_/C _1470_/C vdd gnd AOI21X1
X_1362_ _1461_/C _1431_/B _1431_/A _1368_/B vdd gnd AOI21X1
X_1293_ _983_/A _1396_/D _1294_/D vdd gnd NAND2X1
XFILL_0__1636_ vdd gnd FILL
XFILL_0__1705_ vdd gnd FILL
XFILL_0__1567_ vdd gnd FILL
XFILL_3__1345_ vdd gnd FILL
XFILL_3__1414_ vdd gnd FILL
XFILL_3__1276_ vdd gnd FILL
XFILL_0__1498_ vdd gnd FILL
X_1629_ _1646_/A _1637_/B _1637_/A _1633_/A vdd gnd NAND3X1
XFILL_1__1676_ vdd gnd FILL
XFILL_4__1454_ vdd gnd FILL
XFILL_1__1745_ vdd gnd FILL
XFILL_1__1814_ vdd gnd FILL
XFILL_4__1385_ vdd gnd FILL
XFILL_2__1021_ vdd gnd FILL
XFILL_2__998_ vdd gnd FILL
XFILL_2__1785_ vdd gnd FILL
XFILL_0__1421_ vdd gnd FILL
XFILL_3__1130_ vdd gnd FILL
XFILL_0__1352_ vdd gnd FILL
XFILL_3__1061_ vdd gnd FILL
XFILL_0__1283_ vdd gnd FILL
XFILL_2__1219_ vdd gnd FILL
XFILL_1__1530_ vdd gnd FILL
X_1345_ _1450_/A _1352_/B _1352_/A _1460_/A vdd gnd NAND3X1
X_1414_ _1418_/B _1418_/C _1418_/A _1427_/B vdd gnd AOI21X1
X_1276_ _1382_/A _1382_/B _1285_/C _1289_/A vdd gnd NAND3X1
XFILL_0__1619_ vdd gnd FILL
XFILL_1__1461_ vdd gnd FILL
XFILL_3__1328_ vdd gnd FILL
XFILL_1__1392_ vdd gnd FILL
XFILL_4__1170_ vdd gnd FILL
XFILL_3__1259_ vdd gnd FILL
XFILL_1__1659_ vdd gnd FILL
XFILL_1__1728_ vdd gnd FILL
XFILL_2__1570_ vdd gnd FILL
XFILL_2__1004_ vdd gnd FILL
XFILL_2__1768_ vdd gnd FILL
XFILL_2__1699_ vdd gnd FILL
X_987_ _990_/A _987_/B _987_/C _987_/Y vdd gnd OAI21X1
XFILL_2__1837_ vdd gnd FILL
X_1130_ _1130_/A _1130_/B _1130_/C _1196_/B vdd gnd AOI21X1
XFILL_0__1404_ vdd gnd FILL
XFILL_0__1335_ vdd gnd FILL
X_1061_ _976_/B _1216_/A _1098_/C vdd gnd NAND2X1
XFILL_3__1113_ vdd gnd FILL
X_1894_ _1894_/D _1908_/CLK _1894_/Q vdd gnd DFFPOSX1
XFILL_0__1266_ vdd gnd FILL
XFILL_0__1197_ vdd gnd FILL
XFILL_3__1044_ vdd gnd FILL
XFILL_1__1513_ vdd gnd FILL
XFILL_1__1444_ vdd gnd FILL
XFILL_1__999_ vdd gnd FILL
X_1328_ _949_/A Cin[2] _1420_/A _1331_/B vdd gnd NAND3X1
X_1259_ _1263_/A _1263_/B _1360_/C _1269_/A vdd gnd OAI21X1
XFILL_1__1375_ vdd gnd FILL
XFILL_4__1084_ vdd gnd FILL
XFILL_2__1553_ vdd gnd FILL
XFILL_2__1622_ vdd gnd FILL
XFILL_2__1484_ vdd gnd FILL
XFILL_3_BUFX2_insert17 vdd gnd FILL
XFILL_0__1051_ vdd gnd FILL
XFILL_0__1120_ vdd gnd FILL
XFILL_3__1731_ vdd gnd FILL
XFILL_3__1662_ vdd gnd FILL
XFILL_3__1800_ vdd gnd FILL
XFILL_1__922_ vdd gnd FILL
XFILL_3__1593_ vdd gnd FILL
X_1113_ _1173_/C _1113_/B _1113_/C _1130_/B vdd gnd NAND3X1
X_1044_ _1845_/B _1044_/B _1049_/B _1048_/C vdd gnd OAI21X1
XFILL_0__1318_ vdd gnd FILL
XFILL_1__1160_ vdd gnd FILL
XFILL_1__1091_ vdd gnd FILL
X_1877_ _1877_/D _1904_/CLK _988_/A vdd gnd DFFPOSX1
XFILL_3__1027_ vdd gnd FILL
XFILL_0__1249_ vdd gnd FILL
XFILL_1__1427_ vdd gnd FILL
XFILL_1__1358_ vdd gnd FILL
XFILL_0__940_ vdd gnd FILL
XFILL_1__1289_ vdd gnd FILL
XFILL_2__1536_ vdd gnd FILL
XFILL_2__1605_ vdd gnd FILL
XFILL_2__1467_ vdd gnd FILL
X_1800_ _1800_/A _998_/A _1801_/C vdd gnd AND2X2
XFILL_2__1398_ vdd gnd FILL
X_1731_ _1759_/C _1731_/B _1732_/B _1736_/A vdd gnd NAND3X1
X_1662_ _1711_/B _1720_/A _1711_/A _1671_/A vdd gnd OAI21X1
XFILL_0__1103_ vdd gnd FILL
XFILL_0__1034_ vdd gnd FILL
XFILL_3__1645_ vdd gnd FILL
X_1593_ _1601_/A _1601_/B _1600_/C _1599_/C vdd gnd OAI21X1
XFILL_3__1714_ vdd gnd FILL
XFILL_3__1576_ vdd gnd FILL
XFILL_0__1798_ vdd gnd FILL
X_1027_ _1027_/A _1027_/B _1029_/B vdd gnd NAND2X1
XFILL_1__1212_ vdd gnd FILL
XFILL_1__1143_ vdd gnd FILL
XFILL_1__1074_ vdd gnd FILL
XFILL_4__1823_ vdd gnd FILL
XFILL_2__1321_ vdd gnd FILL
XFILL_2__1183_ vdd gnd FILL
XFILL100950x11850 vdd gnd FILL
XFILL_2__1252_ vdd gnd FILL
XFILL100650x46950 vdd gnd FILL
XFILL_0__923_ vdd gnd FILL
XFILL_0__1721_ vdd gnd FILL
XFILL_3__996_ vdd gnd FILL
XFILL_0__1652_ vdd gnd FILL
XFILL_0__1583_ vdd gnd FILL
XFILL_2__1519_ vdd gnd FILL
XFILL_3__1430_ vdd gnd FILL
XFILL_3__1361_ vdd gnd FILL
XFILL_3__1292_ vdd gnd FILL
X_1645_ _1645_/A _1645_/B _1645_/C _1646_/B vdd gnd AOI21X1
X_1576_ _1576_/A _1576_/B _1693_/A vdd gnd NAND2X1
X_1714_ _952_/A Cin[5] _1749_/A vdd gnd NAND2X1
XFILL_1__1830_ vdd gnd FILL
XFILL_0__1017_ vdd gnd FILL
XFILL_3__1628_ vdd gnd FILL
XFILL_1__1692_ vdd gnd FILL
XFILL_3__1559_ vdd gnd FILL
XFILL_1__1761_ vdd gnd FILL
XFILL_0__1919_ vdd gnd FILL
XFILL_1__1126_ vdd gnd FILL
XFILL_1__1057_ vdd gnd FILL
XFILL_4__1668_ vdd gnd FILL
XFILL_4__1737_ vdd gnd FILL
XFILL_2__1304_ vdd gnd FILL
XFILL100950x23550 vdd gnd FILL
XFILL100650x58650 vdd gnd FILL
XFILL_2__1235_ vdd gnd FILL
XFILL_2__1166_ vdd gnd FILL
X_1430_ _1461_/C _1431_/C vdd gnd INVX1
XFILL_2__1097_ vdd gnd FILL
XFILL_0__1704_ vdd gnd FILL
XFILL_3__1413_ vdd gnd FILL
XFILL_3__979_ vdd gnd FILL
X_1361_ _1361_/A _1361_/B _1361_/C _1473_/C vdd gnd OAI21X1
X_1292_ _1395_/B _1292_/B _1292_/C _1396_/D vdd gnd NAND3X1
XFILL_3__1275_ vdd gnd FILL
XFILL_0__1635_ vdd gnd FILL
XFILL_0__1566_ vdd gnd FILL
XFILL_0__1497_ vdd gnd FILL
XFILL_3__1344_ vdd gnd FILL
X_1628_ _1685_/B _1631_/B _1645_/C _1637_/B vdd gnd OAI21X1
X_1559_ _1574_/C _1574_/B _1574_/A _1575_/C vdd gnd NAND3X1
XFILL_4__1522_ vdd gnd FILL
XFILL_1__1813_ vdd gnd FILL
XFILL_1__1675_ vdd gnd FILL
XFILL_1__1744_ vdd gnd FILL
XFILL_2__997_ vdd gnd FILL
XFILL_2__1020_ vdd gnd FILL
XFILL_1__1109_ vdd gnd FILL
XFILL_2__1784_ vdd gnd FILL
XFILL100950x35250 vdd gnd FILL
XFILL_0__1351_ vdd gnd FILL
XFILL_0__1420_ vdd gnd FILL
XFILL_3__1060_ vdd gnd FILL
XFILL_0__1282_ vdd gnd FILL
XFILL_2__1218_ vdd gnd FILL
XFILL_2__1149_ vdd gnd FILL
X_1413_ _1849_/B _1413_/B _1413_/C _1418_/C vdd gnd OAI21X1
X_1275_ _1301_/A _1372_/C _1301_/B _1382_/B vdd gnd NAND3X1
X_1344_ _1897_/Q _1348_/B _1352_/B vdd gnd NAND2X1
XFILL_1__1460_ vdd gnd FILL
XFILL_0__1618_ vdd gnd FILL
XFILL_0__1549_ vdd gnd FILL
XFILL_3__1327_ vdd gnd FILL
XFILL_3__1258_ vdd gnd FILL
XFILL_1__1391_ vdd gnd FILL
XFILL_3__1189_ vdd gnd FILL
XFILL_1__1727_ vdd gnd FILL
XFILL_1__1589_ vdd gnd FILL
XFILL_1__1658_ vdd gnd FILL
XFILL_4__1436_ vdd gnd FILL
XFILL_4__1367_ vdd gnd FILL
XFILL_4__1298_ vdd gnd FILL
XFILL_2__1003_ vdd gnd FILL
XFILL_2__1836_ vdd gnd FILL
XFILL_2__1767_ vdd gnd FILL
XFILL_2__1698_ vdd gnd FILL
X_986_ _986_/A _990_/A _987_/C vdd gnd NAND2X1
X_1060_ _1060_/A _1060_/B _1060_/C _1872_/D vdd gnd OAI21X1
XFILL_0__1334_ vdd gnd FILL
XFILL_0__1403_ vdd gnd FILL
XFILL_3__1112_ vdd gnd FILL
XFILL_3__1043_ vdd gnd FILL
X_1893_ _1893_/D _1897_/CLK _1893_/Q vdd gnd DFFPOSX1
XFILL_0__1196_ vdd gnd FILL
XFILL_0__1265_ vdd gnd FILL
XFILL_1__1512_ vdd gnd FILL
XFILL_1__1443_ vdd gnd FILL
XFILL_1__998_ vdd gnd FILL
X_1327_ _946_/A Cin[3] _1420_/A vdd gnd NAND2X1
X_1258_ _1258_/A _1258_/B _1338_/A _1263_/B vdd gnd AOI21X1
XFILL_4__1221_ vdd gnd FILL
X_1189_ _1193_/A _1193_/B _1266_/C _1198_/A vdd gnd OAI21X1
XFILL_4__1152_ vdd gnd FILL
XFILL_1__1374_ vdd gnd FILL
XFILL_2__1483_ vdd gnd FILL
XFILL_2__1621_ vdd gnd FILL
XFILL_2__1552_ vdd gnd FILL
XFILL100950x4050 vdd gnd FILL
XFILL_3_BUFX2_insert18 vdd gnd FILL
XFILL_0__1050_ vdd gnd FILL
XFILL_3__1730_ vdd gnd FILL
XFILL_3__1661_ vdd gnd FILL
XFILL_3__1592_ vdd gnd FILL
XFILL_2__1819_ vdd gnd FILL
X_969_ _969_/A _971_/B vdd gnd INVX1
X_1112_ _1131_/A _1131_/B _1131_/C _1161_/B vdd gnd NAND3X1
X_1043_ _1068_/B _1050_/B _1049_/B vdd gnd NOR2X1
XFILL_4__994_ vdd gnd FILL
XFILL_0__1248_ vdd gnd FILL
XFILL_0__1317_ vdd gnd FILL
XFILL_3__1026_ vdd gnd FILL
XFILL_1__1090_ vdd gnd FILL
XFILL_4__1770_ vdd gnd FILL
X_1876_ _1876_/D _1904_/CLK _985_/A vdd gnd DFFPOSX1
XFILL_0__1179_ vdd gnd FILL
XFILL_1__1357_ vdd gnd FILL
XFILL_1__1426_ vdd gnd FILL
XFILL_1__1288_ vdd gnd FILL
XFILL_4__1066_ vdd gnd FILL
XFILL_2__1535_ vdd gnd FILL
XFILL_2__1604_ vdd gnd FILL
XFILL_2__1466_ vdd gnd FILL
XFILL_0__1102_ vdd gnd FILL
XFILL_2__1397_ vdd gnd FILL
X_1730_ _1762_/C _1730_/B _1730_/C _1759_/C vdd gnd NAND3X1
X_1661_ _1661_/A _1661_/B _1720_/A vdd gnd NOR2X1
X_1592_ _1592_/A _1592_/B _1592_/C _1600_/C vdd gnd OAI21X1
XFILL_0__999_ vdd gnd FILL
XFILL_0__1033_ vdd gnd FILL
XFILL_3__1575_ vdd gnd FILL
XFILL_3__1713_ vdd gnd FILL
XFILL_3__1644_ vdd gnd FILL
XFILL_0__1797_ vdd gnd FILL
X_1026_ _1036_/C _1026_/B _1026_/C _1027_/A vdd gnd NAND3X1
XFILL_1__1211_ vdd gnd FILL
XFILL_3__1009_ vdd gnd FILL
X_1859_ _983_/Y _1904_/CLK _981_/A vdd gnd DFFPOSX1
XFILL_1__1142_ vdd gnd FILL
XFILL_1__1073_ vdd gnd FILL
XFILL_2__1320_ vdd gnd FILL
XFILL_1__1409_ vdd gnd FILL
XFILL_0__922_ vdd gnd FILL
XFILL_2__1182_ vdd gnd FILL
XFILL_2__1251_ vdd gnd FILL
XFILL_0__1651_ vdd gnd FILL
XFILL_0__1720_ vdd gnd FILL
XFILL_3__995_ vdd gnd FILL
XFILL_0__1582_ vdd gnd FILL
XFILL_2__1518_ vdd gnd FILL
XFILL_2__1449_ vdd gnd FILL
XFILL_3__1360_ vdd gnd FILL
XFILL_3__1291_ vdd gnd FILL
X_1713_ _955_/A Cin[5] _1794_/B _1749_/D vdd gnd AOI21X1
X_1575_ _1575_/A _1575_/B _1575_/C _1633_/C vdd gnd OAI21X1
XFILL_1__1760_ vdd gnd FILL
X_1644_ _1703_/B _1644_/B _1705_/B _1699_/B vdd gnd OAI21X1
XFILL_0__1016_ vdd gnd FILL
XFILL_3__1627_ vdd gnd FILL
XFILL_1__1691_ vdd gnd FILL
XFILL_3__1558_ vdd gnd FILL
XFILL_0__1918_ vdd gnd FILL
XFILL_0__1849_ vdd gnd FILL
XFILL_3__1489_ vdd gnd FILL
X_1009_ _943_/B _1801_/A _1010_/C vdd gnd NAND2X1
XFILL_4__1805_ vdd gnd FILL
XFILL_1__1125_ vdd gnd FILL
XFILL_1__1056_ vdd gnd FILL
XFILL101250x70350 vdd gnd FILL
XFILL_2__1303_ vdd gnd FILL
XFILL_2__1234_ vdd gnd FILL
XFILL_2__1096_ vdd gnd FILL
XFILL_2__1165_ vdd gnd FILL
X_1360_ _1360_/A _1360_/B _1360_/C _1361_/B vdd gnd AOI21X1
XFILL_0__1634_ vdd gnd FILL
XFILL_0__1703_ vdd gnd FILL
XFILL_3__1343_ vdd gnd FILL
XFILL_3__1412_ vdd gnd FILL
XFILL_3__978_ vdd gnd FILL
X_1291_ _1292_/C _1395_/B _1292_/B _1294_/C vdd gnd AOI21X1
XFILL_0__1496_ vdd gnd FILL
XFILL_0__1565_ vdd gnd FILL
XFILL_3__1274_ vdd gnd FILL
X_1627_ _1687_/A _1687_/B _1685_/B vdd gnd NOR2X1
XFILL_1__1743_ vdd gnd FILL
X_1558_ _1564_/A _1564_/B _1575_/A _1562_/A vdd gnd AOI21X1
X_1489_ _1704_/C _1572_/B _1490_/B vdd gnd XOR2X1
XFILL_1__1812_ vdd gnd FILL
XFILL_2_BUFX2_insert20 vdd gnd FILL
XFILL_1__1674_ vdd gnd FILL
XFILL_2__996_ vdd gnd FILL
XFILL_1__1108_ vdd gnd FILL
XFILL101250x82050 vdd gnd FILL
XFILL_1__1039_ vdd gnd FILL
XFILL_4__1719_ vdd gnd FILL
XFILL_2__1783_ vdd gnd FILL
XFILL_0__1350_ vdd gnd FILL
XFILL_0__1281_ vdd gnd FILL
XFILL_2__1217_ vdd gnd FILL
XFILL_2__1079_ vdd gnd FILL
XFILL_2__1148_ vdd gnd FILL
X_1343_ _955_/A _1449_/B _1348_/B vdd gnd NAND2X1
X_1412_ _1847_/B _1778_/B _1507_/A _1418_/B vdd gnd OAI21X1
XFILL_0__1617_ vdd gnd FILL
XFILL_3__1326_ vdd gnd FILL
XFILL_1__1390_ vdd gnd FILL
X_1274_ _1274_/A _1274_/B _1274_/C _1301_/B vdd gnd OAI21X1
XFILL_0__1548_ vdd gnd FILL
XFILL_0__1479_ vdd gnd FILL
XFILL_3__1257_ vdd gnd FILL
XFILL_3__1188_ vdd gnd FILL
XFILL_1__1726_ vdd gnd FILL
XFILL_4__1504_ vdd gnd FILL
XFILL_1__1588_ vdd gnd FILL
XFILL_1__1657_ vdd gnd FILL
XFILL_2__1002_ vdd gnd FILL
XFILL_2__979_ vdd gnd FILL
X_985_ _985_/A _987_/B vdd gnd INVX1
XFILL_2__1835_ vdd gnd FILL
XFILL100350x150 vdd gnd FILL
XFILL_2__1697_ vdd gnd FILL
XFILL_2__1766_ vdd gnd FILL
X_1892_ _1892_/D _1897_/CLK _1892_/Q vdd gnd DFFPOSX1
XFILL_0__1333_ vdd gnd FILL
XFILL_0__1402_ vdd gnd FILL
XFILL_3__1111_ vdd gnd FILL
XFILL_3__1042_ vdd gnd FILL
XFILL_0__1264_ vdd gnd FILL
XFILL_0__1195_ vdd gnd FILL
XFILL_1__1511_ vdd gnd FILL
XFILL_1__997_ vdd gnd FILL
X_1326_ _956_/B Cin[4] _1416_/A vdd gnd NAND2X1
XFILL_1__1373_ vdd gnd FILL
XFILL_1__1442_ vdd gnd FILL
XFILL_3__1309_ vdd gnd FILL
X_1257_ _963_/A _1257_/B _1896_/Q _1258_/A vdd gnd OAI21X1
X_1188_ _1188_/A _1188_/B _1243_/A _1193_/B vdd gnd AOI21X1
XFILL_2__1620_ vdd gnd FILL
XFILL_1__1709_ vdd gnd FILL
XFILL_2__1551_ vdd gnd FILL
XFILL_2__1482_ vdd gnd FILL
XFILL_4__1418_ vdd gnd FILL
XFILL_4__1349_ vdd gnd FILL
XFILL_3_BUFX2_insert19 vdd gnd FILL
XFILL_3__1660_ vdd gnd FILL
XFILL_3__1591_ vdd gnd FILL
XFILL_2__1749_ vdd gnd FILL
XFILL_2__1818_ vdd gnd FILL
X_968_ _977_/A _968_/B _968_/C _968_/Y vdd gnd OAI21X1
X_1111_ _1173_/B _1114_/B _1113_/B _1131_/B vdd gnd OAI21X1
X_1042_ _1068_/C _1050_/B vdd gnd INVX1
XFILL_0__1316_ vdd gnd FILL
X_1875_ _1875_/D _1903_/CLK _982_/B vdd gnd DFFPOSX1
XFILL_3__1025_ vdd gnd FILL
XFILL_0__1247_ vdd gnd FILL
XFILL_0__1178_ vdd gnd FILL
XFILL_3__1789_ vdd gnd FILL
X_1309_ Cin[6] _1778_/B vdd gnd INVX1
XFILL_1__1356_ vdd gnd FILL
XFILL_1__1425_ vdd gnd FILL
XFILL_1__1287_ vdd gnd FILL
XFILL_4__1203_ vdd gnd FILL
XFILL_4__1134_ vdd gnd FILL
XFILL_2__1603_ vdd gnd FILL
XFILL_2__1534_ vdd gnd FILL
XFILL_2__1465_ vdd gnd FILL
XFILL_2__1396_ vdd gnd FILL
XFILL_0__998_ vdd gnd FILL
XFILL_0__1032_ vdd gnd FILL
XFILL_0__1101_ vdd gnd FILL
X_1660_ _952_/A Cin[6] _1661_/B vdd gnd NAND2X1
X_1591_ _1611_/A _1596_/B _1592_/B vdd gnd NOR2X1
XFILL_3__1712_ vdd gnd FILL
XFILL_3__1574_ vdd gnd FILL
XFILL_0__1796_ vdd gnd FILL
XFILL_3__1643_ vdd gnd FILL
XFILL_4__976_ vdd gnd FILL
XFILL_1__1210_ vdd gnd FILL
XFILL_1__1141_ vdd gnd FILL
X_1025_ _1036_/A _1026_/B vdd gnd INVX1
XFILL_3__1008_ vdd gnd FILL
X_1858_ _980_/Y _1880_/CLK _978_/A vdd gnd DFFPOSX1
XFILL_1__1072_ vdd gnd FILL
XFILL_4__1683_ vdd gnd FILL
X_1789_ _1789_/A _1791_/C _1790_/B vdd gnd XOR2X1
XFILL_4__1752_ vdd gnd FILL
XFILL_2__1250_ vdd gnd FILL
XFILL_1__1339_ vdd gnd FILL
XFILL_1__1408_ vdd gnd FILL
XFILL_4__1117_ vdd gnd FILL
XFILL_4__1048_ vdd gnd FILL
XFILL_2__1181_ vdd gnd FILL
XFILL_0__1650_ vdd gnd FILL
XFILL_3__994_ vdd gnd FILL
XFILL_2__1517_ vdd gnd FILL
XFILL_0__1581_ vdd gnd FILL
XFILL_2__1448_ vdd gnd FILL
XFILL_2__1379_ vdd gnd FILL
XFILL_3__1290_ vdd gnd FILL
X_1712_ _949_/A Cin[7] _1749_/C vdd gnd NAND2X1
X_1643_ _997_/B _1701_/B vdd gnd INVX1
XFILL_0__1015_ vdd gnd FILL
X_1574_ _1574_/A _1574_/B _1574_/C _1575_/B vdd gnd AOI21X1
XFILL_0__1917_ vdd gnd FILL
XFILL_1__1690_ vdd gnd FILL
XFILL_3__1626_ vdd gnd FILL
XFILL_3__1557_ vdd gnd FILL
XFILL_3__1488_ vdd gnd FILL
XFILL_0__1779_ vdd gnd FILL
XFILL_0__1848_ vdd gnd FILL
X_1008_ _1885_/Q _1801_/B vdd gnd INVX1
XFILL_1__1124_ vdd gnd FILL
XFILL_1__1055_ vdd gnd FILL
XFILL101250x89850 vdd gnd FILL
XFILL_4__1597_ vdd gnd FILL
XFILL_2__1302_ vdd gnd FILL
XFILL_2__1233_ vdd gnd FILL
XFILL_2__1095_ vdd gnd FILL
XFILL_2__1164_ vdd gnd FILL
XFILL_3__977_ vdd gnd FILL
XFILL_0__1633_ vdd gnd FILL
XFILL_0__1564_ vdd gnd FILL
XFILL_0__1702_ vdd gnd FILL
XFILL_3__1411_ vdd gnd FILL
XFILL_3__1342_ vdd gnd FILL
X_1290_ _1290_/A _1290_/B _1290_/C _1292_/C vdd gnd OAI21X1
XFILL_0__1495_ vdd gnd FILL
XFILL_3__1273_ vdd gnd FILL
X_1626_ _1649_/A _1649_/B _1626_/C _1631_/B vdd gnd AOI21X1
XFILL_1__1742_ vdd gnd FILL
X_1557_ _1634_/A _1634_/B _1574_/C _1564_/B vdd gnd OAI21X1
XFILL_3__1609_ vdd gnd FILL
XFILL_1__1673_ vdd gnd FILL
X_1488_ _1571_/A _1492_/B _1572_/B vdd gnd NAND2X1
XFILL_4__1451_ vdd gnd FILL
XFILL_1__1811_ vdd gnd FILL
XFILL_2_BUFX2_insert21 vdd gnd FILL
XFILL_4__1382_ vdd gnd FILL
XFILL_2__995_ vdd gnd FILL
XFILL_1__1107_ vdd gnd FILL
XFILL_2__1782_ vdd gnd FILL
XFILL_1__1038_ vdd gnd FILL
XFILL_0__1280_ vdd gnd FILL
XFILL_2__1216_ vdd gnd FILL
XFILL_2__1078_ vdd gnd FILL
XFILL_2__1147_ vdd gnd FILL
X_1411_ _1499_/B _1419_/A _1419_/B _1427_/A vdd gnd AOI21X1
X_1342_ _955_/A _1449_/B _1348_/A _1352_/A vdd gnd NAND3X1
X_1273_ _1371_/B _1371_/C _1371_/A _1372_/C vdd gnd NAND3X1
XFILL_0__1547_ vdd gnd FILL
XFILL_0__1616_ vdd gnd FILL
XFILL_3__1256_ vdd gnd FILL
XFILL_3__1325_ vdd gnd FILL
XFILL_0__1478_ vdd gnd FILL
XFILL_3__1187_ vdd gnd FILL
X_1609_ _952_/A Cin[4] _955_/A Cin[3] _1611_/C vdd gnd AOI22X1
XFILL_1__1725_ vdd gnd FILL
XFILL_1__1656_ vdd gnd FILL
XFILL_1__1587_ vdd gnd FILL
XFILL_2__1001_ vdd gnd FILL
XFILL100350x7950 vdd gnd FILL
XFILL_2__978_ vdd gnd FILL
XFILL_2__1765_ vdd gnd FILL
X_984_ _992_/A _984_/Y vdd gnd INVX8
XFILL_2__1834_ vdd gnd FILL
XFILL_2__1696_ vdd gnd FILL
XFILL_0__1401_ vdd gnd FILL
XFILL_3__1110_ vdd gnd FILL
X_1891_ _1891_/D _1897_/CLK _1891_/Q vdd gnd DFFPOSX1
XFILL_0__1332_ vdd gnd FILL
XFILL_0__1194_ vdd gnd FILL
XFILL_3__1041_ vdd gnd FILL
XFILL_0__1263_ vdd gnd FILL
XFILL_1__1510_ vdd gnd FILL
XFILL_1__996_ vdd gnd FILL
X_1256_ _952_/A _1449_/B _1256_/C _1258_/B vdd gnd NAND3X1
X_1325_ _1325_/A _1325_/B _1325_/C _1368_/C vdd gnd AOI21X1
XFILL_1__1441_ vdd gnd FILL
XFILL_3__1308_ vdd gnd FILL
XFILL_3__1239_ vdd gnd FILL
XFILL_4__1081_ vdd gnd FILL
XFILL_1__1372_ vdd gnd FILL
X_1187_ _961_/A _1257_/B _1895_/Q _1188_/A vdd gnd OAI21X1
XFILL_1__1708_ vdd gnd FILL
XFILL_2__1550_ vdd gnd FILL
XFILL_1__1639_ vdd gnd FILL
XFILL_2__1481_ vdd gnd FILL
XFILL_2__1679_ vdd gnd FILL
XFILL_3__1590_ vdd gnd FILL
XFILL_2__1748_ vdd gnd FILL
XFILL100350x70350 vdd gnd FILL
XFILL_2__1817_ vdd gnd FILL
X_967_ _967_/A _977_/A _968_/C vdd gnd NAND2X1
X_1110_ _1173_/A _1113_/B vdd gnd INVX1
X_1041_ _953_/B _1104_/B _1900_/Q _1068_/C vdd gnd NAND3X1
XFILL_0__1315_ vdd gnd FILL
XFILL_0__1246_ vdd gnd FILL
XFILL_3__1024_ vdd gnd FILL
X_1874_ _1874_/D _1904_/CLK _979_/B vdd gnd DFFPOSX1
XFILL_0__1177_ vdd gnd FILL
XFILL_3__1788_ vdd gnd FILL
XFILL_1__1424_ vdd gnd FILL
X_1308_ _1403_/B _1316_/A _1316_/B _1321_/A vdd gnd AOI21X1
X_1239_ _1239_/A _1334_/A _1313_/C vdd gnd NAND2X1
XFILL_1__979_ vdd gnd FILL
XFILL_1__1355_ vdd gnd FILL
XFILL_1__1286_ vdd gnd FILL
XFILL_2__1602_ vdd gnd FILL
XFILL_2__1533_ vdd gnd FILL
XFILL_2__1464_ vdd gnd FILL
XFILL_2__1395_ vdd gnd FILL
XFILL_0__997_ vdd gnd FILL
XFILL_0__1031_ vdd gnd FILL
XFILL_0__1100_ vdd gnd FILL
X_1590_ _1652_/C _1594_/A _1594_/B _1601_/B vdd gnd AOI21X1
XFILL_3__1711_ vdd gnd FILL
XFILL_3__1642_ vdd gnd FILL
XFILL_3__1573_ vdd gnd FILL
XFILL_0__1795_ vdd gnd FILL
X_1024_ _1036_/B _1026_/C vdd gnd INVX1
XFILL_1__1140_ vdd gnd FILL
XFILL_4__1820_ vdd gnd FILL
X_1788_ _1799_/A _1788_/B _1791_/C vdd gnd AND2X2
XFILL_3__1007_ vdd gnd FILL
X_1857_ _977_/Y _1910_/CLK _975_/A vdd gnd DFFPOSX1
XFILL_1__1071_ vdd gnd FILL
XFILL_0__1229_ vdd gnd FILL
XFILL_1__1407_ vdd gnd FILL
XFILL_2__1180_ vdd gnd FILL
XFILL_1__1338_ vdd gnd FILL
XFILL_1__1269_ vdd gnd FILL
XFILL_3__993_ vdd gnd FILL
XFILL_0__1580_ vdd gnd FILL
XFILL_2__1516_ vdd gnd FILL
XFILL_2__1447_ vdd gnd FILL
XFILL_2__1378_ vdd gnd FILL
X_1711_ _1711_/A _1711_/B _1711_/C _1728_/B vdd gnd OAI21X1
X_1642_ _1642_/A _1642_/B _1642_/C _1880_/D vdd gnd OAI21X1
XFILL_0__1014_ vdd gnd FILL
XFILL_3__1625_ vdd gnd FILL
X_1573_ _1704_/C _1704_/A _1706_/D _1644_/B vdd gnd AOI21X1
XFILL_0__1916_ vdd gnd FILL
XFILL_0__1847_ vdd gnd FILL
XFILL_3__1556_ vdd gnd FILL
XFILL_3__1487_ vdd gnd FILL
XFILL_0__1778_ vdd gnd FILL
X_1007_ _998_/A _1007_/B _1007_/C _1868_/D vdd gnd OAI21X1
X_1909_ _943_/A _1910_/CLK _1910_/D vdd gnd DFFPOSX1
XFILL_4__958_ vdd gnd FILL
XFILL_1__1054_ vdd gnd FILL
XFILL_1__1123_ vdd gnd FILL
XFILL_4__1734_ vdd gnd FILL
XFILL_4__1665_ vdd gnd FILL
XFILL_2__1232_ vdd gnd FILL
XFILL_2__1301_ vdd gnd FILL
XFILL_2__1163_ vdd gnd FILL
XFILL_2__1094_ vdd gnd FILL
XFILL_0__1701_ vdd gnd FILL
XFILL_3__976_ vdd gnd FILL
XFILL_0__1632_ vdd gnd FILL
XFILL_0__1563_ vdd gnd FILL
XFILL_3__1410_ vdd gnd FILL
XFILL_3__1341_ vdd gnd FILL
XFILL_3__1272_ vdd gnd FILL
XFILL_0__1494_ vdd gnd FILL
X_1625_ _1625_/A _1625_/B _1625_/C _1645_/C vdd gnd OAI21X1
X_1556_ _1556_/A _1556_/B _1625_/B _1634_/B vdd gnd AOI21X1
XFILL_1__1810_ vdd gnd FILL
XFILL_2_BUFX2_insert22 vdd gnd FILL
XFILL_1__1672_ vdd gnd FILL
XFILL_1__1741_ vdd gnd FILL
XFILL_3__1608_ vdd gnd FILL
XFILL_3__1539_ vdd gnd FILL
X_1487_ _1487_/A _1565_/D _1487_/C _1492_/B vdd gnd OAI21X1
XFILL_2__994_ vdd gnd FILL
XFILL_1__1037_ vdd gnd FILL
XFILL_1__1106_ vdd gnd FILL
XFILL_2__1781_ vdd gnd FILL
XFILL_4__1579_ vdd gnd FILL
XFILL_2__1146_ vdd gnd FILL
XFILL_2__1215_ vdd gnd FILL
X_1410_ _1847_/B _1778_/B _1502_/A _1419_/A vdd gnd OAI21X1
XFILL_2__1077_ vdd gnd FILL
X_1341_ _1897_/Q _1348_/A vdd gnd INVX1
XFILL_3__959_ vdd gnd FILL
X_1272_ _1299_/B _1299_/A _1301_/A vdd gnd XOR2X1
XFILL_0__1546_ vdd gnd FILL
XFILL_0__1615_ vdd gnd FILL
XFILL_0__1477_ vdd gnd FILL
XFILL_3__1255_ vdd gnd FILL
XFILL_3__1324_ vdd gnd FILL
XFILL_3__1186_ vdd gnd FILL
X_1608_ _1611_/A _1723_/B _1670_/C vdd gnd AND2X2
X_1539_ _1539_/A _1539_/B _1539_/C _1620_/B vdd gnd NAND3X1
XFILL_1__1586_ vdd gnd FILL
XFILL_1__1724_ vdd gnd FILL
XFILL_1__1655_ vdd gnd FILL
XFILL_4__1433_ vdd gnd FILL
XFILL_4__1364_ vdd gnd FILL
XFILL_4__1295_ vdd gnd FILL
XFILL_2__1000_ vdd gnd FILL
XFILL_2__977_ vdd gnd FILL
XFILL_2__1695_ vdd gnd FILL
XFILL_2__1764_ vdd gnd FILL
XFILL_2__1833_ vdd gnd FILL
X_983_ _983_/A _983_/B _983_/C _983_/Y vdd gnd OAI21X1
XFILL_0__1400_ vdd gnd FILL
XFILL_0__1331_ vdd gnd FILL
XFILL_3__1040_ vdd gnd FILL
X_1890_ _1890_/D _1897_/CLK _1890_/Q vdd gnd DFFPOSX1
XFILL_0__1262_ vdd gnd FILL
XFILL_2__1129_ vdd gnd FILL
XFILL_0__1193_ vdd gnd FILL
XFILL_1__1440_ vdd gnd FILL
XFILL_1__995_ vdd gnd FILL
X_1255_ _1896_/Q _1256_/C vdd gnd INVX1
X_1324_ _1361_/C _1325_/C vdd gnd INVX1
X_1186_ _949_/A _1248_/B _1186_/C _1188_/B vdd gnd NAND3X1
XFILL_0__1529_ vdd gnd FILL
XFILL_3__1307_ vdd gnd FILL
XFILL_3__1238_ vdd gnd FILL
XFILL_1__1371_ vdd gnd FILL
XFILL_3__1169_ vdd gnd FILL
XFILL_1__1638_ vdd gnd FILL
XFILL_1__1707_ vdd gnd FILL
XFILL_2__1480_ vdd gnd FILL
XFILL_1__1569_ vdd gnd FILL
XFILL_4__1278_ vdd gnd FILL
XFILL_2__1816_ vdd gnd FILL
XFILL_2__1678_ vdd gnd FILL
XFILL_2__1747_ vdd gnd FILL
X_966_ _966_/A _968_/B vdd gnd INVX1
X_1040_ _953_/B _1106_/B _1900_/Q _1068_/B vdd gnd AOI21X1
XFILL_4__991_ vdd gnd FILL
XFILL_0__1314_ vdd gnd FILL
XFILL_3__1023_ vdd gnd FILL
X_1873_ _1873_/D _1903_/CLK _976_/B vdd gnd DFFPOSX1
XFILL_0__1176_ vdd gnd FILL
XFILL_0__1245_ vdd gnd FILL
XFILL_3__1787_ vdd gnd FILL
XFILL_1__1423_ vdd gnd FILL
X_1307_ _1847_/B _1413_/B _1425_/A _1316_/A vdd gnd OAI21X1
XFILL_1__978_ vdd gnd FILL
X_1238_ _946_/A Cin[3] _1334_/A vdd gnd AND2X2
XFILL_4__1132_ vdd gnd FILL
X_1169_ _1169_/A _1239_/A _1171_/C vdd gnd NAND2X1
XFILL_1__1354_ vdd gnd FILL
XFILL_1__1285_ vdd gnd FILL
XFILL_4__1063_ vdd gnd FILL
XFILL_2__1601_ vdd gnd FILL
XFILL_2__1532_ vdd gnd FILL
XFILL_2__1463_ vdd gnd FILL
XFILL_3_CLKBUF1_insert10 vdd gnd FILL
XFILL100950x31350 vdd gnd FILL
XFILL_2__1394_ vdd gnd FILL
XFILL100650x66450 vdd gnd FILL
XFILL_0__996_ vdd gnd FILL
XFILL_0__1030_ vdd gnd FILL
XFILL_3__1710_ vdd gnd FILL
XFILL_3__1572_ vdd gnd FILL
XFILL_3__1641_ vdd gnd FILL
XFILL_0__1794_ vdd gnd FILL
X_949_ _949_/A _961_/A vdd gnd INVX1
X_1023_ _1036_/B _1023_/B _1036_/A _1027_/B vdd gnd OAI21X1
XFILL_3__1006_ vdd gnd FILL
XFILL_1__1070_ vdd gnd FILL
XFILL_0__1228_ vdd gnd FILL
X_1787_ _1792_/A _1792_/B _1788_/B vdd gnd NAND2X1
X_1856_ _974_/Y _1903_/CLK _972_/A vdd gnd DFFPOSX1
XFILL_0__1159_ vdd gnd FILL
XFILL_3__1839_ vdd gnd FILL
XFILL_1__1337_ vdd gnd FILL
XFILL_1__1406_ vdd gnd FILL
XFILL_1__1199_ vdd gnd FILL
XFILL_1__1268_ vdd gnd FILL
XFILL_3__992_ vdd gnd FILL
XFILL_2__1515_ vdd gnd FILL
XFILL_2__1446_ vdd gnd FILL
XFILL100950x43050 vdd gnd FILL
XFILL100650x78150 vdd gnd FILL
XFILL_2__1377_ vdd gnd FILL
X_1710_ _1710_/A _1710_/B _1733_/B _1731_/B vdd gnd OAI21X1
X_1572_ _1572_/A _1572_/B _1704_/A vdd gnd NOR2X1
X_1641_ _1703_/B _1644_/B _992_/A _1642_/A vdd gnd OAI21X1
XFILL_0__1013_ vdd gnd FILL
XFILL_0__979_ vdd gnd FILL
XFILL_3__1624_ vdd gnd FILL
XFILL_3__1555_ vdd gnd FILL
XFILL_0__1915_ vdd gnd FILL
XFILL_0__1846_ vdd gnd FILL
XFILL_0__1777_ vdd gnd FILL
XFILL_3__1486_ vdd gnd FILL
X_1006_ _998_/A _1884_/Q _1007_/C vdd gnd NAND2X1
X_1908_ _927_/A _1908_/CLK _943_/A vdd gnd DFFPOSX1
X_1839_ _948_/A _1839_/B _1839_/C _1900_/D vdd gnd AOI21X1
XFILL_1__1122_ vdd gnd FILL
XFILL_1__1053_ vdd gnd FILL
XFILL_4__1802_ vdd gnd FILL
XFILL_2__1300_ vdd gnd FILL
XFILL_2__1093_ vdd gnd FILL
XFILL_2__1231_ vdd gnd FILL
XFILL_2__1162_ vdd gnd FILL
XFILL_0__1700_ vdd gnd FILL
XFILL_3__975_ vdd gnd FILL
XFILL_0__1631_ vdd gnd FILL
XFILL_0__1562_ vdd gnd FILL
XFILL_0__1493_ vdd gnd FILL
XFILL_2__1429_ vdd gnd FILL
XFILL_3__1340_ vdd gnd FILL
XFILL_3__1271_ vdd gnd FILL
X_1624_ _1645_/A _1645_/B _1631_/C _1637_/A vdd gnd NAND3X1
XFILL_1__1740_ vdd gnd FILL
X_1555_ _1555_/A _1555_/B _1555_/C _1556_/A vdd gnd OAI21X1
XFILL_2_BUFX2_insert23 vdd gnd FILL
XFILL_2_BUFX2_insert12 vdd gnd FILL
XFILL_1__1671_ vdd gnd FILL
XFILL_3__1538_ vdd gnd FILL
XFILL_3__1607_ vdd gnd FILL
X_1486_ _1486_/A _1486_/B _1486_/C _1565_/D vdd gnd AOI21X1
XFILL_0__1829_ vdd gnd FILL
XFILL_3__1469_ vdd gnd FILL
XFILL_2__993_ vdd gnd FILL
XFILL_1__1105_ vdd gnd FILL
XFILL_1__1036_ vdd gnd FILL
XFILL_4__1647_ vdd gnd FILL
XFILL_2__1780_ vdd gnd FILL
XFILL_4__1716_ vdd gnd FILL
XFILL_2__1076_ vdd gnd FILL
XFILL_2__1145_ vdd gnd FILL
XFILL_2__1214_ vdd gnd FILL
X_1340_ _952_/A Cin[1] _1450_/A vdd gnd NAND2X1
XFILL_0_CLKBUF1_insert5 vdd gnd FILL
XFILL_0__1614_ vdd gnd FILL
XFILL_3__958_ vdd gnd FILL
X_1271_ _1372_/B _1280_/B _1280_/A _1382_/A vdd gnd NAND3X1
XFILL_0__1545_ vdd gnd FILL
XFILL_0__1476_ vdd gnd FILL
XFILL_4_BUFX2_insert2 vdd gnd FILL
XFILL_3__1323_ vdd gnd FILL
XFILL_3__1185_ vdd gnd FILL
XFILL_3__1254_ vdd gnd FILL
X_1538_ _1538_/A _1538_/B _1554_/A vdd gnd NAND2X1
XFILL_4__1501_ vdd gnd FILL
XFILL_1__1723_ vdd gnd FILL
X_1607_ _955_/A Cin[4] _1723_/B vdd gnd AND2X2
X_1469_ _1551_/B _1551_/C _1551_/A _1552_/C vdd gnd NAND3X1
XFILL_1__1585_ vdd gnd FILL
XFILL_1__1654_ vdd gnd FILL
XFILL_2__976_ vdd gnd FILL
XFILL_2__1832_ vdd gnd FILL
XFILL_1__1019_ vdd gnd FILL
XFILL_2__1694_ vdd gnd FILL
XFILL_2__1763_ vdd gnd FILL
X_982_ _983_/A _982_/B _983_/C vdd gnd NAND2X1
XFILL_0__1330_ vdd gnd FILL
XFILL_0__1261_ vdd gnd FILL
XFILL_2__1128_ vdd gnd FILL
XFILL_0__1192_ vdd gnd FILL
XFILL_2__1059_ vdd gnd FILL
XFILL_1__994_ vdd gnd FILL
X_1323_ _1366_/A _1399_/B _1474_/A vdd gnd NAND2X1
XFILL_3__1306_ vdd gnd FILL
XFILL_1__1370_ vdd gnd FILL
X_1185_ _1895_/Q _1186_/C vdd gnd INVX1
X_1254_ _1254_/A _1338_/C _1254_/C _1263_/A vdd gnd AOI21X1
XFILL_0__1528_ vdd gnd FILL
XFILL_0__1459_ vdd gnd FILL
XFILL_3__1237_ vdd gnd FILL
XFILL_3__1168_ vdd gnd FILL
XFILL_3__1099_ vdd gnd FILL
XFILL_1__1706_ vdd gnd FILL
XFILL_4__1415_ vdd gnd FILL
XFILL_1__1637_ vdd gnd FILL
XFILL_4__1346_ vdd gnd FILL
XFILL_1__1568_ vdd gnd FILL
XFILL_1__1499_ vdd gnd FILL
XFILL_2__959_ vdd gnd FILL
XFILL_2__1815_ vdd gnd FILL
X_965_ _965_/A _965_/B _965_/C _965_/Y vdd gnd OAI21X1
XFILL_2__1677_ vdd gnd FILL
XFILL_2__1746_ vdd gnd FILL
XFILL_0__1313_ vdd gnd FILL
XFILL_3__1022_ vdd gnd FILL
XFILL_0__1244_ vdd gnd FILL
X_1872_ _1872_/D _1903_/CLK _973_/B vdd gnd DFFPOSX1
XFILL_0__1175_ vdd gnd FILL
XFILL_3__1786_ vdd gnd FILL
X_1306_ _950_/B Cin[6] _1425_/A vdd gnd NAND2X1
XFILL_1__977_ vdd gnd FILL
XFILL_1__1353_ vdd gnd FILL
XFILL_1__1422_ vdd gnd FILL
X_1237_ _1313_/A _1317_/A vdd gnd INVX1
XFILL_4__1200_ vdd gnd FILL
X_1099_ _979_/B _1216_/A _1151_/C vdd gnd NAND2X1
X_1168_ _1168_/A _1171_/A vdd gnd INVX1
XFILL_1__1284_ vdd gnd FILL
XFILL_2__1600_ vdd gnd FILL
XFILL_2__1531_ vdd gnd FILL
XFILL_2__1462_ vdd gnd FILL
XFILL_3_CLKBUF1_insert11 vdd gnd FILL
XFILL_2__1393_ vdd gnd FILL
XFILL_0__995_ vdd gnd FILL
XFILL_2__1729_ vdd gnd FILL
XFILL_0__1793_ vdd gnd FILL
XFILL_3__1571_ vdd gnd FILL
XFILL_3__1640_ vdd gnd FILL
X_948_ _948_/A _959_/A _948_/C _948_/Y vdd gnd OAI21X1
X_1022_ _947_/B Cin[1] _1036_/A vdd gnd NAND2X1
XFILL_4__973_ vdd gnd FILL
XFILL_3__1005_ vdd gnd FILL
X_1855_ _971_/Y _1880_/CLK _969_/A vdd gnd DFFPOSX1
XFILL_0__1227_ vdd gnd FILL
XFILL_4__1680_ vdd gnd FILL
X_1786_ _1792_/B _1792_/A _1799_/A vdd gnd OR2X2
XFILL_3__1838_ vdd gnd FILL
XFILL_0__1089_ vdd gnd FILL
XFILL_0__1158_ vdd gnd FILL
XFILL_3__1769_ vdd gnd FILL
XFILL_1__1405_ vdd gnd FILL
XFILL_1__1336_ vdd gnd FILL
XFILL_4__1114_ vdd gnd FILL
XFILL_4__1045_ vdd gnd FILL
XFILL_1__1198_ vdd gnd FILL
XFILL_1__1267_ vdd gnd FILL
XFILL_3__991_ vdd gnd FILL
XFILL_2__1514_ vdd gnd FILL
XFILL_2__1445_ vdd gnd FILL
XFILL100950x7950 vdd gnd FILL
XFILL_2__1376_ vdd gnd FILL
XFILL_0__978_ vdd gnd FILL
X_1571_ _1571_/A _1572_/A _1571_/C _1706_/D vdd gnd OAI21X1
X_1640_ _1644_/B _1703_/B _1642_/B vdd gnd AND2X2
XFILL_0__1012_ vdd gnd FILL
XFILL_3__1623_ vdd gnd FILL
XFILL_3__1554_ vdd gnd FILL
XFILL_0__1776_ vdd gnd FILL
XFILL_3__1485_ vdd gnd FILL
XFILL_0__1914_ vdd gnd FILL
XFILL_0__1845_ vdd gnd FILL
X_1005_ _938_/B _1007_/B vdd gnd INVX1
XFILL_1__1121_ vdd gnd FILL
X_1907_ _957_/A _1908_/CLK _927_/A vdd gnd DFFPOSX1
X_1838_ _948_/A _1900_/Q _1839_/C vdd gnd NOR2X1
XFILL_1__1052_ vdd gnd FILL
XFILL_4__1594_ vdd gnd FILL
X_1769_ _1790_/A _1769_/B _1769_/C _1769_/D _1883_/D vdd gnd AOI22X1
XFILL_2__1230_ vdd gnd FILL
XFILL_1__1319_ vdd gnd FILL
XFILL_2__1161_ vdd gnd FILL
XFILL_2__1092_ vdd gnd FILL
XFILL_0__1630_ vdd gnd FILL
XFILL_3__974_ vdd gnd FILL
XFILL_0__1561_ vdd gnd FILL
XFILL_0__1492_ vdd gnd FILL
XFILL_2__1428_ vdd gnd FILL
XFILL_2__1359_ vdd gnd FILL
XFILL_3__1270_ vdd gnd FILL
X_1623_ _1649_/A _1649_/B _1626_/C _1645_/B vdd gnd NAND3X1
X_1554_ _1554_/A _1620_/B _1554_/C _1556_/B vdd gnd NAND3X1
X_1485_ _1494_/B _1493_/A _1494_/A _1487_/A vdd gnd AOI21X1
XFILL_2_BUFX2_insert24 vdd gnd FILL
XFILL_2_BUFX2_insert13 vdd gnd FILL
.ends


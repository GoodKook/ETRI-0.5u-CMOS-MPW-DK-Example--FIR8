VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fir_pe
  CLASS BLOCK ;
  FOREIGN fir_pe ;
  ORIGIN 6.000 6.000 ;
  SIZE 912.000 BY 912.000 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 897.300 909.450 899.700 ;
        RECT 900.450 821.700 909.450 897.300 ;
        RECT 0.600 819.300 909.450 821.700 ;
        RECT 900.450 743.700 909.450 819.300 ;
        RECT 0.600 741.300 909.450 743.700 ;
        RECT 900.450 665.700 909.450 741.300 ;
        RECT 0.600 663.300 909.450 665.700 ;
        RECT 900.450 587.700 909.450 663.300 ;
        RECT 0.600 585.300 909.450 587.700 ;
        RECT 900.450 509.700 909.450 585.300 ;
        RECT 0.600 507.300 909.450 509.700 ;
        RECT 900.450 431.700 909.450 507.300 ;
        RECT 0.600 429.300 909.450 431.700 ;
        RECT 900.450 353.700 909.450 429.300 ;
        RECT 0.600 351.300 909.450 353.700 ;
        RECT 900.450 275.700 909.450 351.300 ;
        RECT 0.600 273.300 909.450 275.700 ;
        RECT 900.450 197.700 909.450 273.300 ;
        RECT 0.600 195.300 909.450 197.700 ;
        RECT 900.450 119.700 909.450 195.300 ;
        RECT 0.600 117.300 909.450 119.700 ;
        RECT 900.450 41.700 909.450 117.300 ;
        RECT 0.600 39.300 909.450 41.700 ;
        RECT 900.450 0.300 909.450 39.300 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -9.450 860.700 -0.450 899.700 ;
        RECT -9.450 858.300 899.400 860.700 ;
        RECT -9.450 782.700 -0.450 858.300 ;
        RECT -9.450 780.300 899.400 782.700 ;
        RECT -9.450 704.700 -0.450 780.300 ;
        RECT -9.450 702.300 899.400 704.700 ;
        RECT -9.450 626.700 -0.450 702.300 ;
        RECT -9.450 624.300 899.400 626.700 ;
        RECT -9.450 548.700 -0.450 624.300 ;
        RECT -9.450 546.300 899.400 548.700 ;
        RECT -9.450 470.700 -0.450 546.300 ;
        RECT -9.450 468.300 899.400 470.700 ;
        RECT -9.450 392.700 -0.450 468.300 ;
        RECT -9.450 390.300 899.400 392.700 ;
        RECT -9.450 314.700 -0.450 390.300 ;
        RECT -9.450 312.300 899.400 314.700 ;
        RECT -9.450 236.700 -0.450 312.300 ;
        RECT -9.450 234.300 899.400 236.700 ;
        RECT -9.450 158.700 -0.450 234.300 ;
        RECT -9.450 156.300 899.400 158.700 ;
        RECT -9.450 80.700 -0.450 156.300 ;
        RECT -9.450 78.300 899.400 80.700 ;
        RECT -9.450 2.700 -0.450 78.300 ;
        RECT -9.450 0.300 899.400 2.700 ;
    END
  END vdd
  PIN Cin[7]
    PORT
      LAYER metal1 ;
        RECT 346.950 375.450 349.050 376.050 ;
        RECT 352.950 375.450 355.050 376.050 ;
        RECT 346.950 374.550 355.050 375.450 ;
        RECT 346.950 373.950 349.050 374.550 ;
        RECT 352.950 373.950 355.050 374.550 ;
        RECT 334.950 342.450 337.050 342.900 ;
        RECT 346.950 342.450 349.050 343.200 ;
        RECT 334.950 341.550 349.050 342.450 ;
        RECT 334.950 340.800 337.050 341.550 ;
        RECT 346.950 341.100 349.050 341.550 ;
      LAYER metal2 ;
        RECT 373.950 494.100 376.050 496.200 ;
        RECT 385.950 494.100 388.050 496.200 ;
        RECT 365.400 489.900 366.600 490.650 ;
        RECT 374.400 490.050 375.450 494.100 ;
        RECT 386.400 493.350 387.600 494.100 ;
        RECT 364.950 487.800 367.050 489.900 ;
        RECT 373.950 487.950 376.050 490.050 ;
        RECT 365.400 466.050 366.450 487.800 ;
        RECT 340.950 463.950 343.050 466.050 ;
        RECT 364.950 463.950 367.050 466.050 ;
        RECT 341.400 450.600 342.450 463.950 ;
        RECT 341.400 448.350 342.600 450.600 ;
        RECT 374.400 394.050 375.450 487.950 ;
        RECT 352.950 391.950 355.050 394.050 ;
        RECT 373.950 391.950 376.050 394.050 ;
        RECT 160.950 382.950 163.050 385.050 ;
        RECT 161.400 376.050 162.450 382.950 ;
        RECT 353.400 376.050 354.450 391.950 ;
        RECT 160.950 372.000 163.050 376.050 ;
        RECT 169.950 373.950 172.050 376.050 ;
        RECT 346.950 373.950 349.050 376.050 ;
        RECT 352.950 373.950 355.050 376.050 ;
        RECT 161.400 370.350 162.600 372.000 ;
        RECT 170.400 352.050 171.450 373.950 ;
        RECT 169.950 349.950 172.050 352.050 ;
        RECT 193.950 349.950 196.050 352.050 ;
        RECT 194.400 313.050 195.450 349.950 ;
        RECT 347.400 343.200 348.450 373.950 ;
        RECT 353.400 372.600 354.450 373.950 ;
        RECT 353.400 370.350 354.600 372.600 ;
        RECT 334.950 340.800 337.050 342.900 ;
        RECT 346.950 341.100 349.050 343.200 ;
        RECT 296.400 332.400 297.600 334.650 ;
        RECT 296.400 322.050 297.450 332.400 ;
        RECT 335.400 322.050 336.450 340.800 ;
        RECT 226.950 319.950 229.050 322.050 ;
        RECT 295.950 319.950 298.050 322.050 ;
        RECT 334.950 319.950 337.050 322.050 ;
        RECT 227.400 313.050 228.450 319.950 ;
        RECT 193.950 310.950 196.050 313.050 ;
        RECT 226.950 310.950 229.050 313.050 ;
        RECT 227.400 295.200 228.450 310.950 ;
        RECT 226.950 293.100 229.050 295.200 ;
        RECT 227.400 292.350 228.600 293.100 ;
        RECT 245.400 288.900 246.600 289.650 ;
        RECT 244.950 286.800 247.050 288.900 ;
      LAYER via2 ;
        RECT 160.950 373.950 163.050 376.050 ;
      LAYER metal3 ;
        RECT 373.950 495.750 376.050 496.200 ;
        RECT 385.950 495.750 388.050 496.200 ;
        RECT 373.950 494.550 388.050 495.750 ;
        RECT 373.950 494.100 376.050 494.550 ;
        RECT 385.950 494.100 388.050 494.550 ;
        RECT 364.950 489.600 367.050 489.900 ;
        RECT 373.950 489.600 376.050 490.050 ;
        RECT 364.950 488.400 376.050 489.600 ;
        RECT 364.950 487.800 367.050 488.400 ;
        RECT 373.950 487.950 376.050 488.400 ;
        RECT 340.950 465.600 343.050 466.050 ;
        RECT 364.950 465.600 367.050 466.050 ;
        RECT 340.950 464.400 367.050 465.600 ;
        RECT 340.950 463.950 343.050 464.400 ;
        RECT 364.950 463.950 367.050 464.400 ;
        RECT 352.950 393.600 355.050 394.050 ;
        RECT 373.950 393.600 376.050 394.050 ;
        RECT 352.950 392.400 376.050 393.600 ;
        RECT 352.950 391.950 355.050 392.400 ;
        RECT 373.950 391.950 376.050 392.400 ;
        RECT 160.950 384.600 163.050 385.050 ;
        RECT -3.600 383.400 163.050 384.600 ;
        RECT 160.950 382.950 163.050 383.400 ;
        RECT 160.950 375.600 163.050 376.050 ;
        RECT 169.950 375.600 172.050 376.050 ;
        RECT 160.950 374.400 172.050 375.600 ;
        RECT 160.950 373.950 163.050 374.400 ;
        RECT 169.950 373.950 172.050 374.400 ;
        RECT 169.950 351.600 172.050 352.050 ;
        RECT 193.950 351.600 196.050 352.050 ;
        RECT 169.950 350.400 196.050 351.600 ;
        RECT 169.950 349.950 172.050 350.400 ;
        RECT 193.950 349.950 196.050 350.400 ;
        RECT 226.950 321.600 229.050 322.050 ;
        RECT 295.950 321.600 298.050 322.050 ;
        RECT 334.950 321.600 337.050 322.050 ;
        RECT 226.950 320.400 337.050 321.600 ;
        RECT 226.950 319.950 229.050 320.400 ;
        RECT 295.950 319.950 298.050 320.400 ;
        RECT 334.950 319.950 337.050 320.400 ;
        RECT 193.950 312.600 196.050 313.050 ;
        RECT 226.950 312.600 229.050 313.050 ;
        RECT 193.950 311.400 229.050 312.600 ;
        RECT 193.950 310.950 196.050 311.400 ;
        RECT 226.950 310.950 229.050 311.400 ;
        RECT 226.950 294.600 229.050 295.200 ;
        RECT 226.950 293.400 246.600 294.600 ;
        RECT 226.950 293.100 229.050 293.400 ;
        RECT 245.400 288.900 246.600 293.400 ;
        RECT 244.950 286.800 247.050 288.900 ;
    END
  END Cin[7]
  PIN Cin[6]
    PORT
      LAYER metal1 ;
        RECT 316.950 375.450 319.050 376.050 ;
        RECT 322.950 375.450 325.050 376.050 ;
        RECT 331.950 375.450 334.050 376.200 ;
        RECT 316.950 374.550 334.050 375.450 ;
        RECT 316.950 373.950 319.050 374.550 ;
        RECT 322.950 373.950 325.050 374.550 ;
        RECT 331.950 374.100 334.050 374.550 ;
      LAYER metal2 ;
        RECT 214.950 494.100 217.050 496.200 ;
        RECT 223.950 494.100 226.050 496.200 ;
        RECT 215.400 493.350 216.600 494.100 ;
        RECT 224.400 490.050 225.450 494.100 ;
        RECT 223.950 487.950 226.050 490.050 ;
        RECT 233.400 489.900 234.600 490.650 ;
        RECT 224.400 463.050 225.450 487.950 ;
        RECT 232.950 487.800 235.050 489.900 ;
        RECT 208.950 460.950 211.050 463.050 ;
        RECT 223.950 460.950 226.050 463.050 ;
        RECT 209.400 444.900 210.450 460.950 ;
        RECT 221.400 444.900 222.600 445.650 ;
        RECT 208.950 442.800 211.050 444.900 ;
        RECT 220.950 442.800 223.050 444.900 ;
        RECT 209.400 418.200 210.450 442.800 ;
        RECT 208.950 416.100 211.050 418.200 ;
        RECT 209.400 415.350 210.600 416.100 ;
        RECT 229.950 415.950 232.050 418.050 ;
        RECT 331.950 416.100 334.050 418.200 ;
        RECT 343.950 416.100 346.050 418.200 ;
        RECT 230.400 382.050 231.450 415.950 ;
        RECT 106.950 379.950 109.050 382.050 ;
        RECT 229.950 379.950 232.050 382.050 ;
        RECT 107.400 376.050 108.450 379.950 ;
        RECT 106.950 373.950 109.050 376.050 ;
        RECT 107.400 372.600 108.450 373.950 ;
        RECT 107.400 370.350 108.600 372.600 ;
        RECT 230.400 358.050 231.450 379.950 ;
        RECT 332.400 376.200 333.450 416.100 ;
        RECT 344.400 415.350 345.600 416.100 ;
        RECT 316.950 372.000 319.050 376.050 ;
        RECT 322.950 373.950 325.050 376.050 ;
        RECT 331.950 374.100 334.050 376.200 ;
        RECT 317.400 370.350 318.600 372.000 ;
        RECT 263.400 365.400 264.600 367.650 ;
        RECT 263.400 358.050 264.450 365.400 ;
        RECT 229.950 355.950 232.050 358.050 ;
        RECT 262.950 357.450 265.050 358.050 ;
        RECT 319.950 357.450 322.050 358.050 ;
        RECT 323.400 357.450 324.450 373.950 ;
        RECT 377.400 365.400 378.600 367.650 ;
        RECT 377.400 358.050 378.450 365.400 ;
        RECT 262.950 356.400 267.450 357.450 ;
        RECT 262.950 355.950 265.050 356.400 ;
        RECT 230.400 333.900 231.600 334.650 ;
        RECT 260.400 333.900 261.600 334.650 ;
        RECT 266.400 333.900 267.450 356.400 ;
        RECT 319.950 356.400 324.450 357.450 ;
        RECT 319.950 355.950 322.050 356.400 ;
        RECT 376.950 355.950 379.050 358.050 ;
        RECT 320.400 339.600 321.450 355.950 ;
        RECT 320.400 337.350 321.600 339.600 ;
        RECT 229.950 331.800 232.050 333.900 ;
        RECT 259.950 331.800 262.050 333.900 ;
        RECT 265.950 331.800 268.050 333.900 ;
      LAYER metal3 ;
        RECT 214.950 495.750 217.050 496.200 ;
        RECT 223.950 495.750 226.050 496.200 ;
        RECT 214.950 494.550 226.050 495.750 ;
        RECT 214.950 494.100 217.050 494.550 ;
        RECT 223.950 494.100 226.050 494.550 ;
        RECT 223.950 489.600 226.050 490.050 ;
        RECT 232.950 489.600 235.050 489.900 ;
        RECT 223.950 488.400 235.050 489.600 ;
        RECT 223.950 487.950 226.050 488.400 ;
        RECT 232.950 487.800 235.050 488.400 ;
        RECT 208.950 462.600 211.050 463.050 ;
        RECT 223.950 462.600 226.050 463.050 ;
        RECT 208.950 461.400 226.050 462.600 ;
        RECT 208.950 460.950 211.050 461.400 ;
        RECT 223.950 460.950 226.050 461.400 ;
        RECT 208.950 444.450 211.050 444.900 ;
        RECT 220.950 444.450 223.050 444.900 ;
        RECT 208.950 443.250 223.050 444.450 ;
        RECT 208.950 442.800 211.050 443.250 ;
        RECT 220.950 442.800 223.050 443.250 ;
        RECT 208.950 417.600 211.050 418.200 ;
        RECT 229.950 417.600 232.050 418.050 ;
        RECT 208.950 416.400 232.050 417.600 ;
        RECT 208.950 416.100 211.050 416.400 ;
        RECT 229.950 415.950 232.050 416.400 ;
        RECT 331.950 417.750 334.050 418.200 ;
        RECT 343.950 417.750 346.050 418.200 ;
        RECT 331.950 416.550 346.050 417.750 ;
        RECT 331.950 416.100 334.050 416.550 ;
        RECT 343.950 416.100 346.050 416.550 ;
        RECT 106.950 381.600 109.050 382.050 ;
        RECT 229.950 381.600 232.050 382.050 ;
        RECT 106.950 380.400 232.050 381.600 ;
        RECT 106.950 379.950 109.050 380.400 ;
        RECT 229.950 379.950 232.050 380.400 ;
        RECT 106.950 375.600 109.050 376.050 ;
        RECT -3.600 374.400 109.050 375.600 ;
        RECT -3.600 371.400 -2.400 374.400 ;
        RECT 106.950 373.950 109.050 374.400 ;
        RECT 229.950 357.600 232.050 358.050 ;
        RECT 262.950 357.600 265.050 358.050 ;
        RECT 319.950 357.600 322.050 358.050 ;
        RECT 376.950 357.600 379.050 358.050 ;
        RECT 229.950 356.400 379.050 357.600 ;
        RECT 229.950 355.950 232.050 356.400 ;
        RECT 262.950 355.950 265.050 356.400 ;
        RECT 319.950 355.950 322.050 356.400 ;
        RECT 376.950 355.950 379.050 356.400 ;
        RECT 230.400 335.400 267.600 336.600 ;
        RECT 230.400 333.900 231.600 335.400 ;
        RECT 266.400 333.900 267.600 335.400 ;
        RECT 229.950 331.800 232.050 333.900 ;
        RECT 259.950 333.450 262.050 333.900 ;
        RECT 265.950 333.450 268.050 333.900 ;
        RECT 259.950 332.250 268.050 333.450 ;
        RECT 259.950 331.800 262.050 332.250 ;
        RECT 265.950 331.800 268.050 332.250 ;
    END
  END Cin[6]
  PIN Cin[5]
    PORT
      LAYER metal2 ;
        RECT 262.950 449.100 265.050 451.200 ;
        RECT 283.950 449.100 286.050 451.200 ;
        RECT 319.950 449.100 322.050 451.200 ;
        RECT 325.950 449.100 328.050 451.200 ;
        RECT 263.400 448.350 264.600 449.100 ;
        RECT 1.950 442.950 4.050 445.050 ;
        RECT 200.400 443.400 201.600 445.650 ;
        RECT 227.400 443.400 228.600 445.650 ;
        RECT 284.400 445.050 285.450 449.100 ;
        RECT 320.400 448.350 321.600 449.100 ;
        RECT 2.400 430.050 3.450 442.950 ;
        RECT 200.400 436.050 201.450 443.400 ;
        RECT 227.400 436.050 228.450 443.400 ;
        RECT 283.950 442.950 286.050 445.050 ;
        RECT 290.400 444.900 291.600 445.650 ;
        RECT 289.950 442.800 292.050 444.900 ;
        RECT 290.400 436.050 291.450 442.800 ;
        RECT 199.950 433.950 202.050 436.050 ;
        RECT 217.950 433.950 220.050 436.050 ;
        RECT 226.950 433.950 229.050 436.050 ;
        RECT 289.950 433.950 292.050 436.050 ;
        RECT 200.400 430.050 201.450 433.950 ;
        RECT 1.950 427.950 4.050 430.050 ;
        RECT 199.950 427.950 202.050 430.050 ;
        RECT 218.400 385.050 219.450 433.950 ;
        RECT 290.400 424.050 291.450 433.950 ;
        RECT 326.400 424.050 327.450 449.100 ;
        RECT 289.950 421.950 292.050 424.050 ;
        RECT 319.950 421.950 322.050 424.050 ;
        RECT 325.950 421.950 328.050 424.050 ;
        RECT 320.400 417.600 321.450 421.950 ;
        RECT 320.400 415.350 321.600 417.600 ;
        RECT 217.950 382.950 220.050 385.050 ;
        RECT 247.950 382.950 250.050 385.050 ;
        RECT 253.950 382.950 256.050 385.050 ;
        RECT 218.400 372.600 219.450 382.950 ;
        RECT 218.400 370.350 219.600 372.600 ;
        RECT 245.400 372.450 246.600 372.600 ;
        RECT 248.400 372.450 249.450 382.950 ;
        RECT 245.400 371.400 249.450 372.450 ;
        RECT 245.400 370.350 246.600 371.400 ;
        RECT 254.400 361.050 255.450 382.950 ;
        RECT 269.400 365.400 270.600 367.650 ;
        RECT 293.400 365.400 294.600 367.650 ;
        RECT 269.400 361.050 270.450 365.400 ;
        RECT 293.400 361.050 294.450 365.400 ;
        RECT 253.950 358.950 256.050 361.050 ;
        RECT 268.950 358.950 271.050 361.050 ;
        RECT 292.950 358.950 295.050 361.050 ;
        RECT 293.400 346.050 294.450 358.950 ;
        RECT 292.950 343.950 295.050 346.050 ;
        RECT 325.950 343.950 328.050 346.050 ;
        RECT 326.400 339.600 327.450 343.950 ;
        RECT 326.400 337.350 327.600 339.600 ;
      LAYER metal3 ;
        RECT 262.950 450.750 265.050 451.200 ;
        RECT 283.950 450.750 286.050 451.200 ;
        RECT 262.950 449.550 286.050 450.750 ;
        RECT 262.950 449.100 265.050 449.550 ;
        RECT 283.950 449.100 286.050 449.550 ;
        RECT 319.950 450.750 322.050 451.200 ;
        RECT 325.950 450.750 328.050 451.200 ;
        RECT 319.950 449.550 328.050 450.750 ;
        RECT 319.950 449.100 322.050 449.550 ;
        RECT 325.950 449.100 328.050 449.550 ;
        RECT 1.950 444.600 4.050 445.050 ;
        RECT -3.600 443.400 4.050 444.600 ;
        RECT 1.950 442.950 4.050 443.400 ;
        RECT 283.950 444.600 286.050 445.050 ;
        RECT 289.950 444.600 292.050 444.900 ;
        RECT 283.950 443.400 292.050 444.600 ;
        RECT 283.950 442.950 286.050 443.400 ;
        RECT 289.950 442.800 292.050 443.400 ;
        RECT 199.950 435.600 202.050 436.050 ;
        RECT 217.950 435.600 220.050 436.050 ;
        RECT 226.950 435.600 229.050 436.050 ;
        RECT 289.950 435.600 292.050 436.050 ;
        RECT 199.950 434.400 292.050 435.600 ;
        RECT 199.950 433.950 202.050 434.400 ;
        RECT 217.950 433.950 220.050 434.400 ;
        RECT 226.950 433.950 229.050 434.400 ;
        RECT 289.950 433.950 292.050 434.400 ;
        RECT 1.950 429.600 4.050 430.050 ;
        RECT 199.950 429.600 202.050 430.050 ;
        RECT 1.950 428.400 202.050 429.600 ;
        RECT 1.950 427.950 4.050 428.400 ;
        RECT 199.950 427.950 202.050 428.400 ;
        RECT 289.950 423.600 292.050 424.050 ;
        RECT 319.950 423.600 322.050 424.050 ;
        RECT 325.950 423.600 328.050 424.050 ;
        RECT 289.950 422.400 328.050 423.600 ;
        RECT 289.950 421.950 292.050 422.400 ;
        RECT 319.950 421.950 322.050 422.400 ;
        RECT 325.950 421.950 328.050 422.400 ;
        RECT 217.950 384.600 220.050 385.050 ;
        RECT 247.950 384.600 250.050 385.050 ;
        RECT 253.950 384.600 256.050 385.050 ;
        RECT 217.950 383.400 256.050 384.600 ;
        RECT 217.950 382.950 220.050 383.400 ;
        RECT 247.950 382.950 250.050 383.400 ;
        RECT 253.950 382.950 256.050 383.400 ;
        RECT 253.950 360.600 256.050 361.050 ;
        RECT 268.950 360.600 271.050 361.050 ;
        RECT 292.950 360.600 295.050 361.050 ;
        RECT 253.950 359.400 295.050 360.600 ;
        RECT 253.950 358.950 256.050 359.400 ;
        RECT 268.950 358.950 271.050 359.400 ;
        RECT 292.950 358.950 295.050 359.400 ;
        RECT 292.950 345.600 295.050 346.050 ;
        RECT 325.950 345.600 328.050 346.050 ;
        RECT 292.950 344.400 328.050 345.600 ;
        RECT 292.950 343.950 295.050 344.400 ;
        RECT 325.950 343.950 328.050 344.400 ;
    END
  END Cin[5]
  PIN Cin[4]
    PORT
      LAYER metal1 ;
        RECT 496.950 450.450 499.050 451.050 ;
        RECT 491.550 450.000 499.050 450.450 ;
        RECT 490.950 449.550 499.050 450.000 ;
        RECT 490.950 445.800 493.050 449.550 ;
        RECT 496.950 448.950 499.050 449.550 ;
      LAYER metal2 ;
        RECT 397.950 610.950 400.050 613.050 ;
        RECT 412.950 610.950 415.050 613.050 ;
        RECT 475.950 610.950 478.050 613.050 ;
        RECT 368.400 567.900 369.600 568.650 ;
        RECT 398.400 567.900 399.450 610.950 ;
        RECT 413.400 606.600 414.450 610.950 ;
        RECT 476.400 607.200 477.450 610.950 ;
        RECT 413.400 604.350 414.600 606.600 ;
        RECT 475.950 605.100 478.050 607.200 ;
        RECT 484.950 605.100 487.050 607.200 ;
        RECT 476.400 604.350 477.600 605.100 ;
        RECT 367.950 565.800 370.050 567.900 ;
        RECT 397.950 565.800 400.050 567.900 ;
        RECT 485.400 532.050 486.450 605.100 ;
        RECT 484.950 531.450 487.050 532.050 ;
        RECT 482.400 530.400 487.050 531.450 ;
        RECT 482.400 502.050 483.450 530.400 ;
        RECT 484.950 529.950 487.050 530.400 ;
        RECT 583.950 528.000 586.050 532.050 ;
        RECT 584.400 526.350 585.600 528.000 ;
        RECT 481.950 499.950 484.050 502.050 ;
        RECT 496.950 499.950 499.050 502.050 ;
        RECT 497.400 451.050 498.450 499.950 ;
        RECT 496.950 448.950 499.050 451.050 ;
        RECT 490.950 445.800 493.050 447.900 ;
        RECT 491.400 426.450 492.450 445.800 ;
        RECT 491.400 425.400 495.450 426.450 ;
        RECT 494.400 385.050 495.450 425.400 ;
        RECT 493.950 382.950 496.050 385.050 ;
        RECT 559.950 382.950 562.050 385.050 ;
        RECT 560.400 340.050 561.450 382.950 ;
        RECT 559.800 337.950 561.900 340.050 ;
        RECT 599.400 333.900 600.600 334.650 ;
        RECT 598.950 331.800 601.050 333.900 ;
        RECT 599.400 295.050 600.450 331.800 ;
        RECT 598.950 292.950 601.050 295.050 ;
        RECT 604.950 292.950 607.050 295.050 ;
        RECT 605.400 261.450 606.450 292.950 ;
        RECT 602.400 260.400 606.450 261.450 ;
        RECT 368.400 255.900 369.600 256.650 ;
        RECT 367.950 253.800 370.050 255.900 ;
        RECT 421.950 253.800 424.050 255.900 ;
        RECT 545.400 254.400 546.600 256.650 ;
        RECT 368.400 223.050 369.450 253.800 ;
        RECT 422.400 244.050 423.450 253.800 ;
        RECT 545.400 247.050 546.450 254.400 ;
        RECT 602.400 247.050 603.450 260.400 ;
        RECT 544.950 244.950 547.050 247.050 ;
        RECT 601.950 244.950 604.050 247.050 ;
        RECT 421.950 241.950 424.050 244.050 ;
        RECT 331.950 220.950 334.050 223.050 ;
        RECT 367.950 220.950 370.050 223.050 ;
        RECT 332.400 177.450 333.450 220.950 ;
        RECT 335.400 177.450 336.600 178.650 ;
        RECT 332.400 176.400 336.600 177.450 ;
        RECT 335.400 142.050 336.450 176.400 ;
        RECT 334.950 139.950 337.050 142.050 ;
        RECT 355.950 139.950 358.050 142.050 ;
        RECT 356.400 64.050 357.450 139.950 ;
        RECT 355.950 61.950 358.050 64.050 ;
        RECT 361.950 61.950 364.050 64.050 ;
        RECT 362.400 37.050 363.450 61.950 ;
        RECT 331.950 34.950 334.050 37.050 ;
        RECT 361.950 34.950 364.050 37.050 ;
        RECT 332.400 -3.600 333.450 34.950 ;
      LAYER via2 ;
        RECT 583.950 529.950 586.050 532.050 ;
      LAYER metal3 ;
        RECT 397.950 612.600 400.050 613.050 ;
        RECT 412.950 612.600 415.050 613.050 ;
        RECT 475.950 612.600 478.050 613.050 ;
        RECT 397.950 611.400 478.050 612.600 ;
        RECT 397.950 610.950 400.050 611.400 ;
        RECT 412.950 610.950 415.050 611.400 ;
        RECT 475.950 610.950 478.050 611.400 ;
        RECT 475.950 606.750 478.050 607.200 ;
        RECT 484.950 606.750 487.050 607.200 ;
        RECT 475.950 605.550 487.050 606.750 ;
        RECT 475.950 605.100 478.050 605.550 ;
        RECT 484.950 605.100 487.050 605.550 ;
        RECT 367.950 567.450 370.050 567.900 ;
        RECT 397.950 567.450 400.050 567.900 ;
        RECT 367.950 566.250 400.050 567.450 ;
        RECT 367.950 565.800 370.050 566.250 ;
        RECT 397.950 565.800 400.050 566.250 ;
        RECT 484.950 531.600 487.050 532.050 ;
        RECT 583.950 531.600 586.050 532.050 ;
        RECT 484.950 530.400 586.050 531.600 ;
        RECT 484.950 529.950 487.050 530.400 ;
        RECT 583.950 529.950 586.050 530.400 ;
        RECT 481.950 501.600 484.050 502.050 ;
        RECT 496.950 501.600 499.050 502.050 ;
        RECT 481.950 500.400 499.050 501.600 ;
        RECT 481.950 499.950 484.050 500.400 ;
        RECT 496.950 499.950 499.050 500.400 ;
        RECT 493.950 384.600 496.050 385.050 ;
        RECT 559.950 384.600 562.050 385.050 ;
        RECT 493.950 383.400 562.050 384.600 ;
        RECT 493.950 382.950 496.050 383.400 ;
        RECT 559.950 382.950 562.050 383.400 ;
        RECT 559.800 339.000 561.900 340.050 ;
        RECT 559.800 337.950 562.050 339.000 ;
        RECT 559.950 336.600 562.050 337.950 ;
        RECT 559.950 336.000 600.600 336.600 ;
        RECT 560.400 335.400 600.600 336.000 ;
        RECT 599.400 333.900 600.600 335.400 ;
        RECT 598.950 331.800 601.050 333.900 ;
        RECT 598.950 294.600 601.050 295.050 ;
        RECT 604.950 294.600 607.050 295.050 ;
        RECT 598.950 293.400 607.050 294.600 ;
        RECT 598.950 292.950 601.050 293.400 ;
        RECT 604.950 292.950 607.050 293.400 ;
        RECT 367.950 255.450 370.050 255.900 ;
        RECT 421.950 255.450 424.050 255.900 ;
        RECT 367.950 254.250 424.050 255.450 ;
        RECT 367.950 253.800 370.050 254.250 ;
        RECT 421.950 253.800 424.050 254.250 ;
        RECT 544.950 246.600 547.050 247.050 ;
        RECT 601.950 246.600 604.050 247.050 ;
        RECT 506.400 245.400 604.050 246.600 ;
        RECT 421.950 243.600 424.050 244.050 ;
        RECT 506.400 243.600 507.600 245.400 ;
        RECT 544.950 244.950 547.050 245.400 ;
        RECT 601.950 244.950 604.050 245.400 ;
        RECT 421.950 242.400 507.600 243.600 ;
        RECT 421.950 241.950 424.050 242.400 ;
        RECT 331.950 222.600 334.050 223.050 ;
        RECT 367.950 222.600 370.050 223.050 ;
        RECT 331.950 221.400 370.050 222.600 ;
        RECT 331.950 220.950 334.050 221.400 ;
        RECT 367.950 220.950 370.050 221.400 ;
        RECT 334.950 141.600 337.050 142.050 ;
        RECT 355.950 141.600 358.050 142.050 ;
        RECT 334.950 140.400 358.050 141.600 ;
        RECT 334.950 139.950 337.050 140.400 ;
        RECT 355.950 139.950 358.050 140.400 ;
        RECT 355.950 63.600 358.050 64.050 ;
        RECT 361.950 63.600 364.050 64.050 ;
        RECT 355.950 62.400 364.050 63.600 ;
        RECT 355.950 61.950 358.050 62.400 ;
        RECT 361.950 61.950 364.050 62.400 ;
        RECT 331.950 36.600 334.050 37.050 ;
        RECT 361.950 36.600 364.050 37.050 ;
        RECT 331.950 35.400 364.050 36.600 ;
        RECT 331.950 34.950 334.050 35.400 ;
        RECT 361.950 34.950 364.050 35.400 ;
    END
  END Cin[4]
  PIN Cin[3]
    PORT
      LAYER metal1 ;
        RECT 490.950 267.450 493.050 268.050 ;
        RECT 496.950 267.450 499.050 267.900 ;
        RECT 490.950 266.550 499.050 267.450 ;
        RECT 490.950 265.950 493.050 266.550 ;
        RECT 496.950 265.800 499.050 266.550 ;
      LAYER metal2 ;
        RECT 460.950 650.100 463.050 652.200 ;
        RECT 469.950 650.100 472.050 652.200 ;
        RECT 461.400 649.350 462.600 650.100 ;
        RECT 317.400 645.000 318.600 646.650 ;
        RECT 316.950 642.450 319.050 645.000 ;
        RECT 314.400 641.400 319.050 642.450 ;
        RECT 314.400 583.050 315.450 641.400 ;
        RECT 316.950 640.950 319.050 641.400 ;
        RECT 361.950 640.950 364.050 643.050 ;
        RECT 362.400 622.050 363.450 640.950 ;
        RECT 470.400 628.050 471.450 650.100 ;
        RECT 530.400 644.400 531.600 646.650 ;
        RECT 530.400 628.050 531.450 644.400 ;
        RECT 469.950 625.950 472.050 628.050 ;
        RECT 499.950 625.950 502.050 628.050 ;
        RECT 529.950 625.950 532.050 628.050 ;
        RECT 598.950 625.950 601.050 628.050 ;
        RECT 470.400 622.050 471.450 625.950 ;
        RECT 361.950 619.950 364.050 622.050 ;
        RECT 469.950 619.950 472.050 622.050 ;
        RECT 362.400 606.600 363.450 619.950 ;
        RECT 362.400 604.350 363.600 606.600 ;
        RECT 295.950 580.950 298.050 583.050 ;
        RECT 313.950 580.950 316.050 583.050 ;
        RECT 296.400 573.600 297.450 580.950 ;
        RECT 500.400 576.450 501.450 625.950 ;
        RECT 497.400 575.400 501.450 576.450 ;
        RECT 497.400 573.600 498.450 575.400 ;
        RECT 296.400 571.350 297.600 573.600 ;
        RECT 497.400 571.350 498.600 573.600 ;
        RECT 599.400 565.050 600.450 625.950 ;
        RECT 650.400 566.400 651.600 568.650 ;
        RECT 650.400 565.050 651.450 566.400 ;
        RECT 598.950 562.950 601.050 565.050 ;
        RECT 649.950 562.950 652.050 565.050 ;
        RECT 650.400 550.050 651.450 562.950 ;
        RECT 649.950 547.950 652.050 550.050 ;
        RECT 685.950 547.950 688.050 550.050 ;
        RECT 686.400 514.050 687.450 547.950 ;
        RECT 685.950 511.950 688.050 514.050 ;
        RECT 683.400 489.450 684.600 490.650 ;
        RECT 686.400 489.450 687.450 511.950 ;
        RECT 683.400 488.400 687.450 489.450 ;
        RECT 686.400 376.050 687.450 488.400 ;
        RECT 670.950 373.950 673.050 376.050 ;
        RECT 685.950 373.950 688.050 376.050 ;
        RECT 671.400 343.050 672.450 373.950 ;
        RECT 658.950 340.950 661.050 343.050 ;
        RECT 670.950 340.950 673.050 343.050 ;
        RECT 659.400 333.900 660.450 340.950 ;
        RECT 677.400 333.900 678.600 334.650 ;
        RECT 658.950 331.800 661.050 333.900 ;
        RECT 676.950 331.800 679.050 333.900 ;
        RECT 659.400 298.050 660.450 331.800 ;
        RECT 652.950 295.950 655.050 298.050 ;
        RECT 658.950 295.950 661.050 298.050 ;
        RECT 445.950 293.100 448.050 295.200 ;
        RECT 446.400 292.350 447.600 293.100 ;
        RECT 415.950 289.950 418.050 292.050 ;
        RECT 356.400 254.400 357.600 256.650 ;
        RECT 356.400 250.050 357.450 254.400 ;
        RECT 416.400 253.050 417.450 289.950 ;
        RECT 490.950 286.950 493.050 289.050 ;
        RECT 491.400 268.050 492.450 286.950 ;
        RECT 653.400 268.050 654.450 295.950 ;
        RECT 659.400 294.600 660.450 295.950 ;
        RECT 659.400 292.350 660.600 294.600 ;
        RECT 490.950 265.950 493.050 268.050 ;
        RECT 498.000 267.900 501.000 268.050 ;
        RECT 496.950 265.950 502.050 267.900 ;
        RECT 532.950 265.950 535.050 268.050 ;
        RECT 598.950 265.950 601.050 268.050 ;
        RECT 652.950 265.950 655.050 268.050 ;
        RECT 496.950 265.800 499.050 265.950 ;
        RECT 499.950 265.800 502.050 265.950 ;
        RECT 533.400 259.050 534.450 265.950 ;
        RECT 599.400 259.050 600.450 265.950 ;
        RECT 532.950 256.950 535.050 259.050 ;
        RECT 598.950 256.950 601.050 259.050 ;
        RECT 527.400 255.000 528.600 256.650 ;
        RECT 415.950 250.950 418.050 253.050 ;
        RECT 526.950 250.950 529.050 255.000 ;
        RECT 533.400 253.050 534.450 256.950 ;
        RECT 532.950 250.950 535.050 253.050 ;
        RECT 355.950 247.950 358.050 250.050 ;
      LAYER metal3 ;
        RECT 460.950 651.750 463.050 652.200 ;
        RECT 469.950 651.750 472.050 652.200 ;
        RECT 460.950 650.550 472.050 651.750 ;
        RECT 460.950 650.100 463.050 650.550 ;
        RECT 469.950 650.100 472.050 650.550 ;
        RECT 316.950 642.600 319.050 643.050 ;
        RECT 361.950 642.600 364.050 643.050 ;
        RECT 316.950 641.400 364.050 642.600 ;
        RECT 316.950 640.950 319.050 641.400 ;
        RECT 361.950 640.950 364.050 641.400 ;
        RECT 469.950 627.600 472.050 628.050 ;
        RECT 499.950 627.600 502.050 628.050 ;
        RECT 529.950 627.600 532.050 628.050 ;
        RECT 598.950 627.600 601.050 628.050 ;
        RECT 469.950 626.400 601.050 627.600 ;
        RECT 469.950 625.950 472.050 626.400 ;
        RECT 499.950 625.950 502.050 626.400 ;
        RECT 529.950 625.950 532.050 626.400 ;
        RECT 598.950 625.950 601.050 626.400 ;
        RECT 361.950 621.600 364.050 622.050 ;
        RECT 469.950 621.600 472.050 622.050 ;
        RECT 361.950 620.400 472.050 621.600 ;
        RECT 361.950 619.950 364.050 620.400 ;
        RECT 469.950 619.950 472.050 620.400 ;
        RECT 295.950 582.600 298.050 583.050 ;
        RECT 313.950 582.600 316.050 583.050 ;
        RECT 295.950 581.400 316.050 582.600 ;
        RECT 295.950 580.950 298.050 581.400 ;
        RECT 313.950 580.950 316.050 581.400 ;
        RECT 598.950 564.600 601.050 565.050 ;
        RECT 649.950 564.600 652.050 565.050 ;
        RECT 598.950 563.400 652.050 564.600 ;
        RECT 598.950 562.950 601.050 563.400 ;
        RECT 649.950 562.950 652.050 563.400 ;
        RECT 649.950 549.600 652.050 550.050 ;
        RECT 685.950 549.600 688.050 550.050 ;
        RECT 649.950 548.400 688.050 549.600 ;
        RECT 649.950 547.950 652.050 548.400 ;
        RECT 685.950 547.950 688.050 548.400 ;
        RECT 905.400 516.600 906.600 528.600 ;
        RECT 848.400 515.400 906.600 516.600 ;
        RECT 685.950 513.600 688.050 514.050 ;
        RECT 848.400 513.600 849.600 515.400 ;
        RECT 685.950 512.400 849.600 513.600 ;
        RECT 685.950 511.950 688.050 512.400 ;
        RECT 670.950 375.600 673.050 376.050 ;
        RECT 685.950 375.600 688.050 376.050 ;
        RECT 670.950 374.400 688.050 375.600 ;
        RECT 670.950 373.950 673.050 374.400 ;
        RECT 685.950 373.950 688.050 374.400 ;
        RECT 658.950 342.600 661.050 343.050 ;
        RECT 670.950 342.600 673.050 343.050 ;
        RECT 658.950 341.400 673.050 342.600 ;
        RECT 658.950 340.950 661.050 341.400 ;
        RECT 670.950 340.950 673.050 341.400 ;
        RECT 658.950 333.450 661.050 333.900 ;
        RECT 676.950 333.450 679.050 333.900 ;
        RECT 658.950 332.250 679.050 333.450 ;
        RECT 658.950 331.800 661.050 332.250 ;
        RECT 676.950 331.800 679.050 332.250 ;
        RECT 652.950 297.600 655.050 298.050 ;
        RECT 658.950 297.600 661.050 298.050 ;
        RECT 652.950 296.400 661.050 297.600 ;
        RECT 652.950 295.950 655.050 296.400 ;
        RECT 658.950 295.950 661.050 296.400 ;
        RECT 445.950 293.100 448.050 295.200 ;
        RECT 415.950 291.600 418.050 292.050 ;
        RECT 446.400 291.600 447.600 293.100 ;
        RECT 415.950 290.400 447.600 291.600 ;
        RECT 415.950 289.950 418.050 290.400 ;
        RECT 446.400 288.600 447.600 290.400 ;
        RECT 490.950 288.600 493.050 289.050 ;
        RECT 446.400 287.400 493.050 288.600 ;
        RECT 490.950 286.950 493.050 287.400 ;
        RECT 499.950 267.600 502.050 267.900 ;
        RECT 532.950 267.600 535.050 268.050 ;
        RECT 499.950 266.400 535.050 267.600 ;
        RECT 499.950 265.800 502.050 266.400 ;
        RECT 532.950 265.950 535.050 266.400 ;
        RECT 598.950 267.600 601.050 268.050 ;
        RECT 652.950 267.600 655.050 268.050 ;
        RECT 598.950 266.400 655.050 267.600 ;
        RECT 598.950 265.950 601.050 266.400 ;
        RECT 652.950 265.950 655.050 266.400 ;
        RECT 532.950 258.600 535.050 259.050 ;
        RECT 598.950 258.600 601.050 259.050 ;
        RECT 532.950 257.400 601.050 258.600 ;
        RECT 532.950 256.950 535.050 257.400 ;
        RECT 598.950 256.950 601.050 257.400 ;
        RECT 415.950 252.600 418.050 253.050 ;
        RECT 371.400 251.400 418.050 252.600 ;
        RECT 355.950 249.600 358.050 250.050 ;
        RECT 371.400 249.600 372.600 251.400 ;
        RECT 415.950 250.950 418.050 251.400 ;
        RECT 526.950 252.600 529.050 253.050 ;
        RECT 532.950 252.600 535.050 253.050 ;
        RECT 526.950 251.400 535.050 252.600 ;
        RECT 526.950 250.950 529.050 251.400 ;
        RECT 532.950 250.950 535.050 251.400 ;
        RECT 355.950 248.400 372.600 249.600 ;
        RECT 355.950 247.950 358.050 248.400 ;
    END
  END Cin[3]
  PIN Cin[2]
    PORT
      LAYER metal1 ;
        RECT 346.950 717.450 349.050 718.050 ;
        RECT 358.950 717.450 361.050 718.050 ;
        RECT 346.950 716.550 361.050 717.450 ;
        RECT 346.950 715.950 349.050 716.550 ;
        RECT 358.950 715.950 361.050 716.550 ;
        RECT 661.950 564.450 664.050 565.050 ;
        RECT 679.950 564.450 682.050 565.050 ;
        RECT 661.950 563.550 682.050 564.450 ;
        RECT 661.950 562.950 664.050 563.550 ;
        RECT 679.950 562.950 682.050 563.550 ;
        RECT 433.950 252.450 436.050 253.050 ;
        RECT 442.950 252.450 445.050 253.050 ;
        RECT 433.950 251.550 445.050 252.450 ;
        RECT 433.950 250.950 436.050 251.550 ;
        RECT 442.950 250.950 445.050 251.550 ;
      LAYER metal2 ;
        RECT 344.400 895.050 345.450 906.450 ;
        RECT 343.950 892.950 346.050 895.050 ;
        RECT 355.950 892.950 358.050 895.050 ;
        RECT 356.400 862.050 357.450 892.950 ;
        RECT 355.950 859.950 358.050 862.050 ;
        RECT 367.950 859.950 370.050 862.050 ;
        RECT 368.400 823.050 369.450 859.950 ;
        RECT 361.950 820.950 364.050 823.050 ;
        RECT 367.950 820.950 370.050 823.050 ;
        RECT 362.400 784.050 363.450 820.950 ;
        RECT 361.950 781.950 364.050 784.050 ;
        RECT 370.950 781.950 373.050 784.050 ;
        RECT 371.400 745.050 372.450 781.950 ;
        RECT 358.950 742.950 361.050 745.050 ;
        RECT 370.950 742.950 373.050 745.050 ;
        RECT 359.400 718.050 360.450 742.950 ;
        RECT 346.950 715.950 349.050 718.050 ;
        RECT 358.950 715.950 361.050 718.050 ;
        RECT 347.400 688.050 348.450 715.950 ;
        RECT 346.950 684.000 349.050 688.050 ;
        RECT 373.950 685.950 376.050 688.050 ;
        RECT 347.400 682.350 348.600 684.000 ;
        RECT 374.400 631.050 375.450 685.950 ;
        RECT 407.400 644.400 408.600 646.650 ;
        RECT 485.400 644.400 486.600 646.650 ;
        RECT 407.400 640.050 408.450 644.400 ;
        RECT 406.950 637.950 409.050 640.050 ;
        RECT 436.950 637.950 439.050 640.050 ;
        RECT 407.400 631.050 408.450 637.950 ;
        RECT 373.950 628.950 376.050 631.050 ;
        RECT 406.950 628.950 409.050 631.050 ;
        RECT 437.400 574.200 438.450 637.950 ;
        RECT 485.400 637.050 486.450 644.400 ;
        RECT 484.950 634.950 487.050 637.050 ;
        RECT 430.950 572.100 433.050 574.200 ;
        RECT 436.950 572.100 439.050 574.200 ;
        RECT 431.400 571.350 432.600 572.100 ;
        RECT 437.400 565.050 438.450 572.100 ;
        RECT 476.400 566.400 477.600 568.650 ;
        RECT 662.400 567.000 663.600 568.650 ;
        RECT 680.400 567.000 681.600 568.650 ;
        RECT 476.400 565.050 477.450 566.400 ;
        RECT 436.950 562.950 439.050 565.050 ;
        RECT 475.950 562.950 478.050 565.050 ;
        RECT 661.950 562.950 664.050 567.000 ;
        RECT 679.950 562.950 682.050 567.000 ;
        RECT 476.400 547.050 477.450 562.950 ;
        RECT 475.950 544.950 478.050 547.050 ;
        RECT 505.950 544.950 508.050 547.050 ;
        RECT 506.400 516.450 507.450 544.950 ;
        RECT 547.950 541.950 550.050 544.050 ;
        RECT 586.950 541.950 589.050 544.050 ;
        RECT 503.400 515.400 507.450 516.450 ;
        RECT 503.400 478.050 504.450 515.400 ;
        RECT 548.400 495.450 549.450 541.950 ;
        RECT 587.400 535.050 588.450 541.950 ;
        RECT 662.400 535.050 663.450 562.950 ;
        RECT 586.950 532.950 589.050 535.050 ;
        RECT 646.950 532.950 649.050 535.050 ;
        RECT 661.950 532.950 664.050 535.050 ;
        RECT 647.400 528.600 648.450 532.950 ;
        RECT 647.400 526.350 648.600 528.600 ;
        RECT 548.400 494.400 552.450 495.450 ;
        RECT 509.400 488.400 510.600 490.650 ;
        RECT 509.400 478.050 510.450 488.400 ;
        RECT 551.400 478.050 552.450 494.400 ;
        RECT 502.950 475.950 505.050 478.050 ;
        RECT 508.950 475.950 511.050 478.050 ;
        RECT 550.950 475.950 553.050 478.050 ;
        RECT 556.950 475.950 559.050 478.050 ;
        RECT 557.400 421.050 558.450 475.950 ;
        RECT 556.950 418.950 559.050 421.050 ;
        RECT 568.950 418.950 571.050 421.050 ;
        RECT 538.950 388.950 541.050 391.050 ;
        RECT 539.400 382.050 540.450 388.950 ;
        RECT 569.400 388.050 570.450 418.950 ;
        RECT 568.950 385.950 571.050 388.050 ;
        RECT 607.950 385.950 610.050 388.050 ;
        RECT 508.950 379.950 511.050 382.050 ;
        RECT 538.950 379.950 541.050 382.050 ;
        RECT 509.400 352.050 510.450 379.950 ;
        RECT 608.400 352.050 609.450 385.950 ;
        RECT 487.950 349.950 490.050 352.050 ;
        RECT 508.950 349.950 511.050 352.050 ;
        RECT 607.950 349.950 610.050 352.050 ;
        RECT 634.950 349.950 637.050 352.050 ;
        RECT 488.400 307.050 489.450 349.950 ;
        RECT 632.400 333.450 633.600 334.650 ;
        RECT 635.400 333.450 636.450 349.950 ;
        RECT 632.400 332.400 636.450 333.450 ;
        RECT 635.400 310.050 636.450 332.400 ;
        RECT 634.950 307.950 637.050 310.050 ;
        RECT 682.950 307.950 685.050 310.050 ;
        RECT 460.950 304.950 463.050 307.050 ;
        RECT 487.950 304.950 490.050 307.050 ;
        RECT 461.400 274.050 462.450 304.950 ;
        RECT 635.400 294.450 636.450 307.950 ;
        RECT 683.400 294.600 684.450 307.950 ;
        RECT 638.400 294.450 639.600 294.600 ;
        RECT 635.400 293.400 639.600 294.450 ;
        RECT 638.400 292.350 639.600 293.400 ;
        RECT 683.400 292.350 684.600 294.600 ;
        RECT 445.950 271.950 448.050 274.050 ;
        RECT 460.950 271.950 463.050 274.050 ;
        RECT 446.400 261.450 447.450 271.950 ;
        RECT 443.400 260.400 447.450 261.450 ;
        RECT 434.400 255.000 435.600 256.650 ;
        RECT 433.950 250.950 436.050 255.000 ;
        RECT 443.400 253.050 444.450 260.400 ;
        RECT 442.950 250.950 445.050 253.050 ;
      LAYER via2 ;
        RECT 346.950 685.950 349.050 688.050 ;
      LAYER metal3 ;
        RECT 343.950 894.600 346.050 895.050 ;
        RECT 355.950 894.600 358.050 895.050 ;
        RECT 343.950 893.400 358.050 894.600 ;
        RECT 343.950 892.950 346.050 893.400 ;
        RECT 355.950 892.950 358.050 893.400 ;
        RECT 355.950 861.600 358.050 862.050 ;
        RECT 367.950 861.600 370.050 862.050 ;
        RECT 355.950 860.400 370.050 861.600 ;
        RECT 355.950 859.950 358.050 860.400 ;
        RECT 367.950 859.950 370.050 860.400 ;
        RECT 361.950 822.600 364.050 823.050 ;
        RECT 367.950 822.600 370.050 823.050 ;
        RECT 361.950 821.400 370.050 822.600 ;
        RECT 361.950 820.950 364.050 821.400 ;
        RECT 367.950 820.950 370.050 821.400 ;
        RECT 361.950 783.600 364.050 784.050 ;
        RECT 370.950 783.600 373.050 784.050 ;
        RECT 361.950 782.400 373.050 783.600 ;
        RECT 361.950 781.950 364.050 782.400 ;
        RECT 370.950 781.950 373.050 782.400 ;
        RECT 358.950 744.600 361.050 745.050 ;
        RECT 370.950 744.600 373.050 745.050 ;
        RECT 358.950 743.400 373.050 744.600 ;
        RECT 358.950 742.950 361.050 743.400 ;
        RECT 370.950 742.950 373.050 743.400 ;
        RECT 346.950 687.600 349.050 688.050 ;
        RECT 373.950 687.600 376.050 688.050 ;
        RECT 346.950 686.400 376.050 687.600 ;
        RECT 346.950 685.950 349.050 686.400 ;
        RECT 373.950 685.950 376.050 686.400 ;
        RECT 406.950 639.600 409.050 640.050 ;
        RECT 436.950 639.600 439.050 640.050 ;
        RECT 406.950 638.400 439.050 639.600 ;
        RECT 406.950 637.950 409.050 638.400 ;
        RECT 436.950 637.950 439.050 638.400 ;
        RECT 437.400 636.600 438.600 637.950 ;
        RECT 484.950 636.600 487.050 637.050 ;
        RECT 437.400 635.400 487.050 636.600 ;
        RECT 484.950 634.950 487.050 635.400 ;
        RECT 373.950 630.600 376.050 631.050 ;
        RECT 406.950 630.600 409.050 631.050 ;
        RECT 373.950 629.400 409.050 630.600 ;
        RECT 373.950 628.950 376.050 629.400 ;
        RECT 406.950 628.950 409.050 629.400 ;
        RECT 430.950 573.750 433.050 574.200 ;
        RECT 436.950 573.750 439.050 574.200 ;
        RECT 430.950 572.550 439.050 573.750 ;
        RECT 430.950 572.100 433.050 572.550 ;
        RECT 436.950 572.100 439.050 572.550 ;
        RECT 436.950 564.600 439.050 565.050 ;
        RECT 475.950 564.600 478.050 565.050 ;
        RECT 436.950 563.400 478.050 564.600 ;
        RECT 436.950 562.950 439.050 563.400 ;
        RECT 475.950 562.950 478.050 563.400 ;
        RECT 475.950 546.600 478.050 547.050 ;
        RECT 505.950 546.600 508.050 547.050 ;
        RECT 475.950 545.400 508.050 546.600 ;
        RECT 475.950 544.950 478.050 545.400 ;
        RECT 505.950 544.950 508.050 545.400 ;
        RECT 547.950 543.600 550.050 544.050 ;
        RECT 586.950 543.600 589.050 544.050 ;
        RECT 547.950 542.400 589.050 543.600 ;
        RECT 547.950 541.950 550.050 542.400 ;
        RECT 586.950 541.950 589.050 542.400 ;
        RECT 586.950 534.600 589.050 535.050 ;
        RECT 646.950 534.600 649.050 535.050 ;
        RECT 661.950 534.600 664.050 535.050 ;
        RECT 586.950 533.400 664.050 534.600 ;
        RECT 586.950 532.950 589.050 533.400 ;
        RECT 646.950 532.950 649.050 533.400 ;
        RECT 661.950 532.950 664.050 533.400 ;
        RECT 502.950 477.600 505.050 478.050 ;
        RECT 508.950 477.600 511.050 478.050 ;
        RECT 550.950 477.600 553.050 478.050 ;
        RECT 556.950 477.600 559.050 478.050 ;
        RECT 502.950 476.400 559.050 477.600 ;
        RECT 502.950 475.950 505.050 476.400 ;
        RECT 508.950 475.950 511.050 476.400 ;
        RECT 550.950 475.950 553.050 476.400 ;
        RECT 556.950 475.950 559.050 476.400 ;
        RECT 556.950 420.600 559.050 421.050 ;
        RECT 568.950 420.600 571.050 421.050 ;
        RECT 556.950 419.400 571.050 420.600 ;
        RECT 556.950 418.950 559.050 419.400 ;
        RECT 568.950 418.950 571.050 419.400 ;
        RECT 538.950 390.600 541.050 391.050 ;
        RECT 538.950 389.400 570.600 390.600 ;
        RECT 538.950 388.950 541.050 389.400 ;
        RECT 569.400 388.050 570.600 389.400 ;
        RECT 568.950 387.600 571.050 388.050 ;
        RECT 607.950 387.600 610.050 388.050 ;
        RECT 568.950 386.400 610.050 387.600 ;
        RECT 568.950 385.950 571.050 386.400 ;
        RECT 607.950 385.950 610.050 386.400 ;
        RECT 508.950 381.600 511.050 382.050 ;
        RECT 538.950 381.600 541.050 382.050 ;
        RECT 508.950 380.400 541.050 381.600 ;
        RECT 508.950 379.950 511.050 380.400 ;
        RECT 538.950 379.950 541.050 380.400 ;
        RECT 487.950 351.600 490.050 352.050 ;
        RECT 508.950 351.600 511.050 352.050 ;
        RECT 487.950 350.400 511.050 351.600 ;
        RECT 487.950 349.950 490.050 350.400 ;
        RECT 508.950 349.950 511.050 350.400 ;
        RECT 607.950 351.600 610.050 352.050 ;
        RECT 634.950 351.600 637.050 352.050 ;
        RECT 607.950 350.400 637.050 351.600 ;
        RECT 607.950 349.950 610.050 350.400 ;
        RECT 634.950 349.950 637.050 350.400 ;
        RECT 634.950 309.600 637.050 310.050 ;
        RECT 682.950 309.600 685.050 310.050 ;
        RECT 634.950 308.400 685.050 309.600 ;
        RECT 634.950 307.950 637.050 308.400 ;
        RECT 682.950 307.950 685.050 308.400 ;
        RECT 460.950 306.600 463.050 307.050 ;
        RECT 487.950 306.600 490.050 307.050 ;
        RECT 460.950 305.400 490.050 306.600 ;
        RECT 460.950 304.950 463.050 305.400 ;
        RECT 487.950 304.950 490.050 305.400 ;
        RECT 445.950 273.600 448.050 274.050 ;
        RECT 460.950 273.600 463.050 274.050 ;
        RECT 445.950 272.400 463.050 273.600 ;
        RECT 445.950 271.950 448.050 272.400 ;
        RECT 460.950 271.950 463.050 272.400 ;
    END
  END Cin[2]
  PIN Cin[1]
    PORT
      LAYER metal1 ;
        RECT 790.950 363.450 793.050 364.050 ;
        RECT 799.950 363.450 802.050 364.050 ;
        RECT 790.950 362.550 802.050 363.450 ;
        RECT 790.950 361.950 793.050 362.550 ;
        RECT 799.950 361.950 802.050 362.550 ;
      LAYER metal2 ;
        RECT 395.400 801.450 396.600 802.650 ;
        RECT 395.400 800.400 399.450 801.450 ;
        RECT 398.400 796.050 399.450 800.400 ;
        RECT 692.400 800.400 693.600 802.650 ;
        RECT 773.400 800.400 774.600 802.650 ;
        RECT 397.950 793.950 400.050 796.050 ;
        RECT 415.950 793.950 418.050 796.050 ;
        RECT 175.950 790.950 178.050 793.050 ;
        RECT 226.950 790.950 229.050 793.050 ;
        RECT 292.950 790.950 295.050 793.050 ;
        RECT 364.950 790.950 367.050 793.050 ;
        RECT 176.400 787.050 177.450 790.950 ;
        RECT 133.950 784.950 136.050 787.050 ;
        RECT 175.950 784.950 178.050 787.050 ;
        RECT 128.400 723.900 129.600 724.650 ;
        RECT 134.400 723.900 135.450 784.950 ;
        RECT 227.400 775.050 228.450 790.950 ;
        RECT 293.400 775.050 294.450 790.950 ;
        RECT 226.950 772.950 229.050 775.050 ;
        RECT 292.950 772.950 295.050 775.050 ;
        RECT 365.400 769.050 366.450 790.950 ;
        RECT 398.400 769.050 399.450 793.950 ;
        RECT 416.400 775.050 417.450 793.950 ;
        RECT 692.400 793.050 693.450 800.400 ;
        RECT 773.400 793.050 774.450 800.400 ;
        RECT 691.950 790.950 694.050 793.050 ;
        RECT 772.950 790.950 775.050 793.050 ;
        RECT 692.400 781.050 693.450 790.950 ;
        RECT 691.950 778.950 694.050 781.050 ;
        RECT 415.950 772.950 418.050 775.050 ;
        RECT 364.950 766.950 367.050 769.050 ;
        RECT 397.950 766.950 400.050 769.050 ;
        RECT 773.400 748.050 774.450 790.950 ;
        RECT 760.950 745.950 763.050 748.050 ;
        RECT 772.950 745.950 775.050 748.050 ;
        RECT 127.950 721.800 130.050 723.900 ;
        RECT 133.950 721.800 136.050 723.900 ;
        RECT 128.400 694.050 129.450 721.800 ;
        RECT 761.400 703.050 762.450 745.950 ;
        RECT 718.950 700.950 721.050 703.050 ;
        RECT 760.950 700.950 763.050 703.050 ;
        RECT 70.950 691.950 73.050 694.050 ;
        RECT 76.950 691.950 79.050 694.050 ;
        RECT 127.950 691.950 130.050 694.050 ;
        RECT 71.400 684.600 72.450 691.950 ;
        RECT 71.400 682.350 72.600 684.600 ;
        RECT 77.400 651.450 78.450 691.950 ;
        RECT 719.400 676.050 720.450 700.950 ;
        RECT 718.950 673.950 721.050 676.050 ;
        RECT 727.950 673.950 730.050 676.050 ;
        RECT 74.400 650.400 78.450 651.450 ;
        RECT 74.400 616.050 75.450 650.400 ;
        RECT 728.400 637.050 729.450 673.950 ;
        RECT 721.950 634.950 724.050 637.050 ;
        RECT 727.950 634.950 730.050 637.050 ;
        RECT 73.950 613.950 76.050 616.050 ;
        RECT 82.950 613.950 85.050 616.050 ;
        RECT 83.400 592.050 84.450 613.950 ;
        RECT 82.950 589.950 85.050 592.050 ;
        RECT 94.950 589.950 97.050 592.050 ;
        RECT 95.400 508.050 96.450 589.950 ;
        RECT 722.400 556.050 723.450 634.950 ;
        RECT 721.950 553.950 724.050 556.050 ;
        RECT 781.950 553.950 784.050 556.050 ;
        RECT 94.950 505.950 97.050 508.050 ;
        RECT 178.950 505.950 181.050 508.050 ;
        RECT 179.400 450.600 180.450 505.950 ;
        RECT 782.400 484.050 783.450 553.950 ;
        RECT 775.950 481.950 778.050 484.050 ;
        RECT 781.950 481.950 784.050 484.050 ;
        RECT 179.400 448.350 180.600 450.600 ;
        RECT 776.400 439.050 777.450 481.950 ;
        RECT 775.950 436.950 778.050 439.050 ;
        RECT 784.950 436.950 787.050 439.050 ;
        RECT 785.400 406.050 786.450 436.950 ;
        RECT 784.950 403.950 787.050 406.050 ;
        RECT 790.950 403.950 793.050 406.050 ;
        RECT 791.400 364.050 792.450 403.950 ;
        RECT 790.950 361.950 793.050 364.050 ;
        RECT 799.950 361.950 802.050 364.050 ;
        RECT 800.400 316.050 801.450 361.950 ;
        RECT 815.400 332.400 816.600 334.650 ;
        RECT 815.400 316.050 816.450 332.400 ;
        RECT 799.950 313.950 802.050 316.050 ;
        RECT 814.950 313.950 817.050 316.050 ;
        RECT 853.950 313.950 856.050 316.050 ;
        RECT 889.950 313.950 892.050 316.050 ;
        RECT 854.400 294.600 855.450 313.950 ;
        RECT 890.400 301.050 891.450 313.950 ;
        RECT 889.950 298.950 892.050 301.050 ;
        RECT 854.400 292.350 855.600 294.600 ;
        RECT 886.950 292.950 889.050 295.050 ;
        RECT 887.400 292.350 888.600 292.950 ;
      LAYER metal3 ;
        RECT 397.950 795.600 400.050 796.050 ;
        RECT 415.950 795.600 418.050 796.050 ;
        RECT 397.950 794.400 418.050 795.600 ;
        RECT 397.950 793.950 400.050 794.400 ;
        RECT 415.950 793.950 418.050 794.400 ;
        RECT 175.950 792.600 178.050 793.050 ;
        RECT 226.950 792.600 229.050 793.050 ;
        RECT 175.950 791.400 229.050 792.600 ;
        RECT 175.950 790.950 178.050 791.400 ;
        RECT 226.950 790.950 229.050 791.400 ;
        RECT 292.950 792.600 295.050 793.050 ;
        RECT 364.950 792.600 367.050 793.050 ;
        RECT 292.950 791.400 367.050 792.600 ;
        RECT 292.950 790.950 295.050 791.400 ;
        RECT 364.950 790.950 367.050 791.400 ;
        RECT 691.950 792.600 694.050 793.050 ;
        RECT 772.950 792.600 775.050 793.050 ;
        RECT 691.950 791.400 775.050 792.600 ;
        RECT 691.950 790.950 694.050 791.400 ;
        RECT 772.950 790.950 775.050 791.400 ;
        RECT 133.950 786.600 136.050 787.050 ;
        RECT 175.950 786.600 178.050 787.050 ;
        RECT 133.950 785.400 178.050 786.600 ;
        RECT 133.950 784.950 136.050 785.400 ;
        RECT 175.950 784.950 178.050 785.400 ;
        RECT 691.950 780.600 694.050 781.050 ;
        RECT 611.400 779.400 694.050 780.600 ;
        RECT 611.400 777.600 612.600 779.400 ;
        RECT 691.950 778.950 694.050 779.400 ;
        RECT 434.400 776.400 612.600 777.600 ;
        RECT 226.950 774.600 229.050 775.050 ;
        RECT 292.950 774.600 295.050 775.050 ;
        RECT 226.950 773.400 295.050 774.600 ;
        RECT 226.950 772.950 229.050 773.400 ;
        RECT 292.950 772.950 295.050 773.400 ;
        RECT 415.950 774.600 418.050 775.050 ;
        RECT 434.400 774.600 435.600 776.400 ;
        RECT 415.950 773.400 435.600 774.600 ;
        RECT 415.950 772.950 418.050 773.400 ;
        RECT 364.950 768.600 367.050 769.050 ;
        RECT 397.950 768.600 400.050 769.050 ;
        RECT 364.950 767.400 400.050 768.600 ;
        RECT 364.950 766.950 367.050 767.400 ;
        RECT 397.950 766.950 400.050 767.400 ;
        RECT 760.950 747.600 763.050 748.050 ;
        RECT 772.950 747.600 775.050 748.050 ;
        RECT 760.950 746.400 775.050 747.600 ;
        RECT 760.950 745.950 763.050 746.400 ;
        RECT 772.950 745.950 775.050 746.400 ;
        RECT 127.950 723.450 130.050 723.900 ;
        RECT 133.950 723.450 136.050 723.900 ;
        RECT 127.950 722.250 136.050 723.450 ;
        RECT 127.950 721.800 130.050 722.250 ;
        RECT 133.950 721.800 136.050 722.250 ;
        RECT 718.950 702.600 721.050 703.050 ;
        RECT 760.950 702.600 763.050 703.050 ;
        RECT 718.950 701.400 763.050 702.600 ;
        RECT 718.950 700.950 721.050 701.400 ;
        RECT 760.950 700.950 763.050 701.400 ;
        RECT 70.950 693.600 73.050 694.050 ;
        RECT 76.950 693.600 79.050 694.050 ;
        RECT 127.950 693.600 130.050 694.050 ;
        RECT 70.950 692.400 130.050 693.600 ;
        RECT 70.950 691.950 73.050 692.400 ;
        RECT 76.950 691.950 79.050 692.400 ;
        RECT 127.950 691.950 130.050 692.400 ;
        RECT 718.950 675.600 721.050 676.050 ;
        RECT 727.950 675.600 730.050 676.050 ;
        RECT 718.950 674.400 730.050 675.600 ;
        RECT 718.950 673.950 721.050 674.400 ;
        RECT 727.950 673.950 730.050 674.400 ;
        RECT 721.950 636.600 724.050 637.050 ;
        RECT 727.950 636.600 730.050 637.050 ;
        RECT 721.950 635.400 730.050 636.600 ;
        RECT 721.950 634.950 724.050 635.400 ;
        RECT 727.950 634.950 730.050 635.400 ;
        RECT 73.950 615.600 76.050 616.050 ;
        RECT 82.950 615.600 85.050 616.050 ;
        RECT 73.950 614.400 85.050 615.600 ;
        RECT 73.950 613.950 76.050 614.400 ;
        RECT 82.950 613.950 85.050 614.400 ;
        RECT 82.950 591.600 85.050 592.050 ;
        RECT 94.950 591.600 97.050 592.050 ;
        RECT 82.950 590.400 97.050 591.600 ;
        RECT 82.950 589.950 85.050 590.400 ;
        RECT 94.950 589.950 97.050 590.400 ;
        RECT 721.950 555.600 724.050 556.050 ;
        RECT 781.950 555.600 784.050 556.050 ;
        RECT 721.950 554.400 784.050 555.600 ;
        RECT 721.950 553.950 724.050 554.400 ;
        RECT 781.950 553.950 784.050 554.400 ;
        RECT 94.950 507.600 97.050 508.050 ;
        RECT 178.950 507.600 181.050 508.050 ;
        RECT 94.950 506.400 181.050 507.600 ;
        RECT 94.950 505.950 97.050 506.400 ;
        RECT 178.950 505.950 181.050 506.400 ;
        RECT 775.950 483.600 778.050 484.050 ;
        RECT 781.950 483.600 784.050 484.050 ;
        RECT 775.950 482.400 784.050 483.600 ;
        RECT 775.950 481.950 778.050 482.400 ;
        RECT 781.950 481.950 784.050 482.400 ;
        RECT 775.950 438.600 778.050 439.050 ;
        RECT 784.950 438.600 787.050 439.050 ;
        RECT 775.950 437.400 787.050 438.600 ;
        RECT 775.950 436.950 778.050 437.400 ;
        RECT 784.950 436.950 787.050 437.400 ;
        RECT 784.950 405.600 787.050 406.050 ;
        RECT 790.950 405.600 793.050 406.050 ;
        RECT 784.950 404.400 793.050 405.600 ;
        RECT 784.950 403.950 787.050 404.400 ;
        RECT 790.950 403.950 793.050 404.400 ;
        RECT 799.950 315.600 802.050 316.050 ;
        RECT 814.950 315.600 817.050 316.050 ;
        RECT 853.950 315.600 856.050 316.050 ;
        RECT 889.950 315.600 892.050 316.050 ;
        RECT 799.950 314.400 892.050 315.600 ;
        RECT 799.950 313.950 802.050 314.400 ;
        RECT 814.950 313.950 817.050 314.400 ;
        RECT 853.950 313.950 856.050 314.400 ;
        RECT 889.950 313.950 892.050 314.400 ;
        RECT 889.950 300.600 894.000 301.050 ;
        RECT 889.950 298.950 894.600 300.600 ;
        RECT 893.400 297.600 894.600 298.950 ;
        RECT 893.400 296.400 906.600 297.600 ;
        RECT 886.950 294.600 889.050 295.050 ;
        RECT 905.400 294.600 906.600 296.400 ;
        RECT 886.950 293.400 906.600 294.600 ;
        RECT 886.950 292.950 889.050 293.400 ;
    END
  END Cin[1]
  PIN Cin[0]
    PORT
      LAYER metal1 ;
        RECT 700.950 720.450 703.050 721.050 ;
        RECT 706.950 720.450 709.050 721.050 ;
        RECT 700.950 719.550 709.050 720.450 ;
        RECT 700.950 718.950 703.050 719.550 ;
        RECT 706.950 718.950 709.050 719.550 ;
        RECT 694.950 684.450 697.050 685.050 ;
        RECT 700.950 684.450 703.050 685.050 ;
        RECT 694.950 683.550 703.050 684.450 ;
        RECT 694.950 682.950 697.050 683.550 ;
        RECT 700.950 682.950 703.050 683.550 ;
        RECT 694.950 678.450 697.050 679.050 ;
        RECT 700.950 678.450 703.050 679.050 ;
        RECT 694.950 677.550 703.050 678.450 ;
        RECT 694.950 676.950 697.050 677.550 ;
        RECT 700.950 676.950 703.050 677.550 ;
        RECT 694.950 645.450 697.050 646.050 ;
        RECT 700.950 645.450 703.050 646.050 ;
        RECT 694.950 644.550 703.050 645.450 ;
        RECT 694.950 643.950 697.050 644.550 ;
        RECT 700.950 643.950 703.050 644.550 ;
        RECT 712.950 363.450 715.050 364.050 ;
        RECT 718.950 363.450 721.050 364.050 ;
        RECT 712.950 362.550 721.050 363.450 ;
        RECT 712.950 361.950 715.050 362.550 ;
        RECT 718.950 361.950 721.050 362.550 ;
      LAYER metal2 ;
        RECT 478.950 895.950 481.050 898.050 ;
        RECT 484.950 895.950 487.050 898.050 ;
        RECT 766.950 895.950 769.050 898.050 ;
        RECT 479.400 885.600 480.450 895.950 ;
        RECT 479.400 883.350 480.600 885.600 ;
        RECT 482.400 807.450 483.600 807.600 ;
        RECT 485.400 807.450 486.450 895.950 ;
        RECT 767.400 885.450 768.450 895.950 ;
        RECT 770.400 885.450 771.600 885.600 ;
        RECT 767.400 884.400 771.600 885.450 ;
        RECT 767.400 844.050 768.450 884.400 ;
        RECT 770.400 883.350 771.600 884.400 ;
        RECT 742.950 841.950 745.050 844.050 ;
        RECT 766.950 841.950 769.050 844.050 ;
        RECT 482.400 806.400 486.450 807.450 ;
        RECT 482.400 805.350 483.600 806.400 ;
        RECT 743.400 790.050 744.450 841.950 ;
        RECT 703.950 787.950 706.050 790.050 ;
        RECT 742.950 787.950 745.050 790.050 ;
        RECT 704.400 756.450 705.450 787.950 ;
        RECT 704.400 755.400 708.450 756.450 ;
        RECT 707.400 721.050 708.450 755.400 ;
        RECT 700.950 718.950 703.050 721.050 ;
        RECT 706.950 718.950 709.050 721.050 ;
        RECT 701.400 685.050 702.450 718.950 ;
        RECT 694.950 682.950 697.050 685.050 ;
        RECT 700.950 682.950 703.050 685.050 ;
        RECT 695.400 679.050 696.450 682.950 ;
        RECT 694.950 676.950 697.050 679.050 ;
        RECT 700.950 676.950 703.050 679.050 ;
        RECT 701.400 646.050 702.450 676.950 ;
        RECT 694.950 643.950 697.050 646.050 ;
        RECT 700.950 643.950 703.050 646.050 ;
        RECT 695.400 550.050 696.450 643.950 ;
        RECT 694.950 547.950 697.050 550.050 ;
        RECT 700.950 547.950 703.050 550.050 ;
        RECT 701.400 517.050 702.450 547.950 ;
        RECT 700.950 514.950 703.050 517.050 ;
        RECT 712.950 514.950 715.050 517.050 ;
        RECT 713.400 489.450 714.450 514.950 ;
        RECT 710.400 488.400 714.450 489.450 ;
        RECT 710.400 409.050 711.450 488.400 ;
        RECT 709.950 406.950 712.050 409.050 ;
        RECT 718.950 406.950 721.050 409.050 ;
        RECT 719.400 364.050 720.450 406.950 ;
        RECT 712.950 361.950 715.050 364.050 ;
        RECT 718.950 361.950 721.050 364.050 ;
        RECT 713.400 328.050 714.450 361.950 ;
        RECT 712.950 325.950 715.050 328.050 ;
        RECT 721.950 325.950 724.050 328.050 ;
        RECT 722.400 265.050 723.450 325.950 ;
        RECT 721.950 262.950 724.050 265.050 ;
        RECT 736.950 259.950 739.050 262.050 ;
        RECT 737.400 247.050 738.450 259.950 ;
        RECT 736.950 244.950 739.050 247.050 ;
        RECT 784.950 244.950 787.050 247.050 ;
        RECT 785.400 232.050 786.450 244.950 ;
        RECT 784.950 229.950 787.050 232.050 ;
        RECT 889.950 229.950 892.050 232.050 ;
        RECT 890.400 169.050 891.450 229.950 ;
        RECT 877.950 166.950 880.050 169.050 ;
        RECT 889.950 166.950 892.050 169.050 ;
        RECT 878.400 127.050 879.450 166.950 ;
        RECT 877.950 124.950 880.050 127.050 ;
        RECT 886.950 124.950 889.050 127.050 ;
        RECT 887.400 28.200 888.450 124.950 ;
        RECT 886.950 26.100 889.050 28.200 ;
        RECT 887.400 25.350 888.600 26.100 ;
      LAYER metal3 ;
        RECT 478.950 897.600 481.050 898.050 ;
        RECT 484.950 897.600 487.050 898.050 ;
        RECT 766.950 897.600 769.050 898.050 ;
        RECT 478.950 896.400 769.050 897.600 ;
        RECT 478.950 895.950 481.050 896.400 ;
        RECT 484.950 895.950 487.050 896.400 ;
        RECT 766.950 895.950 769.050 896.400 ;
        RECT 742.950 843.600 745.050 844.050 ;
        RECT 766.950 843.600 769.050 844.050 ;
        RECT 742.950 842.400 769.050 843.600 ;
        RECT 742.950 841.950 745.050 842.400 ;
        RECT 766.950 841.950 769.050 842.400 ;
        RECT 703.950 789.600 706.050 790.050 ;
        RECT 742.950 789.600 745.050 790.050 ;
        RECT 703.950 788.400 745.050 789.600 ;
        RECT 703.950 787.950 706.050 788.400 ;
        RECT 742.950 787.950 745.050 788.400 ;
        RECT 694.950 549.600 697.050 550.050 ;
        RECT 700.950 549.600 703.050 550.050 ;
        RECT 694.950 548.400 703.050 549.600 ;
        RECT 694.950 547.950 697.050 548.400 ;
        RECT 700.950 547.950 703.050 548.400 ;
        RECT 700.950 516.600 703.050 517.050 ;
        RECT 712.950 516.600 715.050 517.050 ;
        RECT 700.950 515.400 715.050 516.600 ;
        RECT 700.950 514.950 703.050 515.400 ;
        RECT 712.950 514.950 715.050 515.400 ;
        RECT 709.950 408.600 712.050 409.050 ;
        RECT 718.950 408.600 721.050 409.050 ;
        RECT 709.950 407.400 721.050 408.600 ;
        RECT 709.950 406.950 712.050 407.400 ;
        RECT 718.950 406.950 721.050 407.400 ;
        RECT 712.950 327.600 715.050 328.050 ;
        RECT 721.950 327.600 724.050 328.050 ;
        RECT 712.950 326.400 724.050 327.600 ;
        RECT 712.950 325.950 715.050 326.400 ;
        RECT 721.950 325.950 724.050 326.400 ;
        RECT 721.950 261.600 724.050 265.050 ;
        RECT 736.950 261.600 739.050 262.050 ;
        RECT 721.950 261.000 739.050 261.600 ;
        RECT 722.400 260.400 739.050 261.000 ;
        RECT 736.950 259.950 739.050 260.400 ;
        RECT 736.950 246.600 739.050 247.050 ;
        RECT 784.950 246.600 787.050 247.050 ;
        RECT 736.950 245.400 787.050 246.600 ;
        RECT 736.950 244.950 739.050 245.400 ;
        RECT 784.950 244.950 787.050 245.400 ;
        RECT 784.950 231.600 787.050 232.050 ;
        RECT 889.950 231.600 892.050 232.050 ;
        RECT 784.950 230.400 892.050 231.600 ;
        RECT 784.950 229.950 787.050 230.400 ;
        RECT 889.950 229.950 892.050 230.400 ;
        RECT 877.950 168.600 880.050 169.050 ;
        RECT 889.950 168.600 892.050 169.050 ;
        RECT 877.950 167.400 892.050 168.600 ;
        RECT 877.950 166.950 880.050 167.400 ;
        RECT 889.950 166.950 892.050 167.400 ;
        RECT 877.950 126.600 880.050 127.050 ;
        RECT 886.950 126.600 889.050 127.050 ;
        RECT 877.950 125.400 889.050 126.600 ;
        RECT 877.950 124.950 880.050 125.400 ;
        RECT 886.950 124.950 889.050 125.400 ;
        RECT 886.950 27.600 889.050 28.200 ;
        RECT 886.950 26.400 906.600 27.600 ;
        RECT 886.950 26.100 889.050 26.400 ;
    END
  END Cin[0]
  PIN Xin[7]
    PORT
      LAYER metal1 ;
        RECT 112.950 375.450 115.050 376.050 ;
        RECT 118.950 375.450 121.050 376.050 ;
        RECT 112.950 374.550 121.050 375.450 ;
        RECT 112.950 373.950 115.050 374.550 ;
        RECT 118.950 373.950 121.050 374.550 ;
        RECT 880.950 141.450 883.050 142.050 ;
        RECT 886.950 141.450 889.050 142.050 ;
        RECT 880.950 140.550 889.050 141.450 ;
        RECT 880.950 139.950 883.050 140.550 ;
        RECT 886.950 139.950 889.050 140.550 ;
      LAYER metal2 ;
        RECT 850.950 416.100 853.050 418.200 ;
        RECT 859.950 416.100 862.050 418.200 ;
        RECT 86.400 411.000 87.600 412.650 ;
        RECT 85.950 406.950 88.050 411.000 ;
        RECT 851.400 409.050 852.450 416.100 ;
        RECT 860.400 415.350 861.600 416.100 ;
        RECT 112.950 406.950 115.050 409.050 ;
        RECT 850.950 406.950 853.050 409.050 ;
        RECT 859.950 406.950 862.050 409.050 ;
        RECT 113.400 376.050 114.450 406.950 ;
        RECT 112.950 372.000 115.050 376.050 ;
        RECT 118.950 373.950 121.050 376.050 ;
        RECT 113.400 370.350 114.600 372.000 ;
        RECT 119.400 352.050 120.450 373.950 ;
        RECT 118.950 349.950 121.050 352.050 ;
        RECT 139.950 349.950 142.050 352.050 ;
        RECT 140.400 277.050 141.450 349.950 ;
        RECT 860.400 343.050 861.450 406.950 ;
        RECT 844.950 340.950 847.050 343.050 ;
        RECT 845.400 304.050 846.450 340.950 ;
        RECT 859.950 339.000 862.050 343.050 ;
        RECT 883.950 339.000 886.050 343.050 ;
        RECT 895.950 340.950 898.050 343.050 ;
        RECT 860.400 337.350 861.600 339.000 ;
        RECT 884.400 337.350 885.600 339.000 ;
        RECT 896.400 307.050 897.450 340.950 ;
        RECT 895.950 304.950 898.050 307.050 ;
        RECT 436.950 301.950 439.050 304.050 ;
        RECT 844.950 301.950 847.050 304.050 ;
        RECT 139.950 274.950 142.050 277.050 ;
        RECT 160.950 274.950 163.050 277.050 ;
        RECT 161.400 262.200 162.450 274.950 ;
        RECT 437.400 274.050 438.450 301.950 ;
        RECT 845.400 288.900 846.450 301.950 ;
        RECT 857.400 288.900 858.600 289.650 ;
        RECT 844.950 286.800 847.050 288.900 ;
        RECT 856.950 286.800 859.050 288.900 ;
        RECT 884.400 287.400 885.600 289.650 ;
        RECT 845.400 283.050 846.450 286.800 ;
        RECT 884.400 283.050 885.450 287.400 ;
        RECT 844.950 280.950 847.050 283.050 ;
        RECT 883.950 282.450 886.050 283.050 ;
        RECT 883.950 281.400 888.450 282.450 ;
        RECT 883.950 280.950 886.050 281.400 ;
        RECT 349.950 271.950 352.050 274.050 ;
        RECT 358.950 271.950 361.050 274.050 ;
        RECT 436.950 271.950 439.050 274.050 ;
        RECT 160.950 260.100 163.050 262.200 ;
        RECT 169.950 260.100 172.050 262.200 ;
        RECT 161.400 244.050 162.450 260.100 ;
        RECT 170.400 259.350 171.600 260.100 ;
        RECT 160.950 241.950 163.050 244.050 ;
        RECT 350.400 241.050 351.450 271.950 ;
        RECT 359.400 261.600 360.450 271.950 ;
        RECT 437.400 262.200 438.450 271.950 ;
        RECT 359.400 259.350 360.600 261.600 ;
        RECT 427.950 260.100 430.050 262.200 ;
        RECT 436.950 260.100 439.050 262.200 ;
        RECT 428.400 259.350 429.600 260.100 ;
        RECT 349.950 238.950 352.050 241.050 ;
        RECT 350.400 184.200 351.450 238.950 ;
        RECT 340.950 182.100 343.050 184.200 ;
        RECT 349.950 182.100 352.050 184.200 ;
        RECT 341.400 181.350 342.600 182.100 ;
        RECT 887.400 142.050 888.450 281.400 ;
        RECT 880.950 139.950 883.050 142.050 ;
        RECT 886.950 139.950 889.050 142.050 ;
        RECT 881.400 106.050 882.450 139.950 ;
        RECT 880.950 103.950 883.050 106.050 ;
        RECT 889.950 103.950 892.050 106.050 ;
        RECT 839.400 20.400 840.600 22.650 ;
        RECT 839.400 10.050 840.450 20.400 ;
        RECT 890.400 10.050 891.450 103.950 ;
        RECT 838.950 7.950 841.050 10.050 ;
        RECT 889.950 7.950 892.050 10.050 ;
      LAYER via2 ;
        RECT 859.950 340.950 862.050 343.050 ;
        RECT 883.950 340.950 886.050 343.050 ;
      LAYER metal3 ;
        RECT 850.950 417.750 853.050 418.200 ;
        RECT 859.950 417.750 862.050 418.200 ;
        RECT 850.950 416.550 862.050 417.750 ;
        RECT 850.950 416.100 853.050 416.550 ;
        RECT 859.950 416.100 862.050 416.550 ;
        RECT 85.950 408.600 88.050 409.050 ;
        RECT 112.950 408.600 115.050 409.050 ;
        RECT 85.950 407.400 115.050 408.600 ;
        RECT 85.950 406.950 88.050 407.400 ;
        RECT 112.950 406.950 115.050 407.400 ;
        RECT 850.950 408.600 853.050 409.050 ;
        RECT 859.950 408.600 862.050 409.050 ;
        RECT 850.950 407.400 862.050 408.600 ;
        RECT 850.950 406.950 853.050 407.400 ;
        RECT 859.950 406.950 862.050 407.400 ;
        RECT 118.950 351.600 121.050 352.050 ;
        RECT 139.950 351.600 142.050 352.050 ;
        RECT 118.950 350.400 142.050 351.600 ;
        RECT 118.950 349.950 121.050 350.400 ;
        RECT 139.950 349.950 142.050 350.400 ;
        RECT 844.950 342.600 847.050 343.050 ;
        RECT 859.950 342.600 862.050 343.050 ;
        RECT 883.950 342.600 886.050 343.050 ;
        RECT 895.950 342.600 898.050 343.050 ;
        RECT 844.950 341.400 898.050 342.600 ;
        RECT 844.950 340.950 847.050 341.400 ;
        RECT 859.950 340.950 862.050 341.400 ;
        RECT 883.950 340.950 886.050 341.400 ;
        RECT 895.950 340.950 898.050 341.400 ;
        RECT 895.950 306.600 898.050 307.050 ;
        RECT 895.950 305.400 906.600 306.600 ;
        RECT 895.950 304.950 898.050 305.400 ;
        RECT 436.950 303.600 439.050 304.050 ;
        RECT 844.950 303.600 847.050 304.050 ;
        RECT 436.950 302.400 847.050 303.600 ;
        RECT 436.950 301.950 439.050 302.400 ;
        RECT 844.950 301.950 847.050 302.400 ;
        RECT 844.950 288.450 847.050 288.900 ;
        RECT 856.950 288.450 859.050 288.900 ;
        RECT 844.950 287.250 859.050 288.450 ;
        RECT 844.950 286.800 847.050 287.250 ;
        RECT 856.950 286.800 859.050 287.250 ;
        RECT 844.950 282.600 847.050 283.050 ;
        RECT 883.950 282.600 886.050 283.050 ;
        RECT 844.950 281.400 886.050 282.600 ;
        RECT 844.950 280.950 847.050 281.400 ;
        RECT 883.950 280.950 886.050 281.400 ;
        RECT 139.950 276.600 142.050 277.050 ;
        RECT 160.950 276.600 163.050 277.050 ;
        RECT 139.950 275.400 163.050 276.600 ;
        RECT 139.950 274.950 142.050 275.400 ;
        RECT 160.950 274.950 163.050 275.400 ;
        RECT 349.950 273.600 352.050 274.050 ;
        RECT 358.950 273.600 361.050 274.050 ;
        RECT 436.950 273.600 439.050 274.050 ;
        RECT 349.950 272.400 439.050 273.600 ;
        RECT 349.950 271.950 352.050 272.400 ;
        RECT 358.950 271.950 361.050 272.400 ;
        RECT 436.950 271.950 439.050 272.400 ;
        RECT 160.950 261.750 163.050 262.200 ;
        RECT 169.950 261.750 172.050 262.200 ;
        RECT 160.950 260.550 172.050 261.750 ;
        RECT 160.950 260.100 163.050 260.550 ;
        RECT 169.950 260.100 172.050 260.550 ;
        RECT 427.950 261.750 430.050 262.200 ;
        RECT 436.950 261.750 439.050 262.200 ;
        RECT 427.950 260.550 439.050 261.750 ;
        RECT 427.950 260.100 430.050 260.550 ;
        RECT 436.950 260.100 439.050 260.550 ;
        RECT 160.950 240.600 163.050 244.050 ;
        RECT 349.950 240.600 352.050 241.050 ;
        RECT 160.950 240.000 352.050 240.600 ;
        RECT 161.400 239.400 352.050 240.000 ;
        RECT 349.950 238.950 352.050 239.400 ;
        RECT 340.950 183.750 343.050 184.200 ;
        RECT 349.950 183.750 352.050 184.200 ;
        RECT 340.950 182.550 352.050 183.750 ;
        RECT 340.950 182.100 343.050 182.550 ;
        RECT 349.950 182.100 352.050 182.550 ;
        RECT 880.950 105.600 883.050 106.050 ;
        RECT 889.950 105.600 892.050 106.050 ;
        RECT 880.950 104.400 892.050 105.600 ;
        RECT 880.950 103.950 883.050 104.400 ;
        RECT 889.950 103.950 892.050 104.400 ;
        RECT 838.950 9.600 841.050 10.050 ;
        RECT 889.950 9.600 892.050 10.050 ;
        RECT 838.950 8.400 892.050 9.600 ;
        RECT 838.950 7.950 841.050 8.400 ;
        RECT 889.950 7.950 892.050 8.400 ;
    END
  END Xin[7]
  PIN Xin[6]
    PORT
      LAYER metal1 ;
        RECT 163.950 630.450 166.050 631.050 ;
        RECT 172.950 630.450 175.050 631.050 ;
        RECT 163.950 629.550 175.050 630.450 ;
        RECT 163.950 628.950 166.050 629.550 ;
        RECT 172.950 628.950 175.050 629.550 ;
        RECT 223.950 378.450 226.050 379.050 ;
        RECT 235.950 378.450 238.050 379.050 ;
        RECT 223.950 377.550 238.050 378.450 ;
        RECT 223.950 376.950 226.050 377.550 ;
        RECT 235.950 376.950 238.050 377.550 ;
      LAYER metal2 ;
        RECT 785.400 901.050 786.450 906.450 ;
        RECT 607.950 898.950 610.050 901.050 ;
        RECT 784.950 898.950 787.050 901.050 ;
        RECT 185.400 879.450 186.600 880.650 ;
        RECT 182.400 878.400 186.600 879.450 ;
        RECT 182.400 871.050 183.450 878.400 ;
        RECT 181.950 868.950 184.050 871.050 ;
        RECT 193.950 868.950 196.050 871.050 ;
        RECT 409.950 868.950 412.050 871.050 ;
        RECT 194.400 781.050 195.450 868.950 ;
        RECT 410.400 865.050 411.450 868.950 ;
        RECT 608.400 865.050 609.450 898.950 ;
        RECT 785.400 880.050 786.450 898.950 ;
        RECT 784.950 877.950 787.050 880.050 ;
        RECT 791.400 879.900 792.600 880.650 ;
        RECT 790.950 877.800 793.050 879.900 ;
        RECT 409.950 862.950 412.050 865.050 ;
        RECT 607.950 862.950 610.050 865.050 ;
        RECT 791.400 864.450 792.450 877.800 ;
        RECT 791.400 863.400 795.450 864.450 ;
        RECT 794.400 832.050 795.450 863.400 ;
        RECT 830.400 834.900 831.600 835.650 ;
        RECT 851.400 834.900 852.600 835.650 ;
        RECT 793.950 829.950 796.050 832.050 ;
        RECT 829.950 829.950 832.050 834.900 ;
        RECT 850.950 832.800 853.050 834.900 ;
        RECT 851.400 831.450 852.450 832.800 ;
        RECT 848.400 830.400 852.450 831.450 ;
        RECT 848.400 807.600 849.450 830.400 ;
        RECT 848.400 805.350 849.600 807.600 ;
        RECT 172.950 778.950 175.050 781.050 ;
        RECT 193.950 778.950 196.050 781.050 ;
        RECT 173.400 733.050 174.450 778.950 ;
        RECT 163.950 730.950 166.050 733.050 ;
        RECT 172.950 730.950 175.050 733.050 ;
        RECT 164.400 631.050 165.450 730.950 ;
        RECT 163.950 628.950 166.050 631.050 ;
        RECT 172.950 628.950 175.050 631.050 ;
        RECT 173.400 625.050 174.450 628.950 ;
        RECT 172.950 622.950 175.050 625.050 ;
        RECT 196.950 622.950 199.050 625.050 ;
        RECT 197.400 504.450 198.450 622.950 ;
        RECT 197.400 503.400 201.450 504.450 ;
        RECT 200.400 472.050 201.450 503.400 ;
        RECT 199.950 469.950 202.050 472.050 ;
        RECT 235.950 469.950 238.050 472.050 ;
        RECT 236.400 379.050 237.450 469.950 ;
        RECT 223.950 376.950 226.050 379.050 ;
        RECT 235.950 378.450 238.050 379.050 ;
        RECT 233.400 377.400 238.050 378.450 ;
        RECT 224.400 372.600 225.450 376.950 ;
        RECT 224.400 370.350 225.600 372.600 ;
        RECT 233.400 346.050 234.450 377.400 ;
        RECT 235.950 376.950 238.050 377.400 ;
        RECT 220.950 343.950 223.050 346.050 ;
        RECT 232.950 343.950 235.050 346.050 ;
        RECT 221.400 328.050 222.450 343.950 ;
        RECT 236.400 332.400 237.600 334.650 ;
        RECT 809.400 333.000 810.600 334.650 ;
        RECT 236.400 328.050 237.450 332.400 ;
        RECT 682.950 328.950 685.050 331.050 ;
        RECT 808.950 328.950 811.050 333.000 ;
        RECT 220.950 325.950 223.050 328.050 ;
        RECT 235.950 325.950 238.050 328.050 ;
        RECT 236.400 265.050 237.450 325.950 ;
        RECT 550.950 322.950 553.050 325.050 ;
        RECT 643.950 322.950 646.050 325.050 ;
        RECT 551.400 319.050 552.450 322.950 ;
        RECT 644.400 319.050 645.450 322.950 ;
        RECT 683.400 319.050 684.450 328.950 ;
        RECT 523.950 316.950 526.050 319.050 ;
        RECT 550.950 316.950 553.050 319.050 ;
        RECT 643.950 316.950 646.050 319.050 ;
        RECT 682.950 316.950 685.050 319.050 ;
        RECT 457.950 313.950 460.050 316.050 ;
        RECT 452.400 288.000 453.600 289.650 ;
        RECT 364.950 283.950 367.050 286.050 ;
        RECT 451.950 283.950 454.050 288.000 ;
        RECT 458.400 286.050 459.450 313.950 ;
        RECT 524.400 313.050 525.450 316.950 ;
        RECT 523.950 310.950 526.050 313.050 ;
        RECT 644.400 295.200 645.450 316.950 ;
        RECT 631.950 292.950 634.050 295.050 ;
        RECT 643.950 293.100 646.050 295.200 ;
        RECT 632.400 286.050 633.450 292.950 ;
        RECT 644.400 292.350 645.600 293.100 ;
        RECT 686.400 288.000 687.600 289.650 ;
        RECT 457.950 283.950 460.050 286.050 ;
        RECT 631.950 283.950 634.050 286.050 ;
        RECT 685.950 283.950 688.050 288.000 ;
        RECT 365.400 277.050 366.450 283.950 ;
        RECT 364.950 274.950 367.050 277.050 ;
        RECT 274.950 271.950 277.050 274.050 ;
        RECT 275.400 265.050 276.450 271.950 ;
        RECT 235.950 262.950 238.050 265.050 ;
        RECT 253.950 261.000 256.050 265.050 ;
        RECT 274.950 262.950 277.050 265.050 ;
        RECT 365.400 261.600 366.450 274.950 ;
        RECT 254.400 259.350 255.600 261.000 ;
        RECT 365.400 259.350 366.600 261.600 ;
      LAYER via2 ;
        RECT 829.950 832.800 832.050 834.900 ;
        RECT 253.950 262.950 256.050 265.050 ;
      LAYER metal3 ;
        RECT 607.950 900.600 610.050 901.050 ;
        RECT 784.950 900.600 787.050 901.050 ;
        RECT 607.950 899.400 787.050 900.600 ;
        RECT 607.950 898.950 610.050 899.400 ;
        RECT 784.950 898.950 787.050 899.400 ;
        RECT 784.950 879.600 787.050 880.050 ;
        RECT 790.950 879.600 793.050 879.900 ;
        RECT 784.950 878.400 793.050 879.600 ;
        RECT 784.950 877.950 787.050 878.400 ;
        RECT 790.950 877.800 793.050 878.400 ;
        RECT 181.950 870.600 184.050 871.050 ;
        RECT 193.950 870.600 196.050 871.050 ;
        RECT 409.950 870.600 412.050 871.050 ;
        RECT 181.950 869.400 412.050 870.600 ;
        RECT 181.950 868.950 184.050 869.400 ;
        RECT 193.950 868.950 196.050 869.400 ;
        RECT 409.950 868.950 412.050 869.400 ;
        RECT 409.950 864.600 412.050 865.050 ;
        RECT 607.950 864.600 610.050 865.050 ;
        RECT 409.950 863.400 610.050 864.600 ;
        RECT 409.950 862.950 412.050 863.400 ;
        RECT 607.950 862.950 610.050 863.400 ;
        RECT 829.950 834.600 832.050 834.900 ;
        RECT 850.950 834.600 853.050 834.900 ;
        RECT 829.950 833.400 853.050 834.600 ;
        RECT 829.950 832.800 832.050 833.400 ;
        RECT 850.950 832.800 853.050 833.400 ;
        RECT 793.950 831.600 796.050 832.050 ;
        RECT 829.950 831.600 832.050 832.050 ;
        RECT 793.950 830.400 832.050 831.600 ;
        RECT 793.950 829.950 796.050 830.400 ;
        RECT 829.950 829.950 832.050 830.400 ;
        RECT 172.950 780.600 175.050 781.050 ;
        RECT 193.950 780.600 196.050 781.050 ;
        RECT 172.950 779.400 196.050 780.600 ;
        RECT 172.950 778.950 175.050 779.400 ;
        RECT 193.950 778.950 196.050 779.400 ;
        RECT 163.950 732.600 166.050 733.050 ;
        RECT 172.950 732.600 175.050 733.050 ;
        RECT 163.950 731.400 175.050 732.600 ;
        RECT 163.950 730.950 166.050 731.400 ;
        RECT 172.950 730.950 175.050 731.400 ;
        RECT 172.950 624.600 175.050 625.050 ;
        RECT 196.950 624.600 199.050 625.050 ;
        RECT 172.950 623.400 199.050 624.600 ;
        RECT 172.950 622.950 175.050 623.400 ;
        RECT 196.950 622.950 199.050 623.400 ;
        RECT 199.950 471.600 202.050 472.050 ;
        RECT 235.950 471.600 238.050 472.050 ;
        RECT 199.950 470.400 238.050 471.600 ;
        RECT 199.950 469.950 202.050 470.400 ;
        RECT 235.950 469.950 238.050 470.400 ;
        RECT 220.950 345.600 223.050 346.050 ;
        RECT 232.950 345.600 235.050 346.050 ;
        RECT 220.950 344.400 235.050 345.600 ;
        RECT 220.950 343.950 223.050 344.400 ;
        RECT 232.950 343.950 235.050 344.400 ;
        RECT 682.950 330.600 685.050 331.050 ;
        RECT 808.950 330.600 811.050 331.050 ;
        RECT 682.950 329.400 811.050 330.600 ;
        RECT 682.950 328.950 685.050 329.400 ;
        RECT 808.950 328.950 811.050 329.400 ;
        RECT 220.950 327.600 223.050 328.050 ;
        RECT 235.950 327.600 238.050 328.050 ;
        RECT 220.950 326.400 238.050 327.600 ;
        RECT 220.950 325.950 223.050 326.400 ;
        RECT 235.950 325.950 238.050 326.400 ;
        RECT 550.950 324.600 553.050 325.050 ;
        RECT 643.950 324.600 646.050 325.050 ;
        RECT 550.950 323.400 646.050 324.600 ;
        RECT 550.950 322.950 553.050 323.400 ;
        RECT 643.950 322.950 646.050 323.400 ;
        RECT 523.950 318.600 526.050 319.050 ;
        RECT 550.950 318.600 553.050 319.050 ;
        RECT 523.950 317.400 553.050 318.600 ;
        RECT 523.950 316.950 526.050 317.400 ;
        RECT 550.950 316.950 553.050 317.400 ;
        RECT 643.950 318.600 646.050 319.050 ;
        RECT 682.950 318.600 685.050 319.050 ;
        RECT 643.950 317.400 685.050 318.600 ;
        RECT 643.950 316.950 646.050 317.400 ;
        RECT 682.950 316.950 685.050 317.400 ;
        RECT 457.950 315.600 460.050 316.050 ;
        RECT 457.950 314.400 504.600 315.600 ;
        RECT 457.950 313.950 460.050 314.400 ;
        RECT 503.400 312.600 504.600 314.400 ;
        RECT 523.950 312.600 526.050 313.050 ;
        RECT 503.400 311.400 526.050 312.600 ;
        RECT 523.950 310.950 526.050 311.400 ;
        RECT 631.950 294.600 634.050 295.050 ;
        RECT 643.950 294.600 646.050 295.200 ;
        RECT 631.950 293.400 646.050 294.600 ;
        RECT 631.950 292.950 634.050 293.400 ;
        RECT 643.950 293.100 646.050 293.400 ;
        RECT 364.950 285.600 367.050 286.050 ;
        RECT 451.950 285.600 454.050 286.050 ;
        RECT 457.950 285.600 460.050 286.050 ;
        RECT 364.950 284.400 460.050 285.600 ;
        RECT 364.950 283.950 367.050 284.400 ;
        RECT 451.950 283.950 454.050 284.400 ;
        RECT 457.950 283.950 460.050 284.400 ;
        RECT 631.950 285.600 634.050 286.050 ;
        RECT 685.950 285.600 688.050 286.050 ;
        RECT 631.950 284.400 688.050 285.600 ;
        RECT 631.950 283.950 634.050 284.400 ;
        RECT 685.950 283.950 688.050 284.400 ;
        RECT 364.950 276.600 367.050 277.050 ;
        RECT 329.400 275.400 367.050 276.600 ;
        RECT 274.950 273.600 277.050 274.050 ;
        RECT 329.400 273.600 330.600 275.400 ;
        RECT 364.950 274.950 367.050 275.400 ;
        RECT 274.950 272.400 330.600 273.600 ;
        RECT 274.950 271.950 277.050 272.400 ;
        RECT 235.950 264.600 238.050 265.050 ;
        RECT 253.950 264.600 256.050 265.050 ;
        RECT 274.950 264.600 277.050 265.050 ;
        RECT 235.950 263.400 277.050 264.600 ;
        RECT 235.950 262.950 238.050 263.400 ;
        RECT 253.950 262.950 256.050 263.400 ;
        RECT 274.950 262.950 277.050 263.400 ;
    END
  END Xin[6]
  PIN Xin[5]
    PORT
      LAYER metal1 ;
        RECT 583.950 453.450 586.050 454.050 ;
        RECT 592.950 453.450 595.050 454.200 ;
        RECT 583.950 452.550 595.050 453.450 ;
        RECT 583.950 451.950 586.050 452.550 ;
        RECT 592.950 452.100 595.050 452.550 ;
      LAYER metal2 ;
        RECT 614.400 889.050 615.450 906.450 ;
        RECT 577.950 886.950 580.050 889.050 ;
        RECT 613.950 886.950 616.050 889.050 ;
        RECT 578.400 811.050 579.450 886.950 ;
        RECT 619.950 884.100 622.050 889.050 ;
        RECT 637.950 884.100 640.050 886.200 ;
        RECT 620.400 883.350 621.600 884.100 ;
        RECT 638.400 883.350 639.600 884.100 ;
        RECT 577.950 808.950 580.050 811.050 ;
        RECT 586.950 808.950 589.050 811.050 ;
        RECT 587.400 733.050 588.450 808.950 ;
        RECT 586.950 730.950 589.050 733.050 ;
        RECT 592.950 730.950 595.050 733.050 ;
        RECT 593.400 574.050 594.450 730.950 ;
        RECT 592.950 571.950 595.050 574.050 ;
        RECT 592.950 565.950 595.050 568.050 ;
        RECT 593.400 454.200 594.450 565.950 ;
        RECT 583.950 451.950 586.050 454.050 ;
        RECT 592.950 452.100 595.050 454.200 ;
        RECT 584.400 421.050 585.450 451.950 ;
        RECT 583.950 418.950 586.050 421.050 ;
        RECT 592.950 418.950 595.050 421.050 ;
        RECT 593.400 376.050 594.450 418.950 ;
        RECT 586.950 373.950 589.050 376.050 ;
        RECT 592.950 373.950 595.050 376.050 ;
        RECT 425.400 365.400 426.600 367.650 ;
        RECT 425.400 358.050 426.450 365.400 ;
        RECT 587.400 358.050 588.450 373.950 ;
        RECT 424.950 355.950 427.050 358.050 ;
        RECT 586.950 355.950 589.050 358.050 ;
        RECT 587.400 343.050 588.450 355.950 ;
        RECT 586.950 340.950 589.050 343.050 ;
        RECT 646.950 339.000 649.050 343.050 ;
        RECT 647.400 337.350 648.600 339.000 ;
      LAYER via2 ;
        RECT 619.950 886.950 622.050 889.050 ;
        RECT 646.950 340.950 649.050 343.050 ;
      LAYER metal3 ;
        RECT 577.950 888.600 580.050 889.050 ;
        RECT 613.950 888.600 616.050 889.050 ;
        RECT 619.950 888.600 622.050 889.050 ;
        RECT 577.950 887.400 622.050 888.600 ;
        RECT 577.950 886.950 580.050 887.400 ;
        RECT 613.950 886.950 616.050 887.400 ;
        RECT 619.950 886.950 622.050 887.400 ;
        RECT 619.950 885.600 622.050 886.200 ;
        RECT 637.950 885.600 640.050 886.200 ;
        RECT 619.950 884.400 640.050 885.600 ;
        RECT 619.950 884.100 622.050 884.400 ;
        RECT 637.950 884.100 640.050 884.400 ;
        RECT 577.950 810.600 580.050 811.050 ;
        RECT 586.950 810.600 589.050 811.050 ;
        RECT 577.950 809.400 589.050 810.600 ;
        RECT 577.950 808.950 580.050 809.400 ;
        RECT 586.950 808.950 589.050 809.400 ;
        RECT 586.950 732.600 589.050 733.050 ;
        RECT 592.950 732.600 595.050 733.050 ;
        RECT 586.950 731.400 595.050 732.600 ;
        RECT 586.950 730.950 589.050 731.400 ;
        RECT 592.950 730.950 595.050 731.400 ;
        RECT 592.950 571.950 595.050 574.050 ;
        RECT 593.400 568.050 594.600 571.950 ;
        RECT 592.950 565.950 595.050 568.050 ;
        RECT 583.950 420.600 586.050 421.050 ;
        RECT 592.950 420.600 595.050 421.050 ;
        RECT 583.950 419.400 595.050 420.600 ;
        RECT 583.950 418.950 586.050 419.400 ;
        RECT 592.950 418.950 595.050 419.400 ;
        RECT 586.950 375.600 589.050 376.050 ;
        RECT 592.950 375.600 595.050 376.050 ;
        RECT 586.950 374.400 595.050 375.600 ;
        RECT 586.950 373.950 589.050 374.400 ;
        RECT 592.950 373.950 595.050 374.400 ;
        RECT 424.950 357.600 427.050 358.050 ;
        RECT 586.950 357.600 589.050 358.050 ;
        RECT 424.950 356.400 589.050 357.600 ;
        RECT 424.950 355.950 427.050 356.400 ;
        RECT 586.950 355.950 589.050 356.400 ;
        RECT 586.950 342.600 589.050 343.050 ;
        RECT 646.950 342.600 649.050 343.050 ;
        RECT 586.950 341.400 649.050 342.600 ;
        RECT 586.950 340.950 589.050 341.400 ;
        RECT 646.950 340.950 649.050 341.400 ;
    END
  END Xin[5]
  PIN Xin[4]
    PORT
      LAYER metal2 ;
        RECT 395.400 905.400 399.450 906.450 ;
        RECT 373.950 885.000 376.050 889.050 ;
        RECT 398.400 886.200 399.450 905.400 ;
        RECT 374.400 883.350 375.600 885.000 ;
        RECT 397.950 884.100 400.050 886.200 ;
        RECT 406.950 884.100 409.050 886.200 ;
        RECT 398.400 883.350 399.600 884.100 ;
        RECT 407.400 862.050 408.450 884.100 ;
        RECT 406.950 859.950 409.050 862.050 ;
        RECT 628.950 859.950 631.050 862.050 ;
        RECT 629.400 799.050 630.450 859.950 ;
        RECT 686.400 801.000 687.600 802.650 ;
        RECT 628.950 796.950 631.050 799.050 ;
        RECT 679.950 796.950 682.050 799.050 ;
        RECT 685.950 796.950 688.050 801.000 ;
        RECT 680.400 742.050 681.450 796.950 ;
        RECT 661.950 739.950 664.050 742.050 ;
        RECT 679.950 739.950 682.050 742.050 ;
        RECT 662.400 715.050 663.450 739.950 ;
        RECT 661.950 712.950 664.050 715.050 ;
        RECT 670.950 712.950 673.050 715.050 ;
        RECT 671.400 678.450 672.450 712.950 ;
        RECT 671.400 677.400 675.450 678.450 ;
        RECT 674.400 634.050 675.450 677.400 ;
        RECT 646.950 631.950 649.050 634.050 ;
        RECT 673.950 631.950 676.050 634.050 ;
        RECT 647.400 574.050 648.450 631.950 ;
        RECT 646.950 571.950 649.050 574.050 ;
        RECT 652.950 572.100 655.050 574.200 ;
        RECT 673.950 572.100 676.050 574.200 ;
        RECT 653.400 571.350 654.600 572.100 ;
        RECT 674.400 568.050 675.450 572.100 ;
        RECT 673.950 565.950 676.050 568.050 ;
        RECT 686.400 567.900 687.600 568.650 ;
        RECT 685.950 565.800 688.050 567.900 ;
        RECT 686.400 556.050 687.450 565.800 ;
        RECT 679.950 553.950 682.050 556.050 ;
        RECT 685.950 553.950 688.050 556.050 ;
        RECT 680.400 498.450 681.450 553.950 ;
        RECT 677.400 497.400 681.450 498.450 ;
        RECT 677.400 496.200 678.450 497.400 ;
        RECT 499.950 494.100 502.050 496.200 ;
        RECT 514.950 494.100 517.050 496.200 ;
        RECT 320.400 488.400 321.600 490.650 ;
        RECT 320.400 484.050 321.450 488.400 ;
        RECT 319.950 481.950 322.050 484.050 ;
        RECT 328.950 481.950 331.050 484.050 ;
        RECT 122.400 411.000 123.600 412.650 ;
        RECT 121.950 406.950 124.050 411.000 ;
        RECT 259.950 403.950 262.050 406.050 ;
        RECT 260.400 376.050 261.450 403.950 ;
        RECT 329.400 376.050 330.450 481.950 ;
        RECT 500.400 469.050 501.450 494.100 ;
        RECT 515.400 493.350 516.600 494.100 ;
        RECT 667.950 493.950 670.050 496.050 ;
        RECT 676.950 494.100 679.050 496.200 ;
        RECT 668.400 469.050 669.450 493.950 ;
        RECT 677.400 493.350 678.600 494.100 ;
        RECT 499.950 466.950 502.050 469.050 ;
        RECT 637.950 466.950 640.050 469.050 ;
        RECT 667.950 466.950 670.050 469.050 ;
        RECT 500.400 463.050 501.450 466.950 ;
        RECT 469.950 460.950 472.050 463.050 ;
        RECT 499.950 460.950 502.050 463.050 ;
        RECT 382.950 382.950 385.050 385.050 ;
        RECT 383.400 376.050 384.450 382.950 ;
        RECT 470.400 382.050 471.450 460.950 ;
        RECT 638.400 421.050 639.450 466.950 ;
        RECT 637.950 418.950 640.050 421.050 ;
        RECT 643.950 418.950 646.050 421.050 ;
        RECT 469.950 379.950 472.050 382.050 ;
        RECT 644.400 376.050 645.450 418.950 ;
        RECT 259.950 372.000 262.050 376.050 ;
        RECT 328.950 373.950 331.050 376.050 ;
        RECT 364.950 373.950 367.050 376.050 ;
        RECT 382.950 373.950 385.050 376.050 ;
        RECT 628.950 373.950 631.050 376.050 ;
        RECT 643.950 373.950 646.050 376.050 ;
        RECT 260.400 370.350 261.600 372.000 ;
        RECT 365.400 339.450 366.450 373.950 ;
        RECT 383.400 372.600 384.450 373.950 ;
        RECT 383.400 370.350 384.600 372.600 ;
        RECT 629.400 355.050 630.450 373.950 ;
        RECT 613.950 352.950 616.050 355.050 ;
        RECT 628.950 352.950 631.050 355.050 ;
        RECT 362.400 338.400 366.450 339.450 ;
        RECT 254.400 333.000 255.600 334.650 ;
        RECT 329.400 333.000 330.600 334.650 ;
        RECT 253.950 328.950 256.050 333.000 ;
        RECT 328.950 328.950 331.050 333.000 ;
        RECT 362.400 331.050 363.450 338.400 ;
        RECT 605.400 333.900 606.600 334.650 ;
        RECT 614.400 333.900 615.450 352.950 ;
        RECT 604.950 331.800 607.050 333.900 ;
        RECT 613.950 331.800 616.050 333.900 ;
        RECT 361.950 328.950 364.050 331.050 ;
        RECT 254.400 316.050 255.450 328.950 ;
        RECT 220.950 313.950 223.050 316.050 ;
        RECT 253.950 313.950 256.050 316.050 ;
        RECT 221.400 294.600 222.450 313.950 ;
        RECT 221.400 292.350 222.600 294.600 ;
      LAYER via2 ;
        RECT 373.950 886.950 376.050 889.050 ;
        RECT 259.950 373.950 262.050 376.050 ;
      LAYER metal3 ;
        RECT 373.950 888.600 376.050 889.050 ;
        RECT 373.950 887.400 399.600 888.600 ;
        RECT 373.950 886.950 376.050 887.400 ;
        RECT 398.400 886.200 399.600 887.400 ;
        RECT 397.950 885.750 400.050 886.200 ;
        RECT 406.950 885.750 409.050 886.200 ;
        RECT 397.950 884.550 409.050 885.750 ;
        RECT 397.950 884.100 400.050 884.550 ;
        RECT 406.950 884.100 409.050 884.550 ;
        RECT 406.950 861.600 409.050 862.050 ;
        RECT 628.950 861.600 631.050 862.050 ;
        RECT 406.950 860.400 631.050 861.600 ;
        RECT 406.950 859.950 409.050 860.400 ;
        RECT 628.950 859.950 631.050 860.400 ;
        RECT 628.950 798.600 631.050 799.050 ;
        RECT 679.950 798.600 682.050 799.050 ;
        RECT 685.950 798.600 688.050 799.050 ;
        RECT 628.950 797.400 688.050 798.600 ;
        RECT 628.950 796.950 631.050 797.400 ;
        RECT 679.950 796.950 682.050 797.400 ;
        RECT 685.950 796.950 688.050 797.400 ;
        RECT 661.950 741.600 664.050 742.050 ;
        RECT 679.950 741.600 682.050 742.050 ;
        RECT 661.950 740.400 682.050 741.600 ;
        RECT 661.950 739.950 664.050 740.400 ;
        RECT 679.950 739.950 682.050 740.400 ;
        RECT 661.950 714.600 664.050 715.050 ;
        RECT 670.950 714.600 673.050 715.050 ;
        RECT 661.950 713.400 673.050 714.600 ;
        RECT 661.950 712.950 664.050 713.400 ;
        RECT 670.950 712.950 673.050 713.400 ;
        RECT 646.950 633.600 649.050 634.050 ;
        RECT 673.950 633.600 676.050 634.050 ;
        RECT 646.950 632.400 676.050 633.600 ;
        RECT 646.950 631.950 649.050 632.400 ;
        RECT 673.950 631.950 676.050 632.400 ;
        RECT 646.950 573.600 649.050 574.050 ;
        RECT 652.950 573.750 655.050 574.200 ;
        RECT 673.950 573.750 676.050 574.200 ;
        RECT 652.950 573.600 676.050 573.750 ;
        RECT 646.950 572.550 676.050 573.600 ;
        RECT 646.950 572.400 655.050 572.550 ;
        RECT 646.950 571.950 649.050 572.400 ;
        RECT 652.950 572.100 655.050 572.400 ;
        RECT 673.950 572.100 676.050 572.550 ;
        RECT 673.950 567.600 676.050 568.050 ;
        RECT 685.950 567.600 688.050 567.900 ;
        RECT 673.950 566.400 688.050 567.600 ;
        RECT 673.950 565.950 676.050 566.400 ;
        RECT 685.950 565.800 688.050 566.400 ;
        RECT 679.950 555.600 682.050 556.050 ;
        RECT 685.950 555.600 688.050 556.050 ;
        RECT 679.950 554.400 688.050 555.600 ;
        RECT 679.950 553.950 682.050 554.400 ;
        RECT 685.950 553.950 688.050 554.400 ;
        RECT 499.950 495.750 502.050 496.200 ;
        RECT 514.950 495.750 517.050 496.200 ;
        RECT 499.950 494.550 517.050 495.750 ;
        RECT 499.950 494.100 502.050 494.550 ;
        RECT 514.950 494.100 517.050 494.550 ;
        RECT 667.950 495.600 670.050 496.050 ;
        RECT 676.950 495.600 679.050 496.200 ;
        RECT 667.950 494.400 679.050 495.600 ;
        RECT 667.950 493.950 670.050 494.400 ;
        RECT 676.950 494.100 679.050 494.400 ;
        RECT 319.950 483.600 322.050 484.050 ;
        RECT 328.950 483.600 331.050 484.050 ;
        RECT 319.950 482.400 331.050 483.600 ;
        RECT 319.950 481.950 322.050 482.400 ;
        RECT 328.950 481.950 331.050 482.400 ;
        RECT 499.950 468.600 502.050 469.050 ;
        RECT 637.950 468.600 640.050 469.050 ;
        RECT 667.950 468.600 670.050 469.050 ;
        RECT 499.950 467.400 670.050 468.600 ;
        RECT 499.950 466.950 502.050 467.400 ;
        RECT 637.950 466.950 640.050 467.400 ;
        RECT 667.950 466.950 670.050 467.400 ;
        RECT 469.950 462.600 472.050 463.050 ;
        RECT 499.950 462.600 502.050 463.050 ;
        RECT 469.950 461.400 502.050 462.600 ;
        RECT 469.950 460.950 472.050 461.400 ;
        RECT 499.950 460.950 502.050 461.400 ;
        RECT 637.950 420.600 640.050 421.050 ;
        RECT 643.950 420.600 646.050 421.050 ;
        RECT 637.950 419.400 646.050 420.600 ;
        RECT 637.950 418.950 640.050 419.400 ;
        RECT 643.950 418.950 646.050 419.400 ;
        RECT 121.950 405.600 124.050 409.050 ;
        RECT 259.950 405.600 262.050 406.050 ;
        RECT 121.950 405.000 262.050 405.600 ;
        RECT 122.400 404.400 262.050 405.000 ;
        RECT 259.950 403.950 262.050 404.400 ;
        RECT 382.950 384.600 385.050 385.050 ;
        RECT 382.950 383.400 405.600 384.600 ;
        RECT 382.950 382.950 385.050 383.400 ;
        RECT 404.400 381.600 405.600 383.400 ;
        RECT 469.950 381.600 472.050 382.050 ;
        RECT 404.400 380.400 472.050 381.600 ;
        RECT 469.950 379.950 472.050 380.400 ;
        RECT 259.950 375.600 262.050 376.050 ;
        RECT 328.950 375.600 331.050 376.050 ;
        RECT 364.950 375.600 367.050 376.050 ;
        RECT 382.950 375.600 385.050 376.050 ;
        RECT 259.950 374.400 385.050 375.600 ;
        RECT 259.950 373.950 262.050 374.400 ;
        RECT 328.950 373.950 331.050 374.400 ;
        RECT 364.950 373.950 367.050 374.400 ;
        RECT 382.950 373.950 385.050 374.400 ;
        RECT 628.950 375.600 631.050 376.050 ;
        RECT 643.950 375.600 646.050 376.050 ;
        RECT 628.950 374.400 646.050 375.600 ;
        RECT 628.950 373.950 631.050 374.400 ;
        RECT 643.950 373.950 646.050 374.400 ;
        RECT 613.950 354.600 616.050 355.050 ;
        RECT 628.950 354.600 631.050 355.050 ;
        RECT 613.950 353.400 631.050 354.600 ;
        RECT 613.950 352.950 616.050 353.400 ;
        RECT 628.950 352.950 631.050 353.400 ;
        RECT 604.950 333.450 607.050 333.900 ;
        RECT 613.950 333.450 616.050 333.900 ;
        RECT 604.950 332.250 616.050 333.450 ;
        RECT 604.950 331.800 607.050 332.250 ;
        RECT 613.950 331.800 616.050 332.250 ;
        RECT 253.950 330.600 256.050 331.050 ;
        RECT 328.950 330.600 331.050 331.050 ;
        RECT 361.950 330.600 364.050 331.050 ;
        RECT 253.950 329.400 364.050 330.600 ;
        RECT 253.950 328.950 256.050 329.400 ;
        RECT 328.950 328.950 331.050 329.400 ;
        RECT 361.950 328.950 364.050 329.400 ;
        RECT 220.950 315.600 223.050 316.050 ;
        RECT 253.950 315.600 256.050 316.050 ;
        RECT 220.950 314.400 256.050 315.600 ;
        RECT 220.950 313.950 223.050 314.400 ;
        RECT 253.950 313.950 256.050 314.400 ;
    END
  END Xin[4]
  PIN Xin[3]
    PORT
      LAYER metal2 ;
        RECT 20.400 905.400 24.450 906.450 ;
        RECT 23.400 892.050 24.450 905.400 ;
        RECT 22.950 889.950 25.050 892.050 ;
        RECT 220.950 889.950 223.050 892.050 ;
        RECT 23.400 885.600 24.450 889.950 ;
        RECT 23.400 883.350 24.600 885.600 ;
        RECT 221.400 787.050 222.450 889.950 ;
        RECT 220.950 784.950 223.050 787.050 ;
        RECT 247.950 784.950 250.050 787.050 ;
        RECT 248.400 742.050 249.450 784.950 ;
        RECT 247.950 739.950 250.050 742.050 ;
        RECT 259.950 739.950 262.050 742.050 ;
        RECT 260.400 684.450 261.450 739.950 ;
        RECT 260.400 683.400 264.450 684.450 ;
        RECT 263.400 676.050 264.450 683.400 ;
        RECT 272.400 678.000 273.600 679.650 ;
        RECT 241.950 673.950 244.050 676.050 ;
        RECT 262.950 673.950 265.050 676.050 ;
        RECT 271.950 673.950 274.050 678.000 ;
        RECT 242.400 613.050 243.450 673.950 ;
        RECT 241.950 610.950 244.050 613.050 ;
        RECT 259.950 610.950 262.050 613.050 ;
        RECT 260.400 565.050 261.450 610.950 ;
        RECT 244.950 562.950 247.050 565.050 ;
        RECT 259.950 562.950 262.050 565.050 ;
        RECT 236.400 522.900 237.600 523.650 ;
        RECT 245.400 522.900 246.450 562.950 ;
        RECT 235.950 520.800 238.050 522.900 ;
        RECT 244.950 520.800 247.050 522.900 ;
        RECT 253.950 520.950 256.050 523.050 ;
        RECT 254.400 495.600 255.450 520.950 ;
        RECT 254.400 493.350 255.600 495.600 ;
      LAYER metal3 ;
        RECT 22.950 891.600 25.050 892.050 ;
        RECT 220.950 891.600 223.050 892.050 ;
        RECT 22.950 890.400 223.050 891.600 ;
        RECT 22.950 889.950 25.050 890.400 ;
        RECT 220.950 889.950 223.050 890.400 ;
        RECT 220.950 786.600 223.050 787.050 ;
        RECT 247.950 786.600 250.050 787.050 ;
        RECT 220.950 785.400 250.050 786.600 ;
        RECT 220.950 784.950 223.050 785.400 ;
        RECT 247.950 784.950 250.050 785.400 ;
        RECT 247.950 741.600 250.050 742.050 ;
        RECT 259.950 741.600 262.050 742.050 ;
        RECT 247.950 740.400 262.050 741.600 ;
        RECT 247.950 739.950 250.050 740.400 ;
        RECT 259.950 739.950 262.050 740.400 ;
        RECT 241.950 675.600 244.050 676.050 ;
        RECT 262.950 675.600 265.050 676.050 ;
        RECT 271.950 675.600 274.050 676.050 ;
        RECT 241.950 674.400 274.050 675.600 ;
        RECT 241.950 673.950 244.050 674.400 ;
        RECT 262.950 673.950 265.050 674.400 ;
        RECT 271.950 673.950 274.050 674.400 ;
        RECT 241.950 612.600 244.050 613.050 ;
        RECT 259.950 612.600 262.050 613.050 ;
        RECT 241.950 611.400 262.050 612.600 ;
        RECT 241.950 610.950 244.050 611.400 ;
        RECT 259.950 610.950 262.050 611.400 ;
        RECT 244.950 564.600 247.050 565.050 ;
        RECT 259.950 564.600 262.050 565.050 ;
        RECT 244.950 563.400 262.050 564.600 ;
        RECT 244.950 562.950 247.050 563.400 ;
        RECT 259.950 562.950 262.050 563.400 ;
        RECT 235.950 522.450 238.050 522.900 ;
        RECT 244.950 522.600 247.050 522.900 ;
        RECT 253.950 522.600 256.050 523.050 ;
        RECT 244.950 522.450 256.050 522.600 ;
        RECT 235.950 521.400 256.050 522.450 ;
        RECT 235.950 521.250 247.050 521.400 ;
        RECT 235.950 520.800 238.050 521.250 ;
        RECT 244.950 520.800 247.050 521.250 ;
        RECT 253.950 520.950 256.050 521.400 ;
    END
  END Xin[3]
  PIN Xin[2]
    PORT
      LAYER metal1 ;
        RECT 166.950 615.450 169.050 616.050 ;
        RECT 178.950 615.450 181.050 616.050 ;
        RECT 166.950 614.550 181.050 615.450 ;
        RECT 166.950 613.950 169.050 614.550 ;
        RECT 178.950 613.950 181.050 614.550 ;
      LAYER metal2 ;
        RECT 44.400 723.000 45.600 724.650 ;
        RECT 122.400 723.000 123.600 724.650 ;
        RECT 43.950 718.950 46.050 723.000 ;
        RECT 115.950 718.950 118.050 721.050 ;
        RECT 121.950 718.950 124.050 723.000 ;
        RECT 17.400 678.900 18.600 679.650 ;
        RECT 16.950 673.950 19.050 678.900 ;
        RECT 116.400 676.050 117.450 718.950 ;
        RECT 115.950 673.950 118.050 676.050 ;
        RECT 17.400 651.600 18.450 673.950 ;
        RECT 17.400 649.350 18.600 651.600 ;
        RECT 116.400 628.050 117.450 673.950 ;
        RECT 464.400 644.400 465.600 646.650 ;
        RECT 115.950 625.950 118.050 628.050 ;
        RECT 166.950 625.950 169.050 628.050 ;
        RECT 167.400 616.050 168.450 625.950 ;
        RECT 166.950 613.950 169.050 616.050 ;
        RECT 178.950 613.950 184.050 616.050 ;
        RECT 352.950 610.950 355.050 613.050 ;
        RECT 367.950 610.950 370.050 613.050 ;
        RECT 353.400 565.050 354.450 610.950 ;
        RECT 368.400 606.600 369.450 610.950 ;
        RECT 464.400 607.200 465.450 644.400 ;
        RECT 368.400 604.350 369.600 606.600 ;
        RECT 463.950 605.100 466.050 607.200 ;
        RECT 469.950 605.100 472.050 607.200 ;
        RECT 425.400 567.450 426.600 568.650 ;
        RECT 422.400 567.000 426.600 567.450 ;
        RECT 421.950 566.400 426.600 567.000 ;
        RECT 352.950 562.950 355.050 565.050 ;
        RECT 421.950 562.950 424.050 566.400 ;
        RECT 353.400 553.050 354.450 562.950 ;
        RECT 425.400 562.050 426.450 566.400 ;
        RECT 464.400 562.050 465.450 605.100 ;
        RECT 470.400 604.350 471.600 605.100 ;
        RECT 424.950 559.950 427.050 562.050 ;
        RECT 463.950 559.950 466.050 562.050 ;
        RECT 313.950 550.950 316.050 553.050 ;
        RECT 352.800 550.950 354.900 553.050 ;
        RECT 247.950 450.000 250.050 454.050 ;
        RECT 248.400 448.350 249.600 450.000 ;
        RECT 295.950 449.100 298.050 454.050 ;
        RECT 314.400 451.200 315.450 550.950 ;
        RECT 296.400 448.350 297.600 449.100 ;
        RECT 307.950 448.950 310.050 451.050 ;
        RECT 313.950 449.100 316.050 451.200 ;
        RECT 308.400 403.050 309.450 448.950 ;
        RECT 314.400 448.350 315.600 449.100 ;
        RECT 338.400 410.400 339.600 412.650 ;
        RECT 338.400 403.050 339.450 410.400 ;
        RECT 307.950 400.950 310.050 403.050 ;
        RECT 337.950 400.950 340.050 403.050 ;
        RECT 338.400 385.050 339.450 400.950 ;
        RECT 337.950 382.950 340.050 385.050 ;
        RECT 358.950 382.950 361.050 385.050 ;
        RECT 359.400 372.600 360.450 382.950 ;
        RECT 359.400 370.350 360.600 372.600 ;
      LAYER via2 ;
        RECT 16.950 676.800 19.050 678.900 ;
        RECT 181.950 613.950 184.050 616.050 ;
        RECT 247.950 451.950 250.050 454.050 ;
        RECT 295.950 451.950 298.050 454.050 ;
      LAYER metal3 ;
        RECT 43.950 720.600 46.050 721.050 ;
        RECT 115.950 720.600 118.050 721.050 ;
        RECT 121.950 720.600 124.050 721.050 ;
        RECT 43.950 719.400 124.050 720.600 ;
        RECT 43.950 718.950 46.050 719.400 ;
        RECT 115.950 718.950 118.050 719.400 ;
        RECT 121.950 718.950 124.050 719.400 ;
        RECT 16.950 678.600 19.050 678.900 ;
        RECT -3.600 677.400 19.050 678.600 ;
        RECT 16.950 676.800 19.050 677.400 ;
        RECT 16.950 675.600 19.050 676.050 ;
        RECT 115.950 675.600 118.050 676.050 ;
        RECT 16.950 674.400 118.050 675.600 ;
        RECT 16.950 673.950 19.050 674.400 ;
        RECT 115.950 673.950 118.050 674.400 ;
        RECT 115.950 627.600 118.050 628.050 ;
        RECT 166.950 627.600 169.050 628.050 ;
        RECT 115.950 626.400 169.050 627.600 ;
        RECT 115.950 625.950 118.050 626.400 ;
        RECT 166.950 625.950 169.050 626.400 ;
        RECT 181.950 615.600 184.050 616.050 ;
        RECT 181.950 614.400 354.600 615.600 ;
        RECT 181.950 613.950 184.050 614.400 ;
        RECT 353.400 613.050 354.600 614.400 ;
        RECT 352.950 612.600 355.050 613.050 ;
        RECT 367.950 612.600 370.050 613.050 ;
        RECT 352.950 611.400 370.050 612.600 ;
        RECT 352.950 610.950 355.050 611.400 ;
        RECT 367.950 610.950 370.050 611.400 ;
        RECT 463.950 606.750 466.050 607.200 ;
        RECT 469.950 606.750 472.050 607.200 ;
        RECT 463.950 605.550 472.050 606.750 ;
        RECT 463.950 605.100 466.050 605.550 ;
        RECT 469.950 605.100 472.050 605.550 ;
        RECT 352.950 564.600 355.050 565.050 ;
        RECT 421.950 564.600 424.050 565.050 ;
        RECT 352.950 563.400 424.050 564.600 ;
        RECT 352.950 562.950 355.050 563.400 ;
        RECT 421.950 562.950 424.050 563.400 ;
        RECT 424.950 561.600 427.050 562.050 ;
        RECT 463.950 561.600 466.050 562.050 ;
        RECT 424.950 560.400 466.050 561.600 ;
        RECT 424.950 559.950 427.050 560.400 ;
        RECT 463.950 559.950 466.050 560.400 ;
        RECT 313.950 552.600 316.050 553.050 ;
        RECT 352.800 552.600 354.900 553.050 ;
        RECT 313.950 551.400 354.900 552.600 ;
        RECT 313.950 550.950 316.050 551.400 ;
        RECT 352.800 550.950 354.900 551.400 ;
        RECT 247.950 453.600 250.050 454.050 ;
        RECT 295.950 453.600 298.050 454.050 ;
        RECT 247.950 452.400 298.050 453.600 ;
        RECT 247.950 451.950 250.050 452.400 ;
        RECT 295.950 451.950 298.050 452.400 ;
        RECT 295.950 450.600 298.050 451.200 ;
        RECT 307.950 450.600 310.050 451.050 ;
        RECT 313.950 450.600 316.050 451.200 ;
        RECT 295.950 449.400 316.050 450.600 ;
        RECT 295.950 449.100 298.050 449.400 ;
        RECT 307.950 448.950 310.050 449.400 ;
        RECT 313.950 449.100 316.050 449.400 ;
        RECT 307.950 402.600 310.050 403.050 ;
        RECT 337.950 402.600 340.050 403.050 ;
        RECT 307.950 401.400 340.050 402.600 ;
        RECT 307.950 400.950 310.050 401.400 ;
        RECT 337.950 400.950 340.050 401.400 ;
        RECT 337.950 384.600 340.050 385.050 ;
        RECT 358.950 384.600 361.050 385.050 ;
        RECT 337.950 383.400 361.050 384.600 ;
        RECT 337.950 382.950 340.050 383.400 ;
        RECT 358.950 382.950 361.050 383.400 ;
    END
  END Xin[2]
  PIN Xin[1]
    PORT
      LAYER metal1 ;
        RECT 394.950 609.450 397.050 610.050 ;
        RECT 406.950 609.450 409.050 610.050 ;
        RECT 394.950 608.550 409.050 609.450 ;
        RECT 394.950 607.950 397.050 608.550 ;
        RECT 406.950 607.950 409.050 608.550 ;
      LAYER metal2 ;
        RECT 28.950 688.950 31.050 691.050 ;
        RECT 64.950 688.950 67.050 691.050 ;
        RECT 29.400 640.050 30.450 688.950 ;
        RECT 65.400 684.600 66.450 688.950 ;
        RECT 65.400 682.350 66.600 684.600 ;
        RECT 331.950 683.100 334.050 685.200 ;
        RECT 340.950 683.100 343.050 685.200 ;
        RECT 332.400 673.050 333.450 683.100 ;
        RECT 341.400 682.350 342.600 683.100 ;
        RECT 325.950 670.950 328.050 673.050 ;
        RECT 331.950 670.950 334.050 673.050 ;
        RECT 311.400 644.400 312.600 646.650 ;
        RECT 311.400 640.050 312.450 644.400 ;
        RECT 326.400 640.050 327.450 670.950 ;
        RECT 1.950 637.950 4.050 640.050 ;
        RECT 28.950 637.950 31.050 640.050 ;
        RECT 310.950 637.950 313.050 640.050 ;
        RECT 325.950 637.950 328.050 640.050 ;
        RECT 2.400 616.050 3.450 637.950 ;
        RECT 1.950 613.950 4.050 616.050 ;
        RECT 2.400 502.050 3.450 613.950 ;
        RECT 311.400 600.450 312.450 637.950 ;
        RECT 326.400 628.050 327.450 637.950 ;
        RECT 325.950 625.950 328.050 628.050 ;
        RECT 394.950 625.950 397.050 628.050 ;
        RECT 395.400 610.050 396.450 625.950 ;
        RECT 394.950 607.950 397.050 610.050 ;
        RECT 406.950 605.100 409.050 610.050 ;
        RECT 407.400 604.350 408.600 605.100 ;
        RECT 308.400 599.400 312.450 600.450 ;
        RECT 290.400 566.400 291.600 568.650 ;
        RECT 290.400 559.050 291.450 566.400 ;
        RECT 308.400 559.050 309.450 599.400 ;
        RECT 406.950 595.950 409.050 598.050 ;
        RECT 407.400 573.600 408.450 595.950 ;
        RECT 407.400 571.350 408.600 573.600 ;
        RECT 289.950 556.950 292.050 559.050 ;
        RECT 307.950 556.950 310.050 559.050 ;
        RECT 1.950 499.950 4.050 502.050 ;
        RECT 64.950 499.950 67.050 502.050 ;
        RECT 79.950 499.950 82.050 502.050 ;
        RECT 100.950 499.950 103.050 502.050 ;
        RECT 196.950 499.950 199.050 502.050 ;
        RECT 65.400 454.050 66.450 499.950 ;
        RECT 80.400 495.600 81.450 499.950 ;
        RECT 101.400 495.600 102.450 499.950 ;
        RECT 80.400 493.350 81.600 495.600 ;
        RECT 101.400 493.350 102.600 495.600 ;
        RECT 197.400 487.050 198.450 499.950 ;
        RECT 209.400 489.000 210.600 490.650 ;
        RECT 239.400 489.000 240.600 490.650 ;
        RECT 196.950 484.950 199.050 487.050 ;
        RECT 208.950 484.950 211.050 489.000 ;
        RECT 229.950 484.950 232.050 487.050 ;
        RECT 238.950 484.950 241.050 489.000 ;
        RECT 230.400 466.050 231.450 484.950 ;
        RECT 290.400 466.050 291.450 556.950 ;
        RECT 229.950 463.950 232.050 466.050 ;
        RECT 289.950 463.950 292.050 466.050 ;
        RECT 334.950 463.950 337.050 466.050 ;
        RECT 64.950 451.950 67.050 454.050 ;
        RECT 82.950 450.000 85.050 454.050 ;
        RECT 230.400 450.600 231.450 463.950 ;
        RECT 335.400 450.600 336.450 463.950 ;
        RECT 83.400 448.350 84.600 450.000 ;
        RECT 230.400 448.350 231.600 450.600 ;
        RECT 335.400 448.350 336.600 450.600 ;
      LAYER via2 ;
        RECT 82.950 451.950 85.050 454.050 ;
      LAYER metal3 ;
        RECT 28.950 690.600 31.050 691.050 ;
        RECT 64.950 690.600 67.050 691.050 ;
        RECT 28.950 689.400 67.050 690.600 ;
        RECT 28.950 688.950 31.050 689.400 ;
        RECT 64.950 688.950 67.050 689.400 ;
        RECT 331.950 684.750 334.050 685.200 ;
        RECT 340.950 684.750 343.050 685.200 ;
        RECT 331.950 683.550 343.050 684.750 ;
        RECT 331.950 683.100 334.050 683.550 ;
        RECT 340.950 683.100 343.050 683.550 ;
        RECT 325.950 672.600 328.050 673.050 ;
        RECT 331.950 672.600 334.050 673.050 ;
        RECT 325.950 671.400 334.050 672.600 ;
        RECT 325.950 670.950 328.050 671.400 ;
        RECT 331.950 670.950 334.050 671.400 ;
        RECT 1.950 639.600 4.050 640.050 ;
        RECT 28.950 639.600 31.050 640.050 ;
        RECT 1.950 638.400 31.050 639.600 ;
        RECT 1.950 637.950 4.050 638.400 ;
        RECT 28.950 637.950 31.050 638.400 ;
        RECT 310.950 639.600 313.050 640.050 ;
        RECT 325.950 639.600 328.050 640.050 ;
        RECT 310.950 638.400 328.050 639.600 ;
        RECT 310.950 637.950 313.050 638.400 ;
        RECT 325.950 637.950 328.050 638.400 ;
        RECT 325.950 627.600 328.050 628.050 ;
        RECT 394.950 627.600 397.050 628.050 ;
        RECT 325.950 626.400 397.050 627.600 ;
        RECT 325.950 625.950 328.050 626.400 ;
        RECT 394.950 625.950 397.050 626.400 ;
        RECT 1.950 615.600 4.050 616.050 ;
        RECT -3.600 614.400 4.050 615.600 ;
        RECT 1.950 613.950 4.050 614.400 ;
        RECT 406.950 605.100 409.050 607.200 ;
        RECT 407.400 598.050 408.600 605.100 ;
        RECT 406.950 595.950 409.050 598.050 ;
        RECT 289.950 558.600 292.050 559.050 ;
        RECT 307.950 558.600 310.050 559.050 ;
        RECT 289.950 557.400 310.050 558.600 ;
        RECT 289.950 556.950 292.050 557.400 ;
        RECT 307.950 556.950 310.050 557.400 ;
        RECT 1.950 501.600 4.050 502.050 ;
        RECT 64.950 501.600 67.050 502.050 ;
        RECT 79.950 501.600 82.050 502.050 ;
        RECT 100.950 501.600 103.050 502.050 ;
        RECT 196.950 501.600 199.050 502.050 ;
        RECT 1.950 500.400 199.050 501.600 ;
        RECT 1.950 499.950 4.050 500.400 ;
        RECT 64.950 499.950 67.050 500.400 ;
        RECT 79.950 499.950 82.050 500.400 ;
        RECT 100.950 499.950 103.050 500.400 ;
        RECT 196.950 499.950 199.050 500.400 ;
        RECT 196.950 486.600 199.050 487.050 ;
        RECT 208.950 486.600 211.050 487.050 ;
        RECT 229.950 486.600 232.050 487.050 ;
        RECT 238.950 486.600 241.050 487.050 ;
        RECT 196.950 485.400 241.050 486.600 ;
        RECT 196.950 484.950 199.050 485.400 ;
        RECT 208.950 484.950 211.050 485.400 ;
        RECT 229.950 484.950 232.050 485.400 ;
        RECT 238.950 484.950 241.050 485.400 ;
        RECT 229.950 465.600 232.050 466.050 ;
        RECT 289.950 465.600 292.050 466.050 ;
        RECT 334.950 465.600 337.050 466.050 ;
        RECT 229.950 464.400 337.050 465.600 ;
        RECT 229.950 463.950 232.050 464.400 ;
        RECT 289.950 463.950 292.050 464.400 ;
        RECT 334.950 463.950 337.050 464.400 ;
        RECT 64.950 453.600 67.050 454.050 ;
        RECT 82.950 453.600 85.050 454.050 ;
        RECT 64.950 452.400 85.050 453.600 ;
        RECT 64.950 451.950 67.050 452.400 ;
        RECT 82.950 451.950 85.050 452.400 ;
    END
  END Xin[1]
  PIN Xin[0]
    PORT
      LAYER metal2 ;
        RECT 362.400 566.400 363.600 568.650 ;
        RECT 362.400 561.450 363.450 566.400 ;
        RECT 359.400 560.400 363.450 561.450 ;
        RECT 359.400 535.050 360.450 560.400 ;
        RECT 286.950 532.950 289.050 535.050 ;
        RECT 358.950 532.950 361.050 535.050 ;
        RECT 257.400 521.400 258.600 523.650 ;
        RECT 257.400 517.050 258.450 521.400 ;
        RECT 287.400 517.050 288.450 532.950 ;
        RECT 247.950 514.950 250.050 517.050 ;
        RECT 256.950 514.950 259.050 517.050 ;
        RECT 286.950 514.950 289.050 517.050 ;
        RECT 248.400 475.050 249.450 514.950 ;
        RECT 359.400 505.050 360.450 532.950 ;
        RECT 352.950 502.950 355.050 505.050 ;
        RECT 358.800 502.950 360.900 505.050 ;
        RECT 353.400 484.050 354.450 502.950 ;
        RECT 359.400 488.400 360.600 490.650 ;
        RECT 383.400 488.400 384.600 490.650 ;
        RECT 359.400 484.050 360.450 488.400 ;
        RECT 383.400 484.050 384.450 488.400 ;
        RECT 352.950 481.950 355.050 484.050 ;
        RECT 358.950 481.950 361.050 484.050 ;
        RECT 382.950 481.950 385.050 484.050 ;
        RECT 43.950 472.950 46.050 475.050 ;
        RECT 217.950 472.950 220.050 475.050 ;
        RECT 247.950 472.950 250.050 475.050 ;
        RECT 44.400 460.050 45.450 472.950 ;
        RECT 43.950 457.950 46.050 460.050 ;
        RECT 44.400 450.450 45.450 457.950 ;
        RECT 218.400 451.200 219.450 472.950 ;
        RECT 47.400 450.450 48.600 450.600 ;
        RECT 44.400 449.400 48.600 450.450 ;
        RECT 47.400 448.350 48.600 449.400 ;
        RECT 184.950 449.100 187.050 451.200 ;
        RECT 217.950 449.100 220.050 451.200 ;
        RECT 185.400 448.350 186.600 449.100 ;
        RECT 218.400 448.350 219.600 449.100 ;
      LAYER metal3 ;
        RECT 286.950 534.600 289.050 535.050 ;
        RECT 358.950 534.600 361.050 535.050 ;
        RECT 286.950 533.400 361.050 534.600 ;
        RECT 286.950 532.950 289.050 533.400 ;
        RECT 358.950 532.950 361.050 533.400 ;
        RECT 247.950 516.600 250.050 517.050 ;
        RECT 256.950 516.600 259.050 517.050 ;
        RECT 286.950 516.600 289.050 517.050 ;
        RECT 247.950 515.400 289.050 516.600 ;
        RECT 247.950 514.950 250.050 515.400 ;
        RECT 256.950 514.950 259.050 515.400 ;
        RECT 286.950 514.950 289.050 515.400 ;
        RECT 352.950 504.600 355.050 505.050 ;
        RECT 358.800 504.600 360.900 505.050 ;
        RECT 352.950 503.400 360.900 504.600 ;
        RECT 352.950 502.950 355.050 503.400 ;
        RECT 358.800 502.950 360.900 503.400 ;
        RECT 352.950 483.600 355.050 484.050 ;
        RECT 358.950 483.600 361.050 484.050 ;
        RECT 382.950 483.600 385.050 484.050 ;
        RECT 352.950 482.400 385.050 483.600 ;
        RECT 352.950 481.950 355.050 482.400 ;
        RECT 358.950 481.950 361.050 482.400 ;
        RECT 382.950 481.950 385.050 482.400 ;
        RECT 43.950 474.600 46.050 475.050 ;
        RECT 217.950 474.600 220.050 475.050 ;
        RECT 247.950 474.600 250.050 475.050 ;
        RECT 43.950 473.400 250.050 474.600 ;
        RECT 43.950 472.950 46.050 473.400 ;
        RECT 217.950 472.950 220.050 473.400 ;
        RECT 247.950 472.950 250.050 473.400 ;
        RECT 43.950 459.600 46.050 460.050 ;
        RECT -3.600 458.400 46.050 459.600 ;
        RECT 43.950 457.950 46.050 458.400 ;
        RECT 184.950 450.600 187.050 451.200 ;
        RECT 217.950 450.600 220.050 451.200 ;
        RECT 184.950 449.400 220.050 450.600 ;
        RECT 184.950 449.100 187.050 449.400 ;
        RECT 217.950 449.100 220.050 449.400 ;
    END
  END Xin[0]
  PIN Xout[7]
    PORT
      LAYER metal2 ;
        RECT 10.950 415.950 13.050 418.050 ;
        RECT 11.400 411.450 12.450 415.950 ;
        RECT 14.400 411.450 15.600 412.650 ;
        RECT 11.400 410.400 15.600 411.450 ;
      LAYER metal3 ;
        RECT 10.950 417.600 13.050 418.050 ;
        RECT -3.600 416.400 13.050 417.600 ;
        RECT 10.950 415.950 13.050 416.400 ;
    END
  END Xout[7]
  PIN Xout[6]
    PORT
      LAYER metal2 ;
        RECT 158.400 898.050 159.450 906.450 ;
        RECT 151.950 895.950 154.050 898.050 ;
        RECT 157.950 895.950 160.050 898.050 ;
        RECT 152.400 879.450 153.450 895.950 ;
        RECT 155.400 879.450 156.600 880.650 ;
        RECT 152.400 878.400 156.600 879.450 ;
      LAYER metal3 ;
        RECT 151.950 897.600 154.050 898.050 ;
        RECT 157.950 897.600 160.050 898.050 ;
        RECT 151.950 896.400 160.050 897.600 ;
        RECT 151.950 895.950 154.050 896.400 ;
        RECT 157.950 895.950 160.050 896.400 ;
    END
  END Xout[6]
  PIN Xout[5]
    PORT
      LAYER metal2 ;
        RECT 596.400 901.050 597.450 906.450 ;
        RECT 595.950 898.950 598.050 901.050 ;
        RECT 601.950 898.950 604.050 901.050 ;
        RECT 599.400 879.450 600.600 880.650 ;
        RECT 602.400 879.450 603.450 898.950 ;
        RECT 599.400 878.400 603.450 879.450 ;
      LAYER metal3 ;
        RECT 595.950 900.600 598.050 901.050 ;
        RECT 601.950 900.600 604.050 901.050 ;
        RECT 595.950 899.400 604.050 900.600 ;
        RECT 595.950 898.950 598.050 899.400 ;
        RECT 601.950 898.950 604.050 899.400 ;
    END
  END Xout[5]
  PIN Xout[4]
    PORT
      LAYER metal2 ;
        RECT 1.950 421.950 4.050 424.050 ;
        RECT 2.400 412.050 3.450 421.950 ;
        RECT 1.950 409.950 4.050 412.050 ;
        RECT 56.400 411.900 57.600 412.650 ;
        RECT 55.950 409.800 58.050 411.900 ;
      LAYER metal3 ;
        RECT 1.950 423.600 4.050 424.050 ;
        RECT -3.600 422.400 4.050 423.600 ;
        RECT 1.950 421.950 4.050 422.400 ;
        RECT 1.950 411.600 4.050 412.050 ;
        RECT 55.950 411.600 58.050 411.900 ;
        RECT 1.950 410.400 58.050 411.600 ;
        RECT 1.950 409.950 4.050 410.400 ;
        RECT 55.950 409.800 58.050 410.400 ;
    END
  END Xout[4]
  PIN Xout[3]
    PORT
      LAYER metal2 ;
        RECT 14.400 567.900 15.600 568.650 ;
        RECT 13.950 565.800 16.050 567.900 ;
      LAYER metal3 ;
        RECT 13.950 567.600 16.050 567.900 ;
        RECT -3.600 566.400 16.050 567.600 ;
        RECT 13.950 565.800 16.050 566.400 ;
    END
  END Xout[3]
  PIN Xout[2]
    PORT
      LAYER metal2 ;
        RECT 14.400 723.900 15.600 724.650 ;
        RECT 13.950 721.800 16.050 723.900 ;
      LAYER metal3 ;
        RECT 13.950 723.600 16.050 723.900 ;
        RECT -3.600 722.400 16.050 723.600 ;
        RECT 13.950 721.800 16.050 722.400 ;
    END
  END Xout[2]
  PIN Xout[1]
    PORT
      LAYER metal2 ;
        RECT 35.400 411.000 36.600 412.650 ;
        RECT 34.950 406.950 37.050 411.000 ;
      LAYER metal3 ;
        RECT -3.600 408.600 -2.400 411.600 ;
        RECT 34.950 408.600 37.050 409.050 ;
        RECT -3.600 407.400 37.050 408.600 ;
        RECT 34.950 406.950 37.050 407.400 ;
    END
  END Xout[1]
  PIN Xout[0]
    PORT
      LAYER metal2 ;
        RECT 16.950 449.100 19.050 451.200 ;
        RECT 17.400 448.350 18.600 449.100 ;
      LAYER metal3 ;
        RECT 16.950 450.600 19.050 451.200 ;
        RECT -3.600 449.400 19.050 450.600 ;
        RECT 16.950 449.100 19.050 449.400 ;
    END
  END Xout[0]
  PIN Yin[15]
    PORT
      LAYER metal2 ;
        RECT 14.400 210.900 15.600 211.650 ;
        RECT 13.950 208.800 16.050 210.900 ;
      LAYER metal3 ;
        RECT -3.600 210.600 -2.400 216.600 ;
        RECT 13.950 210.600 16.050 210.900 ;
        RECT -3.600 209.400 16.050 210.600 ;
        RECT 13.950 208.800 16.050 209.400 ;
    END
  END Yin[15]
  PIN Yin[14]
    PORT
      LAYER metal2 ;
        RECT 7.950 268.950 10.050 271.050 ;
        RECT 16.950 268.950 19.050 271.050 ;
        RECT 88.950 268.950 91.050 271.050 ;
        RECT 8.400 256.050 9.450 268.950 ;
        RECT 17.400 261.600 18.450 268.950 ;
        RECT 89.400 262.200 90.450 268.950 ;
        RECT 17.400 259.350 18.600 261.600 ;
        RECT 88.950 260.100 91.050 262.200 ;
        RECT 94.950 260.100 97.050 262.200 ;
        RECT 89.400 259.350 90.600 260.100 ;
        RECT 95.400 256.050 96.450 260.100 ;
        RECT 7.950 253.950 10.050 256.050 ;
        RECT 94.950 253.950 97.050 256.050 ;
        RECT 104.400 255.900 105.600 256.650 ;
        RECT 103.950 253.800 106.050 255.900 ;
      LAYER metal3 ;
        RECT 7.950 270.600 10.050 271.050 ;
        RECT 16.950 270.600 19.050 271.050 ;
        RECT 88.950 270.600 91.050 271.050 ;
        RECT 7.950 269.400 91.050 270.600 ;
        RECT 7.950 268.950 10.050 269.400 ;
        RECT 16.950 268.950 19.050 269.400 ;
        RECT 88.950 268.950 91.050 269.400 ;
        RECT 88.950 261.750 91.050 262.200 ;
        RECT 94.950 261.750 97.050 262.200 ;
        RECT 88.950 260.550 97.050 261.750 ;
        RECT 88.950 260.100 91.050 260.550 ;
        RECT 94.950 260.100 97.050 260.550 ;
        RECT 7.950 255.600 10.050 256.050 ;
        RECT -3.600 254.400 10.050 255.600 ;
        RECT 7.950 253.950 10.050 254.400 ;
        RECT 94.950 255.600 97.050 256.050 ;
        RECT 103.950 255.600 106.050 255.900 ;
        RECT 94.950 254.400 106.050 255.600 ;
        RECT 94.950 253.950 97.050 254.400 ;
        RECT 103.950 253.800 106.050 254.400 ;
    END
  END Yin[14]
  PIN Yin[13]
    PORT
      LAYER metal2 ;
        RECT 14.400 176.400 15.600 178.650 ;
        RECT 14.400 171.450 15.450 176.400 ;
        RECT 11.400 170.400 15.450 171.450 ;
        RECT 11.400 139.050 12.450 170.400 ;
        RECT 10.950 136.950 13.050 139.050 ;
        RECT 11.400 132.450 12.450 136.950 ;
        RECT 14.400 132.450 15.600 133.650 ;
        RECT 11.400 131.400 15.600 132.450 ;
      LAYER metal3 ;
        RECT 10.950 138.600 13.050 139.050 ;
        RECT -3.600 137.400 13.050 138.600 ;
        RECT 10.950 136.950 13.050 137.400 ;
    END
  END Yin[13]
  PIN Yin[12]
    PORT
      LAYER metal2 ;
        RECT 16.950 26.100 19.050 28.200 ;
        RECT 17.400 25.350 18.600 26.100 ;
      LAYER metal3 ;
        RECT 16.950 27.600 19.050 28.200 ;
        RECT -3.600 26.400 19.050 27.600 ;
        RECT -3.600 20.400 -2.400 26.400 ;
        RECT 16.950 26.100 19.050 26.400 ;
    END
  END Yin[12]
  PIN Yin[11]
    PORT
      LAYER metal1 ;
        RECT 391.950 9.450 394.050 10.050 ;
        RECT 397.950 9.450 400.050 10.050 ;
        RECT 391.950 8.550 400.050 9.450 ;
        RECT 391.950 7.950 394.050 8.550 ;
        RECT 397.950 7.950 400.050 8.550 ;
      LAYER metal2 ;
        RECT 379.950 59.100 382.050 61.200 ;
        RECT 380.400 58.350 381.600 59.100 ;
        RECT 391.950 52.950 394.050 55.050 ;
        RECT 410.400 54.900 411.600 55.650 ;
        RECT 392.400 10.050 393.450 52.950 ;
        RECT 409.950 52.800 412.050 54.900 ;
        RECT 391.950 7.950 394.050 10.050 ;
        RECT 397.950 7.950 400.050 10.050 ;
        RECT 398.400 -3.600 399.450 7.950 ;
      LAYER metal3 ;
        RECT 379.950 59.100 382.050 61.200 ;
        RECT 380.400 54.600 381.600 59.100 ;
        RECT 391.950 54.600 394.050 55.050 ;
        RECT 409.950 54.600 412.050 54.900 ;
        RECT 380.400 53.400 412.050 54.600 ;
        RECT 391.950 52.950 394.050 53.400 ;
        RECT 409.950 52.800 412.050 53.400 ;
    END
  END Yin[11]
  PIN Yin[10]
    PORT
      LAYER metal2 ;
        RECT 389.400 132.000 390.600 133.650 ;
        RECT 388.950 127.950 391.050 132.000 ;
        RECT 448.950 127.950 451.050 130.050 ;
        RECT 449.400 82.050 450.450 127.950 ;
        RECT 448.950 79.950 451.050 82.050 ;
        RECT 460.950 79.950 463.050 82.050 ;
        RECT 461.400 4.050 462.450 79.950 ;
        RECT 476.400 20.400 477.600 22.650 ;
        RECT 476.400 4.050 477.450 20.400 ;
        RECT 460.950 1.950 463.050 4.050 ;
        RECT 466.950 1.950 469.050 4.050 ;
        RECT 475.950 1.950 478.050 4.050 ;
        RECT 467.400 -3.600 468.450 1.950 ;
      LAYER metal3 ;
        RECT 388.950 129.600 391.050 130.050 ;
        RECT 448.950 129.600 451.050 130.050 ;
        RECT 388.950 128.400 451.050 129.600 ;
        RECT 388.950 127.950 391.050 128.400 ;
        RECT 448.950 127.950 451.050 128.400 ;
        RECT 448.950 81.600 451.050 82.050 ;
        RECT 460.950 81.600 463.050 82.050 ;
        RECT 448.950 80.400 463.050 81.600 ;
        RECT 448.950 79.950 451.050 80.400 ;
        RECT 460.950 79.950 463.050 80.400 ;
        RECT 460.950 3.600 463.050 4.050 ;
        RECT 466.950 3.600 469.050 4.050 ;
        RECT 475.950 3.600 478.050 4.050 ;
        RECT 460.950 2.400 478.050 3.600 ;
        RECT 460.950 1.950 463.050 2.400 ;
        RECT 466.950 1.950 469.050 2.400 ;
        RECT 475.950 1.950 478.050 2.400 ;
    END
  END Yin[10]
  PIN Yin[9]
    PORT
      LAYER metal2 ;
        RECT 866.400 183.450 867.600 183.600 ;
        RECT 863.400 182.400 867.600 183.450 ;
        RECT 851.400 177.900 852.600 178.650 ;
        RECT 863.400 177.900 864.450 182.400 ;
        RECT 866.400 181.350 867.600 182.400 ;
        RECT 850.950 175.800 853.050 177.900 ;
        RECT 862.950 175.800 865.050 177.900 ;
      LAYER metal3 ;
        RECT 850.950 177.450 853.050 177.900 ;
        RECT 862.950 177.600 865.050 177.900 ;
        RECT 862.950 177.450 882.600 177.600 ;
        RECT 850.950 176.400 882.600 177.450 ;
        RECT 850.950 176.250 865.050 176.400 ;
        RECT 850.950 175.800 853.050 176.250 ;
        RECT 862.950 175.800 865.050 176.250 ;
        RECT 881.400 174.600 882.600 176.400 ;
        RECT 896.400 176.400 906.600 177.600 ;
        RECT 896.400 174.600 897.600 176.400 ;
        RECT 881.400 173.400 897.600 174.600 ;
    END
  END Yin[9]
  PIN Yin[8]
    PORT
      LAYER metal1 ;
        RECT 880.950 300.450 883.050 301.050 ;
        RECT 892.950 300.450 895.050 301.050 ;
        RECT 880.950 299.550 895.050 300.450 ;
        RECT 880.950 298.950 883.050 299.550 ;
        RECT 892.950 298.950 895.050 299.550 ;
      LAYER metal2 ;
        RECT 859.950 298.950 862.050 301.050 ;
        RECT 880.950 298.950 883.050 301.050 ;
        RECT 892.950 298.950 898.050 301.050 ;
        RECT 860.400 294.600 861.450 298.950 ;
        RECT 881.400 294.600 882.450 298.950 ;
        RECT 860.400 292.350 861.600 294.600 ;
        RECT 881.400 292.350 882.600 294.600 ;
      LAYER via2 ;
        RECT 895.950 298.950 898.050 301.050 ;
      LAYER metal3 ;
        RECT 859.950 300.600 862.050 301.050 ;
        RECT 880.950 300.600 883.050 301.050 ;
        RECT 859.950 299.400 883.050 300.600 ;
        RECT 859.950 298.950 862.050 299.400 ;
        RECT 880.950 298.950 883.050 299.400 ;
        RECT 895.950 300.600 898.050 301.050 ;
        RECT 895.950 299.400 906.600 300.600 ;
        RECT 895.950 298.950 898.050 299.400 ;
    END
  END Yin[8]
  PIN Yin[7]
    PORT
      LAYER metal2 ;
        RECT 865.950 371.100 868.050 373.200 ;
        RECT 871.950 371.100 874.050 373.200 ;
        RECT 854.400 365.400 855.600 367.650 ;
        RECT 854.400 358.050 855.450 365.400 ;
        RECT 866.400 358.050 867.450 371.100 ;
        RECT 872.400 370.350 873.600 371.100 ;
        RECT 853.950 355.950 856.050 358.050 ;
        RECT 865.950 355.950 868.050 358.050 ;
        RECT 871.950 355.950 874.050 358.050 ;
        RECT 857.400 333.900 858.600 334.650 ;
        RECT 856.950 331.800 859.050 333.900 ;
        RECT 872.400 331.050 873.450 355.950 ;
        RECT 881.400 333.900 882.600 334.650 ;
        RECT 871.950 328.950 874.050 331.050 ;
        RECT 880.950 328.950 883.050 333.900 ;
      LAYER via2 ;
        RECT 880.950 331.800 883.050 333.900 ;
      LAYER metal3 ;
        RECT 865.950 372.750 868.050 373.200 ;
        RECT 871.950 372.750 874.050 373.200 ;
        RECT 865.950 371.550 874.050 372.750 ;
        RECT 865.950 371.100 868.050 371.550 ;
        RECT 871.950 371.100 874.050 371.550 ;
        RECT 853.950 357.600 856.050 358.050 ;
        RECT 865.950 357.600 868.050 358.050 ;
        RECT 871.950 357.600 874.050 358.050 ;
        RECT 853.950 356.400 874.050 357.600 ;
        RECT 853.950 355.950 856.050 356.400 ;
        RECT 865.950 355.950 868.050 356.400 ;
        RECT 871.950 355.950 874.050 356.400 ;
        RECT 856.950 333.600 859.050 333.900 ;
        RECT 880.950 333.600 883.050 333.900 ;
        RECT 856.950 332.400 861.600 333.600 ;
        RECT 856.950 331.800 859.050 332.400 ;
        RECT 860.400 330.600 861.600 332.400 ;
        RECT 880.950 332.400 906.600 333.600 ;
        RECT 880.950 331.800 883.050 332.400 ;
        RECT 871.950 330.600 874.050 331.050 ;
        RECT 880.950 330.600 883.050 331.050 ;
        RECT 860.400 329.400 883.050 330.600 ;
        RECT 871.950 328.950 874.050 329.400 ;
        RECT 880.950 328.950 883.050 329.400 ;
    END
  END Yin[7]
  PIN Yin[6]
    PORT
      LAYER metal2 ;
        RECT 821.400 878.400 822.600 880.650 ;
        RECT 821.400 850.050 822.450 878.400 ;
        RECT 820.950 847.950 823.050 850.050 ;
        RECT 853.800 847.950 855.900 850.050 ;
        RECT 854.400 841.200 855.450 847.950 ;
        RECT 853.950 839.100 856.050 841.200 ;
        RECT 854.400 838.350 855.600 839.100 ;
        RECT 859.950 832.950 862.050 835.050 ;
        RECT 896.400 834.900 897.600 835.650 ;
        RECT 851.400 801.900 852.600 802.650 ;
        RECT 860.400 802.050 861.450 832.950 ;
        RECT 895.950 832.800 898.050 834.900 ;
        RECT 850.950 799.800 853.050 801.900 ;
        RECT 856.950 800.400 861.450 802.050 ;
        RECT 856.950 799.950 861.000 800.400 ;
      LAYER metal3 ;
        RECT 820.950 849.600 823.050 850.050 ;
        RECT 853.800 849.600 855.900 850.050 ;
        RECT 820.950 848.400 855.900 849.600 ;
        RECT 820.950 847.950 823.050 848.400 ;
        RECT 853.800 847.950 855.900 848.400 ;
        RECT 853.950 839.100 856.050 841.200 ;
        RECT 854.400 837.600 855.600 839.100 ;
        RECT 854.400 836.400 858.600 837.600 ;
        RECT 857.400 834.600 858.600 836.400 ;
        RECT 859.950 834.600 862.050 835.050 ;
        RECT 895.950 834.600 898.050 834.900 ;
        RECT 857.400 833.400 906.600 834.600 ;
        RECT 859.950 832.950 862.050 833.400 ;
        RECT 895.950 832.800 898.050 833.400 ;
        RECT 850.950 801.600 853.050 801.900 ;
        RECT 856.950 801.600 859.050 802.050 ;
        RECT 850.950 800.400 859.050 801.600 ;
        RECT 850.950 799.800 853.050 800.400 ;
        RECT 856.950 799.950 859.050 800.400 ;
    END
  END Yin[6]
  PIN Yin[5]
    PORT
      LAYER metal2 ;
        RECT 689.400 905.400 693.450 906.450 ;
        RECT 692.400 886.200 693.450 905.400 ;
        RECT 691.950 884.100 694.050 886.200 ;
        RECT 718.950 884.100 721.050 886.200 ;
        RECT 692.400 883.350 693.600 884.100 ;
        RECT 719.400 874.050 720.450 884.100 ;
        RECT 734.400 878.400 735.600 880.650 ;
        RECT 734.400 874.050 735.450 878.400 ;
        RECT 718.950 871.950 721.050 874.050 ;
        RECT 733.950 871.950 736.050 874.050 ;
        RECT 734.400 850.050 735.450 871.950 ;
        RECT 733.950 847.950 736.050 850.050 ;
        RECT 778.950 847.950 781.050 850.050 ;
        RECT 802.950 847.950 805.050 850.050 ;
        RECT 779.400 840.600 780.450 847.950 ;
        RECT 803.400 840.600 804.450 847.950 ;
        RECT 779.400 838.350 780.600 840.600 ;
        RECT 803.400 838.350 804.600 840.600 ;
      LAYER metal3 ;
        RECT 691.950 885.750 694.050 886.200 ;
        RECT 718.950 885.750 721.050 886.200 ;
        RECT 691.950 884.550 721.050 885.750 ;
        RECT 691.950 884.100 694.050 884.550 ;
        RECT 718.950 884.100 721.050 884.550 ;
        RECT 718.950 873.600 721.050 874.050 ;
        RECT 733.950 873.600 736.050 874.050 ;
        RECT 718.950 872.400 736.050 873.600 ;
        RECT 718.950 871.950 721.050 872.400 ;
        RECT 733.950 871.950 736.050 872.400 ;
        RECT 733.950 849.600 736.050 850.050 ;
        RECT 778.950 849.600 781.050 850.050 ;
        RECT 802.950 849.600 805.050 850.050 ;
        RECT 733.950 848.400 805.050 849.600 ;
        RECT 733.950 847.950 736.050 848.400 ;
        RECT 778.950 847.950 781.050 848.400 ;
        RECT 802.950 847.950 805.050 848.400 ;
    END
  END Yin[5]
  PIN Yin[4]
    PORT
      LAYER metal1 ;
        RECT 370.950 876.450 373.050 877.050 ;
        RECT 379.950 876.450 382.050 877.050 ;
        RECT 370.950 875.550 382.050 876.450 ;
        RECT 370.950 874.950 373.050 875.550 ;
        RECT 379.950 874.950 382.050 875.550 ;
      LAYER metal2 ;
        RECT 386.400 905.400 390.450 906.450 ;
        RECT 371.400 879.000 372.600 880.650 ;
        RECT 386.400 880.050 387.450 905.400 ;
        RECT 370.950 874.950 373.050 879.000 ;
        RECT 379.950 874.950 382.050 879.900 ;
        RECT 385.950 877.950 388.050 880.050 ;
        RECT 395.400 879.900 396.600 880.650 ;
        RECT 394.950 877.800 397.050 879.900 ;
      LAYER via2 ;
        RECT 379.950 877.800 382.050 879.900 ;
      LAYER metal3 ;
        RECT 379.950 879.450 382.050 879.900 ;
        RECT 385.950 879.450 388.050 880.050 ;
        RECT 394.950 879.450 397.050 879.900 ;
        RECT 379.950 878.250 397.050 879.450 ;
        RECT 379.950 877.800 382.050 878.250 ;
        RECT 385.950 877.950 388.050 878.250 ;
        RECT 394.950 877.800 397.050 878.250 ;
    END
  END Yin[4]
  PIN Yin[3]
    PORT
      LAYER metal2 ;
        RECT 61.950 839.100 64.050 841.200 ;
        RECT 62.400 838.350 63.600 839.100 ;
        RECT 67.950 838.950 70.050 841.050 ;
        RECT 82.950 839.100 85.050 841.200 ;
        RECT 106.950 839.100 109.050 841.200 ;
        RECT 1.950 835.950 4.050 838.050 ;
        RECT 2.400 832.050 3.450 835.950 ;
        RECT 14.400 834.000 15.600 835.650 ;
        RECT 1.950 829.950 4.050 832.050 ;
        RECT 13.950 829.950 16.050 834.000 ;
        RECT 68.400 832.050 69.450 838.950 ;
        RECT 83.400 838.350 84.600 839.100 ;
        RECT 107.400 838.350 108.600 839.100 ;
        RECT 67.950 829.950 70.050 832.050 ;
      LAYER metal3 ;
        RECT 61.950 840.600 64.050 841.200 ;
        RECT 67.950 840.600 70.050 841.050 ;
        RECT 82.950 840.600 85.050 841.200 ;
        RECT 106.950 840.600 109.050 841.200 ;
        RECT -3.600 837.600 -2.400 840.600 ;
        RECT 61.950 839.400 109.050 840.600 ;
        RECT 61.950 839.100 64.050 839.400 ;
        RECT 67.950 838.950 70.050 839.400 ;
        RECT 82.950 839.100 85.050 839.400 ;
        RECT 106.950 839.100 109.050 839.400 ;
        RECT 1.950 837.600 4.050 838.050 ;
        RECT -3.600 836.400 4.050 837.600 ;
        RECT 1.950 835.950 4.050 836.400 ;
        RECT 1.950 831.600 4.050 832.050 ;
        RECT 13.950 831.600 16.050 832.050 ;
        RECT 67.950 831.600 70.050 832.050 ;
        RECT 1.950 830.400 70.050 831.600 ;
        RECT 1.950 829.950 4.050 830.400 ;
        RECT 13.950 829.950 16.050 830.400 ;
        RECT 67.950 829.950 70.050 830.400 ;
    END
  END Yin[3]
  PIN Yin[2]
    PORT
      LAYER metal1 ;
        RECT 1.950 687.450 4.050 688.050 ;
        RECT 19.950 687.450 22.050 688.050 ;
        RECT 1.950 686.550 22.050 687.450 ;
        RECT 1.950 685.950 4.050 686.550 ;
        RECT 19.950 685.950 22.050 686.550 ;
      LAYER metal2 ;
        RECT 1.950 682.950 4.050 688.050 ;
        RECT 19.950 684.000 22.050 688.050 ;
        RECT 2.400 646.050 3.450 682.950 ;
        RECT 20.400 682.350 21.600 684.000 ;
        RECT 1.950 643.950 4.050 646.050 ;
        RECT 20.400 645.900 21.600 646.650 ;
        RECT 19.950 643.800 22.050 645.900 ;
      LAYER metal3 ;
        RECT 1.950 684.600 4.050 685.050 ;
        RECT -3.600 683.400 4.050 684.600 ;
        RECT 1.950 682.950 4.050 683.400 ;
        RECT 1.950 645.600 4.050 646.050 ;
        RECT 19.950 645.600 22.050 645.900 ;
        RECT 1.950 644.400 22.050 645.600 ;
        RECT 1.950 643.950 4.050 644.400 ;
        RECT 19.950 643.800 22.050 644.400 ;
    END
  END Yin[2]
  PIN Yin[1]
    PORT
      LAYER metal1 ;
        RECT 76.950 486.450 79.050 487.050 ;
        RECT 103.950 486.450 106.050 487.050 ;
        RECT 76.950 485.550 106.050 486.450 ;
        RECT 76.950 484.950 79.050 485.550 ;
        RECT 103.950 484.950 106.050 485.550 ;
      LAYER metal2 ;
        RECT 1.950 487.950 4.050 490.050 ;
        RECT 77.400 489.000 78.600 490.650 ;
        RECT 104.400 489.000 105.600 490.650 ;
        RECT 2.400 484.050 3.450 487.950 ;
        RECT 1.950 481.950 4.050 484.050 ;
        RECT 76.950 481.950 79.050 489.000 ;
        RECT 103.950 484.950 106.050 489.000 ;
      LAYER metal3 ;
        RECT 1.950 489.600 4.050 490.050 ;
        RECT -3.600 488.400 4.050 489.600 ;
        RECT 1.950 487.950 4.050 488.400 ;
        RECT 1.950 483.600 4.050 484.050 ;
        RECT 76.950 483.600 79.050 484.050 ;
        RECT 1.950 482.400 79.050 483.600 ;
        RECT 1.950 481.950 4.050 482.400 ;
        RECT 76.950 481.950 79.050 482.400 ;
    END
  END Yin[1]
  PIN Yin[0]
    PORT
      LAYER metal2 ;
        RECT 85.950 604.950 88.050 607.050 ;
        RECT 91.950 605.100 94.050 607.200 ;
        RECT 71.400 600.900 72.600 601.650 ;
        RECT 86.400 600.900 87.450 604.950 ;
        RECT 92.400 604.350 93.600 605.100 ;
        RECT 70.950 598.800 73.050 600.900 ;
        RECT 85.950 598.800 88.050 600.900 ;
      LAYER metal3 ;
        RECT 85.950 606.600 88.050 607.050 ;
        RECT 91.950 606.600 94.050 607.200 ;
        RECT 85.950 605.400 94.050 606.600 ;
        RECT 85.950 604.950 88.050 605.400 ;
        RECT 91.950 605.100 94.050 605.400 ;
        RECT 70.950 600.600 73.050 600.900 ;
        RECT -3.600 600.450 73.050 600.600 ;
        RECT 85.950 600.450 88.050 600.900 ;
        RECT -3.600 599.400 88.050 600.450 ;
        RECT 70.950 599.250 88.050 599.400 ;
        RECT 70.950 598.800 73.050 599.250 ;
        RECT 85.950 598.800 88.050 599.250 ;
    END
  END Yin[0]
  PIN Yout[15]
    PORT
      LAYER metal2 ;
        RECT 1.950 337.950 4.050 340.050 ;
        RECT 2.400 328.050 3.450 337.950 ;
        RECT 38.400 332.400 39.600 334.650 ;
        RECT 38.400 328.050 39.450 332.400 ;
        RECT 1.950 325.950 4.050 328.050 ;
        RECT 37.950 325.950 40.050 328.050 ;
      LAYER metal3 ;
        RECT 1.950 339.600 4.050 340.050 ;
        RECT -3.600 338.400 4.050 339.600 ;
        RECT 1.950 337.950 4.050 338.400 ;
        RECT 1.950 327.600 4.050 328.050 ;
        RECT 37.950 327.600 40.050 328.050 ;
        RECT 1.950 326.400 40.050 327.600 ;
        RECT 1.950 325.950 4.050 326.400 ;
        RECT 37.950 325.950 40.050 326.400 ;
    END
  END Yout[15]
  PIN Yout[14]
    PORT
      LAYER metal2 ;
        RECT 17.400 333.900 18.600 334.650 ;
        RECT 16.950 331.800 19.050 333.900 ;
      LAYER metal3 ;
        RECT 16.950 333.600 19.050 333.900 ;
        RECT -3.600 332.400 19.050 333.600 ;
        RECT 16.950 331.800 19.050 332.400 ;
    END
  END Yout[14]
  PIN Yout[13]
    PORT
      LAYER metal2 ;
        RECT 341.400 20.400 342.600 22.650 ;
        RECT 341.400 -2.550 342.450 20.400 ;
        RECT 338.400 -3.600 342.450 -2.550 ;
    END
  END Yout[13]
  PIN Yout[12]
    PORT
      LAYER metal2 ;
        RECT 356.400 20.400 357.600 22.650 ;
        RECT 356.400 -2.550 357.450 20.400 ;
        RECT 356.400 -3.600 360.450 -2.550 ;
    END
  END Yout[12]
  PIN Yout[11]
    PORT
      LAYER metal2 ;
        RECT 779.400 20.400 780.600 22.650 ;
        RECT 779.400 -2.550 780.450 20.400 ;
        RECT 776.400 -3.600 780.450 -2.550 ;
    END
  END Yout[11]
  PIN Yout[10]
    PORT
      LAYER metal1 ;
        RECT 553.950 63.450 556.050 64.050 ;
        RECT 565.950 63.450 568.050 64.050 ;
        RECT 553.950 62.550 568.050 63.450 ;
        RECT 553.950 61.950 556.050 62.550 ;
        RECT 565.950 61.950 568.050 62.550 ;
      LAYER metal2 ;
        RECT 553.950 214.950 556.050 217.050 ;
        RECT 562.950 215.100 565.050 217.200 ;
        RECT 554.400 142.050 555.450 214.950 ;
        RECT 563.400 214.350 564.600 215.100 ;
        RECT 553.950 139.950 556.050 142.050 ;
        RECT 562.950 139.950 565.050 142.050 ;
        RECT 563.400 105.450 564.450 139.950 ;
        RECT 563.400 104.400 567.450 105.450 ;
        RECT 566.400 64.050 567.450 104.400 ;
        RECT 553.950 61.950 556.050 64.050 ;
        RECT 565.950 61.950 568.050 64.050 ;
        RECT 554.400 4.050 555.450 61.950 ;
        RECT 553.950 1.950 556.050 4.050 ;
        RECT 565.950 1.950 568.050 4.050 ;
        RECT 566.400 -3.600 567.450 1.950 ;
      LAYER metal3 ;
        RECT 553.950 216.600 556.050 217.050 ;
        RECT 562.950 216.600 565.050 217.200 ;
        RECT 553.950 215.400 565.050 216.600 ;
        RECT 553.950 214.950 556.050 215.400 ;
        RECT 562.950 215.100 565.050 215.400 ;
        RECT 553.950 141.600 556.050 142.050 ;
        RECT 562.950 141.600 565.050 142.050 ;
        RECT 553.950 140.400 565.050 141.600 ;
        RECT 553.950 139.950 556.050 140.400 ;
        RECT 562.950 139.950 565.050 140.400 ;
        RECT 553.950 3.600 556.050 4.050 ;
        RECT 565.950 3.600 568.050 4.050 ;
        RECT 553.950 2.400 568.050 3.600 ;
        RECT 553.950 1.950 556.050 2.400 ;
        RECT 565.950 1.950 568.050 2.400 ;
    END
  END Yout[10]
  PIN Yout[9]
    PORT
      LAYER metal2 ;
        RECT 500.400 901.050 501.450 906.450 ;
        RECT 493.950 898.950 496.050 901.050 ;
        RECT 499.950 898.950 502.050 901.050 ;
        RECT 494.400 879.450 495.450 898.950 ;
        RECT 497.400 879.450 498.600 880.650 ;
        RECT 494.400 878.400 498.600 879.450 ;
      LAYER metal3 ;
        RECT 493.950 900.600 496.050 901.050 ;
        RECT 499.950 900.600 502.050 901.050 ;
        RECT 493.950 899.400 502.050 900.600 ;
        RECT 493.950 898.950 496.050 899.400 ;
        RECT 499.950 898.950 502.050 899.400 ;
    END
  END Yout[9]
  PIN Yout[8]
    PORT
      LAYER metal2 ;
        RECT 13.950 376.950 16.050 379.050 ;
        RECT 14.400 372.600 15.450 376.950 ;
        RECT 14.400 370.350 15.600 372.600 ;
      LAYER metal3 ;
        RECT 13.950 378.600 16.050 379.050 ;
        RECT -3.600 377.400 16.050 378.600 ;
        RECT 13.950 376.950 16.050 377.400 ;
    END
  END Yout[8]
  PIN Yout[7]
    PORT
      LAYER metal1 ;
        RECT 451.950 729.450 454.050 730.050 ;
        RECT 457.950 729.450 460.050 729.900 ;
        RECT 451.950 728.550 460.050 729.450 ;
        RECT 451.950 727.950 454.050 728.550 ;
        RECT 457.950 727.800 460.050 728.550 ;
      LAYER metal2 ;
        RECT 470.400 802.050 471.450 906.450 ;
        RECT 442.950 799.950 445.050 802.050 ;
        RECT 469.950 799.950 472.050 802.050 ;
        RECT 443.400 751.050 444.450 799.950 ;
        RECT 442.950 748.950 445.050 751.050 ;
        RECT 451.950 748.950 454.050 751.050 ;
        RECT 452.400 730.050 453.450 748.950 ;
        RECT 451.950 727.950 454.050 730.050 ;
        RECT 457.950 727.800 460.050 729.900 ;
        RECT 458.400 715.050 459.450 727.800 ;
        RECT 457.950 712.950 460.050 715.050 ;
        RECT 466.950 712.950 469.050 715.050 ;
        RECT 467.400 684.600 468.450 712.950 ;
        RECT 467.400 682.350 468.600 684.600 ;
      LAYER metal3 ;
        RECT 442.950 801.600 445.050 802.050 ;
        RECT 469.950 801.600 472.050 802.050 ;
        RECT 442.950 800.400 472.050 801.600 ;
        RECT 442.950 799.950 445.050 800.400 ;
        RECT 469.950 799.950 472.050 800.400 ;
        RECT 442.950 750.600 445.050 751.050 ;
        RECT 451.950 750.600 454.050 751.050 ;
        RECT 442.950 749.400 454.050 750.600 ;
        RECT 442.950 748.950 445.050 749.400 ;
        RECT 451.950 748.950 454.050 749.400 ;
        RECT 457.950 714.600 460.050 715.050 ;
        RECT 466.950 714.600 469.050 715.050 ;
        RECT 457.950 713.400 469.050 714.600 ;
        RECT 457.950 712.950 460.050 713.400 ;
        RECT 466.950 712.950 469.050 713.400 ;
    END
  END Yout[7]
  PIN Yout[6]
    PORT
      LAYER metal2 ;
        RECT 419.400 898.050 420.450 906.450 ;
        RECT 412.950 895.950 415.050 898.050 ;
        RECT 418.950 895.950 421.050 898.050 ;
        RECT 413.400 879.450 414.450 895.950 ;
        RECT 416.400 879.450 417.600 880.650 ;
        RECT 413.400 878.400 417.600 879.450 ;
      LAYER metal3 ;
        RECT 412.950 897.600 415.050 898.050 ;
        RECT 418.950 897.600 421.050 898.050 ;
        RECT 412.950 896.400 421.050 897.600 ;
        RECT 412.950 895.950 415.050 896.400 ;
        RECT 418.950 895.950 421.050 896.400 ;
    END
  END Yout[6]
  PIN Yout[5]
    PORT
      LAYER metal2 ;
        RECT 350.400 905.400 354.450 906.450 ;
        RECT 350.400 879.450 351.600 880.650 ;
        RECT 353.400 879.450 354.450 905.400 ;
        RECT 350.400 878.400 354.450 879.450 ;
    END
  END Yout[5]
  PIN Yout[4]
    PORT
      LAYER metal2 ;
        RECT 251.400 889.050 252.450 906.450 ;
        RECT 250.950 886.950 253.050 889.050 ;
        RECT 254.400 879.900 255.600 880.650 ;
        RECT 253.950 877.800 256.050 879.900 ;
      LAYER metal3 ;
        RECT 250.950 886.950 253.050 889.050 ;
        RECT 251.400 879.600 252.600 886.950 ;
        RECT 253.950 879.600 256.050 879.900 ;
        RECT 251.400 878.400 256.050 879.600 ;
        RECT 253.950 877.800 256.050 878.400 ;
    END
  END Yout[4]
  PIN Yout[3]
    PORT
      LAYER metal2 ;
        RECT 62.400 901.050 63.450 906.450 ;
        RECT 55.950 898.950 58.050 901.050 ;
        RECT 61.950 898.950 64.050 901.050 ;
        RECT 56.400 879.450 57.450 898.950 ;
        RECT 59.400 879.450 60.600 880.650 ;
        RECT 56.400 878.400 60.600 879.450 ;
      LAYER metal3 ;
        RECT 55.950 900.600 58.050 901.050 ;
        RECT 61.950 900.600 64.050 901.050 ;
        RECT 55.950 899.400 64.050 900.600 ;
        RECT 55.950 898.950 58.050 899.400 ;
        RECT 61.950 898.950 64.050 899.400 ;
    END
  END Yout[3]
  PIN Yout[2]
    PORT
      LAYER metal2 ;
        RECT 10.950 493.950 13.050 496.050 ;
        RECT 11.400 489.450 12.450 493.950 ;
        RECT 14.400 489.450 15.600 490.650 ;
        RECT 11.400 488.400 15.600 489.450 ;
      LAYER metal3 ;
        RECT 10.950 495.600 13.050 496.050 ;
        RECT -3.600 494.400 13.050 495.600 ;
        RECT 10.950 493.950 13.050 494.400 ;
    END
  END Yout[2]
  PIN Yout[1]
    PORT
      LAYER metal2 ;
        RECT 13.950 527.100 16.050 529.200 ;
        RECT 14.400 526.350 15.600 527.100 ;
      LAYER metal3 ;
        RECT 13.950 528.600 16.050 529.200 ;
        RECT -3.600 527.400 16.050 528.600 ;
        RECT 13.950 527.100 16.050 527.400 ;
    END
  END Yout[1]
  PIN Yout[0]
    PORT
      LAYER metal2 ;
        RECT 13.950 605.100 16.050 607.200 ;
        RECT 14.400 604.350 15.600 605.100 ;
      LAYER metal3 ;
        RECT 13.950 606.600 16.050 607.200 ;
        RECT -3.600 605.400 16.050 606.600 ;
        RECT 13.950 605.100 16.050 605.400 ;
    END
  END Yout[0]
  PIN clk
    PORT
      LAYER metal2 ;
        RECT 131.400 901.050 132.450 906.450 ;
        RECT 130.950 898.950 133.050 901.050 ;
        RECT 178.950 898.950 181.050 901.050 ;
        RECT 463.950 898.950 466.050 901.050 ;
        RECT 131.400 879.900 132.450 898.950 ;
        RECT 137.400 879.900 138.600 880.650 ;
        RECT 130.950 877.800 133.050 879.900 ;
        RECT 136.950 877.800 139.050 879.900 ;
        RECT 179.400 856.050 180.450 898.950 ;
        RECT 178.950 853.950 181.050 856.050 ;
        RECT 196.950 853.950 199.050 856.050 ;
        RECT 197.400 742.050 198.450 853.950 ;
        RECT 464.400 840.600 465.450 898.950 ;
        RECT 464.400 838.350 465.600 840.600 ;
        RECT 187.950 739.950 190.050 742.050 ;
        RECT 196.950 739.950 199.050 742.050 ;
        RECT 188.400 676.050 189.450 739.950 ;
        RECT 187.950 673.950 190.050 676.050 ;
        RECT 235.950 673.950 238.050 676.050 ;
        RECT 236.400 532.050 237.450 673.950 ;
        RECT 193.950 529.950 196.050 532.050 ;
        RECT 188.400 489.900 189.600 490.650 ;
        RECT 194.400 489.900 195.450 529.950 ;
        RECT 217.950 528.000 220.050 532.050 ;
        RECT 235.950 529.950 238.050 532.050 ;
        RECT 218.400 526.350 219.600 528.000 ;
        RECT 187.950 487.800 190.050 489.900 ;
        RECT 193.950 487.800 196.050 489.900 ;
        RECT 188.400 411.900 189.600 412.650 ;
        RECT 194.400 411.900 195.450 487.800 ;
        RECT 227.400 411.900 228.600 412.650 ;
        RECT 187.950 409.800 190.050 411.900 ;
        RECT 193.950 409.800 196.050 411.900 ;
        RECT 226.950 409.800 229.050 411.900 ;
      LAYER via2 ;
        RECT 217.950 529.950 220.050 532.050 ;
      LAYER metal3 ;
        RECT 130.950 900.600 133.050 901.050 ;
        RECT 178.950 900.600 181.050 901.050 ;
        RECT 463.950 900.600 466.050 901.050 ;
        RECT 130.950 899.400 466.050 900.600 ;
        RECT 130.950 898.950 133.050 899.400 ;
        RECT 178.950 898.950 181.050 899.400 ;
        RECT 463.950 898.950 466.050 899.400 ;
        RECT 130.950 879.450 133.050 879.900 ;
        RECT 136.950 879.450 139.050 879.900 ;
        RECT 130.950 878.250 139.050 879.450 ;
        RECT 130.950 877.800 133.050 878.250 ;
        RECT 136.950 877.800 139.050 878.250 ;
        RECT 178.950 855.600 181.050 856.050 ;
        RECT 196.950 855.600 199.050 856.050 ;
        RECT 178.950 854.400 199.050 855.600 ;
        RECT 178.950 853.950 181.050 854.400 ;
        RECT 196.950 853.950 199.050 854.400 ;
        RECT 187.950 741.600 190.050 742.050 ;
        RECT 196.950 741.600 199.050 742.050 ;
        RECT 187.950 740.400 199.050 741.600 ;
        RECT 187.950 739.950 190.050 740.400 ;
        RECT 196.950 739.950 199.050 740.400 ;
        RECT 187.950 675.600 190.050 676.050 ;
        RECT 235.950 675.600 238.050 676.050 ;
        RECT 187.950 674.400 238.050 675.600 ;
        RECT 187.950 673.950 190.050 674.400 ;
        RECT 235.950 673.950 238.050 674.400 ;
        RECT 193.950 531.600 196.050 532.050 ;
        RECT 217.950 531.600 220.050 532.050 ;
        RECT 235.950 531.600 238.050 532.050 ;
        RECT 193.950 530.400 238.050 531.600 ;
        RECT 193.950 529.950 196.050 530.400 ;
        RECT 217.950 529.950 220.050 530.400 ;
        RECT 235.950 529.950 238.050 530.400 ;
        RECT 187.950 489.450 190.050 489.900 ;
        RECT 193.950 489.450 196.050 489.900 ;
        RECT 187.950 488.250 196.050 489.450 ;
        RECT 187.950 487.800 190.050 488.250 ;
        RECT 193.950 487.800 196.050 488.250 ;
        RECT 187.950 411.450 190.050 411.900 ;
        RECT 193.950 411.600 196.050 411.900 ;
        RECT 226.950 411.600 229.050 411.900 ;
        RECT 193.950 411.450 229.050 411.600 ;
        RECT 187.950 410.400 229.050 411.450 ;
        RECT 187.950 410.250 196.050 410.400 ;
        RECT 187.950 409.800 190.050 410.250 ;
        RECT 193.950 409.800 196.050 410.250 ;
        RECT 226.950 409.800 229.050 410.400 ;
    END
  END clk
  OBS
      LAYER metal1 ;
        RECT 17.100 890.400 18.900 896.400 ;
        RECT 20.100 890.400 21.900 897.000 ;
        RECT 23.100 893.400 24.900 896.400 ;
        RECT 17.100 883.050 18.300 890.400 ;
        RECT 23.700 889.500 24.900 893.400 ;
        RECT 19.200 888.600 24.900 889.500 ;
        RECT 38.700 889.200 40.500 896.400 ;
        RECT 43.800 890.400 45.600 897.000 ;
        RECT 59.100 890.400 60.900 896.400 ;
        RECT 62.100 890.400 63.900 897.000 ;
        RECT 65.100 893.400 66.900 896.400 ;
        RECT 19.200 887.700 21.000 888.600 ;
        RECT 38.700 888.300 42.900 889.200 ;
        RECT 17.100 880.950 19.200 883.050 ;
        RECT 17.100 873.600 18.300 880.950 ;
        RECT 20.100 876.300 21.000 887.700 ;
        RECT 38.100 883.050 39.900 884.850 ;
        RECT 41.700 883.050 42.900 888.300 ;
        RECT 43.950 883.050 45.750 884.850 ;
        RECT 59.100 883.050 60.300 890.400 ;
        RECT 65.700 889.500 66.900 893.400 ;
        RECT 61.200 888.600 66.900 889.500 ;
        RECT 68.550 890.400 70.350 896.400 ;
        RECT 71.850 890.400 73.650 897.000 ;
        RECT 76.950 893.400 78.750 896.400 ;
        RECT 81.450 893.400 83.250 897.000 ;
        RECT 84.450 893.400 86.250 896.400 ;
        RECT 87.750 893.400 89.550 897.000 ;
        RECT 92.250 894.300 94.050 896.400 ;
        RECT 92.250 893.400 95.850 894.300 ;
        RECT 76.350 891.300 78.750 893.400 ;
        RECT 85.200 892.500 86.250 893.400 ;
        RECT 92.250 892.800 96.150 893.400 ;
        RECT 85.200 891.450 90.150 892.500 ;
        RECT 88.350 890.700 90.150 891.450 ;
        RECT 61.200 887.700 63.000 888.600 ;
        RECT 22.500 880.950 24.600 883.050 ;
        RECT 37.950 880.950 40.050 883.050 ;
        RECT 40.950 880.950 43.050 883.050 ;
        RECT 43.950 880.950 46.050 883.050 ;
        RECT 59.100 880.950 61.200 883.050 ;
        RECT 22.800 879.150 24.600 880.950 ;
        RECT 19.200 875.400 21.000 876.300 ;
        RECT 19.200 874.500 24.900 875.400 ;
        RECT 17.100 861.600 18.900 873.600 ;
        RECT 20.100 861.000 21.900 871.800 ;
        RECT 23.700 867.600 24.900 874.500 ;
        RECT 41.700 867.600 42.900 880.950 ;
        RECT 59.100 873.600 60.300 880.950 ;
        RECT 62.100 876.300 63.000 887.700 ;
        RECT 68.550 883.050 69.750 890.400 ;
        RECT 91.350 889.800 93.150 891.600 ;
        RECT 94.050 891.300 96.150 892.800 ;
        RECT 97.050 890.400 98.850 897.000 ;
        RECT 100.050 892.200 101.850 896.400 ;
        RECT 100.050 890.400 102.450 892.200 ;
        RECT 116.100 890.400 117.900 897.000 ;
        RECT 81.150 888.000 82.950 888.600 ;
        RECT 92.100 888.000 93.150 889.800 ;
        RECT 81.150 886.800 93.150 888.000 ;
        RECT 64.500 880.950 66.600 883.050 ;
        RECT 64.800 879.150 66.600 880.950 ;
        RECT 68.550 881.250 74.850 883.050 ;
        RECT 68.550 880.950 73.050 881.250 ;
        RECT 61.200 875.400 63.000 876.300 ;
        RECT 61.200 874.500 66.900 875.400 ;
        RECT 23.100 861.600 24.900 867.600 ;
        RECT 38.100 861.000 39.900 867.600 ;
        RECT 41.100 861.600 42.900 867.600 ;
        RECT 44.100 861.000 45.900 867.600 ;
        RECT 59.100 861.600 60.900 873.600 ;
        RECT 62.100 861.000 63.900 871.800 ;
        RECT 65.700 867.600 66.900 874.500 ;
        RECT 65.100 861.600 66.900 867.600 ;
        RECT 68.550 873.600 69.750 880.950 ;
        RECT 70.650 878.100 72.450 878.250 ;
        RECT 76.350 878.100 78.450 878.400 ;
        RECT 70.650 876.900 78.450 878.100 ;
        RECT 70.650 876.450 72.450 876.900 ;
        RECT 76.350 876.300 78.450 876.900 ;
        RECT 81.150 874.200 82.050 886.800 ;
        RECT 92.100 885.600 100.050 886.800 ;
        RECT 92.100 885.000 93.900 885.600 ;
        RECT 95.100 883.800 96.900 884.400 ;
        RECT 88.800 882.600 96.900 883.800 ;
        RECT 98.250 883.050 100.050 885.600 ;
        RECT 88.800 880.950 90.900 882.600 ;
        RECT 97.950 880.950 100.050 883.050 ;
        RECT 90.750 875.700 92.550 876.000 ;
        RECT 101.550 875.700 102.450 890.400 ;
        RECT 119.100 889.500 120.900 896.400 ;
        RECT 122.100 890.400 123.900 897.000 ;
        RECT 125.100 889.500 126.900 896.400 ;
        RECT 128.100 890.400 129.900 897.000 ;
        RECT 131.100 889.500 132.900 896.400 ;
        RECT 134.100 890.400 135.900 897.000 ;
        RECT 137.100 889.500 138.900 896.400 ;
        RECT 140.100 890.400 141.900 897.000 ;
        RECT 155.100 890.400 156.900 896.400 ;
        RECT 158.100 890.400 159.900 897.000 ;
        RECT 161.100 893.400 162.900 896.400 ;
        RECT 90.750 875.100 102.450 875.700 ;
        RECT 68.550 861.600 70.350 873.600 ;
        RECT 71.550 861.000 73.350 873.600 ;
        RECT 77.250 873.300 82.050 874.200 ;
        RECT 84.150 874.500 102.450 875.100 ;
        RECT 118.050 888.300 120.900 889.500 ;
        RECT 123.000 888.300 126.900 889.500 ;
        RECT 129.000 888.300 132.900 889.500 ;
        RECT 135.000 888.300 138.900 889.500 ;
        RECT 118.050 883.050 119.100 888.300 ;
        RECT 123.000 887.400 124.200 888.300 ;
        RECT 129.000 887.400 130.200 888.300 ;
        RECT 135.000 887.400 136.200 888.300 ;
        RECT 120.000 886.200 124.200 887.400 ;
        RECT 120.000 885.600 121.800 886.200 ;
        RECT 118.050 880.950 121.200 883.050 ;
        RECT 118.050 875.700 119.100 880.950 ;
        RECT 123.000 875.700 124.200 886.200 ;
        RECT 126.000 886.200 130.200 887.400 ;
        RECT 126.000 885.600 127.800 886.200 ;
        RECT 129.000 875.700 130.200 886.200 ;
        RECT 132.000 886.200 136.200 887.400 ;
        RECT 132.000 885.600 133.800 886.200 ;
        RECT 135.000 875.700 136.200 886.200 ;
        RECT 137.400 883.050 139.200 884.850 ;
        RECT 137.100 880.950 139.200 883.050 ;
        RECT 155.100 883.050 156.300 890.400 ;
        RECT 161.700 889.500 162.900 893.400 ;
        RECT 157.200 888.600 162.900 889.500 ;
        RECT 164.550 890.400 166.350 896.400 ;
        RECT 167.850 890.400 169.650 897.000 ;
        RECT 172.950 893.400 174.750 896.400 ;
        RECT 177.450 893.400 179.250 897.000 ;
        RECT 180.450 893.400 182.250 896.400 ;
        RECT 183.750 893.400 185.550 897.000 ;
        RECT 188.250 894.300 190.050 896.400 ;
        RECT 188.250 893.400 191.850 894.300 ;
        RECT 172.350 891.300 174.750 893.400 ;
        RECT 181.200 892.500 182.250 893.400 ;
        RECT 188.250 892.800 192.150 893.400 ;
        RECT 181.200 891.450 186.150 892.500 ;
        RECT 184.350 890.700 186.150 891.450 ;
        RECT 157.200 887.700 159.000 888.600 ;
        RECT 155.100 880.950 157.200 883.050 ;
        RECT 118.050 874.500 120.900 875.700 ;
        RECT 123.000 874.500 126.900 875.700 ;
        RECT 129.000 874.500 132.900 875.700 ;
        RECT 135.000 874.500 138.900 875.700 ;
        RECT 84.150 874.200 92.550 874.500 ;
        RECT 77.250 872.400 78.450 873.300 ;
        RECT 75.450 870.600 78.450 872.400 ;
        RECT 79.350 872.100 81.150 872.400 ;
        RECT 84.150 872.100 85.050 874.200 ;
        RECT 101.550 873.600 102.450 874.500 ;
        RECT 79.350 871.200 85.050 872.100 ;
        RECT 85.950 872.700 87.750 873.300 ;
        RECT 85.950 871.500 93.750 872.700 ;
        RECT 79.350 870.600 81.150 871.200 ;
        RECT 91.650 870.600 93.750 871.500 ;
        RECT 76.350 867.600 78.450 869.700 ;
        RECT 82.950 869.550 84.750 870.300 ;
        RECT 87.750 869.550 89.550 870.300 ;
        RECT 82.950 868.500 89.550 869.550 ;
        RECT 76.350 861.600 78.150 867.600 ;
        RECT 80.850 861.000 82.650 867.600 ;
        RECT 83.850 861.600 85.650 868.500 ;
        RECT 86.850 861.000 88.650 867.600 ;
        RECT 91.650 861.600 93.450 870.600 ;
        RECT 97.050 861.000 98.850 873.600 ;
        RECT 100.050 871.800 102.450 873.600 ;
        RECT 100.050 861.600 101.850 871.800 ;
        RECT 116.100 861.000 117.900 873.600 ;
        RECT 119.100 861.600 120.900 874.500 ;
        RECT 122.100 861.000 123.900 873.600 ;
        RECT 125.100 861.600 126.900 874.500 ;
        RECT 128.100 861.000 129.900 873.600 ;
        RECT 131.100 861.600 132.900 874.500 ;
        RECT 134.100 861.000 135.900 873.600 ;
        RECT 137.100 861.600 138.900 874.500 ;
        RECT 155.100 873.600 156.300 880.950 ;
        RECT 158.100 876.300 159.000 887.700 ;
        RECT 164.550 883.050 165.750 890.400 ;
        RECT 187.350 889.800 189.150 891.600 ;
        RECT 190.050 891.300 192.150 892.800 ;
        RECT 193.050 890.400 194.850 897.000 ;
        RECT 196.050 892.200 197.850 896.400 ;
        RECT 201.150 892.200 202.950 896.400 ;
        RECT 196.050 890.400 198.450 892.200 ;
        RECT 177.150 888.000 178.950 888.600 ;
        RECT 188.100 888.000 189.150 889.800 ;
        RECT 177.150 886.800 189.150 888.000 ;
        RECT 160.500 880.950 162.600 883.050 ;
        RECT 160.800 879.150 162.600 880.950 ;
        RECT 164.550 881.250 170.850 883.050 ;
        RECT 164.550 880.950 169.050 881.250 ;
        RECT 157.200 875.400 159.000 876.300 ;
        RECT 157.200 874.500 162.900 875.400 ;
        RECT 140.100 861.000 141.900 873.600 ;
        RECT 155.100 861.600 156.900 873.600 ;
        RECT 158.100 861.000 159.900 871.800 ;
        RECT 161.700 867.600 162.900 874.500 ;
        RECT 161.100 861.600 162.900 867.600 ;
        RECT 164.550 873.600 165.750 880.950 ;
        RECT 166.650 878.100 168.450 878.250 ;
        RECT 172.350 878.100 174.450 878.400 ;
        RECT 166.650 876.900 174.450 878.100 ;
        RECT 166.650 876.450 168.450 876.900 ;
        RECT 172.350 876.300 174.450 876.900 ;
        RECT 177.150 874.200 178.050 886.800 ;
        RECT 188.100 885.600 196.050 886.800 ;
        RECT 188.100 885.000 189.900 885.600 ;
        RECT 191.100 883.800 192.900 884.400 ;
        RECT 184.800 882.600 192.900 883.800 ;
        RECT 194.250 883.050 196.050 885.600 ;
        RECT 184.800 880.950 186.900 882.600 ;
        RECT 193.950 880.950 196.050 883.050 ;
        RECT 186.750 875.700 188.550 876.000 ;
        RECT 197.550 875.700 198.450 890.400 ;
        RECT 186.750 875.100 198.450 875.700 ;
        RECT 164.550 861.600 166.350 873.600 ;
        RECT 167.550 861.000 169.350 873.600 ;
        RECT 173.250 873.300 178.050 874.200 ;
        RECT 180.150 874.500 198.450 875.100 ;
        RECT 180.150 874.200 188.550 874.500 ;
        RECT 173.250 872.400 174.450 873.300 ;
        RECT 171.450 870.600 174.450 872.400 ;
        RECT 175.350 872.100 177.150 872.400 ;
        RECT 180.150 872.100 181.050 874.200 ;
        RECT 197.550 873.600 198.450 874.500 ;
        RECT 175.350 871.200 181.050 872.100 ;
        RECT 181.950 872.700 183.750 873.300 ;
        RECT 181.950 871.500 189.750 872.700 ;
        RECT 175.350 870.600 177.150 871.200 ;
        RECT 187.650 870.600 189.750 871.500 ;
        RECT 172.350 867.600 174.450 869.700 ;
        RECT 178.950 869.550 180.750 870.300 ;
        RECT 183.750 869.550 185.550 870.300 ;
        RECT 178.950 868.500 185.550 869.550 ;
        RECT 172.350 861.600 174.150 867.600 ;
        RECT 176.850 861.000 178.650 867.600 ;
        RECT 179.850 861.600 181.650 868.500 ;
        RECT 182.850 861.000 184.650 867.600 ;
        RECT 187.650 861.600 189.450 870.600 ;
        RECT 193.050 861.000 194.850 873.600 ;
        RECT 196.050 871.800 198.450 873.600 ;
        RECT 200.550 890.400 202.950 892.200 ;
        RECT 204.150 890.400 205.950 897.000 ;
        RECT 208.950 894.300 210.750 896.400 ;
        RECT 207.150 893.400 210.750 894.300 ;
        RECT 213.450 893.400 215.250 897.000 ;
        RECT 216.750 893.400 218.550 896.400 ;
        RECT 219.750 893.400 221.550 897.000 ;
        RECT 224.250 893.400 226.050 896.400 ;
        RECT 206.850 892.800 210.750 893.400 ;
        RECT 206.850 891.300 208.950 892.800 ;
        RECT 216.750 892.500 217.800 893.400 ;
        RECT 200.550 875.700 201.450 890.400 ;
        RECT 209.850 889.800 211.650 891.600 ;
        RECT 212.850 891.450 217.800 892.500 ;
        RECT 212.850 890.700 214.650 891.450 ;
        RECT 224.250 891.300 226.650 893.400 ;
        RECT 229.350 890.400 231.150 897.000 ;
        RECT 232.650 890.400 234.450 896.400 ;
        RECT 209.850 888.000 210.900 889.800 ;
        RECT 220.050 888.000 221.850 888.600 ;
        RECT 209.850 886.800 221.850 888.000 ;
        RECT 202.950 885.600 210.900 886.800 ;
        RECT 202.950 883.050 204.750 885.600 ;
        RECT 209.100 885.000 210.900 885.600 ;
        RECT 206.100 883.800 207.900 884.400 ;
        RECT 202.950 880.950 205.050 883.050 ;
        RECT 206.100 882.600 214.200 883.800 ;
        RECT 212.100 880.950 214.200 882.600 ;
        RECT 210.450 875.700 212.250 876.000 ;
        RECT 200.550 875.100 212.250 875.700 ;
        RECT 200.550 874.500 218.850 875.100 ;
        RECT 200.550 873.600 201.450 874.500 ;
        RECT 210.450 874.200 218.850 874.500 ;
        RECT 200.550 871.800 202.950 873.600 ;
        RECT 196.050 861.600 197.850 871.800 ;
        RECT 201.150 861.600 202.950 871.800 ;
        RECT 204.150 861.000 205.950 873.600 ;
        RECT 215.250 872.700 217.050 873.300 ;
        RECT 209.250 871.500 217.050 872.700 ;
        RECT 217.950 872.100 218.850 874.200 ;
        RECT 220.950 874.200 221.850 886.800 ;
        RECT 233.250 883.050 234.450 890.400 ;
        RECT 248.100 893.400 249.900 896.400 ;
        RECT 248.100 889.500 249.300 893.400 ;
        RECT 251.100 890.400 252.900 897.000 ;
        RECT 254.100 890.400 255.900 896.400 ;
        RECT 269.100 893.400 270.900 896.400 ;
        RECT 272.100 893.400 273.900 897.000 ;
        RECT 287.100 893.400 288.900 897.000 ;
        RECT 290.100 893.400 291.900 896.400 ;
        RECT 248.100 888.600 253.800 889.500 ;
        RECT 252.000 887.700 253.800 888.600 ;
        RECT 228.150 881.250 234.450 883.050 ;
        RECT 229.950 880.950 234.450 881.250 ;
        RECT 224.550 878.100 226.650 878.400 ;
        RECT 230.550 878.100 232.350 878.250 ;
        RECT 224.550 876.900 232.350 878.100 ;
        RECT 224.550 876.300 226.650 876.900 ;
        RECT 230.550 876.450 232.350 876.900 ;
        RECT 220.950 873.300 225.750 874.200 ;
        RECT 233.250 873.600 234.450 880.950 ;
        RECT 248.400 880.950 250.500 883.050 ;
        RECT 248.400 879.150 250.200 880.950 ;
        RECT 252.000 876.300 252.900 887.700 ;
        RECT 254.700 883.050 255.900 890.400 ;
        RECT 269.700 883.050 270.900 893.400 ;
        RECT 290.100 883.050 291.300 893.400 ;
        RECT 294.150 892.200 295.950 896.400 ;
        RECT 293.550 890.400 295.950 892.200 ;
        RECT 297.150 890.400 298.950 897.000 ;
        RECT 301.950 894.300 303.750 896.400 ;
        RECT 300.150 893.400 303.750 894.300 ;
        RECT 306.450 893.400 308.250 897.000 ;
        RECT 309.750 893.400 311.550 896.400 ;
        RECT 312.750 893.400 314.550 897.000 ;
        RECT 317.250 893.400 319.050 896.400 ;
        RECT 299.850 892.800 303.750 893.400 ;
        RECT 299.850 891.300 301.950 892.800 ;
        RECT 309.750 892.500 310.800 893.400 ;
        RECT 253.800 880.950 255.900 883.050 ;
        RECT 268.950 880.950 271.050 883.050 ;
        RECT 271.950 880.950 274.050 883.050 ;
        RECT 286.950 880.950 289.050 883.050 ;
        RECT 289.950 880.950 292.050 883.050 ;
        RECT 252.000 875.400 253.800 876.300 ;
        RECT 224.550 872.400 225.750 873.300 ;
        RECT 221.850 872.100 223.650 872.400 ;
        RECT 209.250 870.600 211.350 871.500 ;
        RECT 217.950 871.200 223.650 872.100 ;
        RECT 221.850 870.600 223.650 871.200 ;
        RECT 224.550 870.600 227.550 872.400 ;
        RECT 209.550 861.600 211.350 870.600 ;
        RECT 213.450 869.550 215.250 870.300 ;
        RECT 218.250 869.550 220.050 870.300 ;
        RECT 213.450 868.500 220.050 869.550 ;
        RECT 214.350 861.000 216.150 867.600 ;
        RECT 217.350 861.600 219.150 868.500 ;
        RECT 224.550 867.600 226.650 869.700 ;
        RECT 220.350 861.000 222.150 867.600 ;
        RECT 224.850 861.600 226.650 867.600 ;
        RECT 229.650 861.000 231.450 873.600 ;
        RECT 232.650 861.600 234.450 873.600 ;
        RECT 248.100 874.500 253.800 875.400 ;
        RECT 248.100 867.600 249.300 874.500 ;
        RECT 254.700 873.600 255.900 880.950 ;
        RECT 248.100 861.600 249.900 867.600 ;
        RECT 251.100 861.000 252.900 871.800 ;
        RECT 254.100 861.600 255.900 873.600 ;
        RECT 269.700 867.600 270.900 880.950 ;
        RECT 272.100 879.150 273.900 880.950 ;
        RECT 287.100 879.150 288.900 880.950 ;
        RECT 290.100 867.600 291.300 880.950 ;
        RECT 293.550 875.700 294.450 890.400 ;
        RECT 302.850 889.800 304.650 891.600 ;
        RECT 305.850 891.450 310.800 892.500 ;
        RECT 305.850 890.700 307.650 891.450 ;
        RECT 317.250 891.300 319.650 893.400 ;
        RECT 322.350 890.400 324.150 897.000 ;
        RECT 325.650 890.400 327.450 896.400 ;
        RECT 302.850 888.000 303.900 889.800 ;
        RECT 313.050 888.000 314.850 888.600 ;
        RECT 302.850 886.800 314.850 888.000 ;
        RECT 295.950 885.600 303.900 886.800 ;
        RECT 295.950 883.050 297.750 885.600 ;
        RECT 302.100 885.000 303.900 885.600 ;
        RECT 299.100 883.800 300.900 884.400 ;
        RECT 295.950 880.950 298.050 883.050 ;
        RECT 299.100 882.600 307.200 883.800 ;
        RECT 305.100 880.950 307.200 882.600 ;
        RECT 303.450 875.700 305.250 876.000 ;
        RECT 293.550 875.100 305.250 875.700 ;
        RECT 293.550 874.500 311.850 875.100 ;
        RECT 293.550 873.600 294.450 874.500 ;
        RECT 303.450 874.200 311.850 874.500 ;
        RECT 293.550 871.800 295.950 873.600 ;
        RECT 269.100 861.600 270.900 867.600 ;
        RECT 272.100 861.000 273.900 867.600 ;
        RECT 287.100 861.000 288.900 867.600 ;
        RECT 290.100 861.600 291.900 867.600 ;
        RECT 294.150 861.600 295.950 871.800 ;
        RECT 297.150 861.000 298.950 873.600 ;
        RECT 308.250 872.700 310.050 873.300 ;
        RECT 302.250 871.500 310.050 872.700 ;
        RECT 310.950 872.100 311.850 874.200 ;
        RECT 313.950 874.200 314.850 886.800 ;
        RECT 326.250 883.050 327.450 890.400 ;
        RECT 344.100 893.400 345.900 896.400 ;
        RECT 344.100 889.500 345.300 893.400 ;
        RECT 347.100 890.400 348.900 897.000 ;
        RECT 350.100 890.400 351.900 896.400 ;
        RECT 344.100 888.600 349.800 889.500 ;
        RECT 348.000 887.700 349.800 888.600 ;
        RECT 321.150 881.250 327.450 883.050 ;
        RECT 322.950 880.950 327.450 881.250 ;
        RECT 317.550 878.100 319.650 878.400 ;
        RECT 323.550 878.100 325.350 878.250 ;
        RECT 317.550 876.900 325.350 878.100 ;
        RECT 317.550 876.300 319.650 876.900 ;
        RECT 323.550 876.450 325.350 876.900 ;
        RECT 313.950 873.300 318.750 874.200 ;
        RECT 326.250 873.600 327.450 880.950 ;
        RECT 344.400 880.950 346.500 883.050 ;
        RECT 344.400 879.150 346.200 880.950 ;
        RECT 348.000 876.300 348.900 887.700 ;
        RECT 350.700 883.050 351.900 890.400 ;
        RECT 370.500 888.000 372.300 896.400 ;
        RECT 369.000 886.800 372.300 888.000 ;
        RECT 377.100 887.400 378.900 897.000 ;
        RECT 392.700 893.400 394.500 897.000 ;
        RECT 395.700 891.600 397.500 896.400 ;
        RECT 392.400 890.400 397.500 891.600 ;
        RECT 400.200 890.400 402.000 897.000 ;
        RECT 416.100 890.400 417.900 896.400 ;
        RECT 419.100 890.400 420.900 897.000 ;
        RECT 422.100 893.400 423.900 896.400 ;
        RECT 369.000 883.050 369.900 886.800 ;
        RECT 371.100 883.050 372.900 884.850 ;
        RECT 377.100 883.050 378.900 884.850 ;
        RECT 392.400 883.050 393.300 890.400 ;
        RECT 394.950 883.050 396.750 884.850 ;
        RECT 401.100 883.050 402.900 884.850 ;
        RECT 416.100 883.050 417.300 890.400 ;
        RECT 422.700 889.500 423.900 893.400 ;
        RECT 418.200 888.600 423.900 889.500 ;
        RECT 425.550 890.400 427.350 896.400 ;
        RECT 428.850 890.400 430.650 897.000 ;
        RECT 433.950 893.400 435.750 896.400 ;
        RECT 438.450 893.400 440.250 897.000 ;
        RECT 441.450 893.400 443.250 896.400 ;
        RECT 444.750 893.400 446.550 897.000 ;
        RECT 449.250 894.300 451.050 896.400 ;
        RECT 449.250 893.400 452.850 894.300 ;
        RECT 433.350 891.300 435.750 893.400 ;
        RECT 442.200 892.500 443.250 893.400 ;
        RECT 449.250 892.800 453.150 893.400 ;
        RECT 442.200 891.450 447.150 892.500 ;
        RECT 445.350 890.700 447.150 891.450 ;
        RECT 418.200 887.700 420.000 888.600 ;
        RECT 349.800 880.950 351.900 883.050 ;
        RECT 367.950 880.950 370.050 883.050 ;
        RECT 370.950 880.950 373.050 883.050 ;
        RECT 373.950 880.950 376.050 883.050 ;
        RECT 376.950 880.950 379.050 883.050 ;
        RECT 391.950 880.950 394.050 883.050 ;
        RECT 394.950 880.950 397.050 883.050 ;
        RECT 397.950 880.950 400.050 883.050 ;
        RECT 400.950 880.950 403.050 883.050 ;
        RECT 416.100 880.950 418.200 883.050 ;
        RECT 348.000 875.400 349.800 876.300 ;
        RECT 317.550 872.400 318.750 873.300 ;
        RECT 314.850 872.100 316.650 872.400 ;
        RECT 302.250 870.600 304.350 871.500 ;
        RECT 310.950 871.200 316.650 872.100 ;
        RECT 314.850 870.600 316.650 871.200 ;
        RECT 317.550 870.600 320.550 872.400 ;
        RECT 302.550 861.600 304.350 870.600 ;
        RECT 306.450 869.550 308.250 870.300 ;
        RECT 311.250 869.550 313.050 870.300 ;
        RECT 306.450 868.500 313.050 869.550 ;
        RECT 307.350 861.000 309.150 867.600 ;
        RECT 310.350 861.600 312.150 868.500 ;
        RECT 317.550 867.600 319.650 869.700 ;
        RECT 313.350 861.000 315.150 867.600 ;
        RECT 317.850 861.600 319.650 867.600 ;
        RECT 322.650 861.000 324.450 873.600 ;
        RECT 325.650 861.600 327.450 873.600 ;
        RECT 344.100 874.500 349.800 875.400 ;
        RECT 344.100 867.600 345.300 874.500 ;
        RECT 350.700 873.600 351.900 880.950 ;
        RECT 344.100 861.600 345.900 867.600 ;
        RECT 347.100 861.000 348.900 871.800 ;
        RECT 350.100 861.600 351.900 873.600 ;
        RECT 369.000 868.800 369.900 880.950 ;
        RECT 374.100 879.150 375.900 880.950 ;
        RECT 392.400 873.600 393.300 880.950 ;
        RECT 397.950 879.150 399.750 880.950 ;
        RECT 416.100 873.600 417.300 880.950 ;
        RECT 419.100 876.300 420.000 887.700 ;
        RECT 425.550 883.050 426.750 890.400 ;
        RECT 448.350 889.800 450.150 891.600 ;
        RECT 451.050 891.300 453.150 892.800 ;
        RECT 454.050 890.400 455.850 897.000 ;
        RECT 457.050 892.200 458.850 896.400 ;
        RECT 457.050 890.400 459.450 892.200 ;
        RECT 438.150 888.000 439.950 888.600 ;
        RECT 449.100 888.000 450.150 889.800 ;
        RECT 438.150 886.800 450.150 888.000 ;
        RECT 421.500 880.950 423.600 883.050 ;
        RECT 421.800 879.150 423.600 880.950 ;
        RECT 425.550 881.250 431.850 883.050 ;
        RECT 425.550 880.950 430.050 881.250 ;
        RECT 418.200 875.400 420.000 876.300 ;
        RECT 418.200 874.500 423.900 875.400 ;
        RECT 369.000 867.900 375.600 868.800 ;
        RECT 369.000 867.600 369.900 867.900 ;
        RECT 368.100 861.600 369.900 867.600 ;
        RECT 374.100 867.600 375.600 867.900 ;
        RECT 371.100 861.000 372.900 867.000 ;
        RECT 374.100 861.600 375.900 867.600 ;
        RECT 377.100 861.000 378.900 867.600 ;
        RECT 392.100 861.600 393.900 873.600 ;
        RECT 395.100 872.700 402.900 873.600 ;
        RECT 395.100 861.600 396.900 872.700 ;
        RECT 398.100 861.000 399.900 871.800 ;
        RECT 401.100 861.600 402.900 872.700 ;
        RECT 416.100 861.600 417.900 873.600 ;
        RECT 419.100 861.000 420.900 871.800 ;
        RECT 422.700 867.600 423.900 874.500 ;
        RECT 422.100 861.600 423.900 867.600 ;
        RECT 425.550 873.600 426.750 880.950 ;
        RECT 427.650 878.100 429.450 878.250 ;
        RECT 433.350 878.100 435.450 878.400 ;
        RECT 427.650 876.900 435.450 878.100 ;
        RECT 427.650 876.450 429.450 876.900 ;
        RECT 433.350 876.300 435.450 876.900 ;
        RECT 438.150 874.200 439.050 886.800 ;
        RECT 449.100 885.600 457.050 886.800 ;
        RECT 449.100 885.000 450.900 885.600 ;
        RECT 452.100 883.800 453.900 884.400 ;
        RECT 445.800 882.600 453.900 883.800 ;
        RECT 455.250 883.050 457.050 885.600 ;
        RECT 445.800 880.950 447.900 882.600 ;
        RECT 454.950 880.950 457.050 883.050 ;
        RECT 447.750 875.700 449.550 876.000 ;
        RECT 458.550 875.700 459.450 890.400 ;
        RECT 447.750 875.100 459.450 875.700 ;
        RECT 425.550 861.600 427.350 873.600 ;
        RECT 428.550 861.000 430.350 873.600 ;
        RECT 434.250 873.300 439.050 874.200 ;
        RECT 441.150 874.500 459.450 875.100 ;
        RECT 441.150 874.200 449.550 874.500 ;
        RECT 434.250 872.400 435.450 873.300 ;
        RECT 432.450 870.600 435.450 872.400 ;
        RECT 436.350 872.100 438.150 872.400 ;
        RECT 441.150 872.100 442.050 874.200 ;
        RECT 458.550 873.600 459.450 874.500 ;
        RECT 436.350 871.200 442.050 872.100 ;
        RECT 442.950 872.700 444.750 873.300 ;
        RECT 442.950 871.500 450.750 872.700 ;
        RECT 436.350 870.600 438.150 871.200 ;
        RECT 448.650 870.600 450.750 871.500 ;
        RECT 433.350 867.600 435.450 869.700 ;
        RECT 439.950 869.550 441.750 870.300 ;
        RECT 444.750 869.550 446.550 870.300 ;
        RECT 439.950 868.500 446.550 869.550 ;
        RECT 433.350 861.600 435.150 867.600 ;
        RECT 437.850 861.000 439.650 867.600 ;
        RECT 440.850 861.600 442.650 868.500 ;
        RECT 443.850 861.000 445.650 867.600 ;
        RECT 448.650 861.600 450.450 870.600 ;
        RECT 454.050 861.000 455.850 873.600 ;
        RECT 457.050 871.800 459.450 873.600 ;
        RECT 473.100 890.400 474.900 896.400 ;
        RECT 476.100 890.400 477.900 897.000 ;
        RECT 479.100 893.400 480.900 896.400 ;
        RECT 473.100 883.050 474.300 890.400 ;
        RECT 479.700 889.500 480.900 893.400 ;
        RECT 475.200 888.600 480.900 889.500 ;
        RECT 497.100 890.400 498.900 896.400 ;
        RECT 500.100 890.400 501.900 897.000 ;
        RECT 503.100 893.400 504.900 896.400 ;
        RECT 475.200 887.700 477.000 888.600 ;
        RECT 473.100 880.950 475.200 883.050 ;
        RECT 473.100 873.600 474.300 880.950 ;
        RECT 476.100 876.300 477.000 887.700 ;
        RECT 497.100 883.050 498.300 890.400 ;
        RECT 503.700 889.500 504.900 893.400 ;
        RECT 499.200 888.600 504.900 889.500 ;
        RECT 506.550 890.400 508.350 896.400 ;
        RECT 509.850 890.400 511.650 897.000 ;
        RECT 514.950 893.400 516.750 896.400 ;
        RECT 519.450 893.400 521.250 897.000 ;
        RECT 522.450 893.400 524.250 896.400 ;
        RECT 525.750 893.400 527.550 897.000 ;
        RECT 530.250 894.300 532.050 896.400 ;
        RECT 530.250 893.400 533.850 894.300 ;
        RECT 514.350 891.300 516.750 893.400 ;
        RECT 523.200 892.500 524.250 893.400 ;
        RECT 530.250 892.800 534.150 893.400 ;
        RECT 523.200 891.450 528.150 892.500 ;
        RECT 526.350 890.700 528.150 891.450 ;
        RECT 499.200 887.700 501.000 888.600 ;
        RECT 478.500 880.950 480.600 883.050 ;
        RECT 478.800 879.150 480.600 880.950 ;
        RECT 497.100 880.950 499.200 883.050 ;
        RECT 475.200 875.400 477.000 876.300 ;
        RECT 475.200 874.500 480.900 875.400 ;
        RECT 457.050 861.600 458.850 871.800 ;
        RECT 473.100 861.600 474.900 873.600 ;
        RECT 476.100 861.000 477.900 871.800 ;
        RECT 479.700 867.600 480.900 874.500 ;
        RECT 479.100 861.600 480.900 867.600 ;
        RECT 497.100 873.600 498.300 880.950 ;
        RECT 500.100 876.300 501.000 887.700 ;
        RECT 506.550 883.050 507.750 890.400 ;
        RECT 529.350 889.800 531.150 891.600 ;
        RECT 532.050 891.300 534.150 892.800 ;
        RECT 535.050 890.400 536.850 897.000 ;
        RECT 538.050 892.200 539.850 896.400 ;
        RECT 543.150 892.200 544.950 896.400 ;
        RECT 538.050 890.400 540.450 892.200 ;
        RECT 519.150 888.000 520.950 888.600 ;
        RECT 530.100 888.000 531.150 889.800 ;
        RECT 519.150 886.800 531.150 888.000 ;
        RECT 502.500 880.950 504.600 883.050 ;
        RECT 502.800 879.150 504.600 880.950 ;
        RECT 506.550 881.250 512.850 883.050 ;
        RECT 506.550 880.950 511.050 881.250 ;
        RECT 499.200 875.400 501.000 876.300 ;
        RECT 499.200 874.500 504.900 875.400 ;
        RECT 497.100 861.600 498.900 873.600 ;
        RECT 500.100 861.000 501.900 871.800 ;
        RECT 503.700 867.600 504.900 874.500 ;
        RECT 503.100 861.600 504.900 867.600 ;
        RECT 506.550 873.600 507.750 880.950 ;
        RECT 508.650 878.100 510.450 878.250 ;
        RECT 514.350 878.100 516.450 878.400 ;
        RECT 508.650 876.900 516.450 878.100 ;
        RECT 508.650 876.450 510.450 876.900 ;
        RECT 514.350 876.300 516.450 876.900 ;
        RECT 519.150 874.200 520.050 886.800 ;
        RECT 530.100 885.600 538.050 886.800 ;
        RECT 530.100 885.000 531.900 885.600 ;
        RECT 533.100 883.800 534.900 884.400 ;
        RECT 526.800 882.600 534.900 883.800 ;
        RECT 536.250 883.050 538.050 885.600 ;
        RECT 526.800 880.950 528.900 882.600 ;
        RECT 535.950 880.950 538.050 883.050 ;
        RECT 528.750 875.700 530.550 876.000 ;
        RECT 539.550 875.700 540.450 890.400 ;
        RECT 528.750 875.100 540.450 875.700 ;
        RECT 506.550 861.600 508.350 873.600 ;
        RECT 509.550 861.000 511.350 873.600 ;
        RECT 515.250 873.300 520.050 874.200 ;
        RECT 522.150 874.500 540.450 875.100 ;
        RECT 522.150 874.200 530.550 874.500 ;
        RECT 515.250 872.400 516.450 873.300 ;
        RECT 513.450 870.600 516.450 872.400 ;
        RECT 517.350 872.100 519.150 872.400 ;
        RECT 522.150 872.100 523.050 874.200 ;
        RECT 539.550 873.600 540.450 874.500 ;
        RECT 517.350 871.200 523.050 872.100 ;
        RECT 523.950 872.700 525.750 873.300 ;
        RECT 523.950 871.500 531.750 872.700 ;
        RECT 517.350 870.600 519.150 871.200 ;
        RECT 529.650 870.600 531.750 871.500 ;
        RECT 514.350 867.600 516.450 869.700 ;
        RECT 520.950 869.550 522.750 870.300 ;
        RECT 525.750 869.550 527.550 870.300 ;
        RECT 520.950 868.500 527.550 869.550 ;
        RECT 514.350 861.600 516.150 867.600 ;
        RECT 518.850 861.000 520.650 867.600 ;
        RECT 521.850 861.600 523.650 868.500 ;
        RECT 524.850 861.000 526.650 867.600 ;
        RECT 529.650 861.600 531.450 870.600 ;
        RECT 535.050 861.000 536.850 873.600 ;
        RECT 538.050 871.800 540.450 873.600 ;
        RECT 542.550 890.400 544.950 892.200 ;
        RECT 546.150 890.400 547.950 897.000 ;
        RECT 550.950 894.300 552.750 896.400 ;
        RECT 549.150 893.400 552.750 894.300 ;
        RECT 555.450 893.400 557.250 897.000 ;
        RECT 558.750 893.400 560.550 896.400 ;
        RECT 561.750 893.400 563.550 897.000 ;
        RECT 566.250 893.400 568.050 896.400 ;
        RECT 548.850 892.800 552.750 893.400 ;
        RECT 548.850 891.300 550.950 892.800 ;
        RECT 558.750 892.500 559.800 893.400 ;
        RECT 542.550 875.700 543.450 890.400 ;
        RECT 551.850 889.800 553.650 891.600 ;
        RECT 554.850 891.450 559.800 892.500 ;
        RECT 554.850 890.700 556.650 891.450 ;
        RECT 566.250 891.300 568.650 893.400 ;
        RECT 571.350 890.400 573.150 897.000 ;
        RECT 574.650 890.400 576.450 896.400 ;
        RECT 551.850 888.000 552.900 889.800 ;
        RECT 562.050 888.000 563.850 888.600 ;
        RECT 551.850 886.800 563.850 888.000 ;
        RECT 544.950 885.600 552.900 886.800 ;
        RECT 544.950 883.050 546.750 885.600 ;
        RECT 551.100 885.000 552.900 885.600 ;
        RECT 548.100 883.800 549.900 884.400 ;
        RECT 544.950 880.950 547.050 883.050 ;
        RECT 548.100 882.600 556.200 883.800 ;
        RECT 554.100 880.950 556.200 882.600 ;
        RECT 552.450 875.700 554.250 876.000 ;
        RECT 542.550 875.100 554.250 875.700 ;
        RECT 542.550 874.500 560.850 875.100 ;
        RECT 542.550 873.600 543.450 874.500 ;
        RECT 552.450 874.200 560.850 874.500 ;
        RECT 542.550 871.800 544.950 873.600 ;
        RECT 538.050 861.600 539.850 871.800 ;
        RECT 543.150 861.600 544.950 871.800 ;
        RECT 546.150 861.000 547.950 873.600 ;
        RECT 557.250 872.700 559.050 873.300 ;
        RECT 551.250 871.500 559.050 872.700 ;
        RECT 559.950 872.100 560.850 874.200 ;
        RECT 562.950 874.200 563.850 886.800 ;
        RECT 575.250 883.050 576.450 890.400 ;
        RECT 593.100 893.400 594.900 896.400 ;
        RECT 593.100 889.500 594.300 893.400 ;
        RECT 596.100 890.400 597.900 897.000 ;
        RECT 599.100 890.400 600.900 896.400 ;
        RECT 593.100 888.600 598.800 889.500 ;
        RECT 597.000 887.700 598.800 888.600 ;
        RECT 570.150 881.250 576.450 883.050 ;
        RECT 571.950 880.950 576.450 881.250 ;
        RECT 566.550 878.100 568.650 878.400 ;
        RECT 572.550 878.100 574.350 878.250 ;
        RECT 566.550 876.900 574.350 878.100 ;
        RECT 566.550 876.300 568.650 876.900 ;
        RECT 572.550 876.450 574.350 876.900 ;
        RECT 562.950 873.300 567.750 874.200 ;
        RECT 575.250 873.600 576.450 880.950 ;
        RECT 593.400 880.950 595.500 883.050 ;
        RECT 593.400 879.150 595.200 880.950 ;
        RECT 597.000 876.300 597.900 887.700 ;
        RECT 599.700 883.050 600.900 890.400 ;
        RECT 598.800 880.950 600.900 883.050 ;
        RECT 597.000 875.400 598.800 876.300 ;
        RECT 566.550 872.400 567.750 873.300 ;
        RECT 563.850 872.100 565.650 872.400 ;
        RECT 551.250 870.600 553.350 871.500 ;
        RECT 559.950 871.200 565.650 872.100 ;
        RECT 563.850 870.600 565.650 871.200 ;
        RECT 566.550 870.600 569.550 872.400 ;
        RECT 551.550 861.600 553.350 870.600 ;
        RECT 555.450 869.550 557.250 870.300 ;
        RECT 560.250 869.550 562.050 870.300 ;
        RECT 555.450 868.500 562.050 869.550 ;
        RECT 556.350 861.000 558.150 867.600 ;
        RECT 559.350 861.600 561.150 868.500 ;
        RECT 566.550 867.600 568.650 869.700 ;
        RECT 562.350 861.000 564.150 867.600 ;
        RECT 566.850 861.600 568.650 867.600 ;
        RECT 571.650 861.000 573.450 873.600 ;
        RECT 574.650 861.600 576.450 873.600 ;
        RECT 593.100 874.500 598.800 875.400 ;
        RECT 593.100 867.600 594.300 874.500 ;
        RECT 599.700 873.600 600.900 880.950 ;
        RECT 593.100 861.600 594.900 867.600 ;
        RECT 596.100 861.000 597.900 871.800 ;
        RECT 599.100 861.600 600.900 873.600 ;
        RECT 614.100 890.400 615.900 896.400 ;
        RECT 617.100 890.400 618.900 897.000 ;
        RECT 620.100 893.400 621.900 896.400 ;
        RECT 614.100 883.050 615.300 890.400 ;
        RECT 620.700 889.500 621.900 893.400 ;
        RECT 616.200 888.600 621.900 889.500 ;
        RECT 638.100 893.400 639.900 896.400 ;
        RECT 638.100 889.500 639.300 893.400 ;
        RECT 641.100 890.400 642.900 897.000 ;
        RECT 644.100 890.400 645.900 896.400 ;
        RECT 638.100 888.600 643.800 889.500 ;
        RECT 616.200 887.700 618.000 888.600 ;
        RECT 614.100 880.950 616.200 883.050 ;
        RECT 614.100 873.600 615.300 880.950 ;
        RECT 617.100 876.300 618.000 887.700 ;
        RECT 642.000 887.700 643.800 888.600 ;
        RECT 619.500 880.950 621.600 883.050 ;
        RECT 619.800 879.150 621.600 880.950 ;
        RECT 638.400 880.950 640.500 883.050 ;
        RECT 638.400 879.150 640.200 880.950 ;
        RECT 616.200 875.400 618.000 876.300 ;
        RECT 642.000 876.300 642.900 887.700 ;
        RECT 644.700 883.050 645.900 890.400 ;
        RECT 662.100 887.400 663.900 897.000 ;
        RECT 668.700 888.000 670.500 896.400 ;
        RECT 689.100 893.400 690.900 896.400 ;
        RECT 692.100 893.400 693.900 897.000 ;
        RECT 668.700 886.800 672.000 888.000 ;
        RECT 662.100 883.050 663.900 884.850 ;
        RECT 668.100 883.050 669.900 884.850 ;
        RECT 671.100 883.050 672.000 886.800 ;
        RECT 689.700 883.050 690.900 893.400 ;
        RECT 707.400 890.400 709.200 897.000 ;
        RECT 712.500 889.200 714.300 896.400 ;
        RECT 710.100 888.300 714.300 889.200 ;
        RECT 728.700 889.200 730.500 896.400 ;
        RECT 733.800 890.400 735.600 897.000 ;
        RECT 749.700 889.200 751.500 896.400 ;
        RECT 754.800 890.400 756.600 897.000 ;
        RECT 770.100 893.400 771.900 896.400 ;
        RECT 770.100 889.500 771.300 893.400 ;
        RECT 773.100 890.400 774.900 897.000 ;
        RECT 776.100 890.400 777.900 896.400 ;
        RECT 728.700 888.300 732.900 889.200 ;
        RECT 749.700 888.300 753.900 889.200 ;
        RECT 770.100 888.600 775.800 889.500 ;
        RECT 707.250 883.050 709.050 884.850 ;
        RECT 710.100 883.050 711.300 888.300 ;
        RECT 713.100 883.050 714.900 884.850 ;
        RECT 728.100 883.050 729.900 884.850 ;
        RECT 731.700 883.050 732.900 888.300 ;
        RECT 733.950 883.050 735.750 884.850 ;
        RECT 749.100 883.050 750.900 884.850 ;
        RECT 752.700 883.050 753.900 888.300 ;
        RECT 774.000 887.700 775.800 888.600 ;
        RECT 754.950 883.050 756.750 884.850 ;
        RECT 643.800 880.950 645.900 883.050 ;
        RECT 661.950 880.950 664.050 883.050 ;
        RECT 664.950 880.950 667.050 883.050 ;
        RECT 667.950 880.950 670.050 883.050 ;
        RECT 670.950 880.950 673.050 883.050 ;
        RECT 688.950 880.950 691.050 883.050 ;
        RECT 691.950 880.950 694.050 883.050 ;
        RECT 706.950 880.950 709.050 883.050 ;
        RECT 709.950 880.950 712.050 883.050 ;
        RECT 712.950 880.950 715.050 883.050 ;
        RECT 727.950 880.950 730.050 883.050 ;
        RECT 730.950 880.950 733.050 883.050 ;
        RECT 733.950 880.950 736.050 883.050 ;
        RECT 748.950 880.950 751.050 883.050 ;
        RECT 751.950 880.950 754.050 883.050 ;
        RECT 754.950 880.950 757.050 883.050 ;
        RECT 770.400 880.950 772.500 883.050 ;
        RECT 642.000 875.400 643.800 876.300 ;
        RECT 616.200 874.500 621.900 875.400 ;
        RECT 614.100 861.600 615.900 873.600 ;
        RECT 617.100 861.000 618.900 871.800 ;
        RECT 620.700 867.600 621.900 874.500 ;
        RECT 620.100 861.600 621.900 867.600 ;
        RECT 638.100 874.500 643.800 875.400 ;
        RECT 638.100 867.600 639.300 874.500 ;
        RECT 644.700 873.600 645.900 880.950 ;
        RECT 665.100 879.150 666.900 880.950 ;
        RECT 638.100 861.600 639.900 867.600 ;
        RECT 641.100 861.000 642.900 871.800 ;
        RECT 644.100 861.600 645.900 873.600 ;
        RECT 671.100 868.800 672.000 880.950 ;
        RECT 665.400 867.900 672.000 868.800 ;
        RECT 665.400 867.600 666.900 867.900 ;
        RECT 662.100 861.000 663.900 867.600 ;
        RECT 665.100 861.600 666.900 867.600 ;
        RECT 671.100 867.600 672.000 867.900 ;
        RECT 689.700 867.600 690.900 880.950 ;
        RECT 692.100 879.150 693.900 880.950 ;
        RECT 710.100 867.600 711.300 880.950 ;
        RECT 731.700 867.600 732.900 880.950 ;
        RECT 752.700 867.600 753.900 880.950 ;
        RECT 770.400 879.150 772.200 880.950 ;
        RECT 774.000 876.300 774.900 887.700 ;
        RECT 776.700 883.050 777.900 890.400 ;
        RECT 791.700 889.200 793.500 896.400 ;
        RECT 796.800 890.400 798.600 897.000 ;
        RECT 815.700 889.200 817.500 896.400 ;
        RECT 820.800 890.400 822.600 897.000 ;
        RECT 836.100 893.400 837.900 897.000 ;
        RECT 839.100 893.400 840.900 896.400 ;
        RECT 842.100 893.400 843.900 897.000 ;
        RECT 860.100 893.400 861.900 896.400 ;
        RECT 863.100 893.400 864.900 897.000 ;
        RECT 878.100 893.400 879.900 897.000 ;
        RECT 881.100 893.400 882.900 896.400 ;
        RECT 791.700 888.300 795.900 889.200 ;
        RECT 815.700 888.300 819.900 889.200 ;
        RECT 791.100 883.050 792.900 884.850 ;
        RECT 794.700 883.050 795.900 888.300 ;
        RECT 796.950 883.050 798.750 884.850 ;
        RECT 815.100 883.050 816.900 884.850 ;
        RECT 818.700 883.050 819.900 888.300 ;
        RECT 820.950 883.050 822.750 884.850 ;
        RECT 839.700 883.050 840.600 893.400 ;
        RECT 860.700 883.050 861.900 893.400 ;
        RECT 871.950 888.450 874.050 889.050 ;
        RECT 877.950 888.450 880.050 889.050 ;
        RECT 871.950 887.550 880.050 888.450 ;
        RECT 871.950 886.950 874.050 887.550 ;
        RECT 877.950 886.950 880.050 887.550 ;
        RECT 881.100 883.050 882.300 893.400 ;
        RECT 775.800 880.950 777.900 883.050 ;
        RECT 790.950 880.950 793.050 883.050 ;
        RECT 793.950 880.950 796.050 883.050 ;
        RECT 796.950 880.950 799.050 883.050 ;
        RECT 814.950 880.950 817.050 883.050 ;
        RECT 817.950 880.950 820.050 883.050 ;
        RECT 820.950 880.950 823.050 883.050 ;
        RECT 835.950 880.950 838.050 883.050 ;
        RECT 838.950 880.950 841.050 883.050 ;
        RECT 841.950 880.950 844.050 883.050 ;
        RECT 859.950 880.950 862.050 883.050 ;
        RECT 862.950 880.950 865.050 883.050 ;
        RECT 877.950 880.950 880.050 883.050 ;
        RECT 880.950 880.950 883.050 883.050 ;
        RECT 774.000 875.400 775.800 876.300 ;
        RECT 770.100 874.500 775.800 875.400 ;
        RECT 770.100 867.600 771.300 874.500 ;
        RECT 776.700 873.600 777.900 880.950 ;
        RECT 668.100 861.000 669.900 867.000 ;
        RECT 671.100 861.600 672.900 867.600 ;
        RECT 689.100 861.600 690.900 867.600 ;
        RECT 692.100 861.000 693.900 867.600 ;
        RECT 707.100 861.000 708.900 867.600 ;
        RECT 710.100 861.600 711.900 867.600 ;
        RECT 713.100 861.000 714.900 867.600 ;
        RECT 728.100 861.000 729.900 867.600 ;
        RECT 731.100 861.600 732.900 867.600 ;
        RECT 734.100 861.000 735.900 867.600 ;
        RECT 749.100 861.000 750.900 867.600 ;
        RECT 752.100 861.600 753.900 867.600 ;
        RECT 755.100 861.000 756.900 867.600 ;
        RECT 770.100 861.600 771.900 867.600 ;
        RECT 773.100 861.000 774.900 871.800 ;
        RECT 776.100 861.600 777.900 873.600 ;
        RECT 794.700 867.600 795.900 880.950 ;
        RECT 818.700 867.600 819.900 880.950 ;
        RECT 836.100 879.150 837.900 880.950 ;
        RECT 839.700 873.600 840.600 880.950 ;
        RECT 841.950 879.150 843.750 880.950 ;
        RECT 837.000 872.400 840.600 873.600 ;
        RECT 791.100 861.000 792.900 867.600 ;
        RECT 794.100 861.600 795.900 867.600 ;
        RECT 797.100 861.000 798.900 867.600 ;
        RECT 815.100 861.000 816.900 867.600 ;
        RECT 818.100 861.600 819.900 867.600 ;
        RECT 821.100 861.000 822.900 867.600 ;
        RECT 837.000 861.600 838.800 872.400 ;
        RECT 842.100 861.000 843.900 873.600 ;
        RECT 860.700 867.600 861.900 880.950 ;
        RECT 863.100 879.150 864.900 880.950 ;
        RECT 878.100 879.150 879.900 880.950 ;
        RECT 881.100 867.600 882.300 880.950 ;
        RECT 860.100 861.600 861.900 867.600 ;
        RECT 863.100 861.000 864.900 867.600 ;
        RECT 878.100 861.000 879.900 867.600 ;
        RECT 881.100 861.600 882.900 867.600 ;
        RECT 14.100 851.400 15.900 858.000 ;
        RECT 17.100 851.400 18.900 857.400 ;
        RECT 35.100 851.400 36.900 858.000 ;
        RECT 38.100 851.400 39.900 857.400 ;
        RECT 41.100 851.400 42.900 858.000 ;
        RECT 56.100 851.400 57.900 858.000 ;
        RECT 59.100 851.400 60.900 857.400 ;
        RECT 62.100 851.400 63.900 858.000 ;
        RECT 77.100 851.400 78.900 858.000 ;
        RECT 80.100 851.400 81.900 857.400 ;
        RECT 83.100 852.000 84.900 858.000 ;
        RECT 14.100 838.050 15.900 839.850 ;
        RECT 17.100 838.050 18.300 851.400 ;
        RECT 38.100 838.050 39.300 851.400 ;
        RECT 59.700 838.050 60.900 851.400 ;
        RECT 80.400 851.100 81.900 851.400 ;
        RECT 86.100 851.400 87.900 857.400 ;
        RECT 86.100 851.100 87.000 851.400 ;
        RECT 80.400 850.200 87.000 851.100 ;
        RECT 80.100 838.050 81.900 839.850 ;
        RECT 86.100 838.050 87.000 850.200 ;
        RECT 101.100 846.300 102.900 857.400 ;
        RECT 104.100 847.200 105.900 858.000 ;
        RECT 107.100 846.300 108.900 857.400 ;
        RECT 101.100 845.400 108.900 846.300 ;
        RECT 110.100 845.400 111.900 857.400 ;
        RECT 128.100 846.300 129.900 857.400 ;
        RECT 131.100 847.200 132.900 858.000 ;
        RECT 134.100 846.300 135.900 857.400 ;
        RECT 128.100 845.400 135.900 846.300 ;
        RECT 137.100 845.400 138.900 857.400 ;
        RECT 152.100 851.400 153.900 857.400 ;
        RECT 155.100 851.400 156.900 858.000 ;
        RECT 104.250 838.050 106.050 839.850 ;
        RECT 110.700 838.050 111.600 845.400 ;
        RECT 131.250 838.050 133.050 839.850 ;
        RECT 137.700 838.050 138.600 845.400 ;
        RECT 152.700 838.050 153.900 851.400 ;
        RECT 158.550 845.400 160.350 857.400 ;
        RECT 161.550 845.400 163.350 858.000 ;
        RECT 166.350 851.400 168.150 857.400 ;
        RECT 170.850 851.400 172.650 858.000 ;
        RECT 166.350 849.300 168.450 851.400 ;
        RECT 173.850 850.500 175.650 857.400 ;
        RECT 176.850 851.400 178.650 858.000 ;
        RECT 172.950 849.450 179.550 850.500 ;
        RECT 172.950 848.700 174.750 849.450 ;
        RECT 177.750 848.700 179.550 849.450 ;
        RECT 181.650 848.400 183.450 857.400 ;
        RECT 165.450 846.600 168.450 848.400 ;
        RECT 169.350 847.800 171.150 848.400 ;
        RECT 169.350 846.900 175.050 847.800 ;
        RECT 181.650 847.500 183.750 848.400 ;
        RECT 169.350 846.600 171.150 846.900 ;
        RECT 167.250 845.700 168.450 846.600 ;
        RECT 155.100 838.050 156.900 839.850 ;
        RECT 158.550 838.050 159.750 845.400 ;
        RECT 167.250 844.800 172.050 845.700 ;
        RECT 160.650 842.100 162.450 842.550 ;
        RECT 166.350 842.100 168.450 842.700 ;
        RECT 160.650 840.900 168.450 842.100 ;
        RECT 160.650 840.750 162.450 840.900 ;
        RECT 166.350 840.600 168.450 840.900 ;
        RECT 13.950 835.950 16.050 838.050 ;
        RECT 16.950 835.950 19.050 838.050 ;
        RECT 34.950 835.950 37.050 838.050 ;
        RECT 37.950 835.950 40.050 838.050 ;
        RECT 40.950 835.950 43.050 838.050 ;
        RECT 55.950 835.950 58.050 838.050 ;
        RECT 58.950 835.950 61.050 838.050 ;
        RECT 61.950 835.950 64.050 838.050 ;
        RECT 76.950 835.950 79.050 838.050 ;
        RECT 79.950 835.950 82.050 838.050 ;
        RECT 82.950 835.950 85.050 838.050 ;
        RECT 85.950 835.950 88.050 838.050 ;
        RECT 100.950 835.950 103.050 838.050 ;
        RECT 103.950 835.950 106.050 838.050 ;
        RECT 106.950 835.950 109.050 838.050 ;
        RECT 109.950 835.950 112.050 838.050 ;
        RECT 127.950 835.950 130.050 838.050 ;
        RECT 130.950 835.950 133.050 838.050 ;
        RECT 133.950 835.950 136.050 838.050 ;
        RECT 136.950 835.950 139.050 838.050 ;
        RECT 151.950 835.950 154.050 838.050 ;
        RECT 154.950 835.950 157.050 838.050 ;
        RECT 158.550 837.750 163.050 838.050 ;
        RECT 158.550 835.950 164.850 837.750 ;
        RECT 17.100 825.600 18.300 835.950 ;
        RECT 35.250 834.150 37.050 835.950 ;
        RECT 38.100 830.700 39.300 835.950 ;
        RECT 41.100 834.150 42.900 835.950 ;
        RECT 56.100 834.150 57.900 835.950 ;
        RECT 59.700 830.700 60.900 835.950 ;
        RECT 61.950 834.150 63.750 835.950 ;
        RECT 77.100 834.150 78.900 835.950 ;
        RECT 83.100 834.150 84.900 835.950 ;
        RECT 86.100 832.200 87.000 835.950 ;
        RECT 101.100 834.150 102.900 835.950 ;
        RECT 107.250 834.150 109.050 835.950 ;
        RECT 38.100 829.800 42.300 830.700 ;
        RECT 14.100 822.000 15.900 825.600 ;
        RECT 17.100 822.600 18.900 825.600 ;
        RECT 35.400 822.000 37.200 828.600 ;
        RECT 40.500 822.600 42.300 829.800 ;
        RECT 56.700 829.800 60.900 830.700 ;
        RECT 56.700 822.600 58.500 829.800 ;
        RECT 61.800 822.000 63.600 828.600 ;
        RECT 77.100 822.000 78.900 831.600 ;
        RECT 83.700 831.000 87.000 832.200 ;
        RECT 83.700 822.600 85.500 831.000 ;
        RECT 110.700 828.600 111.600 835.950 ;
        RECT 128.100 834.150 129.900 835.950 ;
        RECT 134.250 834.150 136.050 835.950 ;
        RECT 137.700 828.600 138.600 835.950 ;
        RECT 102.000 822.000 103.800 828.600 ;
        RECT 106.500 827.400 111.600 828.600 ;
        RECT 106.500 822.600 108.300 827.400 ;
        RECT 109.500 822.000 111.300 825.600 ;
        RECT 129.000 822.000 130.800 828.600 ;
        RECT 133.500 827.400 138.600 828.600 ;
        RECT 133.500 822.600 135.300 827.400 ;
        RECT 152.700 825.600 153.900 835.950 ;
        RECT 158.550 828.600 159.750 835.950 ;
        RECT 171.150 832.200 172.050 844.800 ;
        RECT 174.150 844.800 175.050 846.900 ;
        RECT 175.950 846.300 183.750 847.500 ;
        RECT 175.950 845.700 177.750 846.300 ;
        RECT 187.050 845.400 188.850 858.000 ;
        RECT 190.050 847.200 191.850 857.400 ;
        RECT 206.100 851.400 207.900 857.400 ;
        RECT 209.100 852.000 210.900 858.000 ;
        RECT 207.000 851.100 207.900 851.400 ;
        RECT 212.100 851.400 213.900 857.400 ;
        RECT 215.100 851.400 216.900 858.000 ;
        RECT 212.100 851.100 213.600 851.400 ;
        RECT 207.000 850.200 213.600 851.100 ;
        RECT 190.050 845.400 192.450 847.200 ;
        RECT 174.150 844.500 182.550 844.800 ;
        RECT 191.550 844.500 192.450 845.400 ;
        RECT 174.150 843.900 192.450 844.500 ;
        RECT 180.750 843.300 192.450 843.900 ;
        RECT 180.750 843.000 182.550 843.300 ;
        RECT 178.800 836.400 180.900 838.050 ;
        RECT 178.800 835.200 186.900 836.400 ;
        RECT 187.950 835.950 190.050 838.050 ;
        RECT 185.100 834.600 186.900 835.200 ;
        RECT 182.100 833.400 183.900 834.000 ;
        RECT 188.250 833.400 190.050 835.950 ;
        RECT 182.100 832.200 190.050 833.400 ;
        RECT 171.150 831.000 183.150 832.200 ;
        RECT 171.150 830.400 172.950 831.000 ;
        RECT 182.100 829.200 183.150 831.000 ;
        RECT 136.500 822.000 138.300 825.600 ;
        RECT 152.100 822.600 153.900 825.600 ;
        RECT 155.100 822.000 156.900 825.600 ;
        RECT 158.550 822.600 160.350 828.600 ;
        RECT 161.850 822.000 163.650 828.600 ;
        RECT 166.350 825.600 168.750 827.700 ;
        RECT 178.350 827.550 180.150 828.300 ;
        RECT 175.200 826.500 180.150 827.550 ;
        RECT 181.350 827.400 183.150 829.200 ;
        RECT 191.550 828.600 192.450 843.300 ;
        RECT 207.000 838.050 207.900 850.200 ;
        RECT 230.100 846.300 231.900 857.400 ;
        RECT 233.100 847.200 234.900 858.000 ;
        RECT 236.100 846.300 237.900 857.400 ;
        RECT 230.100 845.400 237.900 846.300 ;
        RECT 239.100 845.400 240.900 857.400 ;
        RECT 254.100 851.400 255.900 857.400 ;
        RECT 257.100 852.000 258.900 858.000 ;
        RECT 255.000 851.100 255.900 851.400 ;
        RECT 260.100 851.400 261.900 857.400 ;
        RECT 263.100 851.400 264.900 858.000 ;
        RECT 281.100 851.400 282.900 857.400 ;
        RECT 284.100 852.000 285.900 858.000 ;
        RECT 260.100 851.100 261.600 851.400 ;
        RECT 255.000 850.200 261.600 851.100 ;
        RECT 282.000 851.100 282.900 851.400 ;
        RECT 287.100 851.400 288.900 857.400 ;
        RECT 290.100 851.400 291.900 858.000 ;
        RECT 305.700 851.400 307.500 858.000 ;
        RECT 287.100 851.100 288.600 851.400 ;
        RECT 282.000 850.200 288.600 851.100 ;
        RECT 212.100 838.050 213.900 839.850 ;
        RECT 233.250 838.050 235.050 839.850 ;
        RECT 239.700 838.050 240.600 845.400 ;
        RECT 255.000 838.050 255.900 850.200 ;
        RECT 260.100 838.050 261.900 839.850 ;
        RECT 282.000 838.050 282.900 850.200 ;
        RECT 306.000 848.100 307.800 849.900 ;
        RECT 308.700 846.900 310.500 857.400 ;
        RECT 308.100 845.400 310.500 846.900 ;
        RECT 313.800 845.400 315.600 858.000 ;
        RECT 317.550 845.400 319.350 857.400 ;
        RECT 320.550 845.400 322.350 858.000 ;
        RECT 325.350 851.400 327.150 857.400 ;
        RECT 329.850 851.400 331.650 858.000 ;
        RECT 325.350 849.300 327.450 851.400 ;
        RECT 332.850 850.500 334.650 857.400 ;
        RECT 335.850 851.400 337.650 858.000 ;
        RECT 331.950 849.450 338.550 850.500 ;
        RECT 331.950 848.700 333.750 849.450 ;
        RECT 336.750 848.700 338.550 849.450 ;
        RECT 340.650 848.400 342.450 857.400 ;
        RECT 324.450 846.600 327.450 848.400 ;
        RECT 328.350 847.800 330.150 848.400 ;
        RECT 328.350 846.900 334.050 847.800 ;
        RECT 340.650 847.500 342.750 848.400 ;
        RECT 328.350 846.600 330.150 846.900 ;
        RECT 326.250 845.700 327.450 846.600 ;
        RECT 287.100 838.050 288.900 839.850 ;
        RECT 308.100 838.050 309.300 845.400 ;
        RECT 314.100 838.050 315.900 839.850 ;
        RECT 317.550 838.050 318.750 845.400 ;
        RECT 326.250 844.800 331.050 845.700 ;
        RECT 319.650 842.100 321.450 842.550 ;
        RECT 325.350 842.100 327.450 842.700 ;
        RECT 319.650 840.900 327.450 842.100 ;
        RECT 319.650 840.750 321.450 840.900 ;
        RECT 325.350 840.600 327.450 840.900 ;
        RECT 205.950 835.950 208.050 838.050 ;
        RECT 208.950 835.950 211.050 838.050 ;
        RECT 211.950 835.950 214.050 838.050 ;
        RECT 214.950 835.950 217.050 838.050 ;
        RECT 229.950 835.950 232.050 838.050 ;
        RECT 232.950 835.950 235.050 838.050 ;
        RECT 235.950 835.950 238.050 838.050 ;
        RECT 238.950 835.950 241.050 838.050 ;
        RECT 253.950 835.950 256.050 838.050 ;
        RECT 256.950 835.950 259.050 838.050 ;
        RECT 259.950 835.950 262.050 838.050 ;
        RECT 262.950 835.950 265.050 838.050 ;
        RECT 280.950 835.950 283.050 838.050 ;
        RECT 283.950 835.950 286.050 838.050 ;
        RECT 286.950 835.950 289.050 838.050 ;
        RECT 289.950 835.950 292.050 838.050 ;
        RECT 304.950 835.950 307.050 838.050 ;
        RECT 307.950 835.950 310.050 838.050 ;
        RECT 310.950 835.950 313.050 838.050 ;
        RECT 313.950 835.950 316.050 838.050 ;
        RECT 317.550 837.750 322.050 838.050 ;
        RECT 317.550 835.950 323.850 837.750 ;
        RECT 207.000 832.200 207.900 835.950 ;
        RECT 209.100 834.150 210.900 835.950 ;
        RECT 215.100 834.150 216.900 835.950 ;
        RECT 230.100 834.150 231.900 835.950 ;
        RECT 236.250 834.150 238.050 835.950 ;
        RECT 207.000 831.000 210.300 832.200 ;
        RECT 175.200 825.600 176.250 826.500 ;
        RECT 184.050 826.200 186.150 827.700 ;
        RECT 182.250 825.600 186.150 826.200 ;
        RECT 166.950 822.600 168.750 825.600 ;
        RECT 171.450 822.000 173.250 825.600 ;
        RECT 174.450 822.600 176.250 825.600 ;
        RECT 177.750 822.000 179.550 825.600 ;
        RECT 182.250 824.700 185.850 825.600 ;
        RECT 182.250 822.600 184.050 824.700 ;
        RECT 187.050 822.000 188.850 828.600 ;
        RECT 190.050 826.800 192.450 828.600 ;
        RECT 190.050 822.600 191.850 826.800 ;
        RECT 208.500 822.600 210.300 831.000 ;
        RECT 215.100 822.000 216.900 831.600 ;
        RECT 239.700 828.600 240.600 835.950 ;
        RECT 255.000 832.200 255.900 835.950 ;
        RECT 257.100 834.150 258.900 835.950 ;
        RECT 263.100 834.150 264.900 835.950 ;
        RECT 282.000 832.200 282.900 835.950 ;
        RECT 284.100 834.150 285.900 835.950 ;
        RECT 290.100 834.150 291.900 835.950 ;
        RECT 305.100 834.150 306.900 835.950 ;
        RECT 255.000 831.000 258.300 832.200 ;
        RECT 231.000 822.000 232.800 828.600 ;
        RECT 235.500 827.400 240.600 828.600 ;
        RECT 235.500 822.600 237.300 827.400 ;
        RECT 238.500 822.000 240.300 825.600 ;
        RECT 256.500 822.600 258.300 831.000 ;
        RECT 263.100 822.000 264.900 831.600 ;
        RECT 282.000 831.000 285.300 832.200 ;
        RECT 308.100 831.600 309.300 835.950 ;
        RECT 311.100 834.150 312.900 835.950 ;
        RECT 283.500 822.600 285.300 831.000 ;
        RECT 290.100 822.000 291.900 831.600 ;
        RECT 305.700 830.700 309.300 831.600 ;
        RECT 305.700 828.600 306.900 830.700 ;
        RECT 305.100 822.600 306.900 828.600 ;
        RECT 308.100 827.700 315.900 829.050 ;
        RECT 308.100 822.600 309.900 827.700 ;
        RECT 311.100 822.000 312.900 826.800 ;
        RECT 314.100 822.600 315.900 827.700 ;
        RECT 317.550 828.600 318.750 835.950 ;
        RECT 330.150 832.200 331.050 844.800 ;
        RECT 333.150 844.800 334.050 846.900 ;
        RECT 334.950 846.300 342.750 847.500 ;
        RECT 334.950 845.700 336.750 846.300 ;
        RECT 346.050 845.400 347.850 858.000 ;
        RECT 349.050 847.200 350.850 857.400 ;
        RECT 349.050 845.400 351.450 847.200 ;
        RECT 333.150 844.500 341.550 844.800 ;
        RECT 350.550 844.500 351.450 845.400 ;
        RECT 333.150 843.900 351.450 844.500 ;
        RECT 339.750 843.300 351.450 843.900 ;
        RECT 339.750 843.000 341.550 843.300 ;
        RECT 337.800 836.400 339.900 838.050 ;
        RECT 337.800 835.200 345.900 836.400 ;
        RECT 346.950 835.950 349.050 838.050 ;
        RECT 344.100 834.600 345.900 835.200 ;
        RECT 341.100 833.400 342.900 834.000 ;
        RECT 347.250 833.400 349.050 835.950 ;
        RECT 341.100 832.200 349.050 833.400 ;
        RECT 330.150 831.000 342.150 832.200 ;
        RECT 330.150 830.400 331.950 831.000 ;
        RECT 341.100 829.200 342.150 831.000 ;
        RECT 317.550 822.600 319.350 828.600 ;
        RECT 320.850 822.000 322.650 828.600 ;
        RECT 325.350 825.600 327.750 827.700 ;
        RECT 337.350 827.550 339.150 828.300 ;
        RECT 334.200 826.500 339.150 827.550 ;
        RECT 340.350 827.400 342.150 829.200 ;
        RECT 350.550 828.600 351.450 843.300 ;
        RECT 334.200 825.600 335.250 826.500 ;
        RECT 343.050 826.200 345.150 827.700 ;
        RECT 341.250 825.600 345.150 826.200 ;
        RECT 325.950 822.600 327.750 825.600 ;
        RECT 330.450 822.000 332.250 825.600 ;
        RECT 333.450 822.600 335.250 825.600 ;
        RECT 336.750 822.000 338.550 825.600 ;
        RECT 341.250 824.700 344.850 825.600 ;
        RECT 341.250 822.600 343.050 824.700 ;
        RECT 346.050 822.000 347.850 828.600 ;
        RECT 349.050 826.800 351.450 828.600 ;
        RECT 353.550 845.400 355.350 857.400 ;
        RECT 356.550 845.400 358.350 858.000 ;
        RECT 361.350 851.400 363.150 857.400 ;
        RECT 365.850 851.400 367.650 858.000 ;
        RECT 361.350 849.300 363.450 851.400 ;
        RECT 368.850 850.500 370.650 857.400 ;
        RECT 371.850 851.400 373.650 858.000 ;
        RECT 367.950 849.450 374.550 850.500 ;
        RECT 367.950 848.700 369.750 849.450 ;
        RECT 372.750 848.700 374.550 849.450 ;
        RECT 376.650 848.400 378.450 857.400 ;
        RECT 360.450 846.600 363.450 848.400 ;
        RECT 364.350 847.800 366.150 848.400 ;
        RECT 364.350 846.900 370.050 847.800 ;
        RECT 376.650 847.500 378.750 848.400 ;
        RECT 364.350 846.600 366.150 846.900 ;
        RECT 362.250 845.700 363.450 846.600 ;
        RECT 353.550 838.050 354.750 845.400 ;
        RECT 362.250 844.800 367.050 845.700 ;
        RECT 355.650 842.100 357.450 842.550 ;
        RECT 361.350 842.100 363.450 842.700 ;
        RECT 355.650 840.900 363.450 842.100 ;
        RECT 355.650 840.750 357.450 840.900 ;
        RECT 361.350 840.600 363.450 840.900 ;
        RECT 353.550 837.750 358.050 838.050 ;
        RECT 353.550 835.950 359.850 837.750 ;
        RECT 353.550 828.600 354.750 835.950 ;
        RECT 366.150 832.200 367.050 844.800 ;
        RECT 369.150 844.800 370.050 846.900 ;
        RECT 370.950 846.300 378.750 847.500 ;
        RECT 370.950 845.700 372.750 846.300 ;
        RECT 382.050 845.400 383.850 858.000 ;
        RECT 385.050 847.200 386.850 857.400 ;
        RECT 385.050 845.400 387.450 847.200 ;
        RECT 404.400 845.400 406.200 858.000 ;
        RECT 409.500 846.900 411.300 857.400 ;
        RECT 412.500 851.400 414.300 858.000 ;
        RECT 412.200 848.100 414.000 849.900 ;
        RECT 409.500 845.400 411.900 846.900 ;
        RECT 431.100 846.600 432.900 857.400 ;
        RECT 434.100 847.500 435.900 858.000 ;
        RECT 431.100 845.400 435.900 846.600 ;
        RECT 369.150 844.500 377.550 844.800 ;
        RECT 386.550 844.500 387.450 845.400 ;
        RECT 369.150 843.900 387.450 844.500 ;
        RECT 375.750 843.300 387.450 843.900 ;
        RECT 375.750 843.000 377.550 843.300 ;
        RECT 373.800 836.400 375.900 838.050 ;
        RECT 373.800 835.200 381.900 836.400 ;
        RECT 382.950 835.950 385.050 838.050 ;
        RECT 380.100 834.600 381.900 835.200 ;
        RECT 377.100 833.400 378.900 834.000 ;
        RECT 383.250 833.400 385.050 835.950 ;
        RECT 377.100 832.200 385.050 833.400 ;
        RECT 366.150 831.000 378.150 832.200 ;
        RECT 366.150 830.400 367.950 831.000 ;
        RECT 377.100 829.200 378.150 831.000 ;
        RECT 349.050 822.600 350.850 826.800 ;
        RECT 353.550 822.600 355.350 828.600 ;
        RECT 356.850 822.000 358.650 828.600 ;
        RECT 361.350 825.600 363.750 827.700 ;
        RECT 373.350 827.550 375.150 828.300 ;
        RECT 370.200 826.500 375.150 827.550 ;
        RECT 376.350 827.400 378.150 829.200 ;
        RECT 386.550 828.600 387.450 843.300 ;
        RECT 404.100 838.050 405.900 839.850 ;
        RECT 410.700 838.050 411.900 845.400 ;
        RECT 433.800 844.500 435.900 845.400 ;
        RECT 438.600 845.400 440.400 857.400 ;
        RECT 443.100 847.500 444.900 858.000 ;
        RECT 446.100 846.300 447.900 857.400 ;
        RECT 443.400 845.400 447.900 846.300 ;
        RECT 461.100 845.400 462.900 858.000 ;
        RECT 438.600 844.050 439.800 845.400 ;
        RECT 438.300 843.000 439.800 844.050 ;
        RECT 443.400 843.300 445.500 845.400 ;
        RECT 464.100 844.500 465.900 857.400 ;
        RECT 467.100 845.400 468.900 858.000 ;
        RECT 470.100 844.500 471.900 857.400 ;
        RECT 473.100 845.400 474.900 858.000 ;
        RECT 476.100 844.500 477.900 857.400 ;
        RECT 479.100 845.400 480.900 858.000 ;
        RECT 482.100 844.500 483.900 857.400 ;
        RECT 485.100 845.400 486.900 858.000 ;
        RECT 488.550 845.400 490.350 857.400 ;
        RECT 491.550 845.400 493.350 858.000 ;
        RECT 496.350 851.400 498.150 857.400 ;
        RECT 500.850 851.400 502.650 858.000 ;
        RECT 496.350 849.300 498.450 851.400 ;
        RECT 503.850 850.500 505.650 857.400 ;
        RECT 506.850 851.400 508.650 858.000 ;
        RECT 502.950 849.450 509.550 850.500 ;
        RECT 502.950 848.700 504.750 849.450 ;
        RECT 507.750 848.700 509.550 849.450 ;
        RECT 511.650 848.400 513.450 857.400 ;
        RECT 495.450 846.600 498.450 848.400 ;
        RECT 499.350 847.800 501.150 848.400 ;
        RECT 499.350 846.900 505.050 847.800 ;
        RECT 511.650 847.500 513.750 848.400 ;
        RECT 499.350 846.600 501.150 846.900 ;
        RECT 497.250 845.700 498.450 846.600 ;
        RECT 464.100 843.300 468.000 844.500 ;
        RECT 470.100 843.300 474.000 844.500 ;
        RECT 476.100 843.300 480.000 844.500 ;
        RECT 482.100 843.300 484.950 844.500 ;
        RECT 438.300 841.050 439.200 843.000 ;
        RECT 431.400 838.050 433.200 839.850 ;
        RECT 437.100 838.950 439.200 841.050 ;
        RECT 440.100 841.500 442.200 841.800 ;
        RECT 440.100 839.700 444.000 841.500 ;
        RECT 403.950 835.950 406.050 838.050 ;
        RECT 406.950 835.950 409.050 838.050 ;
        RECT 409.950 835.950 412.050 838.050 ;
        RECT 412.950 835.950 415.050 838.050 ;
        RECT 431.100 835.950 433.200 838.050 ;
        RECT 437.700 838.800 439.200 838.950 ;
        RECT 437.700 837.900 440.100 838.800 ;
        RECT 407.100 834.150 408.900 835.950 ;
        RECT 410.700 831.600 411.900 835.950 ;
        RECT 413.100 834.150 414.900 835.950 ;
        RECT 435.900 835.200 437.700 837.000 ;
        RECT 435.900 833.100 438.000 835.200 ;
        RECT 438.900 832.200 440.100 837.900 ;
        RECT 441.000 838.050 442.800 838.500 ;
        RECT 441.000 836.700 447.900 838.050 ;
        RECT 445.800 835.950 447.900 836.700 ;
        RECT 463.800 835.950 465.900 838.050 ;
        RECT 410.700 830.700 414.300 831.600 ;
        RECT 370.200 825.600 371.250 826.500 ;
        RECT 379.050 826.200 381.150 827.700 ;
        RECT 377.250 825.600 381.150 826.200 ;
        RECT 361.950 822.600 363.750 825.600 ;
        RECT 366.450 822.000 368.250 825.600 ;
        RECT 369.450 822.600 371.250 825.600 ;
        RECT 372.750 822.000 374.550 825.600 ;
        RECT 377.250 824.700 380.850 825.600 ;
        RECT 377.250 822.600 379.050 824.700 ;
        RECT 382.050 822.000 383.850 828.600 ;
        RECT 385.050 826.800 387.450 828.600 ;
        RECT 404.100 827.700 411.900 829.050 ;
        RECT 385.050 822.600 386.850 826.800 ;
        RECT 404.100 822.600 405.900 827.700 ;
        RECT 407.100 822.000 408.900 826.800 ;
        RECT 410.100 822.600 411.900 827.700 ;
        RECT 413.100 828.600 414.300 830.700 ;
        RECT 433.800 829.500 435.900 830.700 ;
        RECT 437.100 830.100 440.100 832.200 ;
        RECT 441.000 833.400 442.800 835.200 ;
        RECT 445.800 834.150 447.600 835.950 ;
        RECT 463.800 834.150 465.600 835.950 ;
        RECT 441.000 831.300 443.100 833.400 ;
        RECT 466.800 832.800 468.000 843.300 ;
        RECT 469.200 832.800 471.000 833.400 ;
        RECT 466.800 831.600 471.000 832.800 ;
        RECT 472.800 832.800 474.000 843.300 ;
        RECT 475.200 832.800 477.000 833.400 ;
        RECT 472.800 831.600 477.000 832.800 ;
        RECT 478.800 832.800 480.000 843.300 ;
        RECT 483.900 838.050 484.950 843.300 ;
        RECT 481.800 835.950 484.950 838.050 ;
        RECT 481.200 832.800 483.000 833.400 ;
        RECT 478.800 831.600 483.000 832.800 ;
        RECT 441.000 830.400 447.300 831.300 ;
        RECT 466.800 830.700 468.000 831.600 ;
        RECT 472.800 830.700 474.000 831.600 ;
        RECT 478.800 830.700 480.000 831.600 ;
        RECT 483.900 830.700 484.950 835.950 ;
        RECT 431.100 828.600 435.900 829.500 ;
        RECT 438.900 828.600 440.100 830.100 ;
        RECT 446.100 828.600 447.300 830.400 ;
        RECT 464.100 829.500 468.000 830.700 ;
        RECT 470.100 829.500 474.000 830.700 ;
        RECT 476.100 829.500 480.000 830.700 ;
        RECT 482.100 829.500 484.950 830.700 ;
        RECT 488.550 838.050 489.750 845.400 ;
        RECT 497.250 844.800 502.050 845.700 ;
        RECT 490.650 842.100 492.450 842.550 ;
        RECT 496.350 842.100 498.450 842.700 ;
        RECT 490.650 840.900 498.450 842.100 ;
        RECT 490.650 840.750 492.450 840.900 ;
        RECT 496.350 840.600 498.450 840.900 ;
        RECT 488.550 837.750 493.050 838.050 ;
        RECT 488.550 835.950 494.850 837.750 ;
        RECT 413.100 822.600 414.900 828.600 ;
        RECT 431.100 822.600 432.900 828.600 ;
        RECT 434.100 822.000 435.900 827.700 ;
        RECT 438.600 822.600 440.400 828.600 ;
        RECT 443.100 822.000 444.900 827.700 ;
        RECT 446.100 822.600 447.900 828.600 ;
        RECT 461.100 822.000 462.900 828.600 ;
        RECT 464.100 822.600 465.900 829.500 ;
        RECT 467.100 822.000 468.900 828.600 ;
        RECT 470.100 822.600 471.900 829.500 ;
        RECT 473.100 822.000 474.900 828.600 ;
        RECT 476.100 822.600 477.900 829.500 ;
        RECT 479.100 822.000 480.900 828.600 ;
        RECT 482.100 822.600 483.900 829.500 ;
        RECT 488.550 828.600 489.750 835.950 ;
        RECT 501.150 832.200 502.050 844.800 ;
        RECT 504.150 844.800 505.050 846.900 ;
        RECT 505.950 846.300 513.750 847.500 ;
        RECT 505.950 845.700 507.750 846.300 ;
        RECT 517.050 845.400 518.850 858.000 ;
        RECT 520.050 847.200 521.850 857.400 ;
        RECT 520.050 845.400 522.450 847.200 ;
        RECT 536.100 845.400 537.900 858.000 ;
        RECT 541.200 846.600 543.000 857.400 ;
        RECT 539.400 845.400 543.000 846.600 ;
        RECT 560.100 845.400 561.900 857.400 ;
        RECT 563.100 846.300 564.900 857.400 ;
        RECT 566.100 847.200 567.900 858.000 ;
        RECT 569.100 846.300 570.900 857.400 ;
        RECT 584.100 851.400 585.900 857.400 ;
        RECT 587.100 852.000 588.900 858.000 ;
        RECT 563.100 845.400 570.900 846.300 ;
        RECT 585.000 851.100 585.900 851.400 ;
        RECT 590.100 851.400 591.900 857.400 ;
        RECT 593.100 851.400 594.900 858.000 ;
        RECT 611.700 851.400 613.500 858.000 ;
        RECT 590.100 851.100 591.600 851.400 ;
        RECT 585.000 850.200 591.600 851.100 ;
        RECT 504.150 844.500 512.550 844.800 ;
        RECT 521.550 844.500 522.450 845.400 ;
        RECT 504.150 843.900 522.450 844.500 ;
        RECT 510.750 843.300 522.450 843.900 ;
        RECT 510.750 843.000 512.550 843.300 ;
        RECT 508.800 836.400 510.900 838.050 ;
        RECT 508.800 835.200 516.900 836.400 ;
        RECT 517.950 835.950 520.050 838.050 ;
        RECT 515.100 834.600 516.900 835.200 ;
        RECT 512.100 833.400 513.900 834.000 ;
        RECT 518.250 833.400 520.050 835.950 ;
        RECT 512.100 832.200 520.050 833.400 ;
        RECT 501.150 831.000 513.150 832.200 ;
        RECT 501.150 830.400 502.950 831.000 ;
        RECT 512.100 829.200 513.150 831.000 ;
        RECT 485.100 822.000 486.900 828.600 ;
        RECT 488.550 822.600 490.350 828.600 ;
        RECT 491.850 822.000 493.650 828.600 ;
        RECT 496.350 825.600 498.750 827.700 ;
        RECT 508.350 827.550 510.150 828.300 ;
        RECT 505.200 826.500 510.150 827.550 ;
        RECT 511.350 827.400 513.150 829.200 ;
        RECT 521.550 828.600 522.450 843.300 ;
        RECT 536.250 838.050 538.050 839.850 ;
        RECT 539.400 838.050 540.300 845.400 ;
        RECT 542.100 838.050 543.900 839.850 ;
        RECT 560.400 838.050 561.300 845.400 ;
        RECT 565.950 838.050 567.750 839.850 ;
        RECT 585.000 838.050 585.900 850.200 ;
        RECT 612.000 848.100 613.800 849.900 ;
        RECT 614.700 846.900 616.500 857.400 ;
        RECT 614.100 845.400 616.500 846.900 ;
        RECT 619.800 845.400 621.600 858.000 ;
        RECT 635.400 845.400 637.200 858.000 ;
        RECT 640.500 846.900 642.300 857.400 ;
        RECT 643.500 851.400 645.300 858.000 ;
        RECT 659.100 851.400 660.900 858.000 ;
        RECT 662.100 851.400 663.900 857.400 ;
        RECT 677.100 851.400 678.900 857.400 ;
        RECT 680.100 852.000 681.900 858.000 ;
        RECT 643.200 848.100 645.000 849.900 ;
        RECT 640.500 845.400 642.900 846.900 ;
        RECT 586.950 843.450 589.050 844.050 ;
        RECT 598.950 843.450 601.050 844.050 ;
        RECT 586.950 842.550 601.050 843.450 ;
        RECT 586.950 841.950 589.050 842.550 ;
        RECT 598.950 841.950 601.050 842.550 ;
        RECT 590.100 838.050 591.900 839.850 ;
        RECT 614.100 838.050 615.300 845.400 ;
        RECT 620.100 838.050 621.900 839.850 ;
        RECT 635.100 838.050 636.900 839.850 ;
        RECT 641.700 838.050 642.900 845.400 ;
        RECT 659.100 838.050 660.900 839.850 ;
        RECT 662.100 838.050 663.300 851.400 ;
        RECT 678.000 851.100 678.900 851.400 ;
        RECT 683.100 851.400 684.900 857.400 ;
        RECT 686.100 851.400 687.900 858.000 ;
        RECT 683.100 851.100 684.600 851.400 ;
        RECT 678.000 850.200 684.600 851.100 ;
        RECT 678.000 838.050 678.900 850.200 ;
        RECT 701.100 845.400 702.900 857.400 ;
        RECT 704.100 846.300 705.900 857.400 ;
        RECT 707.100 847.200 708.900 858.000 ;
        RECT 710.100 846.300 711.900 857.400 ;
        RECT 725.100 851.400 726.900 857.400 ;
        RECT 728.100 852.000 729.900 858.000 ;
        RECT 704.100 845.400 711.900 846.300 ;
        RECT 726.000 851.100 726.900 851.400 ;
        RECT 731.100 851.400 732.900 857.400 ;
        RECT 734.100 851.400 735.900 858.000 ;
        RECT 731.100 851.100 732.600 851.400 ;
        RECT 726.000 850.200 732.600 851.100 ;
        RECT 683.100 838.050 684.900 839.850 ;
        RECT 701.400 838.050 702.300 845.400 ;
        RECT 706.950 838.050 708.750 839.850 ;
        RECT 726.000 838.050 726.900 850.200 ;
        RECT 752.100 845.400 753.900 857.400 ;
        RECT 755.100 846.300 756.900 857.400 ;
        RECT 758.100 847.200 759.900 858.000 ;
        RECT 761.100 846.300 762.900 857.400 ;
        RECT 755.100 845.400 762.900 846.300 ;
        RECT 776.100 845.400 777.900 857.400 ;
        RECT 779.100 846.300 780.900 857.400 ;
        RECT 782.100 847.200 783.900 858.000 ;
        RECT 785.100 846.300 786.900 857.400 ;
        RECT 800.100 851.400 801.900 857.400 ;
        RECT 803.100 852.000 804.900 858.000 ;
        RECT 779.100 845.400 786.900 846.300 ;
        RECT 801.000 851.100 801.900 851.400 ;
        RECT 806.100 851.400 807.900 857.400 ;
        RECT 809.100 851.400 810.900 858.000 ;
        RECT 824.100 851.400 825.900 857.400 ;
        RECT 827.100 852.000 828.900 858.000 ;
        RECT 806.100 851.100 807.600 851.400 ;
        RECT 801.000 850.200 807.600 851.100 ;
        RECT 825.000 851.100 825.900 851.400 ;
        RECT 830.100 851.400 831.900 857.400 ;
        RECT 833.100 851.400 834.900 858.000 ;
        RECT 848.100 851.400 849.900 858.000 ;
        RECT 851.100 851.400 852.900 857.400 ;
        RECT 854.100 852.000 855.900 858.000 ;
        RECT 830.100 851.100 831.600 851.400 ;
        RECT 825.000 850.200 831.600 851.100 ;
        RECT 851.400 851.100 852.900 851.400 ;
        RECT 857.100 851.400 858.900 857.400 ;
        RECT 872.100 851.400 873.900 858.000 ;
        RECT 875.100 851.400 876.900 857.400 ;
        RECT 878.100 851.400 879.900 858.000 ;
        RECT 893.100 851.400 894.900 857.400 ;
        RECT 896.100 851.400 897.900 858.000 ;
        RECT 857.100 851.100 858.000 851.400 ;
        RECT 851.400 850.200 858.000 851.100 ;
        RECT 731.100 838.050 732.900 839.850 ;
        RECT 752.400 838.050 753.300 845.400 ;
        RECT 757.950 838.050 759.750 839.850 ;
        RECT 776.400 838.050 777.300 845.400 ;
        RECT 781.950 838.050 783.750 839.850 ;
        RECT 801.000 838.050 801.900 850.200 ;
        RECT 808.950 843.450 811.050 844.200 ;
        RECT 817.950 843.450 820.050 844.050 ;
        RECT 808.950 842.550 820.050 843.450 ;
        RECT 808.950 842.100 811.050 842.550 ;
        RECT 817.950 841.950 820.050 842.550 ;
        RECT 806.100 838.050 807.900 839.850 ;
        RECT 825.000 838.050 825.900 850.200 ;
        RECT 826.950 843.450 829.050 844.050 ;
        RECT 850.950 843.450 853.050 844.050 ;
        RECT 826.950 842.550 853.050 843.450 ;
        RECT 826.950 841.950 829.050 842.550 ;
        RECT 850.950 841.950 853.050 842.550 ;
        RECT 830.100 838.050 831.900 839.850 ;
        RECT 851.100 838.050 852.900 839.850 ;
        RECT 857.100 838.050 858.000 850.200 ;
        RECT 859.950 840.450 862.050 841.050 ;
        RECT 859.950 839.550 867.450 840.450 ;
        RECT 859.950 838.950 862.050 839.550 ;
        RECT 535.950 835.950 538.050 838.050 ;
        RECT 538.950 835.950 541.050 838.050 ;
        RECT 541.950 835.950 544.050 838.050 ;
        RECT 559.950 835.950 562.050 838.050 ;
        RECT 562.950 835.950 565.050 838.050 ;
        RECT 565.950 835.950 568.050 838.050 ;
        RECT 568.950 835.950 571.050 838.050 ;
        RECT 583.950 835.950 586.050 838.050 ;
        RECT 586.950 835.950 589.050 838.050 ;
        RECT 589.950 835.950 592.050 838.050 ;
        RECT 592.950 835.950 595.050 838.050 ;
        RECT 610.950 835.950 613.050 838.050 ;
        RECT 613.950 835.950 616.050 838.050 ;
        RECT 616.950 835.950 619.050 838.050 ;
        RECT 619.950 835.950 622.050 838.050 ;
        RECT 634.950 835.950 637.050 838.050 ;
        RECT 637.950 835.950 640.050 838.050 ;
        RECT 640.950 835.950 643.050 838.050 ;
        RECT 643.950 835.950 646.050 838.050 ;
        RECT 658.950 835.950 661.050 838.050 ;
        RECT 661.950 835.950 664.050 838.050 ;
        RECT 676.950 835.950 679.050 838.050 ;
        RECT 679.950 835.950 682.050 838.050 ;
        RECT 682.950 835.950 685.050 838.050 ;
        RECT 685.950 835.950 688.050 838.050 ;
        RECT 700.950 835.950 703.050 838.050 ;
        RECT 703.950 835.950 706.050 838.050 ;
        RECT 706.950 835.950 709.050 838.050 ;
        RECT 709.950 835.950 712.050 838.050 ;
        RECT 724.950 835.950 727.050 838.050 ;
        RECT 727.950 835.950 730.050 838.050 ;
        RECT 730.950 835.950 733.050 838.050 ;
        RECT 733.950 835.950 736.050 838.050 ;
        RECT 751.950 835.950 754.050 838.050 ;
        RECT 754.950 835.950 757.050 838.050 ;
        RECT 757.950 835.950 760.050 838.050 ;
        RECT 760.950 835.950 763.050 838.050 ;
        RECT 775.950 835.950 778.050 838.050 ;
        RECT 778.950 835.950 781.050 838.050 ;
        RECT 781.950 835.950 784.050 838.050 ;
        RECT 784.950 835.950 787.050 838.050 ;
        RECT 799.950 835.950 802.050 838.050 ;
        RECT 802.950 835.950 805.050 838.050 ;
        RECT 805.950 835.950 808.050 838.050 ;
        RECT 808.950 835.950 811.050 838.050 ;
        RECT 823.950 835.950 826.050 838.050 ;
        RECT 826.950 835.950 829.050 838.050 ;
        RECT 829.950 835.950 832.050 838.050 ;
        RECT 832.950 835.950 835.050 838.050 ;
        RECT 847.950 835.950 850.050 838.050 ;
        RECT 850.950 835.950 853.050 838.050 ;
        RECT 853.950 835.950 856.050 838.050 ;
        RECT 856.950 835.950 859.050 838.050 ;
        RECT 505.200 825.600 506.250 826.500 ;
        RECT 514.050 826.200 516.150 827.700 ;
        RECT 512.250 825.600 516.150 826.200 ;
        RECT 496.950 822.600 498.750 825.600 ;
        RECT 501.450 822.000 503.250 825.600 ;
        RECT 504.450 822.600 506.250 825.600 ;
        RECT 507.750 822.000 509.550 825.600 ;
        RECT 512.250 824.700 515.850 825.600 ;
        RECT 512.250 822.600 514.050 824.700 ;
        RECT 517.050 822.000 518.850 828.600 ;
        RECT 520.050 826.800 522.450 828.600 ;
        RECT 520.050 822.600 521.850 826.800 ;
        RECT 539.400 825.600 540.300 835.950 ;
        RECT 560.400 828.600 561.300 835.950 ;
        RECT 562.950 834.150 564.750 835.950 ;
        RECT 569.100 834.150 570.900 835.950 ;
        RECT 585.000 832.200 585.900 835.950 ;
        RECT 587.100 834.150 588.900 835.950 ;
        RECT 593.100 834.150 594.900 835.950 ;
        RECT 611.100 834.150 612.900 835.950 ;
        RECT 585.000 831.000 588.300 832.200 ;
        RECT 614.100 831.600 615.300 835.950 ;
        RECT 617.100 834.150 618.900 835.950 ;
        RECT 638.100 834.150 639.900 835.950 ;
        RECT 560.400 827.400 565.500 828.600 ;
        RECT 536.100 822.000 537.900 825.600 ;
        RECT 539.100 822.600 540.900 825.600 ;
        RECT 542.100 822.000 543.900 825.600 ;
        RECT 560.700 822.000 562.500 825.600 ;
        RECT 563.700 822.600 565.500 827.400 ;
        RECT 568.200 822.000 570.000 828.600 ;
        RECT 586.500 822.600 588.300 831.000 ;
        RECT 593.100 822.000 594.900 831.600 ;
        RECT 611.700 830.700 615.300 831.600 ;
        RECT 641.700 831.600 642.900 835.950 ;
        RECT 644.100 834.150 645.900 835.950 ;
        RECT 641.700 830.700 645.300 831.600 ;
        RECT 611.700 828.600 612.900 830.700 ;
        RECT 611.100 822.600 612.900 828.600 ;
        RECT 614.100 827.700 621.900 829.050 ;
        RECT 614.100 822.600 615.900 827.700 ;
        RECT 617.100 822.000 618.900 826.800 ;
        RECT 620.100 822.600 621.900 827.700 ;
        RECT 635.100 827.700 642.900 829.050 ;
        RECT 635.100 822.600 636.900 827.700 ;
        RECT 638.100 822.000 639.900 826.800 ;
        RECT 641.100 822.600 642.900 827.700 ;
        RECT 644.100 828.600 645.300 830.700 ;
        RECT 644.100 822.600 645.900 828.600 ;
        RECT 662.100 825.600 663.300 835.950 ;
        RECT 678.000 832.200 678.900 835.950 ;
        RECT 680.100 834.150 681.900 835.950 ;
        RECT 686.100 834.150 687.900 835.950 ;
        RECT 678.000 831.000 681.300 832.200 ;
        RECT 659.100 822.000 660.900 825.600 ;
        RECT 662.100 822.600 663.900 825.600 ;
        RECT 679.500 822.600 681.300 831.000 ;
        RECT 686.100 822.000 687.900 831.600 ;
        RECT 701.400 828.600 702.300 835.950 ;
        RECT 703.950 834.150 705.750 835.950 ;
        RECT 710.100 834.150 711.900 835.950 ;
        RECT 726.000 832.200 726.900 835.950 ;
        RECT 728.100 834.150 729.900 835.950 ;
        RECT 734.100 834.150 735.900 835.950 ;
        RECT 706.950 831.450 709.050 832.050 ;
        RECT 715.950 831.450 718.050 832.050 ;
        RECT 706.950 830.550 718.050 831.450 ;
        RECT 726.000 831.000 729.300 832.200 ;
        RECT 706.950 829.950 709.050 830.550 ;
        RECT 715.950 829.950 718.050 830.550 ;
        RECT 701.400 827.400 706.500 828.600 ;
        RECT 701.700 822.000 703.500 825.600 ;
        RECT 704.700 822.600 706.500 827.400 ;
        RECT 709.200 822.000 711.000 828.600 ;
        RECT 727.500 822.600 729.300 831.000 ;
        RECT 734.100 822.000 735.900 831.600 ;
        RECT 752.400 828.600 753.300 835.950 ;
        RECT 754.950 834.150 756.750 835.950 ;
        RECT 761.100 834.150 762.900 835.950 ;
        RECT 776.400 828.600 777.300 835.950 ;
        RECT 778.950 834.150 780.750 835.950 ;
        RECT 785.100 834.150 786.900 835.950 ;
        RECT 801.000 832.200 801.900 835.950 ;
        RECT 803.100 834.150 804.900 835.950 ;
        RECT 809.100 834.150 810.900 835.950 ;
        RECT 825.000 832.200 825.900 835.950 ;
        RECT 827.100 834.150 828.900 835.950 ;
        RECT 833.100 834.150 834.900 835.950 ;
        RECT 848.100 834.150 849.900 835.950 ;
        RECT 854.100 834.150 855.900 835.950 ;
        RECT 857.100 832.200 858.000 835.950 ;
        RECT 866.550 835.050 867.450 839.550 ;
        RECT 875.700 838.050 876.900 851.400 ;
        RECT 880.950 840.450 883.050 841.050 ;
        RECT 886.950 840.450 889.050 841.050 ;
        RECT 880.950 839.550 889.050 840.450 ;
        RECT 880.950 838.950 883.050 839.550 ;
        RECT 886.950 838.950 889.050 839.550 ;
        RECT 893.700 838.050 894.900 851.400 ;
        RECT 896.100 838.050 897.900 839.850 ;
        RECT 871.950 835.950 874.050 838.050 ;
        RECT 874.950 835.950 877.050 838.050 ;
        RECT 877.950 835.950 880.050 838.050 ;
        RECT 892.950 835.950 895.050 838.050 ;
        RECT 895.950 835.950 898.050 838.050 ;
        RECT 866.550 833.550 871.050 835.050 ;
        RECT 872.100 834.150 873.900 835.950 ;
        RECT 867.000 832.950 871.050 833.550 ;
        RECT 801.000 831.000 804.300 832.200 ;
        RECT 752.400 827.400 757.500 828.600 ;
        RECT 752.700 822.000 754.500 825.600 ;
        RECT 755.700 822.600 757.500 827.400 ;
        RECT 760.200 822.000 762.000 828.600 ;
        RECT 776.400 827.400 781.500 828.600 ;
        RECT 776.700 822.000 778.500 825.600 ;
        RECT 779.700 822.600 781.500 827.400 ;
        RECT 784.200 822.000 786.000 828.600 ;
        RECT 802.500 822.600 804.300 831.000 ;
        RECT 809.100 822.000 810.900 831.600 ;
        RECT 825.000 831.000 828.300 832.200 ;
        RECT 826.500 822.600 828.300 831.000 ;
        RECT 833.100 822.000 834.900 831.600 ;
        RECT 848.100 822.000 849.900 831.600 ;
        RECT 854.700 831.000 858.000 832.200 ;
        RECT 854.700 822.600 856.500 831.000 ;
        RECT 875.700 830.700 876.900 835.950 ;
        RECT 877.950 834.150 879.750 835.950 ;
        RECT 872.700 829.800 876.900 830.700 ;
        RECT 872.700 822.600 874.500 829.800 ;
        RECT 877.800 822.000 879.600 828.600 ;
        RECT 893.700 825.600 894.900 835.950 ;
        RECT 893.100 822.600 894.900 825.600 ;
        RECT 896.100 822.000 897.900 825.600 ;
        RECT 16.500 810.000 18.300 818.400 ;
        RECT 15.000 808.800 18.300 810.000 ;
        RECT 23.100 809.400 24.900 819.000 ;
        RECT 38.700 815.400 40.500 819.000 ;
        RECT 41.700 813.600 43.500 818.400 ;
        RECT 38.400 812.400 43.500 813.600 ;
        RECT 46.200 812.400 48.000 819.000 ;
        RECT 15.000 805.050 15.900 808.800 ;
        RECT 17.100 805.050 18.900 806.850 ;
        RECT 23.100 805.050 24.900 806.850 ;
        RECT 38.400 805.050 39.300 812.400 ;
        RECT 65.100 809.400 66.900 819.000 ;
        RECT 71.700 810.000 73.500 818.400 ;
        RECT 89.700 815.400 91.500 819.000 ;
        RECT 92.700 813.600 94.500 818.400 ;
        RECT 89.400 812.400 94.500 813.600 ;
        RECT 97.200 812.400 99.000 819.000 ;
        RECT 71.700 808.800 75.000 810.000 ;
        RECT 40.950 805.050 42.750 806.850 ;
        RECT 47.100 805.050 48.900 806.850 ;
        RECT 65.100 805.050 66.900 806.850 ;
        RECT 71.100 805.050 72.900 806.850 ;
        RECT 74.100 805.050 75.000 808.800 ;
        RECT 76.950 807.450 79.050 808.050 ;
        RECT 85.950 807.450 88.050 807.900 ;
        RECT 76.950 806.550 88.050 807.450 ;
        RECT 76.950 805.950 79.050 806.550 ;
        RECT 85.950 805.800 88.050 806.550 ;
        RECT 89.400 805.050 90.300 812.400 ;
        RECT 91.950 810.450 94.050 811.050 ;
        RECT 103.950 810.450 106.050 811.050 ;
        RECT 91.950 809.550 106.050 810.450 ;
        RECT 115.500 810.000 117.300 818.400 ;
        RECT 91.950 808.950 94.050 809.550 ;
        RECT 103.950 808.950 106.050 809.550 ;
        RECT 114.000 808.800 117.300 810.000 ;
        RECT 122.100 809.400 123.900 819.000 ;
        RECT 137.100 815.400 138.900 819.000 ;
        RECT 140.100 815.400 141.900 818.400 ;
        RECT 91.950 805.050 93.750 806.850 ;
        RECT 98.100 805.050 99.900 806.850 ;
        RECT 114.000 805.050 114.900 808.800 ;
        RECT 116.100 805.050 117.900 806.850 ;
        RECT 122.100 805.050 123.900 806.850 ;
        RECT 140.100 805.050 141.300 815.400 ;
        RECT 155.100 813.300 156.900 818.400 ;
        RECT 158.100 814.200 159.900 819.000 ;
        RECT 161.100 813.300 162.900 818.400 ;
        RECT 155.100 811.950 162.900 813.300 ;
        RECT 164.100 812.400 165.900 818.400 ;
        RECT 180.600 814.200 182.400 818.400 ;
        RECT 179.700 812.400 182.400 814.200 ;
        RECT 183.600 812.400 185.400 819.000 ;
        RECT 164.100 810.300 165.300 812.400 ;
        RECT 161.700 809.400 165.300 810.300 ;
        RECT 158.100 805.050 159.900 806.850 ;
        RECT 161.700 805.050 162.900 809.400 ;
        RECT 164.100 805.050 165.900 806.850 ;
        RECT 179.700 805.050 180.600 812.400 ;
        RECT 181.500 810.600 183.300 811.500 ;
        RECT 188.100 810.600 189.900 818.400 ;
        RECT 203.100 813.300 204.900 818.400 ;
        RECT 206.100 814.200 207.900 819.000 ;
        RECT 209.100 813.300 210.900 818.400 ;
        RECT 203.100 811.950 210.900 813.300 ;
        RECT 212.100 812.400 213.900 818.400 ;
        RECT 227.100 815.400 228.900 818.400 ;
        RECT 230.100 815.400 231.900 819.000 ;
        RECT 181.500 809.700 189.900 810.600 ;
        RECT 212.100 810.300 213.300 812.400 ;
        RECT 13.950 802.950 16.050 805.050 ;
        RECT 16.950 802.950 19.050 805.050 ;
        RECT 19.950 802.950 22.050 805.050 ;
        RECT 22.950 802.950 25.050 805.050 ;
        RECT 37.950 802.950 40.050 805.050 ;
        RECT 40.950 802.950 43.050 805.050 ;
        RECT 43.950 802.950 46.050 805.050 ;
        RECT 46.950 802.950 49.050 805.050 ;
        RECT 64.950 802.950 67.050 805.050 ;
        RECT 67.950 802.950 70.050 805.050 ;
        RECT 70.950 802.950 73.050 805.050 ;
        RECT 73.950 802.950 76.050 805.050 ;
        RECT 88.950 802.950 91.050 805.050 ;
        RECT 91.950 802.950 94.050 805.050 ;
        RECT 94.950 802.950 97.050 805.050 ;
        RECT 97.950 802.950 100.050 805.050 ;
        RECT 112.950 802.950 115.050 805.050 ;
        RECT 115.950 802.950 118.050 805.050 ;
        RECT 118.950 802.950 121.050 805.050 ;
        RECT 121.950 802.950 124.050 805.050 ;
        RECT 136.950 802.950 139.050 805.050 ;
        RECT 139.950 802.950 142.050 805.050 ;
        RECT 154.950 802.950 157.050 805.050 ;
        RECT 157.950 802.950 160.050 805.050 ;
        RECT 160.950 802.950 163.050 805.050 ;
        RECT 163.950 802.950 166.050 805.050 ;
        RECT 179.100 802.950 181.200 805.050 ;
        RECT 182.400 802.950 184.500 805.050 ;
        RECT 15.000 790.800 15.900 802.950 ;
        RECT 20.100 801.150 21.900 802.950 ;
        RECT 38.400 795.600 39.300 802.950 ;
        RECT 43.950 801.150 45.750 802.950 ;
        RECT 68.100 801.150 69.900 802.950 ;
        RECT 46.950 798.450 49.050 799.050 ;
        RECT 70.950 798.450 73.050 799.050 ;
        RECT 46.950 797.550 73.050 798.450 ;
        RECT 46.950 796.950 49.050 797.550 ;
        RECT 70.950 796.950 73.050 797.550 ;
        RECT 15.000 789.900 21.600 790.800 ;
        RECT 15.000 789.600 15.900 789.900 ;
        RECT 14.100 783.600 15.900 789.600 ;
        RECT 20.100 789.600 21.600 789.900 ;
        RECT 17.100 783.000 18.900 789.000 ;
        RECT 20.100 783.600 21.900 789.600 ;
        RECT 23.100 783.000 24.900 789.600 ;
        RECT 38.100 783.600 39.900 795.600 ;
        RECT 41.100 794.700 48.900 795.600 ;
        RECT 41.100 783.600 42.900 794.700 ;
        RECT 44.100 783.000 45.900 793.800 ;
        RECT 47.100 783.600 48.900 794.700 ;
        RECT 74.100 790.800 75.000 802.950 ;
        RECT 89.400 795.600 90.300 802.950 ;
        RECT 94.950 801.150 96.750 802.950 ;
        RECT 68.400 789.900 75.000 790.800 ;
        RECT 68.400 789.600 69.900 789.900 ;
        RECT 65.100 783.000 66.900 789.600 ;
        RECT 68.100 783.600 69.900 789.600 ;
        RECT 74.100 789.600 75.000 789.900 ;
        RECT 71.100 783.000 72.900 789.000 ;
        RECT 74.100 783.600 75.900 789.600 ;
        RECT 89.100 783.600 90.900 795.600 ;
        RECT 92.100 794.700 99.900 795.600 ;
        RECT 92.100 783.600 93.900 794.700 ;
        RECT 95.100 783.000 96.900 793.800 ;
        RECT 98.100 783.600 99.900 794.700 ;
        RECT 114.000 790.800 114.900 802.950 ;
        RECT 119.100 801.150 120.900 802.950 ;
        RECT 137.100 801.150 138.900 802.950 ;
        RECT 114.000 789.900 120.600 790.800 ;
        RECT 114.000 789.600 114.900 789.900 ;
        RECT 113.100 783.600 114.900 789.600 ;
        RECT 119.100 789.600 120.600 789.900 ;
        RECT 140.100 789.600 141.300 802.950 ;
        RECT 155.100 801.150 156.900 802.950 ;
        RECT 161.700 795.600 162.900 802.950 ;
        RECT 179.700 795.600 180.600 802.950 ;
        RECT 183.000 801.150 184.800 802.950 ;
        RECT 116.100 783.000 117.900 789.000 ;
        RECT 119.100 783.600 120.900 789.600 ;
        RECT 122.100 783.000 123.900 789.600 ;
        RECT 137.100 783.000 138.900 789.600 ;
        RECT 140.100 783.600 141.900 789.600 ;
        RECT 155.400 783.000 157.200 795.600 ;
        RECT 160.500 794.100 162.900 795.600 ;
        RECT 160.500 783.600 162.300 794.100 ;
        RECT 163.200 791.100 165.000 792.900 ;
        RECT 163.500 783.000 165.300 789.600 ;
        RECT 179.100 783.600 180.900 795.600 ;
        RECT 182.100 783.000 183.900 795.000 ;
        RECT 186.000 789.600 186.900 809.700 ;
        RECT 209.700 809.400 213.300 810.300 ;
        RECT 187.950 805.050 189.750 806.850 ;
        RECT 206.100 805.050 207.900 806.850 ;
        RECT 209.700 805.050 210.900 809.400 ;
        RECT 212.100 805.050 213.900 806.850 ;
        RECT 227.700 805.050 228.900 815.400 ;
        RECT 247.500 810.000 249.300 818.400 ;
        RECT 246.000 808.800 249.300 810.000 ;
        RECT 254.100 809.400 255.900 819.000 ;
        RECT 272.700 815.400 274.500 819.000 ;
        RECT 275.700 813.600 277.500 818.400 ;
        RECT 272.400 812.400 277.500 813.600 ;
        RECT 280.200 812.400 282.000 819.000 ;
        RECT 296.100 812.400 297.900 818.400 ;
        RECT 246.000 805.050 246.900 808.800 ;
        RECT 248.100 805.050 249.900 806.850 ;
        RECT 254.100 805.050 255.900 806.850 ;
        RECT 272.400 805.050 273.300 812.400 ;
        RECT 296.700 810.300 297.900 812.400 ;
        RECT 299.100 813.300 300.900 818.400 ;
        RECT 302.100 814.200 303.900 819.000 ;
        RECT 305.100 813.300 306.900 818.400 ;
        RECT 320.100 815.400 321.900 819.000 ;
        RECT 323.100 815.400 324.900 818.400 ;
        RECT 299.100 811.950 306.900 813.300 ;
        RECT 296.700 809.400 300.300 810.300 ;
        RECT 274.950 805.050 276.750 806.850 ;
        RECT 281.100 805.050 282.900 806.850 ;
        RECT 296.100 805.050 297.900 806.850 ;
        RECT 299.100 805.050 300.300 809.400 ;
        RECT 302.100 805.050 303.900 806.850 ;
        RECT 323.100 805.050 324.300 815.400 ;
        RECT 338.100 812.400 339.900 818.400 ;
        RECT 341.100 813.300 342.900 819.000 ;
        RECT 345.600 812.400 347.400 818.400 ;
        RECT 350.100 813.300 351.900 819.000 ;
        RECT 353.100 812.400 354.900 818.400 ;
        RECT 368.400 812.400 370.200 819.000 ;
        RECT 338.700 810.600 339.900 812.400 ;
        RECT 345.900 810.900 347.100 812.400 ;
        RECT 350.100 811.500 354.900 812.400 ;
        RECT 338.700 809.700 345.000 810.600 ;
        RECT 342.900 807.600 345.000 809.700 ;
        RECT 338.400 805.050 340.200 806.850 ;
        RECT 343.200 805.800 345.000 807.600 ;
        RECT 345.900 808.800 348.900 810.900 ;
        RECT 350.100 810.300 352.200 811.500 ;
        RECT 373.500 811.200 375.300 818.400 ;
        RECT 371.100 810.300 375.300 811.200 ;
        RECT 389.700 811.200 391.500 818.400 ;
        RECT 394.800 812.400 396.600 819.000 ;
        RECT 410.100 813.300 411.900 818.400 ;
        RECT 413.100 814.200 414.900 819.000 ;
        RECT 416.100 813.300 417.900 818.400 ;
        RECT 410.100 811.950 417.900 813.300 ;
        RECT 419.100 812.400 420.900 818.400 ;
        RECT 434.400 812.400 436.200 819.000 ;
        RECT 389.700 810.300 393.900 811.200 ;
        RECT 419.100 810.300 420.300 812.400 ;
        RECT 439.500 811.200 441.300 818.400 ;
        RECT 455.100 815.400 456.900 819.000 ;
        RECT 458.100 815.400 459.900 818.400 ;
        RECT 187.800 802.950 189.900 805.050 ;
        RECT 202.950 802.950 205.050 805.050 ;
        RECT 205.950 802.950 208.050 805.050 ;
        RECT 208.950 802.950 211.050 805.050 ;
        RECT 211.950 802.950 214.050 805.050 ;
        RECT 226.950 802.950 229.050 805.050 ;
        RECT 229.950 802.950 232.050 805.050 ;
        RECT 244.950 802.950 247.050 805.050 ;
        RECT 247.950 802.950 250.050 805.050 ;
        RECT 250.950 802.950 253.050 805.050 ;
        RECT 253.950 802.950 256.050 805.050 ;
        RECT 271.950 802.950 274.050 805.050 ;
        RECT 274.950 802.950 277.050 805.050 ;
        RECT 277.950 802.950 280.050 805.050 ;
        RECT 280.950 802.950 283.050 805.050 ;
        RECT 295.950 802.950 298.050 805.050 ;
        RECT 298.950 802.950 301.050 805.050 ;
        RECT 301.950 802.950 304.050 805.050 ;
        RECT 304.950 802.950 307.050 805.050 ;
        RECT 319.950 802.950 322.050 805.050 ;
        RECT 322.950 802.950 325.050 805.050 ;
        RECT 338.100 804.300 340.200 805.050 ;
        RECT 338.100 802.950 345.000 804.300 ;
        RECT 203.100 801.150 204.900 802.950 ;
        RECT 209.700 795.600 210.900 802.950 ;
        RECT 185.100 783.600 186.900 789.600 ;
        RECT 188.100 783.000 189.900 789.600 ;
        RECT 203.400 783.000 205.200 795.600 ;
        RECT 208.500 794.100 210.900 795.600 ;
        RECT 208.500 783.600 210.300 794.100 ;
        RECT 211.200 791.100 213.000 792.900 ;
        RECT 227.700 789.600 228.900 802.950 ;
        RECT 230.100 801.150 231.900 802.950 ;
        RECT 246.000 790.800 246.900 802.950 ;
        RECT 251.100 801.150 252.900 802.950 ;
        RECT 272.400 795.600 273.300 802.950 ;
        RECT 277.950 801.150 279.750 802.950 ;
        RECT 286.950 801.450 289.050 802.050 ;
        RECT 292.950 801.450 295.050 802.050 ;
        RECT 286.950 800.550 295.050 801.450 ;
        RECT 286.950 799.950 289.050 800.550 ;
        RECT 292.950 799.950 295.050 800.550 ;
        RECT 299.100 795.600 300.300 802.950 ;
        RECT 305.100 801.150 306.900 802.950 ;
        RECT 320.100 801.150 321.900 802.950 ;
        RECT 246.000 789.900 252.600 790.800 ;
        RECT 246.000 789.600 246.900 789.900 ;
        RECT 211.500 783.000 213.300 789.600 ;
        RECT 227.100 783.600 228.900 789.600 ;
        RECT 230.100 783.000 231.900 789.600 ;
        RECT 245.100 783.600 246.900 789.600 ;
        RECT 251.100 789.600 252.600 789.900 ;
        RECT 248.100 783.000 249.900 789.000 ;
        RECT 251.100 783.600 252.900 789.600 ;
        RECT 254.100 783.000 255.900 789.600 ;
        RECT 272.100 783.600 273.900 795.600 ;
        RECT 275.100 794.700 282.900 795.600 ;
        RECT 275.100 783.600 276.900 794.700 ;
        RECT 278.100 783.000 279.900 793.800 ;
        RECT 281.100 783.600 282.900 794.700 ;
        RECT 299.100 794.100 301.500 795.600 ;
        RECT 297.000 791.100 298.800 792.900 ;
        RECT 296.700 783.000 298.500 789.600 ;
        RECT 299.700 783.600 301.500 794.100 ;
        RECT 304.800 783.000 306.600 795.600 ;
        RECT 323.100 789.600 324.300 802.950 ;
        RECT 343.200 802.500 345.000 802.950 ;
        RECT 345.900 803.100 347.100 808.800 ;
        RECT 348.000 805.800 350.100 807.900 ;
        RECT 348.300 804.000 350.100 805.800 ;
        RECT 368.250 805.050 370.050 806.850 ;
        RECT 371.100 805.050 372.300 810.300 ;
        RECT 374.100 805.050 375.900 806.850 ;
        RECT 389.100 805.050 390.900 806.850 ;
        RECT 392.700 805.050 393.900 810.300 ;
        RECT 416.700 809.400 420.300 810.300 ;
        RECT 437.100 810.300 441.300 811.200 ;
        RECT 394.950 805.050 396.750 806.850 ;
        RECT 413.100 805.050 414.900 806.850 ;
        RECT 416.700 805.050 417.900 809.400 ;
        RECT 419.100 805.050 420.900 806.850 ;
        RECT 434.250 805.050 436.050 806.850 ;
        RECT 437.100 805.050 438.300 810.300 ;
        RECT 440.100 805.050 441.900 806.850 ;
        RECT 458.100 805.050 459.300 815.400 ;
        RECT 476.100 812.400 477.900 818.400 ;
        RECT 479.100 812.400 480.900 819.000 ;
        RECT 482.100 815.400 483.900 818.400 ;
        RECT 476.100 805.050 477.300 812.400 ;
        RECT 482.700 811.500 483.900 815.400 ;
        RECT 497.100 812.400 498.900 818.400 ;
        RECT 478.200 810.600 483.900 811.500 ;
        RECT 478.200 809.700 480.000 810.600 ;
        RECT 345.900 802.200 348.300 803.100 ;
        RECT 346.800 802.050 348.300 802.200 ;
        RECT 352.800 802.950 354.900 805.050 ;
        RECT 367.950 802.950 370.050 805.050 ;
        RECT 370.950 802.950 373.050 805.050 ;
        RECT 373.950 802.950 376.050 805.050 ;
        RECT 388.950 802.950 391.050 805.050 ;
        RECT 391.950 802.950 394.050 805.050 ;
        RECT 394.950 802.950 397.050 805.050 ;
        RECT 409.950 802.950 412.050 805.050 ;
        RECT 412.950 802.950 415.050 805.050 ;
        RECT 415.950 802.950 418.050 805.050 ;
        RECT 418.950 802.950 421.050 805.050 ;
        RECT 433.950 802.950 436.050 805.050 ;
        RECT 436.950 802.950 439.050 805.050 ;
        RECT 439.950 802.950 442.050 805.050 ;
        RECT 454.950 802.950 457.050 805.050 ;
        RECT 457.950 802.950 460.050 805.050 ;
        RECT 476.100 802.950 478.200 805.050 ;
        RECT 342.000 799.500 345.900 801.300 ;
        RECT 343.800 799.200 345.900 799.500 ;
        RECT 346.800 799.950 348.900 802.050 ;
        RECT 352.800 801.150 354.600 802.950 ;
        RECT 346.800 798.000 347.700 799.950 ;
        RECT 340.500 795.600 342.600 797.700 ;
        RECT 346.200 796.950 347.700 798.000 ;
        RECT 346.200 795.600 347.400 796.950 ;
        RECT 338.100 794.700 342.600 795.600 ;
        RECT 320.100 783.000 321.900 789.600 ;
        RECT 323.100 783.600 324.900 789.600 ;
        RECT 338.100 783.600 339.900 794.700 ;
        RECT 341.100 783.000 342.900 793.500 ;
        RECT 345.600 783.600 347.400 795.600 ;
        RECT 350.100 795.600 352.200 796.500 ;
        RECT 350.100 794.400 354.900 795.600 ;
        RECT 350.100 783.000 351.900 793.500 ;
        RECT 353.100 783.600 354.900 794.400 ;
        RECT 371.100 789.600 372.300 802.950 ;
        RECT 392.700 789.600 393.900 802.950 ;
        RECT 410.100 801.150 411.900 802.950 ;
        RECT 416.700 795.600 417.900 802.950 ;
        RECT 368.100 783.000 369.900 789.600 ;
        RECT 371.100 783.600 372.900 789.600 ;
        RECT 374.100 783.000 375.900 789.600 ;
        RECT 389.100 783.000 390.900 789.600 ;
        RECT 392.100 783.600 393.900 789.600 ;
        RECT 395.100 783.000 396.900 789.600 ;
        RECT 410.400 783.000 412.200 795.600 ;
        RECT 415.500 794.100 417.900 795.600 ;
        RECT 415.500 783.600 417.300 794.100 ;
        RECT 418.200 791.100 420.000 792.900 ;
        RECT 437.100 789.600 438.300 802.950 ;
        RECT 455.100 801.150 456.900 802.950 ;
        RECT 439.950 798.450 442.050 799.050 ;
        RECT 454.950 798.450 457.050 799.050 ;
        RECT 439.950 797.550 457.050 798.450 ;
        RECT 439.950 796.950 442.050 797.550 ;
        RECT 454.950 796.950 457.050 797.550 ;
        RECT 458.100 789.600 459.300 802.950 ;
        RECT 476.100 795.600 477.300 802.950 ;
        RECT 479.100 798.300 480.000 809.700 ;
        RECT 497.700 810.300 498.900 812.400 ;
        RECT 500.100 813.300 501.900 818.400 ;
        RECT 503.100 814.200 504.900 819.000 ;
        RECT 506.100 813.300 507.900 818.400 ;
        RECT 500.100 811.950 507.900 813.300 ;
        RECT 521.100 813.300 522.900 818.400 ;
        RECT 524.100 814.200 525.900 819.000 ;
        RECT 527.100 813.300 528.900 818.400 ;
        RECT 521.100 811.950 528.900 813.300 ;
        RECT 530.100 812.400 531.900 818.400 ;
        RECT 545.400 812.400 547.200 819.000 ;
        RECT 530.100 810.300 531.300 812.400 ;
        RECT 550.500 811.200 552.300 818.400 ;
        RECT 566.700 812.400 568.500 819.000 ;
        RECT 571.200 812.400 573.000 818.400 ;
        RECT 575.700 812.400 577.500 819.000 ;
        RECT 593.100 813.300 594.900 818.400 ;
        RECT 596.100 814.200 597.900 819.000 ;
        RECT 599.100 813.300 600.900 818.400 ;
        RECT 497.700 809.400 501.300 810.300 ;
        RECT 497.100 805.050 498.900 806.850 ;
        RECT 500.100 805.050 501.300 809.400 ;
        RECT 527.700 809.400 531.300 810.300 ;
        RECT 548.100 810.300 552.300 811.200 ;
        RECT 503.100 805.050 504.900 806.850 ;
        RECT 524.100 805.050 525.900 806.850 ;
        RECT 527.700 805.050 528.900 809.400 ;
        RECT 530.100 805.050 531.900 806.850 ;
        RECT 545.250 805.050 547.050 806.850 ;
        RECT 548.100 805.050 549.300 810.300 ;
        RECT 551.100 805.050 552.900 806.850 ;
        RECT 566.250 805.050 568.050 806.850 ;
        RECT 572.100 805.050 573.300 812.400 ;
        RECT 593.100 811.950 600.900 813.300 ;
        RECT 602.100 812.400 603.900 818.400 ;
        RECT 620.100 815.400 621.900 819.000 ;
        RECT 623.100 815.400 624.900 818.400 ;
        RECT 638.700 815.400 640.500 819.000 ;
        RECT 602.100 810.300 603.300 812.400 ;
        RECT 599.700 809.400 603.300 810.300 ;
        RECT 578.100 805.050 579.900 806.850 ;
        RECT 596.100 805.050 597.900 806.850 ;
        RECT 599.700 805.050 600.900 809.400 ;
        RECT 602.100 805.050 603.900 806.850 ;
        RECT 623.100 805.050 624.300 815.400 ;
        RECT 641.700 813.600 643.500 818.400 ;
        RECT 638.400 812.400 643.500 813.600 ;
        RECT 646.200 812.400 648.000 819.000 ;
        RECT 638.400 805.050 639.300 812.400 ;
        RECT 662.100 809.400 663.900 819.000 ;
        RECT 668.700 810.000 670.500 818.400 ;
        RECT 686.700 811.200 688.500 818.400 ;
        RECT 691.800 812.400 693.600 819.000 ;
        RECT 686.700 810.300 690.900 811.200 ;
        RECT 668.700 808.800 672.000 810.000 ;
        RECT 640.950 805.050 642.750 806.850 ;
        RECT 647.100 805.050 648.900 806.850 ;
        RECT 662.100 805.050 663.900 806.850 ;
        RECT 668.100 805.050 669.900 806.850 ;
        RECT 671.100 805.050 672.000 808.800 ;
        RECT 686.100 805.050 687.900 806.850 ;
        RECT 689.700 805.050 690.900 810.300 ;
        RECT 709.500 810.000 711.300 818.400 ;
        RECT 708.000 808.800 711.300 810.000 ;
        RECT 716.100 809.400 717.900 819.000 ;
        RECT 731.100 815.400 732.900 818.400 ;
        RECT 734.100 815.400 735.900 819.000 ;
        RECT 691.950 805.050 693.750 806.850 ;
        RECT 708.000 805.050 708.900 808.800 ;
        RECT 710.100 805.050 711.900 806.850 ;
        RECT 716.100 805.050 717.900 806.850 ;
        RECT 731.700 805.050 732.900 815.400 ;
        RECT 749.100 813.300 750.900 818.400 ;
        RECT 752.100 814.200 753.900 819.000 ;
        RECT 755.100 813.300 756.900 818.400 ;
        RECT 749.100 811.950 756.900 813.300 ;
        RECT 758.100 812.400 759.900 818.400 ;
        RECT 773.400 812.400 775.200 819.000 ;
        RECT 758.100 810.300 759.300 812.400 ;
        RECT 778.500 811.200 780.300 818.400 ;
        RECT 794.700 815.400 796.500 819.000 ;
        RECT 797.700 813.600 799.500 818.400 ;
        RECT 755.700 809.400 759.300 810.300 ;
        RECT 776.100 810.300 780.300 811.200 ;
        RECT 794.400 812.400 799.500 813.600 ;
        RECT 802.200 812.400 804.000 819.000 ;
        RECT 752.100 805.050 753.900 806.850 ;
        RECT 755.700 805.050 756.900 809.400 ;
        RECT 758.100 805.050 759.900 806.850 ;
        RECT 773.250 805.050 775.050 806.850 ;
        RECT 776.100 805.050 777.300 810.300 ;
        RECT 779.100 805.050 780.900 806.850 ;
        RECT 794.400 805.050 795.300 812.400 ;
        RECT 796.950 810.450 799.050 811.050 ;
        RECT 811.950 810.450 814.050 811.050 ;
        RECT 796.950 809.550 814.050 810.450 ;
        RECT 796.950 808.950 799.050 809.550 ;
        RECT 811.950 808.950 814.050 809.550 ;
        RECT 818.100 809.400 819.900 819.000 ;
        RECT 824.700 810.000 826.500 818.400 ;
        RECT 846.000 812.400 847.800 819.000 ;
        RECT 850.500 813.600 852.300 818.400 ;
        RECT 853.500 815.400 855.300 819.000 ;
        RECT 850.500 812.400 855.600 813.600 ;
        RECT 824.700 808.800 828.000 810.000 ;
        RECT 796.950 805.050 798.750 806.850 ;
        RECT 803.100 805.050 804.900 806.850 ;
        RECT 818.100 805.050 819.900 806.850 ;
        RECT 824.100 805.050 825.900 806.850 ;
        RECT 827.100 805.050 828.000 808.800 ;
        RECT 845.100 805.050 846.900 806.850 ;
        RECT 851.250 805.050 853.050 806.850 ;
        RECT 854.700 805.050 855.600 812.400 ;
        RECT 869.100 813.300 870.900 818.400 ;
        RECT 872.100 814.200 873.900 819.000 ;
        RECT 875.100 813.300 876.900 818.400 ;
        RECT 869.100 811.950 876.900 813.300 ;
        RECT 878.100 812.400 879.900 818.400 ;
        RECT 878.100 810.300 879.300 812.400 ;
        RECT 875.700 809.400 879.300 810.300 ;
        RECT 856.950 807.450 861.000 808.050 ;
        RECT 856.950 805.950 861.450 807.450 ;
        RECT 481.500 802.950 483.600 805.050 ;
        RECT 496.950 802.950 499.050 805.050 ;
        RECT 499.950 802.950 502.050 805.050 ;
        RECT 502.950 802.950 505.050 805.050 ;
        RECT 505.950 802.950 508.050 805.050 ;
        RECT 520.950 802.950 523.050 805.050 ;
        RECT 523.950 802.950 526.050 805.050 ;
        RECT 526.950 802.950 529.050 805.050 ;
        RECT 529.950 802.950 532.050 805.050 ;
        RECT 544.950 802.950 547.050 805.050 ;
        RECT 547.950 802.950 550.050 805.050 ;
        RECT 550.950 802.950 553.050 805.050 ;
        RECT 565.950 802.950 568.050 805.050 ;
        RECT 568.950 802.950 571.050 805.050 ;
        RECT 571.950 802.950 574.050 805.050 ;
        RECT 574.950 802.950 577.050 805.050 ;
        RECT 577.950 802.950 580.050 805.050 ;
        RECT 592.950 802.950 595.050 805.050 ;
        RECT 595.950 802.950 598.050 805.050 ;
        RECT 598.950 802.950 601.050 805.050 ;
        RECT 601.950 802.950 604.050 805.050 ;
        RECT 619.950 802.950 622.050 805.050 ;
        RECT 622.950 802.950 625.050 805.050 ;
        RECT 637.950 802.950 640.050 805.050 ;
        RECT 640.950 802.950 643.050 805.050 ;
        RECT 643.950 802.950 646.050 805.050 ;
        RECT 646.950 802.950 649.050 805.050 ;
        RECT 661.950 802.950 664.050 805.050 ;
        RECT 664.950 802.950 667.050 805.050 ;
        RECT 667.950 802.950 670.050 805.050 ;
        RECT 670.950 802.950 673.050 805.050 ;
        RECT 685.950 802.950 688.050 805.050 ;
        RECT 688.950 802.950 691.050 805.050 ;
        RECT 691.950 802.950 694.050 805.050 ;
        RECT 706.950 802.950 709.050 805.050 ;
        RECT 709.950 802.950 712.050 805.050 ;
        RECT 712.950 802.950 715.050 805.050 ;
        RECT 715.950 802.950 718.050 805.050 ;
        RECT 730.950 802.950 733.050 805.050 ;
        RECT 733.950 802.950 736.050 805.050 ;
        RECT 748.950 802.950 751.050 805.050 ;
        RECT 751.950 802.950 754.050 805.050 ;
        RECT 754.950 802.950 757.050 805.050 ;
        RECT 757.950 802.950 760.050 805.050 ;
        RECT 772.950 802.950 775.050 805.050 ;
        RECT 775.950 802.950 778.050 805.050 ;
        RECT 778.950 802.950 781.050 805.050 ;
        RECT 793.950 802.950 796.050 805.050 ;
        RECT 796.950 802.950 799.050 805.050 ;
        RECT 799.950 802.950 802.050 805.050 ;
        RECT 802.950 802.950 805.050 805.050 ;
        RECT 817.950 802.950 820.050 805.050 ;
        RECT 820.950 802.950 823.050 805.050 ;
        RECT 823.950 802.950 826.050 805.050 ;
        RECT 826.950 802.950 829.050 805.050 ;
        RECT 844.950 802.950 847.050 805.050 ;
        RECT 847.950 802.950 850.050 805.050 ;
        RECT 850.950 802.950 853.050 805.050 ;
        RECT 853.950 802.950 856.050 805.050 ;
        RECT 481.800 801.150 483.600 802.950 ;
        RECT 478.200 797.400 480.000 798.300 ;
        RECT 478.200 796.500 483.900 797.400 ;
        RECT 418.500 783.000 420.300 789.600 ;
        RECT 434.100 783.000 435.900 789.600 ;
        RECT 437.100 783.600 438.900 789.600 ;
        RECT 440.100 783.000 441.900 789.600 ;
        RECT 455.100 783.000 456.900 789.600 ;
        RECT 458.100 783.600 459.900 789.600 ;
        RECT 476.100 783.600 477.900 795.600 ;
        RECT 479.100 783.000 480.900 793.800 ;
        RECT 482.700 789.600 483.900 796.500 ;
        RECT 500.100 795.600 501.300 802.950 ;
        RECT 506.100 801.150 507.900 802.950 ;
        RECT 521.100 801.150 522.900 802.950 ;
        RECT 502.950 798.450 505.050 799.050 ;
        RECT 514.950 798.450 517.050 799.050 ;
        RECT 502.950 797.550 517.050 798.450 ;
        RECT 502.950 796.950 505.050 797.550 ;
        RECT 514.950 796.950 517.050 797.550 ;
        RECT 527.700 795.600 528.900 802.950 ;
        RECT 500.100 794.100 502.500 795.600 ;
        RECT 498.000 791.100 499.800 792.900 ;
        RECT 482.100 783.600 483.900 789.600 ;
        RECT 497.700 783.000 499.500 789.600 ;
        RECT 500.700 783.600 502.500 794.100 ;
        RECT 505.800 783.000 507.600 795.600 ;
        RECT 521.400 783.000 523.200 795.600 ;
        RECT 526.500 794.100 528.900 795.600 ;
        RECT 526.500 783.600 528.300 794.100 ;
        RECT 529.200 791.100 531.000 792.900 ;
        RECT 548.100 789.600 549.300 802.950 ;
        RECT 569.250 801.150 571.050 802.950 ;
        RECT 572.100 797.400 573.000 802.950 ;
        RECT 575.100 801.150 576.900 802.950 ;
        RECT 593.100 801.150 594.900 802.950 ;
        RECT 572.100 796.500 576.900 797.400 ;
        RECT 566.100 794.400 573.900 795.300 ;
        RECT 529.500 783.000 531.300 789.600 ;
        RECT 545.100 783.000 546.900 789.600 ;
        RECT 548.100 783.600 549.900 789.600 ;
        RECT 551.100 783.000 552.900 789.600 ;
        RECT 566.100 783.600 567.900 794.400 ;
        RECT 569.100 783.000 570.900 793.500 ;
        RECT 572.100 784.500 573.900 794.400 ;
        RECT 575.100 785.400 576.900 796.500 ;
        RECT 599.700 795.600 600.900 802.950 ;
        RECT 620.100 801.150 621.900 802.950 ;
        RECT 578.100 784.500 579.900 795.600 ;
        RECT 572.100 783.600 579.900 784.500 ;
        RECT 593.400 783.000 595.200 795.600 ;
        RECT 598.500 794.100 600.900 795.600 ;
        RECT 598.500 783.600 600.300 794.100 ;
        RECT 601.200 791.100 603.000 792.900 ;
        RECT 623.100 789.600 624.300 802.950 ;
        RECT 638.400 795.600 639.300 802.950 ;
        RECT 643.950 801.150 645.750 802.950 ;
        RECT 665.100 801.150 666.900 802.950 ;
        RECT 655.950 798.450 658.050 799.050 ;
        RECT 667.950 798.450 670.050 799.050 ;
        RECT 655.950 797.550 670.050 798.450 ;
        RECT 655.950 796.950 658.050 797.550 ;
        RECT 667.950 796.950 670.050 797.550 ;
        RECT 601.500 783.000 603.300 789.600 ;
        RECT 620.100 783.000 621.900 789.600 ;
        RECT 623.100 783.600 624.900 789.600 ;
        RECT 638.100 783.600 639.900 795.600 ;
        RECT 641.100 794.700 648.900 795.600 ;
        RECT 641.100 783.600 642.900 794.700 ;
        RECT 644.100 783.000 645.900 793.800 ;
        RECT 647.100 783.600 648.900 794.700 ;
        RECT 671.100 790.800 672.000 802.950 ;
        RECT 665.400 789.900 672.000 790.800 ;
        RECT 665.400 789.600 666.900 789.900 ;
        RECT 662.100 783.000 663.900 789.600 ;
        RECT 665.100 783.600 666.900 789.600 ;
        RECT 671.100 789.600 672.000 789.900 ;
        RECT 689.700 789.600 690.900 802.950 ;
        RECT 708.000 790.800 708.900 802.950 ;
        RECT 713.100 801.150 714.900 802.950 ;
        RECT 708.000 789.900 714.600 790.800 ;
        RECT 708.000 789.600 708.900 789.900 ;
        RECT 668.100 783.000 669.900 789.000 ;
        RECT 671.100 783.600 672.900 789.600 ;
        RECT 686.100 783.000 687.900 789.600 ;
        RECT 689.100 783.600 690.900 789.600 ;
        RECT 692.100 783.000 693.900 789.600 ;
        RECT 707.100 783.600 708.900 789.600 ;
        RECT 713.100 789.600 714.600 789.900 ;
        RECT 731.700 789.600 732.900 802.950 ;
        RECT 734.100 801.150 735.900 802.950 ;
        RECT 749.100 801.150 750.900 802.950 ;
        RECT 755.700 795.600 756.900 802.950 ;
        RECT 710.100 783.000 711.900 789.000 ;
        RECT 713.100 783.600 714.900 789.600 ;
        RECT 716.100 783.000 717.900 789.600 ;
        RECT 731.100 783.600 732.900 789.600 ;
        RECT 734.100 783.000 735.900 789.600 ;
        RECT 749.400 783.000 751.200 795.600 ;
        RECT 754.500 794.100 756.900 795.600 ;
        RECT 754.500 783.600 756.300 794.100 ;
        RECT 757.200 791.100 759.000 792.900 ;
        RECT 776.100 789.600 777.300 802.950 ;
        RECT 794.400 795.600 795.300 802.950 ;
        RECT 799.950 801.150 801.750 802.950 ;
        RECT 821.100 801.150 822.900 802.950 ;
        RECT 808.950 798.450 811.050 799.050 ;
        RECT 823.950 798.450 826.050 799.050 ;
        RECT 808.950 797.550 826.050 798.450 ;
        RECT 808.950 796.950 811.050 797.550 ;
        RECT 823.950 796.950 826.050 797.550 ;
        RECT 757.500 783.000 759.300 789.600 ;
        RECT 773.100 783.000 774.900 789.600 ;
        RECT 776.100 783.600 777.900 789.600 ;
        RECT 779.100 783.000 780.900 789.600 ;
        RECT 794.100 783.600 795.900 795.600 ;
        RECT 797.100 794.700 804.900 795.600 ;
        RECT 797.100 783.600 798.900 794.700 ;
        RECT 800.100 783.000 801.900 793.800 ;
        RECT 803.100 783.600 804.900 794.700 ;
        RECT 827.100 790.800 828.000 802.950 ;
        RECT 832.950 801.450 835.050 802.050 ;
        RECT 841.950 801.450 844.050 802.050 ;
        RECT 832.950 800.550 844.050 801.450 ;
        RECT 848.250 801.150 850.050 802.950 ;
        RECT 832.950 799.950 835.050 800.550 ;
        RECT 841.950 799.950 844.050 800.550 ;
        RECT 854.700 795.600 855.600 802.950 ;
        RECT 860.550 801.450 861.450 805.950 ;
        RECT 872.100 805.050 873.900 806.850 ;
        RECT 875.700 805.050 876.900 809.400 ;
        RECT 878.100 805.050 879.900 806.850 ;
        RECT 868.950 802.950 871.050 805.050 ;
        RECT 871.950 802.950 874.050 805.050 ;
        RECT 874.950 802.950 877.050 805.050 ;
        RECT 877.950 802.950 880.050 805.050 ;
        RECT 865.950 801.450 868.050 802.050 ;
        RECT 860.550 800.550 868.050 801.450 ;
        RECT 869.100 801.150 870.900 802.950 ;
        RECT 865.950 799.950 868.050 800.550 ;
        RECT 875.700 795.600 876.900 802.950 ;
        RECT 821.400 789.900 828.000 790.800 ;
        RECT 821.400 789.600 822.900 789.900 ;
        RECT 818.100 783.000 819.900 789.600 ;
        RECT 821.100 783.600 822.900 789.600 ;
        RECT 827.100 789.600 828.000 789.900 ;
        RECT 845.100 794.700 852.900 795.600 ;
        RECT 824.100 783.000 825.900 789.000 ;
        RECT 827.100 783.600 828.900 789.600 ;
        RECT 845.100 783.600 846.900 794.700 ;
        RECT 848.100 783.000 849.900 793.800 ;
        RECT 851.100 783.600 852.900 794.700 ;
        RECT 854.100 783.600 855.900 795.600 ;
        RECT 869.400 783.000 871.200 795.600 ;
        RECT 874.500 794.100 876.900 795.600 ;
        RECT 874.500 783.600 876.300 794.100 ;
        RECT 877.200 791.100 879.000 792.900 ;
        RECT 877.500 783.000 879.300 789.600 ;
        RECT 14.100 773.400 15.900 779.400 ;
        RECT 17.100 773.400 18.900 780.000 ;
        RECT 35.700 773.400 37.500 780.000 ;
        RECT 14.700 760.050 15.900 773.400 ;
        RECT 36.000 770.100 37.800 771.900 ;
        RECT 38.700 768.900 40.500 779.400 ;
        RECT 38.100 767.400 40.500 768.900 ;
        RECT 43.800 767.400 45.600 780.000 ;
        RECT 59.100 769.500 60.900 779.400 ;
        RECT 62.100 770.400 63.900 780.000 ;
        RECT 65.100 778.500 72.900 779.400 ;
        RECT 65.100 769.500 66.900 778.500 ;
        RECT 59.100 768.600 66.900 769.500 ;
        RECT 68.100 769.800 69.900 777.600 ;
        RECT 71.100 770.700 72.900 778.500 ;
        RECT 74.100 778.500 81.900 779.400 ;
        RECT 74.100 769.800 75.900 778.500 ;
        RECT 68.100 768.900 75.900 769.800 ;
        RECT 77.100 769.800 78.900 777.600 ;
        RECT 17.100 760.050 18.900 761.850 ;
        RECT 38.100 760.050 39.300 767.400 ;
        RECT 44.100 760.050 45.900 761.850 ;
        RECT 62.100 760.050 63.900 761.850 ;
        RECT 71.250 760.050 73.050 761.850 ;
        RECT 77.100 760.050 78.300 769.800 ;
        RECT 80.100 769.200 81.900 778.500 ;
        RECT 95.400 767.400 97.200 780.000 ;
        RECT 100.500 768.900 102.300 779.400 ;
        RECT 103.500 773.400 105.300 780.000 ;
        RECT 103.200 770.100 105.000 771.900 ;
        RECT 100.500 767.400 102.900 768.900 ;
        RECT 119.100 767.400 120.900 780.000 ;
        RECT 124.200 768.600 126.000 779.400 ;
        RECT 140.100 773.400 141.900 779.400 ;
        RECT 143.100 773.400 144.900 780.000 ;
        RECT 158.100 773.400 159.900 779.400 ;
        RECT 161.100 774.000 162.900 780.000 ;
        RECT 122.400 767.400 126.000 768.600 ;
        RECT 95.100 760.050 96.900 761.850 ;
        RECT 101.700 760.050 102.900 767.400 ;
        RECT 106.950 762.450 109.050 763.050 ;
        RECT 112.950 762.450 115.050 763.050 ;
        RECT 106.950 761.550 115.050 762.450 ;
        RECT 106.950 760.950 109.050 761.550 ;
        RECT 112.950 760.950 115.050 761.550 ;
        RECT 119.250 760.050 121.050 761.850 ;
        RECT 122.400 760.050 123.300 767.400 ;
        RECT 125.100 760.050 126.900 761.850 ;
        RECT 140.700 760.050 141.900 773.400 ;
        RECT 159.000 773.100 159.900 773.400 ;
        RECT 164.100 773.400 165.900 779.400 ;
        RECT 167.100 773.400 168.900 780.000 ;
        RECT 182.100 773.400 183.900 780.000 ;
        RECT 185.100 773.400 186.900 779.400 ;
        RECT 188.100 774.000 189.900 780.000 ;
        RECT 164.100 773.100 165.600 773.400 ;
        RECT 159.000 772.200 165.600 773.100 ;
        RECT 185.400 773.100 186.900 773.400 ;
        RECT 191.100 773.400 192.900 779.400 ;
        RECT 191.100 773.100 192.000 773.400 ;
        RECT 185.400 772.200 192.000 773.100 ;
        RECT 143.100 760.050 144.900 761.850 ;
        RECT 159.000 760.050 159.900 772.200 ;
        RECT 164.100 760.050 165.900 761.850 ;
        RECT 185.100 760.050 186.900 761.850 ;
        RECT 191.100 760.050 192.000 772.200 ;
        RECT 206.100 768.300 207.900 779.400 ;
        RECT 209.100 769.200 210.900 780.000 ;
        RECT 212.100 768.300 213.900 779.400 ;
        RECT 206.100 767.400 213.900 768.300 ;
        RECT 215.100 767.400 216.900 779.400 ;
        RECT 230.400 767.400 232.200 780.000 ;
        RECT 235.500 768.900 237.300 779.400 ;
        RECT 238.500 773.400 240.300 780.000 ;
        RECT 238.200 770.100 240.000 771.900 ;
        RECT 241.950 771.450 244.050 772.050 ;
        RECT 253.950 771.450 256.050 772.050 ;
        RECT 241.950 770.550 256.050 771.450 ;
        RECT 241.950 769.950 244.050 770.550 ;
        RECT 253.950 769.950 256.050 770.550 ;
        RECT 235.500 767.400 237.900 768.900 ;
        RECT 257.100 767.400 258.900 779.400 ;
        RECT 260.100 768.000 261.900 780.000 ;
        RECT 263.100 773.400 264.900 779.400 ;
        RECT 266.100 773.400 267.900 780.000 ;
        RECT 281.100 773.400 282.900 780.000 ;
        RECT 284.100 773.400 285.900 779.400 ;
        RECT 287.100 774.000 288.900 780.000 ;
        RECT 199.950 765.450 202.050 766.050 ;
        RECT 205.950 765.450 208.050 766.200 ;
        RECT 199.950 764.550 208.050 765.450 ;
        RECT 199.950 763.950 202.050 764.550 ;
        RECT 205.950 764.100 208.050 764.550 ;
        RECT 209.250 760.050 211.050 761.850 ;
        RECT 215.700 760.050 216.600 767.400 ;
        RECT 230.100 760.050 231.900 761.850 ;
        RECT 236.700 760.050 237.900 767.400 ;
        RECT 238.950 765.450 241.050 766.050 ;
        RECT 244.950 765.450 247.050 766.050 ;
        RECT 238.950 764.550 247.050 765.450 ;
        RECT 238.950 763.950 241.050 764.550 ;
        RECT 244.950 763.950 247.050 764.550 ;
        RECT 257.700 760.050 258.600 767.400 ;
        RECT 261.000 760.050 262.800 761.850 ;
        RECT 13.950 757.950 16.050 760.050 ;
        RECT 16.950 757.950 19.050 760.050 ;
        RECT 34.950 757.950 37.050 760.050 ;
        RECT 37.950 757.950 40.050 760.050 ;
        RECT 40.950 757.950 43.050 760.050 ;
        RECT 43.950 757.950 46.050 760.050 ;
        RECT 61.800 757.950 63.900 760.050 ;
        RECT 67.950 757.950 70.050 760.050 ;
        RECT 70.950 757.950 73.050 760.050 ;
        RECT 76.500 757.950 78.600 760.050 ;
        RECT 94.950 757.950 97.050 760.050 ;
        RECT 97.950 757.950 100.050 760.050 ;
        RECT 100.950 757.950 103.050 760.050 ;
        RECT 103.950 757.950 106.050 760.050 ;
        RECT 118.950 757.950 121.050 760.050 ;
        RECT 121.950 757.950 124.050 760.050 ;
        RECT 124.950 757.950 127.050 760.050 ;
        RECT 139.950 757.950 142.050 760.050 ;
        RECT 142.950 757.950 145.050 760.050 ;
        RECT 157.950 757.950 160.050 760.050 ;
        RECT 160.950 757.950 163.050 760.050 ;
        RECT 163.950 757.950 166.050 760.050 ;
        RECT 166.950 757.950 169.050 760.050 ;
        RECT 181.950 757.950 184.050 760.050 ;
        RECT 184.950 757.950 187.050 760.050 ;
        RECT 187.950 757.950 190.050 760.050 ;
        RECT 190.950 757.950 193.050 760.050 ;
        RECT 205.950 757.950 208.050 760.050 ;
        RECT 208.950 757.950 211.050 760.050 ;
        RECT 211.950 757.950 214.050 760.050 ;
        RECT 214.950 757.950 217.050 760.050 ;
        RECT 229.950 757.950 232.050 760.050 ;
        RECT 232.950 757.950 235.050 760.050 ;
        RECT 235.950 757.950 238.050 760.050 ;
        RECT 238.950 757.950 241.050 760.050 ;
        RECT 257.100 757.950 259.200 760.050 ;
        RECT 260.400 757.950 262.500 760.050 ;
        RECT 14.700 747.600 15.900 757.950 ;
        RECT 35.100 756.150 36.900 757.950 ;
        RECT 38.100 753.600 39.300 757.950 ;
        RECT 41.100 756.150 42.900 757.950 ;
        RECT 67.950 756.150 69.750 757.950 ;
        RECT 35.700 752.700 39.300 753.600 ;
        RECT 35.700 750.600 36.900 752.700 ;
        RECT 14.100 744.600 15.900 747.600 ;
        RECT 17.100 744.000 18.900 747.600 ;
        RECT 35.100 744.600 36.900 750.600 ;
        RECT 38.100 749.700 45.900 751.050 ;
        RECT 38.100 744.600 39.900 749.700 ;
        RECT 41.100 744.000 42.900 748.800 ;
        RECT 44.100 744.600 45.900 749.700 ;
        RECT 77.100 749.400 78.300 757.950 ;
        RECT 98.100 756.150 99.900 757.950 ;
        RECT 101.700 753.600 102.900 757.950 ;
        RECT 104.100 756.150 105.900 757.950 ;
        RECT 101.700 752.700 105.300 753.600 ;
        RECT 65.700 748.500 78.300 749.400 ;
        RECT 95.100 749.700 102.900 751.050 ;
        RECT 65.700 747.600 66.600 748.500 ;
        RECT 72.900 747.600 73.800 748.500 ;
        RECT 61.800 744.000 63.900 747.600 ;
        RECT 65.100 744.600 66.900 747.600 ;
        RECT 68.100 744.000 69.900 747.600 ;
        RECT 71.100 744.600 73.800 747.600 ;
        RECT 95.100 744.600 96.900 749.700 ;
        RECT 98.100 744.000 99.900 748.800 ;
        RECT 101.100 744.600 102.900 749.700 ;
        RECT 104.100 750.600 105.300 752.700 ;
        RECT 104.100 744.600 105.900 750.600 ;
        RECT 122.400 747.600 123.300 757.950 ;
        RECT 140.700 747.600 141.900 757.950 ;
        RECT 159.000 754.200 159.900 757.950 ;
        RECT 161.100 756.150 162.900 757.950 ;
        RECT 167.100 756.150 168.900 757.950 ;
        RECT 182.100 756.150 183.900 757.950 ;
        RECT 188.100 756.150 189.900 757.950 ;
        RECT 191.100 754.200 192.000 757.950 ;
        RECT 206.100 756.150 207.900 757.950 ;
        RECT 212.250 756.150 214.050 757.950 ;
        RECT 159.000 753.000 162.300 754.200 ;
        RECT 119.100 744.000 120.900 747.600 ;
        RECT 122.100 744.600 123.900 747.600 ;
        RECT 125.100 744.000 126.900 747.600 ;
        RECT 140.100 744.600 141.900 747.600 ;
        RECT 143.100 744.000 144.900 747.600 ;
        RECT 160.500 744.600 162.300 753.000 ;
        RECT 167.100 744.000 168.900 753.600 ;
        RECT 182.100 744.000 183.900 753.600 ;
        RECT 188.700 753.000 192.000 754.200 ;
        RECT 188.700 744.600 190.500 753.000 ;
        RECT 215.700 750.600 216.600 757.950 ;
        RECT 233.100 756.150 234.900 757.950 ;
        RECT 236.700 753.600 237.900 757.950 ;
        RECT 239.100 756.150 240.900 757.950 ;
        RECT 236.700 752.700 240.300 753.600 ;
        RECT 207.000 744.000 208.800 750.600 ;
        RECT 211.500 749.400 216.600 750.600 ;
        RECT 230.100 749.700 237.900 751.050 ;
        RECT 211.500 744.600 213.300 749.400 ;
        RECT 214.500 744.000 216.300 747.600 ;
        RECT 230.100 744.600 231.900 749.700 ;
        RECT 233.100 744.000 234.900 748.800 ;
        RECT 236.100 744.600 237.900 749.700 ;
        RECT 239.100 750.600 240.300 752.700 ;
        RECT 257.700 750.600 258.600 757.950 ;
        RECT 264.000 753.300 264.900 773.400 ;
        RECT 284.400 773.100 285.900 773.400 ;
        RECT 290.100 773.400 291.900 779.400 ;
        RECT 305.100 773.400 306.900 780.000 ;
        RECT 308.100 773.400 309.900 779.400 ;
        RECT 323.100 778.500 330.900 779.400 ;
        RECT 290.100 773.100 291.000 773.400 ;
        RECT 284.400 772.200 291.000 773.100 ;
        RECT 265.950 765.450 268.050 766.050 ;
        RECT 286.950 765.450 289.050 766.050 ;
        RECT 265.950 764.550 289.050 765.450 ;
        RECT 265.950 763.950 268.050 764.550 ;
        RECT 286.950 763.950 289.050 764.550 ;
        RECT 284.100 760.050 285.900 761.850 ;
        RECT 290.100 760.050 291.000 772.200 ;
        RECT 305.100 760.050 306.900 761.850 ;
        RECT 308.100 760.050 309.300 773.400 ;
        RECT 323.100 767.400 324.900 778.500 ;
        RECT 326.100 766.500 327.900 777.600 ;
        RECT 329.100 768.600 330.900 778.500 ;
        RECT 332.100 769.500 333.900 780.000 ;
        RECT 335.100 768.600 336.900 779.400 ;
        RECT 353.100 773.400 354.900 780.000 ;
        RECT 356.100 773.400 357.900 779.400 ;
        RECT 359.100 774.000 360.900 780.000 ;
        RECT 356.400 773.100 357.900 773.400 ;
        RECT 362.100 773.400 363.900 779.400 ;
        RECT 362.100 773.100 363.000 773.400 ;
        RECT 356.400 772.200 363.000 773.100 ;
        RECT 329.100 767.700 336.900 768.600 ;
        RECT 326.100 765.600 330.900 766.500 ;
        RECT 326.100 760.050 327.900 761.850 ;
        RECT 330.000 760.050 330.900 765.600 ;
        RECT 337.950 762.450 340.050 763.050 ;
        RECT 346.950 762.450 349.050 763.050 ;
        RECT 331.950 760.050 333.750 761.850 ;
        RECT 337.950 761.550 349.050 762.450 ;
        RECT 337.950 760.950 340.050 761.550 ;
        RECT 346.950 760.950 349.050 761.550 ;
        RECT 356.100 760.050 357.900 761.850 ;
        RECT 362.100 760.050 363.000 772.200 ;
        RECT 377.100 768.300 378.900 779.400 ;
        RECT 380.100 769.200 381.900 780.000 ;
        RECT 383.100 768.300 384.900 779.400 ;
        RECT 377.100 767.400 384.900 768.300 ;
        RECT 386.100 767.400 387.900 779.400 ;
        RECT 401.100 773.400 402.900 780.000 ;
        RECT 404.100 773.400 405.900 779.400 ;
        RECT 407.100 774.000 408.900 780.000 ;
        RECT 404.400 773.100 405.900 773.400 ;
        RECT 410.100 773.400 411.900 779.400 ;
        RECT 425.100 773.400 426.900 779.400 ;
        RECT 428.100 774.000 429.900 780.000 ;
        RECT 410.100 773.100 411.000 773.400 ;
        RECT 404.400 772.200 411.000 773.100 ;
        RECT 380.250 760.050 382.050 761.850 ;
        RECT 386.700 760.050 387.600 767.400 ;
        RECT 404.100 760.050 405.900 761.850 ;
        RECT 410.100 760.050 411.000 772.200 ;
        RECT 426.000 773.100 426.900 773.400 ;
        RECT 431.100 773.400 432.900 779.400 ;
        RECT 434.100 773.400 435.900 780.000 ;
        RECT 449.100 773.400 450.900 780.000 ;
        RECT 452.100 773.400 453.900 779.400 ;
        RECT 455.100 774.000 456.900 780.000 ;
        RECT 431.100 773.100 432.600 773.400 ;
        RECT 426.000 772.200 432.600 773.100 ;
        RECT 452.400 773.100 453.900 773.400 ;
        RECT 458.100 773.400 459.900 779.400 ;
        RECT 458.100 773.100 459.000 773.400 ;
        RECT 452.400 772.200 459.000 773.100 ;
        RECT 426.000 760.050 426.900 772.200 ;
        RECT 431.100 760.050 432.900 761.850 ;
        RECT 452.100 760.050 453.900 761.850 ;
        RECT 458.100 760.050 459.000 772.200 ;
        RECT 473.100 768.300 474.900 779.400 ;
        RECT 476.100 769.200 477.900 780.000 ;
        RECT 479.100 768.300 480.900 779.400 ;
        RECT 473.100 767.400 480.900 768.300 ;
        RECT 482.100 767.400 483.900 779.400 ;
        RECT 497.100 767.400 498.900 779.400 ;
        RECT 500.100 768.300 501.900 779.400 ;
        RECT 503.100 769.200 504.900 780.000 ;
        RECT 506.100 768.300 507.900 779.400 ;
        RECT 521.100 773.400 522.900 780.000 ;
        RECT 524.100 773.400 525.900 779.400 ;
        RECT 527.100 774.000 528.900 780.000 ;
        RECT 524.400 773.100 525.900 773.400 ;
        RECT 530.100 773.400 531.900 779.400 ;
        RECT 545.100 773.400 546.900 780.000 ;
        RECT 548.100 773.400 549.900 779.400 ;
        RECT 530.100 773.100 531.000 773.400 ;
        RECT 524.400 772.200 531.000 773.100 ;
        RECT 500.100 767.400 507.900 768.300 ;
        RECT 463.950 765.450 466.050 766.050 ;
        RECT 475.950 765.450 478.050 766.050 ;
        RECT 463.950 764.550 478.050 765.450 ;
        RECT 463.950 763.950 466.050 764.550 ;
        RECT 475.950 763.950 478.050 764.550 ;
        RECT 476.250 760.050 478.050 761.850 ;
        RECT 482.700 760.050 483.600 767.400 ;
        RECT 497.400 760.050 498.300 767.400 ;
        RECT 502.950 760.050 504.750 761.850 ;
        RECT 524.100 760.050 525.900 761.850 ;
        RECT 530.100 760.050 531.000 772.200 ;
        RECT 265.800 757.950 267.900 760.050 ;
        RECT 280.950 757.950 283.050 760.050 ;
        RECT 283.950 757.950 286.050 760.050 ;
        RECT 286.950 757.950 289.050 760.050 ;
        RECT 289.950 757.950 292.050 760.050 ;
        RECT 304.950 757.950 307.050 760.050 ;
        RECT 307.950 757.950 310.050 760.050 ;
        RECT 322.950 757.950 325.050 760.050 ;
        RECT 325.950 757.950 328.050 760.050 ;
        RECT 328.950 757.950 331.050 760.050 ;
        RECT 331.950 757.950 334.050 760.050 ;
        RECT 334.950 757.950 337.050 760.050 ;
        RECT 352.950 757.950 355.050 760.050 ;
        RECT 355.950 757.950 358.050 760.050 ;
        RECT 358.950 757.950 361.050 760.050 ;
        RECT 361.950 757.950 364.050 760.050 ;
        RECT 376.950 757.950 379.050 760.050 ;
        RECT 379.950 757.950 382.050 760.050 ;
        RECT 382.950 757.950 385.050 760.050 ;
        RECT 385.950 757.950 388.050 760.050 ;
        RECT 400.950 757.950 403.050 760.050 ;
        RECT 403.950 757.950 406.050 760.050 ;
        RECT 406.950 757.950 409.050 760.050 ;
        RECT 409.950 757.950 412.050 760.050 ;
        RECT 424.950 757.950 427.050 760.050 ;
        RECT 427.950 757.950 430.050 760.050 ;
        RECT 430.950 757.950 433.050 760.050 ;
        RECT 433.950 757.950 436.050 760.050 ;
        RECT 448.950 757.950 451.050 760.050 ;
        RECT 451.950 757.950 454.050 760.050 ;
        RECT 454.950 757.950 457.050 760.050 ;
        RECT 457.950 757.950 460.050 760.050 ;
        RECT 472.950 757.950 475.050 760.050 ;
        RECT 475.950 757.950 478.050 760.050 ;
        RECT 478.950 757.950 481.050 760.050 ;
        RECT 481.950 757.950 484.050 760.050 ;
        RECT 496.950 757.950 499.050 760.050 ;
        RECT 499.950 757.950 502.050 760.050 ;
        RECT 502.950 757.950 505.050 760.050 ;
        RECT 505.950 757.950 508.050 760.050 ;
        RECT 520.950 757.950 523.050 760.050 ;
        RECT 523.950 757.950 526.050 760.050 ;
        RECT 526.950 757.950 529.050 760.050 ;
        RECT 529.950 757.950 532.050 760.050 ;
        RECT 545.100 757.950 547.200 760.050 ;
        RECT 265.950 756.150 267.750 757.950 ;
        RECT 281.100 756.150 282.900 757.950 ;
        RECT 287.100 756.150 288.900 757.950 ;
        RECT 290.100 754.200 291.000 757.950 ;
        RECT 259.500 752.400 267.900 753.300 ;
        RECT 259.500 751.500 261.300 752.400 ;
        RECT 239.100 744.600 240.900 750.600 ;
        RECT 257.700 748.800 260.400 750.600 ;
        RECT 258.600 744.600 260.400 748.800 ;
        RECT 261.600 744.000 263.400 750.600 ;
        RECT 266.100 744.600 267.900 752.400 ;
        RECT 281.100 744.000 282.900 753.600 ;
        RECT 287.700 753.000 291.000 754.200 ;
        RECT 287.700 744.600 289.500 753.000 ;
        RECT 308.100 747.600 309.300 757.950 ;
        RECT 323.100 756.150 324.900 757.950 ;
        RECT 329.700 750.600 330.900 757.950 ;
        RECT 334.950 756.150 336.750 757.950 ;
        RECT 353.100 756.150 354.900 757.950 ;
        RECT 359.100 756.150 360.900 757.950 ;
        RECT 362.100 754.200 363.000 757.950 ;
        RECT 377.100 756.150 378.900 757.950 ;
        RECT 383.250 756.150 385.050 757.950 ;
        RECT 305.100 744.000 306.900 747.600 ;
        RECT 308.100 744.600 309.900 747.600 ;
        RECT 325.500 744.000 327.300 750.600 ;
        RECT 330.000 744.600 331.800 750.600 ;
        RECT 334.500 744.000 336.300 750.600 ;
        RECT 353.100 744.000 354.900 753.600 ;
        RECT 359.700 753.000 363.000 754.200 ;
        RECT 359.700 744.600 361.500 753.000 ;
        RECT 386.700 750.600 387.600 757.950 ;
        RECT 401.100 756.150 402.900 757.950 ;
        RECT 407.100 756.150 408.900 757.950 ;
        RECT 410.100 754.200 411.000 757.950 ;
        RECT 378.000 744.000 379.800 750.600 ;
        RECT 382.500 749.400 387.600 750.600 ;
        RECT 382.500 744.600 384.300 749.400 ;
        RECT 385.500 744.000 387.300 747.600 ;
        RECT 401.100 744.000 402.900 753.600 ;
        RECT 407.700 753.000 411.000 754.200 ;
        RECT 426.000 754.200 426.900 757.950 ;
        RECT 428.100 756.150 429.900 757.950 ;
        RECT 434.100 756.150 435.900 757.950 ;
        RECT 449.100 756.150 450.900 757.950 ;
        RECT 455.100 756.150 456.900 757.950 ;
        RECT 458.100 754.200 459.000 757.950 ;
        RECT 473.100 756.150 474.900 757.950 ;
        RECT 479.250 756.150 481.050 757.950 ;
        RECT 426.000 753.000 429.300 754.200 ;
        RECT 407.700 744.600 409.500 753.000 ;
        RECT 427.500 744.600 429.300 753.000 ;
        RECT 434.100 744.000 435.900 753.600 ;
        RECT 449.100 744.000 450.900 753.600 ;
        RECT 455.700 753.000 459.000 754.200 ;
        RECT 455.700 744.600 457.500 753.000 ;
        RECT 482.700 750.600 483.600 757.950 ;
        RECT 474.000 744.000 475.800 750.600 ;
        RECT 478.500 749.400 483.600 750.600 ;
        RECT 497.400 750.600 498.300 757.950 ;
        RECT 499.950 756.150 501.750 757.950 ;
        RECT 506.100 756.150 507.900 757.950 ;
        RECT 521.100 756.150 522.900 757.950 ;
        RECT 527.100 756.150 528.900 757.950 ;
        RECT 530.100 754.200 531.000 757.950 ;
        RECT 545.250 756.150 547.050 757.950 ;
        RECT 497.400 749.400 502.500 750.600 ;
        RECT 478.500 744.600 480.300 749.400 ;
        RECT 481.500 744.000 483.300 747.600 ;
        RECT 497.700 744.000 499.500 747.600 ;
        RECT 500.700 744.600 502.500 749.400 ;
        RECT 505.200 744.000 507.000 750.600 ;
        RECT 521.100 744.000 522.900 753.600 ;
        RECT 527.700 753.000 531.000 754.200 ;
        RECT 548.100 753.300 549.000 773.400 ;
        RECT 551.100 768.000 552.900 780.000 ;
        RECT 554.100 767.400 555.900 779.400 ;
        RECT 556.950 774.450 559.050 775.050 ;
        RECT 562.950 774.450 565.050 775.050 ;
        RECT 556.950 773.550 565.050 774.450 ;
        RECT 556.950 772.950 559.050 773.550 ;
        RECT 562.950 772.950 565.050 773.550 ;
        RECT 569.100 773.400 570.900 779.400 ;
        RECT 572.100 774.000 573.900 780.000 ;
        RECT 570.000 773.100 570.900 773.400 ;
        RECT 575.100 773.400 576.900 779.400 ;
        RECT 578.100 773.400 579.900 780.000 ;
        RECT 593.100 773.400 594.900 780.000 ;
        RECT 596.100 773.400 597.900 779.400 ;
        RECT 611.100 773.400 612.900 779.400 ;
        RECT 614.100 774.000 615.900 780.000 ;
        RECT 575.100 773.100 576.600 773.400 ;
        RECT 570.000 772.200 576.600 773.100 ;
        RECT 550.200 760.050 552.000 761.850 ;
        RECT 554.400 760.050 555.300 767.400 ;
        RECT 570.000 760.050 570.900 772.200 ;
        RECT 575.100 760.050 576.900 761.850 ;
        RECT 593.100 760.050 594.900 761.850 ;
        RECT 596.100 760.050 597.300 773.400 ;
        RECT 612.000 773.100 612.900 773.400 ;
        RECT 617.100 773.400 618.900 779.400 ;
        RECT 620.100 773.400 621.900 780.000 ;
        RECT 617.100 773.100 618.600 773.400 ;
        RECT 612.000 772.200 618.600 773.100 ;
        RECT 612.000 760.050 612.900 772.200 ;
        RECT 635.100 768.300 636.900 779.400 ;
        RECT 638.100 769.200 639.900 780.000 ;
        RECT 641.100 768.300 642.900 779.400 ;
        RECT 635.100 767.400 642.900 768.300 ;
        RECT 644.100 767.400 645.900 779.400 ;
        RECT 662.100 773.400 663.900 779.400 ;
        RECT 665.100 774.000 666.900 780.000 ;
        RECT 663.000 773.100 663.900 773.400 ;
        RECT 668.100 773.400 669.900 779.400 ;
        RECT 671.100 773.400 672.900 780.000 ;
        RECT 668.100 773.100 669.600 773.400 ;
        RECT 663.000 772.200 669.600 773.100 ;
        RECT 622.950 765.450 625.050 766.050 ;
        RECT 640.950 765.450 643.050 766.050 ;
        RECT 622.950 764.550 643.050 765.450 ;
        RECT 622.950 763.950 625.050 764.550 ;
        RECT 640.950 763.950 643.050 764.550 ;
        RECT 617.100 760.050 618.900 761.850 ;
        RECT 638.250 760.050 640.050 761.850 ;
        RECT 644.700 760.050 645.600 767.400 ;
        RECT 663.000 760.050 663.900 772.200 ;
        RECT 686.100 768.300 687.900 779.400 ;
        RECT 689.100 769.200 690.900 780.000 ;
        RECT 692.100 768.300 693.900 779.400 ;
        RECT 686.100 767.400 693.900 768.300 ;
        RECT 695.100 767.400 696.900 779.400 ;
        RECT 710.100 773.400 711.900 780.000 ;
        RECT 713.100 773.400 714.900 779.400 ;
        RECT 670.950 765.450 673.050 766.050 ;
        RECT 676.950 765.450 679.050 766.050 ;
        RECT 670.950 764.550 679.050 765.450 ;
        RECT 670.950 763.950 673.050 764.550 ;
        RECT 676.950 763.950 679.050 764.550 ;
        RECT 668.100 760.050 669.900 761.850 ;
        RECT 689.250 760.050 691.050 761.850 ;
        RECT 695.700 760.050 696.600 767.400 ;
        RECT 710.100 760.050 711.900 761.850 ;
        RECT 713.100 760.050 714.300 773.400 ;
        RECT 731.100 767.400 732.900 779.400 ;
        RECT 734.100 768.300 735.900 779.400 ;
        RECT 737.100 769.200 738.900 780.000 ;
        RECT 740.100 768.300 741.900 779.400 ;
        RECT 734.100 767.400 741.900 768.300 ;
        RECT 755.100 768.300 756.900 779.400 ;
        RECT 758.100 769.200 759.900 780.000 ;
        RECT 761.100 768.300 762.900 779.400 ;
        RECT 755.100 767.400 762.900 768.300 ;
        RECT 764.100 767.400 765.900 779.400 ;
        RECT 779.100 773.400 780.900 779.400 ;
        RECT 782.100 773.400 783.900 780.000 ;
        RECT 797.100 773.400 798.900 779.400 ;
        RECT 800.100 774.000 801.900 780.000 ;
        RECT 731.400 760.050 732.300 767.400 ;
        RECT 733.950 765.450 736.050 766.050 ;
        RECT 754.950 765.450 757.050 766.050 ;
        RECT 733.950 764.550 757.050 765.450 ;
        RECT 733.950 763.950 736.050 764.550 ;
        RECT 754.950 763.950 757.050 764.550 ;
        RECT 736.950 760.050 738.750 761.850 ;
        RECT 758.250 760.050 760.050 761.850 ;
        RECT 764.700 760.050 765.600 767.400 ;
        RECT 779.700 760.050 780.900 773.400 ;
        RECT 798.000 773.100 798.900 773.400 ;
        RECT 803.100 773.400 804.900 779.400 ;
        RECT 806.100 773.400 807.900 780.000 ;
        RECT 821.700 773.400 823.500 780.000 ;
        RECT 803.100 773.100 804.600 773.400 ;
        RECT 798.000 772.200 804.600 773.100 ;
        RECT 782.100 760.050 783.900 761.850 ;
        RECT 798.000 760.050 798.900 772.200 ;
        RECT 822.000 770.100 823.800 771.900 ;
        RECT 824.700 768.900 826.500 779.400 ;
        RECT 824.100 767.400 826.500 768.900 ;
        RECT 829.800 767.400 831.600 780.000 ;
        RECT 845.100 767.400 846.900 779.400 ;
        RECT 848.100 768.300 849.900 779.400 ;
        RECT 851.100 769.200 852.900 780.000 ;
        RECT 854.100 768.300 855.900 779.400 ;
        RECT 869.100 773.400 870.900 780.000 ;
        RECT 872.100 773.400 873.900 779.400 ;
        RECT 875.100 774.000 876.900 780.000 ;
        RECT 872.400 773.100 873.900 773.400 ;
        RECT 878.100 773.400 879.900 779.400 ;
        RECT 878.100 773.100 879.000 773.400 ;
        RECT 872.400 772.200 879.000 773.100 ;
        RECT 848.100 767.400 855.900 768.300 ;
        RECT 803.100 760.050 804.900 761.850 ;
        RECT 824.100 760.050 825.300 767.400 ;
        RECT 830.100 760.050 831.900 761.850 ;
        RECT 845.400 760.050 846.300 767.400 ;
        RECT 853.950 765.450 856.050 766.050 ;
        RECT 874.950 765.450 877.050 766.050 ;
        RECT 853.950 764.550 877.050 765.450 ;
        RECT 853.950 763.950 856.050 764.550 ;
        RECT 874.950 763.950 877.050 764.550 ;
        RECT 850.950 760.050 852.750 761.850 ;
        RECT 872.100 760.050 873.900 761.850 ;
        RECT 878.100 760.050 879.000 772.200 ;
        RECT 550.500 757.950 552.600 760.050 ;
        RECT 553.800 757.950 555.900 760.050 ;
        RECT 568.950 757.950 571.050 760.050 ;
        RECT 571.950 757.950 574.050 760.050 ;
        RECT 574.950 757.950 577.050 760.050 ;
        RECT 577.950 757.950 580.050 760.050 ;
        RECT 592.950 757.950 595.050 760.050 ;
        RECT 595.950 757.950 598.050 760.050 ;
        RECT 610.950 757.950 613.050 760.050 ;
        RECT 613.950 757.950 616.050 760.050 ;
        RECT 616.950 757.950 619.050 760.050 ;
        RECT 619.950 757.950 622.050 760.050 ;
        RECT 634.950 757.950 637.050 760.050 ;
        RECT 637.950 757.950 640.050 760.050 ;
        RECT 640.950 757.950 643.050 760.050 ;
        RECT 643.950 757.950 646.050 760.050 ;
        RECT 661.950 757.950 664.050 760.050 ;
        RECT 664.950 757.950 667.050 760.050 ;
        RECT 667.950 757.950 670.050 760.050 ;
        RECT 670.950 757.950 673.050 760.050 ;
        RECT 685.950 757.950 688.050 760.050 ;
        RECT 688.950 757.950 691.050 760.050 ;
        RECT 691.950 757.950 694.050 760.050 ;
        RECT 694.950 757.950 697.050 760.050 ;
        RECT 709.950 757.950 712.050 760.050 ;
        RECT 712.950 757.950 715.050 760.050 ;
        RECT 730.950 757.950 733.050 760.050 ;
        RECT 733.950 757.950 736.050 760.050 ;
        RECT 736.950 757.950 739.050 760.050 ;
        RECT 739.950 757.950 742.050 760.050 ;
        RECT 754.950 757.950 757.050 760.050 ;
        RECT 757.950 757.950 760.050 760.050 ;
        RECT 760.950 757.950 763.050 760.050 ;
        RECT 763.950 757.950 766.050 760.050 ;
        RECT 778.950 757.950 781.050 760.050 ;
        RECT 781.950 757.950 784.050 760.050 ;
        RECT 796.950 757.950 799.050 760.050 ;
        RECT 799.950 757.950 802.050 760.050 ;
        RECT 802.950 757.950 805.050 760.050 ;
        RECT 805.950 757.950 808.050 760.050 ;
        RECT 820.950 757.950 823.050 760.050 ;
        RECT 823.950 757.950 826.050 760.050 ;
        RECT 826.950 757.950 829.050 760.050 ;
        RECT 829.950 757.950 832.050 760.050 ;
        RECT 844.950 757.950 847.050 760.050 ;
        RECT 847.950 757.950 850.050 760.050 ;
        RECT 850.950 757.950 853.050 760.050 ;
        RECT 853.950 757.950 856.050 760.050 ;
        RECT 868.950 757.950 871.050 760.050 ;
        RECT 871.950 757.950 874.050 760.050 ;
        RECT 874.950 757.950 877.050 760.050 ;
        RECT 877.950 757.950 880.050 760.050 ;
        RECT 527.700 744.600 529.500 753.000 ;
        RECT 545.100 752.400 553.500 753.300 ;
        RECT 545.100 744.600 546.900 752.400 ;
        RECT 551.700 751.500 553.500 752.400 ;
        RECT 554.400 750.600 555.300 757.950 ;
        RECT 570.000 754.200 570.900 757.950 ;
        RECT 572.100 756.150 573.900 757.950 ;
        RECT 578.100 756.150 579.900 757.950 ;
        RECT 570.000 753.000 573.300 754.200 ;
        RECT 549.600 744.000 551.400 750.600 ;
        RECT 552.600 748.800 555.300 750.600 ;
        RECT 552.600 744.600 554.400 748.800 ;
        RECT 571.500 744.600 573.300 753.000 ;
        RECT 578.100 744.000 579.900 753.600 ;
        RECT 596.100 747.600 597.300 757.950 ;
        RECT 612.000 754.200 612.900 757.950 ;
        RECT 614.100 756.150 615.900 757.950 ;
        RECT 620.100 756.150 621.900 757.950 ;
        RECT 635.100 756.150 636.900 757.950 ;
        RECT 641.250 756.150 643.050 757.950 ;
        RECT 612.000 753.000 615.300 754.200 ;
        RECT 593.100 744.000 594.900 747.600 ;
        RECT 596.100 744.600 597.900 747.600 ;
        RECT 613.500 744.600 615.300 753.000 ;
        RECT 620.100 744.000 621.900 753.600 ;
        RECT 644.700 750.600 645.600 757.950 ;
        RECT 663.000 754.200 663.900 757.950 ;
        RECT 665.100 756.150 666.900 757.950 ;
        RECT 671.100 756.150 672.900 757.950 ;
        RECT 686.100 756.150 687.900 757.950 ;
        RECT 692.250 756.150 694.050 757.950 ;
        RECT 663.000 753.000 666.300 754.200 ;
        RECT 636.000 744.000 637.800 750.600 ;
        RECT 640.500 749.400 645.600 750.600 ;
        RECT 640.500 744.600 642.300 749.400 ;
        RECT 643.500 744.000 645.300 747.600 ;
        RECT 664.500 744.600 666.300 753.000 ;
        RECT 671.100 744.000 672.900 753.600 ;
        RECT 695.700 750.600 696.600 757.950 ;
        RECT 687.000 744.000 688.800 750.600 ;
        RECT 691.500 749.400 696.600 750.600 ;
        RECT 691.500 744.600 693.300 749.400 ;
        RECT 713.100 747.600 714.300 757.950 ;
        RECT 718.950 750.450 721.050 751.050 ;
        RECT 727.950 750.450 730.050 751.050 ;
        RECT 718.950 749.550 730.050 750.450 ;
        RECT 718.950 748.950 721.050 749.550 ;
        RECT 727.950 748.950 730.050 749.550 ;
        RECT 731.400 750.600 732.300 757.950 ;
        RECT 733.950 756.150 735.750 757.950 ;
        RECT 740.100 756.150 741.900 757.950 ;
        RECT 755.100 756.150 756.900 757.950 ;
        RECT 761.250 756.150 763.050 757.950 ;
        RECT 764.700 750.600 765.600 757.950 ;
        RECT 731.400 749.400 736.500 750.600 ;
        RECT 694.500 744.000 696.300 747.600 ;
        RECT 710.100 744.000 711.900 747.600 ;
        RECT 713.100 744.600 714.900 747.600 ;
        RECT 731.700 744.000 733.500 747.600 ;
        RECT 734.700 744.600 736.500 749.400 ;
        RECT 739.200 744.000 741.000 750.600 ;
        RECT 756.000 744.000 757.800 750.600 ;
        RECT 760.500 749.400 765.600 750.600 ;
        RECT 760.500 744.600 762.300 749.400 ;
        RECT 779.700 747.600 780.900 757.950 ;
        RECT 798.000 754.200 798.900 757.950 ;
        RECT 800.100 756.150 801.900 757.950 ;
        RECT 806.100 756.150 807.900 757.950 ;
        RECT 821.100 756.150 822.900 757.950 ;
        RECT 798.000 753.000 801.300 754.200 ;
        RECT 824.100 753.600 825.300 757.950 ;
        RECT 827.100 756.150 828.900 757.950 ;
        RECT 763.500 744.000 765.300 747.600 ;
        RECT 779.100 744.600 780.900 747.600 ;
        RECT 782.100 744.000 783.900 747.600 ;
        RECT 799.500 744.600 801.300 753.000 ;
        RECT 806.100 744.000 807.900 753.600 ;
        RECT 821.700 752.700 825.300 753.600 ;
        RECT 821.700 750.600 822.900 752.700 ;
        RECT 821.100 744.600 822.900 750.600 ;
        RECT 824.100 749.700 831.900 751.050 ;
        RECT 824.100 744.600 825.900 749.700 ;
        RECT 827.100 744.000 828.900 748.800 ;
        RECT 830.100 744.600 831.900 749.700 ;
        RECT 845.400 750.600 846.300 757.950 ;
        RECT 847.950 756.150 849.750 757.950 ;
        RECT 854.100 756.150 855.900 757.950 ;
        RECT 869.100 756.150 870.900 757.950 ;
        RECT 875.100 756.150 876.900 757.950 ;
        RECT 878.100 754.200 879.000 757.950 ;
        RECT 845.400 749.400 850.500 750.600 ;
        RECT 845.700 744.000 847.500 747.600 ;
        RECT 848.700 744.600 850.500 749.400 ;
        RECT 853.200 744.000 855.000 750.600 ;
        RECT 869.100 744.000 870.900 753.600 ;
        RECT 875.700 753.000 879.000 754.200 ;
        RECT 875.700 744.600 877.500 753.000 ;
        RECT 14.100 734.400 15.900 740.400 ;
        RECT 17.100 734.400 18.900 741.000 ;
        RECT 20.100 737.400 21.900 740.400 ;
        RECT 14.100 727.050 15.300 734.400 ;
        RECT 20.700 733.500 21.900 737.400 ;
        RECT 16.200 732.600 21.900 733.500 ;
        RECT 23.550 734.400 25.350 740.400 ;
        RECT 26.850 734.400 28.650 741.000 ;
        RECT 31.950 737.400 33.750 740.400 ;
        RECT 36.450 737.400 38.250 741.000 ;
        RECT 39.450 737.400 41.250 740.400 ;
        RECT 42.750 737.400 44.550 741.000 ;
        RECT 47.250 738.300 49.050 740.400 ;
        RECT 47.250 737.400 50.850 738.300 ;
        RECT 31.350 735.300 33.750 737.400 ;
        RECT 40.200 736.500 41.250 737.400 ;
        RECT 47.250 736.800 51.150 737.400 ;
        RECT 40.200 735.450 45.150 736.500 ;
        RECT 43.350 734.700 45.150 735.450 ;
        RECT 16.200 731.700 18.000 732.600 ;
        RECT 14.100 724.950 16.200 727.050 ;
        RECT 14.100 717.600 15.300 724.950 ;
        RECT 17.100 720.300 18.000 731.700 ;
        RECT 23.550 727.050 24.750 734.400 ;
        RECT 46.350 733.800 48.150 735.600 ;
        RECT 49.050 735.300 51.150 736.800 ;
        RECT 52.050 734.400 53.850 741.000 ;
        RECT 55.050 736.200 56.850 740.400 ;
        RECT 55.050 734.400 57.450 736.200 ;
        RECT 36.150 732.000 37.950 732.600 ;
        RECT 47.100 732.000 48.150 733.800 ;
        RECT 36.150 730.800 48.150 732.000 ;
        RECT 19.500 724.950 21.600 727.050 ;
        RECT 19.800 723.150 21.600 724.950 ;
        RECT 23.550 725.250 29.850 727.050 ;
        RECT 23.550 724.950 28.050 725.250 ;
        RECT 16.200 719.400 18.000 720.300 ;
        RECT 16.200 718.500 21.900 719.400 ;
        RECT 14.100 705.600 15.900 717.600 ;
        RECT 17.100 705.000 18.900 715.800 ;
        RECT 20.700 711.600 21.900 718.500 ;
        RECT 20.100 705.600 21.900 711.600 ;
        RECT 23.550 717.600 24.750 724.950 ;
        RECT 25.650 722.100 27.450 722.250 ;
        RECT 31.350 722.100 33.450 722.400 ;
        RECT 25.650 720.900 33.450 722.100 ;
        RECT 25.650 720.450 27.450 720.900 ;
        RECT 31.350 720.300 33.450 720.900 ;
        RECT 36.150 718.200 37.050 730.800 ;
        RECT 47.100 729.600 55.050 730.800 ;
        RECT 47.100 729.000 48.900 729.600 ;
        RECT 50.100 727.800 51.900 728.400 ;
        RECT 43.800 726.600 51.900 727.800 ;
        RECT 53.250 727.050 55.050 729.600 ;
        RECT 43.800 724.950 45.900 726.600 ;
        RECT 52.950 724.950 55.050 727.050 ;
        RECT 45.750 719.700 47.550 720.000 ;
        RECT 56.550 719.700 57.450 734.400 ;
        RECT 71.100 731.400 72.900 741.000 ;
        RECT 77.700 732.000 79.500 740.400 ;
        RECT 96.000 734.400 97.800 741.000 ;
        RECT 100.500 735.600 102.300 740.400 ;
        RECT 103.500 737.400 105.300 741.000 ;
        RECT 100.500 734.400 105.600 735.600 ;
        RECT 77.700 730.800 81.000 732.000 ;
        RECT 71.100 727.050 72.900 728.850 ;
        RECT 77.100 727.050 78.900 728.850 ;
        RECT 80.100 727.050 81.000 730.800 ;
        RECT 95.100 727.050 96.900 728.850 ;
        RECT 101.250 727.050 103.050 728.850 ;
        RECT 104.700 727.050 105.600 734.400 ;
        RECT 122.700 733.200 124.500 740.400 ;
        RECT 127.800 734.400 129.600 741.000 ;
        RECT 122.700 732.300 126.900 733.200 ;
        RECT 122.100 727.050 123.900 728.850 ;
        RECT 125.700 727.050 126.900 732.300 ;
        RECT 143.100 731.400 144.900 741.000 ;
        RECT 149.700 732.000 151.500 740.400 ;
        RECT 170.700 737.400 172.500 741.000 ;
        RECT 173.700 735.600 175.500 740.400 ;
        RECT 170.400 734.400 175.500 735.600 ;
        RECT 178.200 734.400 180.000 741.000 ;
        RECT 149.700 730.800 153.000 732.000 ;
        RECT 127.950 727.050 129.750 728.850 ;
        RECT 143.100 727.050 144.900 728.850 ;
        RECT 149.100 727.050 150.900 728.850 ;
        RECT 152.100 727.050 153.000 730.800 ;
        RECT 170.400 727.050 171.300 734.400 ;
        RECT 194.700 733.200 196.500 740.400 ;
        RECT 199.800 734.400 201.600 741.000 ;
        RECT 215.700 734.400 217.500 741.000 ;
        RECT 220.200 734.400 222.000 740.400 ;
        RECT 224.700 734.400 226.500 741.000 ;
        RECT 242.100 735.300 243.900 740.400 ;
        RECT 245.100 736.200 246.900 741.000 ;
        RECT 248.100 735.300 249.900 740.400 ;
        RECT 194.700 732.300 198.900 733.200 ;
        RECT 172.950 727.050 174.750 728.850 ;
        RECT 179.100 727.050 180.900 728.850 ;
        RECT 194.100 727.050 195.900 728.850 ;
        RECT 197.700 727.050 198.900 732.300 ;
        RECT 199.950 727.050 201.750 728.850 ;
        RECT 215.250 727.050 217.050 728.850 ;
        RECT 221.100 727.050 222.300 734.400 ;
        RECT 242.100 733.950 249.900 735.300 ;
        RECT 251.100 734.400 252.900 740.400 ;
        RECT 266.100 735.300 267.900 740.400 ;
        RECT 269.100 736.200 270.900 741.000 ;
        RECT 272.100 735.300 273.900 740.400 ;
        RECT 251.100 732.300 252.300 734.400 ;
        RECT 266.100 733.950 273.900 735.300 ;
        RECT 275.100 734.400 276.900 740.400 ;
        RECT 290.100 735.300 291.900 740.400 ;
        RECT 293.100 736.200 294.900 741.000 ;
        RECT 296.100 735.300 297.900 740.400 ;
        RECT 275.100 732.300 276.300 734.400 ;
        RECT 290.100 733.950 297.900 735.300 ;
        RECT 299.100 734.400 300.900 740.400 ;
        RECT 299.100 732.300 300.300 734.400 ;
        RECT 248.700 731.400 252.300 732.300 ;
        RECT 272.700 731.400 276.300 732.300 ;
        RECT 296.700 731.400 300.300 732.300 ;
        RECT 317.100 731.400 318.900 741.000 ;
        RECT 323.700 732.000 325.500 740.400 ;
        RECT 343.500 732.000 345.300 740.400 ;
        RECT 227.100 727.050 228.900 728.850 ;
        RECT 245.100 727.050 246.900 728.850 ;
        RECT 248.700 727.050 249.900 731.400 ;
        RECT 251.100 727.050 252.900 728.850 ;
        RECT 269.100 727.050 270.900 728.850 ;
        RECT 272.700 727.050 273.900 731.400 ;
        RECT 275.100 727.050 276.900 728.850 ;
        RECT 293.100 727.050 294.900 728.850 ;
        RECT 296.700 727.050 297.900 731.400 ;
        RECT 323.700 730.800 327.000 732.000 ;
        RECT 299.100 727.050 300.900 728.850 ;
        RECT 317.100 727.050 318.900 728.850 ;
        RECT 323.100 727.050 324.900 728.850 ;
        RECT 326.100 727.050 327.000 730.800 ;
        RECT 342.000 730.800 345.300 732.000 ;
        RECT 350.100 731.400 351.900 741.000 ;
        RECT 366.000 734.400 367.800 741.000 ;
        RECT 370.500 735.600 372.300 740.400 ;
        RECT 373.500 737.400 375.300 741.000 ;
        RECT 370.500 734.400 375.600 735.600 ;
        RECT 389.100 734.400 390.900 740.400 ;
        RECT 342.000 727.050 342.900 730.800 ;
        RECT 344.100 727.050 345.900 728.850 ;
        RECT 350.100 727.050 351.900 728.850 ;
        RECT 365.100 727.050 366.900 728.850 ;
        RECT 371.250 727.050 373.050 728.850 ;
        RECT 374.700 727.050 375.600 734.400 ;
        RECT 389.700 732.300 390.900 734.400 ;
        RECT 392.100 735.300 393.900 740.400 ;
        RECT 395.100 736.200 396.900 741.000 ;
        RECT 398.100 735.300 399.900 740.400 ;
        RECT 392.100 733.950 399.900 735.300 ;
        RECT 389.700 731.400 393.300 732.300 ;
        RECT 418.500 732.000 420.300 740.400 ;
        RECT 389.100 727.050 390.900 728.850 ;
        RECT 392.100 727.050 393.300 731.400 ;
        RECT 417.000 730.800 420.300 732.000 ;
        RECT 425.100 731.400 426.900 741.000 ;
        RECT 440.700 737.400 442.500 741.000 ;
        RECT 443.700 735.600 445.500 740.400 ;
        RECT 440.400 734.400 445.500 735.600 ;
        RECT 448.200 734.400 450.000 741.000 ;
        RECT 395.100 727.050 396.900 728.850 ;
        RECT 417.000 727.050 417.900 730.800 ;
        RECT 419.100 727.050 420.900 728.850 ;
        RECT 425.100 727.050 426.900 728.850 ;
        RECT 440.400 727.050 441.300 734.400 ;
        RECT 445.950 732.450 448.050 733.200 ;
        RECT 460.950 732.450 463.050 733.050 ;
        RECT 445.950 731.550 463.050 732.450 ;
        RECT 466.500 732.000 468.300 740.400 ;
        RECT 445.950 731.100 448.050 731.550 ;
        RECT 460.950 730.950 463.050 731.550 ;
        RECT 465.000 730.800 468.300 732.000 ;
        RECT 473.100 731.400 474.900 741.000 ;
        RECT 488.100 735.300 489.900 740.400 ;
        RECT 491.100 736.200 492.900 741.000 ;
        RECT 494.100 735.300 495.900 740.400 ;
        RECT 488.100 733.950 495.900 735.300 ;
        RECT 497.100 734.400 498.900 740.400 ;
        RECT 512.100 737.400 513.900 740.400 ;
        RECT 515.100 737.400 516.900 741.000 ;
        RECT 497.100 732.300 498.300 734.400 ;
        RECT 494.700 731.400 498.300 732.300 ;
        RECT 442.950 727.050 444.750 728.850 ;
        RECT 449.100 727.050 450.900 728.850 ;
        RECT 465.000 727.050 465.900 730.800 ;
        RECT 467.100 727.050 468.900 728.850 ;
        RECT 473.100 727.050 474.900 728.850 ;
        RECT 491.100 727.050 492.900 728.850 ;
        RECT 494.700 727.050 495.900 731.400 ;
        RECT 497.100 727.050 498.900 728.850 ;
        RECT 512.700 727.050 513.900 737.400 ;
        RECT 531.000 734.400 532.800 741.000 ;
        RECT 535.500 735.600 537.300 740.400 ;
        RECT 538.500 737.400 540.300 741.000 ;
        RECT 535.500 734.400 540.600 735.600 ;
        RECT 554.100 734.400 555.900 740.400 ;
        RECT 525.000 729.450 529.050 730.050 ;
        RECT 524.550 727.950 529.050 729.450 ;
        RECT 70.950 724.950 73.050 727.050 ;
        RECT 73.950 724.950 76.050 727.050 ;
        RECT 76.950 724.950 79.050 727.050 ;
        RECT 79.950 724.950 82.050 727.050 ;
        RECT 94.950 724.950 97.050 727.050 ;
        RECT 97.950 724.950 100.050 727.050 ;
        RECT 100.950 724.950 103.050 727.050 ;
        RECT 103.950 724.950 106.050 727.050 ;
        RECT 121.950 724.950 124.050 727.050 ;
        RECT 124.950 724.950 127.050 727.050 ;
        RECT 127.950 724.950 130.050 727.050 ;
        RECT 142.950 724.950 145.050 727.050 ;
        RECT 145.950 724.950 148.050 727.050 ;
        RECT 148.950 724.950 151.050 727.050 ;
        RECT 151.950 724.950 154.050 727.050 ;
        RECT 169.950 724.950 172.050 727.050 ;
        RECT 172.950 724.950 175.050 727.050 ;
        RECT 175.950 724.950 178.050 727.050 ;
        RECT 178.950 724.950 181.050 727.050 ;
        RECT 193.950 724.950 196.050 727.050 ;
        RECT 196.950 724.950 199.050 727.050 ;
        RECT 199.950 724.950 202.050 727.050 ;
        RECT 214.950 724.950 217.050 727.050 ;
        RECT 217.950 724.950 220.050 727.050 ;
        RECT 220.950 724.950 223.050 727.050 ;
        RECT 223.950 724.950 226.050 727.050 ;
        RECT 226.950 724.950 229.050 727.050 ;
        RECT 241.950 724.950 244.050 727.050 ;
        RECT 244.950 724.950 247.050 727.050 ;
        RECT 247.950 724.950 250.050 727.050 ;
        RECT 250.950 724.950 253.050 727.050 ;
        RECT 265.950 724.950 268.050 727.050 ;
        RECT 268.950 724.950 271.050 727.050 ;
        RECT 271.950 724.950 274.050 727.050 ;
        RECT 274.950 724.950 277.050 727.050 ;
        RECT 289.950 724.950 292.050 727.050 ;
        RECT 292.950 724.950 295.050 727.050 ;
        RECT 295.950 724.950 298.050 727.050 ;
        RECT 298.950 724.950 301.050 727.050 ;
        RECT 316.950 724.950 319.050 727.050 ;
        RECT 319.950 724.950 322.050 727.050 ;
        RECT 322.950 724.950 325.050 727.050 ;
        RECT 325.950 724.950 328.050 727.050 ;
        RECT 340.950 724.950 343.050 727.050 ;
        RECT 343.950 724.950 346.050 727.050 ;
        RECT 346.950 724.950 349.050 727.050 ;
        RECT 349.950 724.950 352.050 727.050 ;
        RECT 364.950 724.950 367.050 727.050 ;
        RECT 367.950 724.950 370.050 727.050 ;
        RECT 370.950 724.950 373.050 727.050 ;
        RECT 373.950 724.950 376.050 727.050 ;
        RECT 388.950 724.950 391.050 727.050 ;
        RECT 391.950 724.950 394.050 727.050 ;
        RECT 394.950 724.950 397.050 727.050 ;
        RECT 397.950 724.950 400.050 727.050 ;
        RECT 415.950 724.950 418.050 727.050 ;
        RECT 418.950 724.950 421.050 727.050 ;
        RECT 421.950 724.950 424.050 727.050 ;
        RECT 424.950 724.950 427.050 727.050 ;
        RECT 439.950 724.950 442.050 727.050 ;
        RECT 442.950 724.950 445.050 727.050 ;
        RECT 445.950 724.950 448.050 727.050 ;
        RECT 448.950 724.950 451.050 727.050 ;
        RECT 463.950 724.950 466.050 727.050 ;
        RECT 466.950 724.950 469.050 727.050 ;
        RECT 469.950 724.950 472.050 727.050 ;
        RECT 472.950 724.950 475.050 727.050 ;
        RECT 487.950 724.950 490.050 727.050 ;
        RECT 490.950 724.950 493.050 727.050 ;
        RECT 493.950 724.950 496.050 727.050 ;
        RECT 496.950 724.950 499.050 727.050 ;
        RECT 511.950 724.950 514.050 727.050 ;
        RECT 514.950 724.950 517.050 727.050 ;
        RECT 74.100 723.150 75.900 724.950 ;
        RECT 45.750 719.100 57.450 719.700 ;
        RECT 23.550 705.600 25.350 717.600 ;
        RECT 26.550 705.000 28.350 717.600 ;
        RECT 32.250 717.300 37.050 718.200 ;
        RECT 39.150 718.500 57.450 719.100 ;
        RECT 39.150 718.200 47.550 718.500 ;
        RECT 32.250 716.400 33.450 717.300 ;
        RECT 30.450 714.600 33.450 716.400 ;
        RECT 34.350 716.100 36.150 716.400 ;
        RECT 39.150 716.100 40.050 718.200 ;
        RECT 56.550 717.600 57.450 718.500 ;
        RECT 34.350 715.200 40.050 716.100 ;
        RECT 40.950 716.700 42.750 717.300 ;
        RECT 40.950 715.500 48.750 716.700 ;
        RECT 34.350 714.600 36.150 715.200 ;
        RECT 46.650 714.600 48.750 715.500 ;
        RECT 31.350 711.600 33.450 713.700 ;
        RECT 37.950 713.550 39.750 714.300 ;
        RECT 42.750 713.550 44.550 714.300 ;
        RECT 37.950 712.500 44.550 713.550 ;
        RECT 31.350 705.600 33.150 711.600 ;
        RECT 35.850 705.000 37.650 711.600 ;
        RECT 38.850 705.600 40.650 712.500 ;
        RECT 41.850 705.000 43.650 711.600 ;
        RECT 46.650 705.600 48.450 714.600 ;
        RECT 52.050 705.000 53.850 717.600 ;
        RECT 55.050 715.800 57.450 717.600 ;
        RECT 55.050 705.600 56.850 715.800 ;
        RECT 80.100 712.800 81.000 724.950 ;
        RECT 98.250 723.150 100.050 724.950 ;
        RECT 82.950 720.450 85.050 721.050 ;
        RECT 100.950 720.450 103.050 721.050 ;
        RECT 82.950 719.550 103.050 720.450 ;
        RECT 82.950 718.950 85.050 719.550 ;
        RECT 100.950 718.950 103.050 719.550 ;
        RECT 104.700 717.600 105.600 724.950 ;
        RECT 74.400 711.900 81.000 712.800 ;
        RECT 74.400 711.600 75.900 711.900 ;
        RECT 71.100 705.000 72.900 711.600 ;
        RECT 74.100 705.600 75.900 711.600 ;
        RECT 80.100 711.600 81.000 711.900 ;
        RECT 95.100 716.700 102.900 717.600 ;
        RECT 77.100 705.000 78.900 711.000 ;
        RECT 80.100 705.600 81.900 711.600 ;
        RECT 95.100 705.600 96.900 716.700 ;
        RECT 98.100 705.000 99.900 715.800 ;
        RECT 101.100 705.600 102.900 716.700 ;
        RECT 104.100 705.600 105.900 717.600 ;
        RECT 125.700 711.600 126.900 724.950 ;
        RECT 146.100 723.150 147.900 724.950 ;
        RECT 152.100 712.800 153.000 724.950 ;
        RECT 170.400 717.600 171.300 724.950 ;
        RECT 175.950 723.150 177.750 724.950 ;
        RECT 146.400 711.900 153.000 712.800 ;
        RECT 146.400 711.600 147.900 711.900 ;
        RECT 122.100 705.000 123.900 711.600 ;
        RECT 125.100 705.600 126.900 711.600 ;
        RECT 128.100 705.000 129.900 711.600 ;
        RECT 143.100 705.000 144.900 711.600 ;
        RECT 146.100 705.600 147.900 711.600 ;
        RECT 152.100 711.600 153.000 711.900 ;
        RECT 149.100 705.000 150.900 711.000 ;
        RECT 152.100 705.600 153.900 711.600 ;
        RECT 170.100 705.600 171.900 717.600 ;
        RECT 173.100 716.700 180.900 717.600 ;
        RECT 173.100 705.600 174.900 716.700 ;
        RECT 176.100 705.000 177.900 715.800 ;
        RECT 179.100 705.600 180.900 716.700 ;
        RECT 197.700 711.600 198.900 724.950 ;
        RECT 218.250 723.150 220.050 724.950 ;
        RECT 221.100 719.400 222.000 724.950 ;
        RECT 224.100 723.150 225.900 724.950 ;
        RECT 242.100 723.150 243.900 724.950 ;
        RECT 226.950 720.450 229.050 721.050 ;
        RECT 235.950 720.450 238.050 721.050 ;
        RECT 226.950 719.550 238.050 720.450 ;
        RECT 221.100 718.500 225.900 719.400 ;
        RECT 226.950 718.950 229.050 719.550 ;
        RECT 235.950 718.950 238.050 719.550 ;
        RECT 215.100 716.400 222.900 717.300 ;
        RECT 194.100 705.000 195.900 711.600 ;
        RECT 197.100 705.600 198.900 711.600 ;
        RECT 200.100 705.000 201.900 711.600 ;
        RECT 215.100 705.600 216.900 716.400 ;
        RECT 218.100 705.000 219.900 715.500 ;
        RECT 221.100 706.500 222.900 716.400 ;
        RECT 224.100 707.400 225.900 718.500 ;
        RECT 248.700 717.600 249.900 724.950 ;
        RECT 266.100 723.150 267.900 724.950 ;
        RECT 272.700 717.600 273.900 724.950 ;
        RECT 290.100 723.150 291.900 724.950 ;
        RECT 296.700 717.600 297.900 724.950 ;
        RECT 320.100 723.150 321.900 724.950 ;
        RECT 227.100 706.500 228.900 717.600 ;
        RECT 221.100 705.600 228.900 706.500 ;
        RECT 242.400 705.000 244.200 717.600 ;
        RECT 247.500 716.100 249.900 717.600 ;
        RECT 247.500 705.600 249.300 716.100 ;
        RECT 250.200 713.100 252.000 714.900 ;
        RECT 250.500 705.000 252.300 711.600 ;
        RECT 266.400 705.000 268.200 717.600 ;
        RECT 271.500 716.100 273.900 717.600 ;
        RECT 271.500 705.600 273.300 716.100 ;
        RECT 274.200 713.100 276.000 714.900 ;
        RECT 274.500 705.000 276.300 711.600 ;
        RECT 290.400 705.000 292.200 717.600 ;
        RECT 295.500 716.100 297.900 717.600 ;
        RECT 295.500 705.600 297.300 716.100 ;
        RECT 298.200 713.100 300.000 714.900 ;
        RECT 326.100 712.800 327.000 724.950 ;
        RECT 320.400 711.900 327.000 712.800 ;
        RECT 320.400 711.600 321.900 711.900 ;
        RECT 298.500 705.000 300.300 711.600 ;
        RECT 317.100 705.000 318.900 711.600 ;
        RECT 320.100 705.600 321.900 711.600 ;
        RECT 326.100 711.600 327.000 711.900 ;
        RECT 342.000 712.800 342.900 724.950 ;
        RECT 347.100 723.150 348.900 724.950 ;
        RECT 368.250 723.150 370.050 724.950 ;
        RECT 343.950 720.450 346.050 721.050 ;
        RECT 364.950 720.450 367.050 721.050 ;
        RECT 343.950 719.550 367.050 720.450 ;
        RECT 343.950 718.950 346.050 719.550 ;
        RECT 364.950 718.950 367.050 719.550 ;
        RECT 374.700 717.600 375.600 724.950 ;
        RECT 392.100 717.600 393.300 724.950 ;
        RECT 398.100 723.150 399.900 724.950 ;
        RECT 406.950 723.450 409.050 724.050 ;
        RECT 412.950 723.450 415.050 724.050 ;
        RECT 406.950 722.550 415.050 723.450 ;
        RECT 406.950 721.950 409.050 722.550 ;
        RECT 412.950 721.950 415.050 722.550 ;
        RECT 365.100 716.700 372.900 717.600 ;
        RECT 342.000 711.900 348.600 712.800 ;
        RECT 342.000 711.600 342.900 711.900 ;
        RECT 323.100 705.000 324.900 711.000 ;
        RECT 326.100 705.600 327.900 711.600 ;
        RECT 341.100 705.600 342.900 711.600 ;
        RECT 347.100 711.600 348.600 711.900 ;
        RECT 344.100 705.000 345.900 711.000 ;
        RECT 347.100 705.600 348.900 711.600 ;
        RECT 350.100 705.000 351.900 711.600 ;
        RECT 365.100 705.600 366.900 716.700 ;
        RECT 368.100 705.000 369.900 715.800 ;
        RECT 371.100 705.600 372.900 716.700 ;
        RECT 374.100 705.600 375.900 717.600 ;
        RECT 392.100 716.100 394.500 717.600 ;
        RECT 390.000 713.100 391.800 714.900 ;
        RECT 389.700 705.000 391.500 711.600 ;
        RECT 392.700 705.600 394.500 716.100 ;
        RECT 397.800 705.000 399.600 717.600 ;
        RECT 417.000 712.800 417.900 724.950 ;
        RECT 422.100 723.150 423.900 724.950 ;
        RECT 440.400 717.600 441.300 724.950 ;
        RECT 445.950 723.150 447.750 724.950 ;
        RECT 417.000 711.900 423.600 712.800 ;
        RECT 417.000 711.600 417.900 711.900 ;
        RECT 416.100 705.600 417.900 711.600 ;
        RECT 422.100 711.600 423.600 711.900 ;
        RECT 419.100 705.000 420.900 711.000 ;
        RECT 422.100 705.600 423.900 711.600 ;
        RECT 425.100 705.000 426.900 711.600 ;
        RECT 440.100 705.600 441.900 717.600 ;
        RECT 443.100 716.700 450.900 717.600 ;
        RECT 443.100 705.600 444.900 716.700 ;
        RECT 446.100 705.000 447.900 715.800 ;
        RECT 449.100 705.600 450.900 716.700 ;
        RECT 465.000 712.800 465.900 724.950 ;
        RECT 470.100 723.150 471.900 724.950 ;
        RECT 488.100 723.150 489.900 724.950 ;
        RECT 494.700 717.600 495.900 724.950 ;
        RECT 465.000 711.900 471.600 712.800 ;
        RECT 465.000 711.600 465.900 711.900 ;
        RECT 464.100 705.600 465.900 711.600 ;
        RECT 470.100 711.600 471.600 711.900 ;
        RECT 467.100 705.000 468.900 711.000 ;
        RECT 470.100 705.600 471.900 711.600 ;
        RECT 473.100 705.000 474.900 711.600 ;
        RECT 488.400 705.000 490.200 717.600 ;
        RECT 493.500 716.100 495.900 717.600 ;
        RECT 493.500 705.600 495.300 716.100 ;
        RECT 496.200 713.100 498.000 714.900 ;
        RECT 512.700 711.600 513.900 724.950 ;
        RECT 515.100 723.150 516.900 724.950 ;
        RECT 524.550 724.050 525.450 727.950 ;
        RECT 530.100 727.050 531.900 728.850 ;
        RECT 536.250 727.050 538.050 728.850 ;
        RECT 539.700 727.050 540.600 734.400 ;
        RECT 554.700 732.300 555.900 734.400 ;
        RECT 557.100 735.300 558.900 740.400 ;
        RECT 560.100 736.200 561.900 741.000 ;
        RECT 563.100 735.300 564.900 740.400 ;
        RECT 578.700 737.400 580.500 741.000 ;
        RECT 581.700 735.600 583.500 740.400 ;
        RECT 557.100 733.950 564.900 735.300 ;
        RECT 578.400 734.400 583.500 735.600 ;
        RECT 586.200 734.400 588.000 741.000 ;
        RECT 554.700 731.400 558.300 732.300 ;
        RECT 554.100 727.050 555.900 728.850 ;
        RECT 557.100 727.050 558.300 731.400 ;
        RECT 560.100 727.050 561.900 728.850 ;
        RECT 578.400 727.050 579.300 734.400 ;
        RECT 583.950 732.450 586.050 733.050 ;
        RECT 595.950 732.450 598.050 733.050 ;
        RECT 583.950 731.550 598.050 732.450 ;
        RECT 583.950 730.950 586.050 731.550 ;
        RECT 595.950 730.950 598.050 731.550 ;
        RECT 602.100 731.400 603.900 741.000 ;
        RECT 608.700 732.000 610.500 740.400 ;
        RECT 626.100 737.400 627.900 741.000 ;
        RECT 629.100 737.400 630.900 740.400 ;
        RECT 644.700 737.400 646.500 741.000 ;
        RECT 608.700 730.800 612.000 732.000 ;
        RECT 580.950 727.050 582.750 728.850 ;
        RECT 587.100 727.050 588.900 728.850 ;
        RECT 602.100 727.050 603.900 728.850 ;
        RECT 608.100 727.050 609.900 728.850 ;
        RECT 611.100 727.050 612.000 730.800 ;
        RECT 629.100 727.050 630.300 737.400 ;
        RECT 647.700 735.600 649.500 740.400 ;
        RECT 644.400 734.400 649.500 735.600 ;
        RECT 652.200 734.400 654.000 741.000 ;
        RECT 668.100 734.400 669.900 740.400 ;
        RECT 644.400 727.050 645.300 734.400 ;
        RECT 668.700 732.300 669.900 734.400 ;
        RECT 671.100 735.300 672.900 740.400 ;
        RECT 674.100 736.200 675.900 741.000 ;
        RECT 677.100 735.300 678.900 740.400 ;
        RECT 671.100 733.950 678.900 735.300 ;
        RECT 692.100 734.400 693.900 740.400 ;
        RECT 692.700 732.300 693.900 734.400 ;
        RECT 695.100 735.300 696.900 740.400 ;
        RECT 698.100 736.200 699.900 741.000 ;
        RECT 701.100 735.300 702.900 740.400 ;
        RECT 695.100 733.950 702.900 735.300 ;
        RECT 668.700 731.400 672.300 732.300 ;
        RECT 692.700 731.400 696.300 732.300 ;
        RECT 718.500 732.000 720.300 740.400 ;
        RECT 646.950 727.050 648.750 728.850 ;
        RECT 653.100 727.050 654.900 728.850 ;
        RECT 668.100 727.050 669.900 728.850 ;
        RECT 671.100 727.050 672.300 731.400 ;
        RECT 687.000 729.450 691.050 730.050 ;
        RECT 674.100 727.050 675.900 728.850 ;
        RECT 686.550 727.950 691.050 729.450 ;
        RECT 529.950 724.950 532.050 727.050 ;
        RECT 532.950 724.950 535.050 727.050 ;
        RECT 535.950 724.950 538.050 727.050 ;
        RECT 538.950 724.950 541.050 727.050 ;
        RECT 553.950 724.950 556.050 727.050 ;
        RECT 556.950 724.950 559.050 727.050 ;
        RECT 559.950 724.950 562.050 727.050 ;
        RECT 562.950 724.950 565.050 727.050 ;
        RECT 577.950 724.950 580.050 727.050 ;
        RECT 580.950 724.950 583.050 727.050 ;
        RECT 583.950 724.950 586.050 727.050 ;
        RECT 586.950 724.950 589.050 727.050 ;
        RECT 601.950 724.950 604.050 727.050 ;
        RECT 604.950 724.950 607.050 727.050 ;
        RECT 607.950 724.950 610.050 727.050 ;
        RECT 610.950 724.950 613.050 727.050 ;
        RECT 625.950 724.950 628.050 727.050 ;
        RECT 628.950 724.950 631.050 727.050 ;
        RECT 643.950 724.950 646.050 727.050 ;
        RECT 646.950 724.950 649.050 727.050 ;
        RECT 649.950 724.950 652.050 727.050 ;
        RECT 652.950 724.950 655.050 727.050 ;
        RECT 667.950 724.950 670.050 727.050 ;
        RECT 670.950 724.950 673.050 727.050 ;
        RECT 673.950 724.950 676.050 727.050 ;
        RECT 676.950 724.950 679.050 727.050 ;
        RECT 524.550 722.550 529.050 724.050 ;
        RECT 533.250 723.150 535.050 724.950 ;
        RECT 525.000 721.950 529.050 722.550 ;
        RECT 539.700 717.600 540.600 724.950 ;
        RECT 557.100 717.600 558.300 724.950 ;
        RECT 563.100 723.150 564.900 724.950 ;
        RECT 559.950 720.450 562.050 721.050 ;
        RECT 571.950 720.450 574.050 721.050 ;
        RECT 559.950 719.550 574.050 720.450 ;
        RECT 559.950 718.950 562.050 719.550 ;
        RECT 571.950 718.950 574.050 719.550 ;
        RECT 578.400 717.600 579.300 724.950 ;
        RECT 583.950 723.150 585.750 724.950 ;
        RECT 605.100 723.150 606.900 724.950 ;
        RECT 530.100 716.700 537.900 717.600 ;
        RECT 496.500 705.000 498.300 711.600 ;
        RECT 512.100 705.600 513.900 711.600 ;
        RECT 515.100 705.000 516.900 711.600 ;
        RECT 530.100 705.600 531.900 716.700 ;
        RECT 533.100 705.000 534.900 715.800 ;
        RECT 536.100 705.600 537.900 716.700 ;
        RECT 539.100 705.600 540.900 717.600 ;
        RECT 557.100 716.100 559.500 717.600 ;
        RECT 555.000 713.100 556.800 714.900 ;
        RECT 554.700 705.000 556.500 711.600 ;
        RECT 557.700 705.600 559.500 716.100 ;
        RECT 562.800 705.000 564.600 717.600 ;
        RECT 578.100 705.600 579.900 717.600 ;
        RECT 581.100 716.700 588.900 717.600 ;
        RECT 581.100 705.600 582.900 716.700 ;
        RECT 584.100 705.000 585.900 715.800 ;
        RECT 587.100 705.600 588.900 716.700 ;
        RECT 611.100 712.800 612.000 724.950 ;
        RECT 626.100 723.150 627.900 724.950 ;
        RECT 605.400 711.900 612.000 712.800 ;
        RECT 605.400 711.600 606.900 711.900 ;
        RECT 602.100 705.000 603.900 711.600 ;
        RECT 605.100 705.600 606.900 711.600 ;
        RECT 611.100 711.600 612.000 711.900 ;
        RECT 629.100 711.600 630.300 724.950 ;
        RECT 644.400 717.600 645.300 724.950 ;
        RECT 649.950 723.150 651.750 724.950 ;
        RECT 671.100 717.600 672.300 724.950 ;
        RECT 677.100 723.150 678.900 724.950 ;
        RECT 686.550 724.050 687.450 727.950 ;
        RECT 692.100 727.050 693.900 728.850 ;
        RECT 695.100 727.050 696.300 731.400 ;
        RECT 717.000 730.800 720.300 732.000 ;
        RECT 725.100 731.400 726.900 741.000 ;
        RECT 745.500 732.000 747.300 740.400 ;
        RECT 744.000 730.800 747.300 732.000 ;
        RECT 752.100 731.400 753.900 741.000 ;
        RECT 770.100 734.400 771.900 740.400 ;
        RECT 770.700 732.300 771.900 734.400 ;
        RECT 773.100 735.300 774.900 740.400 ;
        RECT 776.100 736.200 777.900 741.000 ;
        RECT 779.100 735.300 780.900 740.400 ;
        RECT 794.700 737.400 796.500 741.000 ;
        RECT 797.700 735.600 799.500 740.400 ;
        RECT 773.100 733.950 780.900 735.300 ;
        RECT 794.400 734.400 799.500 735.600 ;
        RECT 802.200 734.400 804.000 741.000 ;
        RECT 770.700 731.400 774.300 732.300 ;
        RECT 698.100 727.050 699.900 728.850 ;
        RECT 717.000 727.050 717.900 730.800 ;
        RECT 738.000 729.450 742.050 730.050 ;
        RECT 719.100 727.050 720.900 728.850 ;
        RECT 725.100 727.050 726.900 728.850 ;
        RECT 737.550 727.950 742.050 729.450 ;
        RECT 691.950 724.950 694.050 727.050 ;
        RECT 694.950 724.950 697.050 727.050 ;
        RECT 697.950 724.950 700.050 727.050 ;
        RECT 700.950 724.950 703.050 727.050 ;
        RECT 715.950 724.950 718.050 727.050 ;
        RECT 718.950 724.950 721.050 727.050 ;
        RECT 721.950 724.950 724.050 727.050 ;
        RECT 724.950 724.950 727.050 727.050 ;
        RECT 686.550 722.550 691.050 724.050 ;
        RECT 687.000 721.950 691.050 722.550 ;
        RECT 673.950 720.450 676.050 721.050 ;
        RECT 685.950 720.450 688.050 721.050 ;
        RECT 673.950 719.550 688.050 720.450 ;
        RECT 673.950 718.950 676.050 719.550 ;
        RECT 685.950 718.950 688.050 719.550 ;
        RECT 695.100 717.600 696.300 724.950 ;
        RECT 701.100 723.150 702.900 724.950 ;
        RECT 608.100 705.000 609.900 711.000 ;
        RECT 611.100 705.600 612.900 711.600 ;
        RECT 626.100 705.000 627.900 711.600 ;
        RECT 629.100 705.600 630.900 711.600 ;
        RECT 644.100 705.600 645.900 717.600 ;
        RECT 647.100 716.700 654.900 717.600 ;
        RECT 647.100 705.600 648.900 716.700 ;
        RECT 650.100 705.000 651.900 715.800 ;
        RECT 653.100 705.600 654.900 716.700 ;
        RECT 671.100 716.100 673.500 717.600 ;
        RECT 669.000 713.100 670.800 714.900 ;
        RECT 668.700 705.000 670.500 711.600 ;
        RECT 671.700 705.600 673.500 716.100 ;
        RECT 676.800 705.000 678.600 717.600 ;
        RECT 695.100 716.100 697.500 717.600 ;
        RECT 693.000 713.100 694.800 714.900 ;
        RECT 692.700 705.000 694.500 711.600 ;
        RECT 695.700 705.600 697.500 716.100 ;
        RECT 700.800 705.000 702.600 717.600 ;
        RECT 717.000 712.800 717.900 724.950 ;
        RECT 722.100 723.150 723.900 724.950 ;
        RECT 737.550 724.050 738.450 727.950 ;
        RECT 744.000 727.050 744.900 730.800 ;
        RECT 746.100 727.050 747.900 728.850 ;
        RECT 752.100 727.050 753.900 728.850 ;
        RECT 770.100 727.050 771.900 728.850 ;
        RECT 773.100 727.050 774.300 731.400 ;
        RECT 781.950 729.450 784.050 733.050 ;
        RECT 781.950 729.000 786.450 729.450 ;
        RECT 776.100 727.050 777.900 728.850 ;
        RECT 782.550 728.550 786.450 729.000 ;
        RECT 742.950 724.950 745.050 727.050 ;
        RECT 745.950 724.950 748.050 727.050 ;
        RECT 748.950 724.950 751.050 727.050 ;
        RECT 751.950 724.950 754.050 727.050 ;
        RECT 769.950 724.950 772.050 727.050 ;
        RECT 772.950 724.950 775.050 727.050 ;
        RECT 775.950 724.950 778.050 727.050 ;
        RECT 778.950 724.950 781.050 727.050 ;
        RECT 737.550 722.550 742.050 724.050 ;
        RECT 738.000 721.950 742.050 722.550 ;
        RECT 744.000 712.800 744.900 724.950 ;
        RECT 749.100 723.150 750.900 724.950 ;
        RECT 745.950 720.450 748.050 721.050 ;
        RECT 769.950 720.450 772.050 721.050 ;
        RECT 745.950 719.550 772.050 720.450 ;
        RECT 745.950 718.950 748.050 719.550 ;
        RECT 769.950 718.950 772.050 719.550 ;
        RECT 773.100 717.600 774.300 724.950 ;
        RECT 779.100 723.150 780.900 724.950 ;
        RECT 785.550 724.050 786.450 728.550 ;
        RECT 794.400 727.050 795.300 734.400 ;
        RECT 799.950 732.450 802.050 733.050 ;
        RECT 799.950 731.550 807.450 732.450 ;
        RECT 820.500 732.000 822.300 740.400 ;
        RECT 799.950 730.950 802.050 731.550 ;
        RECT 806.550 729.450 807.450 731.550 ;
        RECT 819.000 730.800 822.300 732.000 ;
        RECT 827.100 731.400 828.900 741.000 ;
        RECT 842.100 735.300 843.900 740.400 ;
        RECT 845.100 736.200 846.900 741.000 ;
        RECT 848.100 735.300 849.900 740.400 ;
        RECT 842.100 733.950 849.900 735.300 ;
        RECT 851.100 734.400 852.900 740.400 ;
        RECT 851.100 732.300 852.300 734.400 ;
        RECT 848.700 731.400 852.300 732.300 ;
        RECT 868.500 732.000 870.300 740.400 ;
        RECT 796.950 727.050 798.750 728.850 ;
        RECT 803.100 727.050 804.900 728.850 ;
        RECT 806.550 728.550 810.450 729.450 ;
        RECT 793.950 724.950 796.050 727.050 ;
        RECT 796.950 724.950 799.050 727.050 ;
        RECT 799.950 724.950 802.050 727.050 ;
        RECT 802.950 724.950 805.050 727.050 ;
        RECT 781.950 722.550 786.450 724.050 ;
        RECT 781.950 721.950 786.000 722.550 ;
        RECT 794.400 717.600 795.300 724.950 ;
        RECT 799.950 723.150 801.750 724.950 ;
        RECT 809.550 723.450 810.450 728.550 ;
        RECT 819.000 727.050 819.900 730.800 ;
        RECT 837.000 729.450 841.050 730.050 ;
        RECT 821.100 727.050 822.900 728.850 ;
        RECT 827.100 727.050 828.900 728.850 ;
        RECT 836.550 727.950 841.050 729.450 ;
        RECT 817.950 724.950 820.050 727.050 ;
        RECT 820.950 724.950 823.050 727.050 ;
        RECT 823.950 724.950 826.050 727.050 ;
        RECT 826.950 724.950 829.050 727.050 ;
        RECT 814.950 723.450 817.050 724.050 ;
        RECT 809.550 722.550 817.050 723.450 ;
        RECT 814.950 721.950 817.050 722.550 ;
        RECT 773.100 716.100 775.500 717.600 ;
        RECT 771.000 713.100 772.800 714.900 ;
        RECT 717.000 711.900 723.600 712.800 ;
        RECT 717.000 711.600 717.900 711.900 ;
        RECT 716.100 705.600 717.900 711.600 ;
        RECT 722.100 711.600 723.600 711.900 ;
        RECT 744.000 711.900 750.600 712.800 ;
        RECT 744.000 711.600 744.900 711.900 ;
        RECT 719.100 705.000 720.900 711.000 ;
        RECT 722.100 705.600 723.900 711.600 ;
        RECT 725.100 705.000 726.900 711.600 ;
        RECT 743.100 705.600 744.900 711.600 ;
        RECT 749.100 711.600 750.600 711.900 ;
        RECT 746.100 705.000 747.900 711.000 ;
        RECT 749.100 705.600 750.900 711.600 ;
        RECT 752.100 705.000 753.900 711.600 ;
        RECT 770.700 705.000 772.500 711.600 ;
        RECT 773.700 705.600 775.500 716.100 ;
        RECT 778.800 705.000 780.600 717.600 ;
        RECT 794.100 705.600 795.900 717.600 ;
        RECT 797.100 716.700 804.900 717.600 ;
        RECT 797.100 705.600 798.900 716.700 ;
        RECT 800.100 705.000 801.900 715.800 ;
        RECT 803.100 705.600 804.900 716.700 ;
        RECT 819.000 712.800 819.900 724.950 ;
        RECT 824.100 723.150 825.900 724.950 ;
        RECT 836.550 723.450 837.450 727.950 ;
        RECT 845.100 727.050 846.900 728.850 ;
        RECT 848.700 727.050 849.900 731.400 ;
        RECT 867.000 730.800 870.300 732.000 ;
        RECT 875.100 731.400 876.900 741.000 ;
        RECT 893.100 737.400 894.900 740.400 ;
        RECT 896.100 737.400 897.900 741.000 ;
        RECT 851.100 727.050 852.900 728.850 ;
        RECT 867.000 727.050 867.900 730.800 ;
        RECT 869.100 727.050 870.900 728.850 ;
        RECT 875.100 727.050 876.900 728.850 ;
        RECT 893.700 727.050 894.900 737.400 ;
        RECT 841.950 724.950 844.050 727.050 ;
        RECT 844.950 724.950 847.050 727.050 ;
        RECT 847.950 724.950 850.050 727.050 ;
        RECT 850.950 724.950 853.050 727.050 ;
        RECT 865.950 724.950 868.050 727.050 ;
        RECT 868.950 724.950 871.050 727.050 ;
        RECT 871.950 724.950 874.050 727.050 ;
        RECT 874.950 724.950 877.050 727.050 ;
        RECT 892.950 724.950 895.050 727.050 ;
        RECT 895.950 724.950 898.050 727.050 ;
        RECT 830.550 722.550 837.450 723.450 ;
        RECT 842.100 723.150 843.900 724.950 ;
        RECT 820.950 720.450 823.050 721.050 ;
        RECT 830.550 720.450 831.450 722.550 ;
        RECT 820.950 719.550 831.450 720.450 ;
        RECT 820.950 718.950 823.050 719.550 ;
        RECT 820.950 717.450 823.050 717.900 ;
        RECT 826.950 717.450 829.050 718.050 ;
        RECT 848.700 717.600 849.900 724.950 ;
        RECT 820.950 716.550 829.050 717.450 ;
        RECT 820.950 715.800 823.050 716.550 ;
        RECT 826.950 715.950 829.050 716.550 ;
        RECT 819.000 711.900 825.600 712.800 ;
        RECT 819.000 711.600 819.900 711.900 ;
        RECT 818.100 705.600 819.900 711.600 ;
        RECT 824.100 711.600 825.600 711.900 ;
        RECT 821.100 705.000 822.900 711.000 ;
        RECT 824.100 705.600 825.900 711.600 ;
        RECT 827.100 705.000 828.900 711.600 ;
        RECT 842.400 705.000 844.200 717.600 ;
        RECT 847.500 716.100 849.900 717.600 ;
        RECT 847.500 705.600 849.300 716.100 ;
        RECT 850.200 713.100 852.000 714.900 ;
        RECT 867.000 712.800 867.900 724.950 ;
        RECT 872.100 723.150 873.900 724.950 ;
        RECT 868.950 720.450 871.050 721.050 ;
        RECT 877.950 720.450 880.050 721.050 ;
        RECT 868.950 719.550 880.050 720.450 ;
        RECT 868.950 718.950 871.050 719.550 ;
        RECT 877.950 718.950 880.050 719.550 ;
        RECT 867.000 711.900 873.600 712.800 ;
        RECT 867.000 711.600 867.900 711.900 ;
        RECT 850.500 705.000 852.300 711.600 ;
        RECT 866.100 705.600 867.900 711.600 ;
        RECT 872.100 711.600 873.600 711.900 ;
        RECT 893.700 711.600 894.900 724.950 ;
        RECT 896.100 723.150 897.900 724.950 ;
        RECT 869.100 705.000 870.900 711.000 ;
        RECT 872.100 705.600 873.900 711.600 ;
        RECT 875.100 705.000 876.900 711.600 ;
        RECT 893.100 705.600 894.900 711.600 ;
        RECT 896.100 705.000 897.900 711.600 ;
        RECT 14.100 690.300 15.900 701.400 ;
        RECT 17.100 691.200 18.900 702.000 ;
        RECT 20.100 690.300 21.900 701.400 ;
        RECT 14.100 689.400 21.900 690.300 ;
        RECT 23.100 689.400 24.900 701.400 ;
        RECT 38.700 695.400 40.500 702.000 ;
        RECT 39.000 692.100 40.800 693.900 ;
        RECT 41.700 690.900 43.500 701.400 ;
        RECT 41.100 689.400 43.500 690.900 ;
        RECT 46.800 689.400 48.600 702.000 ;
        RECT 65.100 695.400 66.900 702.000 ;
        RECT 68.100 695.400 69.900 701.400 ;
        RECT 71.100 695.400 72.900 702.000 ;
        RECT 86.100 695.400 87.900 702.000 ;
        RECT 89.100 695.400 90.900 701.400 ;
        RECT 107.100 695.400 108.900 702.000 ;
        RECT 110.100 695.400 111.900 701.400 ;
        RECT 17.250 682.050 19.050 683.850 ;
        RECT 23.700 682.050 24.600 689.400 ;
        RECT 41.100 682.050 42.300 689.400 ;
        RECT 47.100 682.050 48.900 683.850 ;
        RECT 68.100 682.050 69.300 695.400 ;
        RECT 86.100 682.050 87.900 683.850 ;
        RECT 89.100 682.050 90.300 695.400 ;
        RECT 107.100 682.050 108.900 683.850 ;
        RECT 110.100 682.050 111.300 695.400 ;
        RECT 125.100 689.400 126.900 701.400 ;
        RECT 128.100 690.300 129.900 701.400 ;
        RECT 131.100 691.200 132.900 702.000 ;
        RECT 134.100 690.300 135.900 701.400 ;
        RECT 139.950 699.450 142.050 700.050 ;
        RECT 145.950 699.450 148.050 700.050 ;
        RECT 139.950 698.550 148.050 699.450 ;
        RECT 139.950 697.950 142.050 698.550 ;
        RECT 145.950 697.950 148.050 698.550 ;
        RECT 128.100 689.400 135.900 690.300 ;
        RECT 149.400 689.400 151.200 702.000 ;
        RECT 154.500 690.900 156.300 701.400 ;
        RECT 157.500 695.400 159.300 702.000 ;
        RECT 157.200 692.100 159.000 693.900 ;
        RECT 154.500 689.400 156.900 690.900 ;
        RECT 173.400 689.400 175.200 702.000 ;
        RECT 178.500 690.900 180.300 701.400 ;
        RECT 181.500 695.400 183.300 702.000 ;
        RECT 181.200 692.100 183.000 693.900 ;
        RECT 178.500 689.400 180.900 690.900 ;
        RECT 197.100 689.400 198.900 701.400 ;
        RECT 200.100 690.000 201.900 702.000 ;
        RECT 203.100 695.400 204.900 701.400 ;
        RECT 206.100 695.400 207.900 702.000 ;
        RECT 224.100 695.400 225.900 702.000 ;
        RECT 227.100 695.400 228.900 701.400 ;
        RECT 230.100 696.000 231.900 702.000 ;
        RECT 125.400 682.050 126.300 689.400 ;
        RECT 127.950 687.450 130.050 688.050 ;
        RECT 151.950 687.450 154.050 688.050 ;
        RECT 127.950 686.550 154.050 687.450 ;
        RECT 127.950 685.950 130.050 686.550 ;
        RECT 151.950 685.950 154.050 686.550 ;
        RECT 130.950 682.050 132.750 683.850 ;
        RECT 149.100 682.050 150.900 683.850 ;
        RECT 155.700 682.050 156.900 689.400 ;
        RECT 173.100 682.050 174.900 683.850 ;
        RECT 179.700 682.050 180.900 689.400 ;
        RECT 197.700 682.050 198.600 689.400 ;
        RECT 201.000 682.050 202.800 683.850 ;
        RECT 13.950 679.950 16.050 682.050 ;
        RECT 16.950 679.950 19.050 682.050 ;
        RECT 19.950 679.950 22.050 682.050 ;
        RECT 22.950 679.950 25.050 682.050 ;
        RECT 37.950 679.950 40.050 682.050 ;
        RECT 40.950 679.950 43.050 682.050 ;
        RECT 43.950 679.950 46.050 682.050 ;
        RECT 46.950 679.950 49.050 682.050 ;
        RECT 64.950 679.950 67.050 682.050 ;
        RECT 67.950 679.950 70.050 682.050 ;
        RECT 70.950 679.950 73.050 682.050 ;
        RECT 85.950 679.950 88.050 682.050 ;
        RECT 88.950 679.950 91.050 682.050 ;
        RECT 106.950 679.950 109.050 682.050 ;
        RECT 109.950 679.950 112.050 682.050 ;
        RECT 124.950 679.950 127.050 682.050 ;
        RECT 127.950 679.950 130.050 682.050 ;
        RECT 130.950 679.950 133.050 682.050 ;
        RECT 133.950 679.950 136.050 682.050 ;
        RECT 148.950 679.950 151.050 682.050 ;
        RECT 151.950 679.950 154.050 682.050 ;
        RECT 154.950 679.950 157.050 682.050 ;
        RECT 157.950 679.950 160.050 682.050 ;
        RECT 172.950 679.950 175.050 682.050 ;
        RECT 175.950 679.950 178.050 682.050 ;
        RECT 178.950 679.950 181.050 682.050 ;
        RECT 181.950 679.950 184.050 682.050 ;
        RECT 193.950 681.450 196.050 682.050 ;
        RECT 188.550 680.550 196.050 681.450 ;
        RECT 14.100 678.150 15.900 679.950 ;
        RECT 20.250 678.150 22.050 679.950 ;
        RECT 23.700 672.600 24.600 679.950 ;
        RECT 38.100 678.150 39.900 679.950 ;
        RECT 41.100 675.600 42.300 679.950 ;
        RECT 44.100 678.150 45.900 679.950 ;
        RECT 65.250 678.150 67.050 679.950 ;
        RECT 38.700 674.700 42.300 675.600 ;
        RECT 68.100 674.700 69.300 679.950 ;
        RECT 71.100 678.150 72.900 679.950 ;
        RECT 38.700 672.600 39.900 674.700 ;
        RECT 68.100 673.800 72.300 674.700 ;
        RECT 15.000 666.000 16.800 672.600 ;
        RECT 19.500 671.400 24.600 672.600 ;
        RECT 19.500 666.600 21.300 671.400 ;
        RECT 22.500 666.000 24.300 669.600 ;
        RECT 25.950 669.450 28.050 670.050 ;
        RECT 31.950 669.450 34.050 670.050 ;
        RECT 25.950 668.550 34.050 669.450 ;
        RECT 25.950 667.950 28.050 668.550 ;
        RECT 31.950 667.950 34.050 668.550 ;
        RECT 38.100 666.600 39.900 672.600 ;
        RECT 41.100 671.700 48.900 673.050 ;
        RECT 41.100 666.600 42.900 671.700 ;
        RECT 44.100 666.000 45.900 670.800 ;
        RECT 47.100 666.600 48.900 671.700 ;
        RECT 65.400 666.000 67.200 672.600 ;
        RECT 70.500 666.600 72.300 673.800 ;
        RECT 89.100 669.600 90.300 679.950 ;
        RECT 110.100 669.600 111.300 679.950 ;
        RECT 125.400 672.600 126.300 679.950 ;
        RECT 127.950 678.150 129.750 679.950 ;
        RECT 134.100 678.150 135.900 679.950 ;
        RECT 152.100 678.150 153.900 679.950 ;
        RECT 155.700 675.600 156.900 679.950 ;
        RECT 158.100 678.150 159.900 679.950 ;
        RECT 176.100 678.150 177.900 679.950 ;
        RECT 179.700 675.600 180.900 679.950 ;
        RECT 182.100 678.150 183.900 679.950 ;
        RECT 188.550 679.050 189.450 680.550 ;
        RECT 193.950 679.950 196.050 680.550 ;
        RECT 197.100 679.950 199.200 682.050 ;
        RECT 200.400 679.950 202.500 682.050 ;
        RECT 184.950 677.550 189.450 679.050 ;
        RECT 184.950 676.950 189.000 677.550 ;
        RECT 155.700 674.700 159.300 675.600 ;
        RECT 179.700 674.700 183.300 675.600 ;
        RECT 125.400 671.400 130.500 672.600 ;
        RECT 86.100 666.000 87.900 669.600 ;
        RECT 89.100 666.600 90.900 669.600 ;
        RECT 107.100 666.000 108.900 669.600 ;
        RECT 110.100 666.600 111.900 669.600 ;
        RECT 125.700 666.000 127.500 669.600 ;
        RECT 128.700 666.600 130.500 671.400 ;
        RECT 133.200 666.000 135.000 672.600 ;
        RECT 149.100 671.700 156.900 673.050 ;
        RECT 149.100 666.600 150.900 671.700 ;
        RECT 152.100 666.000 153.900 670.800 ;
        RECT 155.100 666.600 156.900 671.700 ;
        RECT 158.100 672.600 159.300 674.700 ;
        RECT 158.100 666.600 159.900 672.600 ;
        RECT 173.100 671.700 180.900 673.050 ;
        RECT 173.100 666.600 174.900 671.700 ;
        RECT 176.100 666.000 177.900 670.800 ;
        RECT 179.100 666.600 180.900 671.700 ;
        RECT 182.100 672.600 183.300 674.700 ;
        RECT 197.700 672.600 198.600 679.950 ;
        RECT 204.000 675.300 204.900 695.400 ;
        RECT 227.400 695.100 228.900 695.400 ;
        RECT 233.100 695.400 234.900 701.400 ;
        RECT 233.100 695.100 234.000 695.400 ;
        RECT 227.400 694.200 234.000 695.100 ;
        RECT 227.100 682.050 228.900 683.850 ;
        RECT 233.100 682.050 234.000 694.200 ;
        RECT 248.100 690.300 249.900 701.400 ;
        RECT 251.100 691.200 252.900 702.000 ;
        RECT 254.100 690.300 255.900 701.400 ;
        RECT 248.100 689.400 255.900 690.300 ;
        RECT 257.100 689.400 258.900 701.400 ;
        RECT 272.100 695.400 273.900 701.400 ;
        RECT 251.250 682.050 253.050 683.850 ;
        RECT 257.700 682.050 258.600 689.400 ;
        RECT 272.100 688.500 273.300 695.400 ;
        RECT 275.100 691.200 276.900 702.000 ;
        RECT 278.100 689.400 279.900 701.400 ;
        RECT 296.700 695.400 298.500 702.000 ;
        RECT 297.000 692.100 298.800 693.900 ;
        RECT 299.700 690.900 301.500 701.400 ;
        RECT 272.100 687.600 277.800 688.500 ;
        RECT 276.000 686.700 277.800 687.600 ;
        RECT 272.400 682.050 274.200 683.850 ;
        RECT 205.800 679.950 207.900 682.050 ;
        RECT 223.950 679.950 226.050 682.050 ;
        RECT 226.950 679.950 229.050 682.050 ;
        RECT 229.950 679.950 232.050 682.050 ;
        RECT 232.950 679.950 235.050 682.050 ;
        RECT 247.950 679.950 250.050 682.050 ;
        RECT 250.950 679.950 253.050 682.050 ;
        RECT 253.950 679.950 256.050 682.050 ;
        RECT 256.950 679.950 259.050 682.050 ;
        RECT 272.400 679.950 274.500 682.050 ;
        RECT 205.950 678.150 207.750 679.950 ;
        RECT 224.100 678.150 225.900 679.950 ;
        RECT 230.100 678.150 231.900 679.950 ;
        RECT 233.100 676.200 234.000 679.950 ;
        RECT 248.100 678.150 249.900 679.950 ;
        RECT 254.250 678.150 256.050 679.950 ;
        RECT 199.500 674.400 207.900 675.300 ;
        RECT 199.500 673.500 201.300 674.400 ;
        RECT 182.100 666.600 183.900 672.600 ;
        RECT 197.700 670.800 200.400 672.600 ;
        RECT 198.600 666.600 200.400 670.800 ;
        RECT 201.600 666.000 203.400 672.600 ;
        RECT 206.100 666.600 207.900 674.400 ;
        RECT 224.100 666.000 225.900 675.600 ;
        RECT 230.700 675.000 234.000 676.200 ;
        RECT 230.700 666.600 232.500 675.000 ;
        RECT 257.700 672.600 258.600 679.950 ;
        RECT 276.000 675.300 276.900 686.700 ;
        RECT 278.700 682.050 279.900 689.400 ;
        RECT 299.100 689.400 301.500 690.900 ;
        RECT 304.800 689.400 306.600 702.000 ;
        RECT 323.100 695.400 324.900 702.000 ;
        RECT 326.100 695.400 327.900 701.400 ;
        RECT 341.100 695.400 342.900 702.000 ;
        RECT 344.100 695.400 345.900 701.400 ;
        RECT 347.100 695.400 348.900 702.000 ;
        RECT 365.100 695.400 366.900 702.000 ;
        RECT 368.100 695.400 369.900 701.400 ;
        RECT 299.100 682.050 300.300 689.400 ;
        RECT 305.100 682.050 306.900 683.850 ;
        RECT 323.100 682.050 324.900 683.850 ;
        RECT 326.100 682.050 327.300 695.400 ;
        RECT 344.100 682.050 345.300 695.400 ;
        RECT 365.100 682.050 366.900 683.850 ;
        RECT 368.100 682.050 369.300 695.400 ;
        RECT 383.100 690.600 384.900 701.400 ;
        RECT 386.100 691.500 387.900 702.000 ;
        RECT 383.100 689.400 387.900 690.600 ;
        RECT 385.800 688.500 387.900 689.400 ;
        RECT 390.600 689.400 392.400 701.400 ;
        RECT 395.100 691.500 396.900 702.000 ;
        RECT 398.100 690.300 399.900 701.400 ;
        RECT 395.400 689.400 399.900 690.300 ;
        RECT 416.100 690.300 417.900 701.400 ;
        RECT 419.100 691.500 420.900 702.000 ;
        RECT 416.100 689.400 420.600 690.300 ;
        RECT 423.600 689.400 425.400 701.400 ;
        RECT 428.100 691.500 429.900 702.000 ;
        RECT 431.100 690.600 432.900 701.400 ;
        RECT 446.100 695.400 447.900 702.000 ;
        RECT 449.100 695.400 450.900 701.400 ;
        RECT 452.100 695.400 453.900 702.000 ;
        RECT 390.600 688.050 391.800 689.400 ;
        RECT 390.300 687.000 391.800 688.050 ;
        RECT 395.400 687.300 397.500 689.400 ;
        RECT 418.500 687.300 420.600 689.400 ;
        RECT 424.200 688.050 425.400 689.400 ;
        RECT 428.100 689.400 432.900 690.600 ;
        RECT 428.100 688.500 430.200 689.400 ;
        RECT 424.200 687.000 425.700 688.050 ;
        RECT 390.300 685.050 391.200 687.000 ;
        RECT 383.400 682.050 385.200 683.850 ;
        RECT 389.100 682.950 391.200 685.050 ;
        RECT 392.100 685.500 394.200 685.800 ;
        RECT 421.800 685.500 423.900 685.800 ;
        RECT 392.100 683.700 396.000 685.500 ;
        RECT 420.000 683.700 423.900 685.500 ;
        RECT 424.800 685.050 425.700 687.000 ;
        RECT 277.800 679.950 279.900 682.050 ;
        RECT 295.950 679.950 298.050 682.050 ;
        RECT 298.950 679.950 301.050 682.050 ;
        RECT 301.950 679.950 304.050 682.050 ;
        RECT 304.950 679.950 307.050 682.050 ;
        RECT 322.950 679.950 325.050 682.050 ;
        RECT 325.950 679.950 328.050 682.050 ;
        RECT 340.950 679.950 343.050 682.050 ;
        RECT 343.950 679.950 346.050 682.050 ;
        RECT 346.950 679.950 349.050 682.050 ;
        RECT 364.950 679.950 367.050 682.050 ;
        RECT 367.950 679.950 370.050 682.050 ;
        RECT 383.100 679.950 385.200 682.050 ;
        RECT 389.700 682.800 391.200 682.950 ;
        RECT 424.800 682.950 426.900 685.050 ;
        RECT 424.800 682.800 426.300 682.950 ;
        RECT 389.700 681.900 392.100 682.800 ;
        RECT 276.000 674.400 277.800 675.300 ;
        RECT 249.000 666.000 250.800 672.600 ;
        RECT 253.500 671.400 258.600 672.600 ;
        RECT 272.100 673.500 277.800 674.400 ;
        RECT 253.500 666.600 255.300 671.400 ;
        RECT 272.100 669.600 273.300 673.500 ;
        RECT 278.700 672.600 279.900 679.950 ;
        RECT 296.100 678.150 297.900 679.950 ;
        RECT 299.100 675.600 300.300 679.950 ;
        RECT 302.100 678.150 303.900 679.950 ;
        RECT 296.700 674.700 300.300 675.600 ;
        RECT 296.700 672.600 297.900 674.700 ;
        RECT 256.500 666.000 258.300 669.600 ;
        RECT 272.100 666.600 273.900 669.600 ;
        RECT 275.100 666.000 276.900 672.600 ;
        RECT 278.100 666.600 279.900 672.600 ;
        RECT 296.100 666.600 297.900 672.600 ;
        RECT 299.100 671.700 306.900 673.050 ;
        RECT 299.100 666.600 300.900 671.700 ;
        RECT 302.100 666.000 303.900 670.800 ;
        RECT 305.100 666.600 306.900 671.700 ;
        RECT 326.100 669.600 327.300 679.950 ;
        RECT 341.250 678.150 343.050 679.950 ;
        RECT 344.100 674.700 345.300 679.950 ;
        RECT 347.100 678.150 348.900 679.950 ;
        RECT 344.100 673.800 348.300 674.700 ;
        RECT 323.100 666.000 324.900 669.600 ;
        RECT 326.100 666.600 327.900 669.600 ;
        RECT 341.400 666.000 343.200 672.600 ;
        RECT 346.500 666.600 348.300 673.800 ;
        RECT 368.100 669.600 369.300 679.950 ;
        RECT 387.900 679.200 389.700 681.000 ;
        RECT 387.900 677.100 390.000 679.200 ;
        RECT 390.900 676.200 392.100 681.900 ;
        RECT 393.000 682.050 394.800 682.500 ;
        RECT 421.200 682.050 423.000 682.500 ;
        RECT 393.000 680.700 399.900 682.050 ;
        RECT 397.800 679.950 399.900 680.700 ;
        RECT 416.100 680.700 423.000 682.050 ;
        RECT 423.900 681.900 426.300 682.800 ;
        RECT 430.800 682.050 432.600 683.850 ;
        RECT 449.700 682.050 450.900 695.400 ;
        RECT 467.100 689.400 468.900 701.400 ;
        RECT 470.100 691.200 471.900 702.000 ;
        RECT 473.100 695.400 474.900 701.400 ;
        RECT 467.100 682.050 468.300 689.400 ;
        RECT 473.700 688.500 474.900 695.400 ;
        RECT 469.200 687.600 474.900 688.500 ;
        RECT 476.550 689.400 478.350 701.400 ;
        RECT 479.550 689.400 481.350 702.000 ;
        RECT 484.350 695.400 486.150 701.400 ;
        RECT 488.850 695.400 490.650 702.000 ;
        RECT 484.350 693.300 486.450 695.400 ;
        RECT 491.850 694.500 493.650 701.400 ;
        RECT 494.850 695.400 496.650 702.000 ;
        RECT 490.950 693.450 497.550 694.500 ;
        RECT 490.950 692.700 492.750 693.450 ;
        RECT 495.750 692.700 497.550 693.450 ;
        RECT 499.650 692.400 501.450 701.400 ;
        RECT 483.450 690.600 486.450 692.400 ;
        RECT 487.350 691.800 489.150 692.400 ;
        RECT 487.350 690.900 493.050 691.800 ;
        RECT 499.650 691.500 501.750 692.400 ;
        RECT 487.350 690.600 489.150 690.900 ;
        RECT 485.250 689.700 486.450 690.600 ;
        RECT 469.200 686.700 471.000 687.600 ;
        RECT 416.100 679.950 418.200 680.700 ;
        RECT 385.800 673.500 387.900 674.700 ;
        RECT 389.100 674.100 392.100 676.200 ;
        RECT 393.000 677.400 394.800 679.200 ;
        RECT 397.800 678.150 399.600 679.950 ;
        RECT 416.400 678.150 418.200 679.950 ;
        RECT 421.200 677.400 423.000 679.200 ;
        RECT 393.000 675.300 395.100 677.400 ;
        RECT 420.900 675.300 423.000 677.400 ;
        RECT 393.000 674.400 399.300 675.300 ;
        RECT 383.100 672.600 387.900 673.500 ;
        RECT 390.900 672.600 392.100 674.100 ;
        RECT 398.100 672.600 399.300 674.400 ;
        RECT 416.700 674.400 423.000 675.300 ;
        RECT 423.900 676.200 425.100 681.900 ;
        RECT 426.300 679.200 428.100 681.000 ;
        RECT 430.800 679.950 432.900 682.050 ;
        RECT 445.950 679.950 448.050 682.050 ;
        RECT 448.950 679.950 451.050 682.050 ;
        RECT 451.950 679.950 454.050 682.050 ;
        RECT 467.100 679.950 469.200 682.050 ;
        RECT 426.000 677.100 428.100 679.200 ;
        RECT 446.100 678.150 447.900 679.950 ;
        RECT 416.700 672.600 417.900 674.400 ;
        RECT 423.900 674.100 426.900 676.200 ;
        RECT 449.700 674.700 450.900 679.950 ;
        RECT 451.950 678.150 453.750 679.950 ;
        RECT 423.900 672.600 425.100 674.100 ;
        RECT 428.100 673.500 430.200 674.700 ;
        RECT 446.700 673.800 450.900 674.700 ;
        RECT 428.100 672.600 432.900 673.500 ;
        RECT 365.100 666.000 366.900 669.600 ;
        RECT 368.100 666.600 369.900 669.600 ;
        RECT 383.100 666.600 384.900 672.600 ;
        RECT 386.100 666.000 387.900 671.700 ;
        RECT 390.600 666.600 392.400 672.600 ;
        RECT 395.100 666.000 396.900 671.700 ;
        RECT 398.100 666.600 399.900 672.600 ;
        RECT 416.100 666.600 417.900 672.600 ;
        RECT 419.100 666.000 420.900 671.700 ;
        RECT 423.600 666.600 425.400 672.600 ;
        RECT 428.100 666.000 429.900 671.700 ;
        RECT 431.100 666.600 432.900 672.600 ;
        RECT 446.700 666.600 448.500 673.800 ;
        RECT 467.100 672.600 468.300 679.950 ;
        RECT 470.100 675.300 471.000 686.700 ;
        RECT 472.800 682.050 474.600 683.850 ;
        RECT 472.500 679.950 474.600 682.050 ;
        RECT 476.550 682.050 477.750 689.400 ;
        RECT 485.250 688.800 490.050 689.700 ;
        RECT 478.650 686.100 480.450 686.550 ;
        RECT 484.350 686.100 486.450 686.700 ;
        RECT 478.650 684.900 486.450 686.100 ;
        RECT 478.650 684.750 480.450 684.900 ;
        RECT 484.350 684.600 486.450 684.900 ;
        RECT 476.550 681.750 481.050 682.050 ;
        RECT 476.550 679.950 482.850 681.750 ;
        RECT 469.200 674.400 471.000 675.300 ;
        RECT 469.200 673.500 474.900 674.400 ;
        RECT 451.800 666.000 453.600 672.600 ;
        RECT 467.100 666.600 468.900 672.600 ;
        RECT 470.100 666.000 471.900 672.600 ;
        RECT 473.700 669.600 474.900 673.500 ;
        RECT 473.100 666.600 474.900 669.600 ;
        RECT 476.550 672.600 477.750 679.950 ;
        RECT 489.150 676.200 490.050 688.800 ;
        RECT 492.150 688.800 493.050 690.900 ;
        RECT 493.950 690.300 501.750 691.500 ;
        RECT 493.950 689.700 495.750 690.300 ;
        RECT 505.050 689.400 506.850 702.000 ;
        RECT 508.050 691.200 509.850 701.400 ;
        RECT 508.050 689.400 510.450 691.200 ;
        RECT 492.150 688.500 500.550 688.800 ;
        RECT 509.550 688.500 510.450 689.400 ;
        RECT 492.150 687.900 510.450 688.500 ;
        RECT 498.750 687.300 510.450 687.900 ;
        RECT 498.750 687.000 500.550 687.300 ;
        RECT 496.800 680.400 498.900 682.050 ;
        RECT 496.800 679.200 504.900 680.400 ;
        RECT 505.950 679.950 508.050 682.050 ;
        RECT 503.100 678.600 504.900 679.200 ;
        RECT 500.100 677.400 501.900 678.000 ;
        RECT 506.250 677.400 508.050 679.950 ;
        RECT 500.100 676.200 508.050 677.400 ;
        RECT 489.150 675.000 501.150 676.200 ;
        RECT 489.150 674.400 490.950 675.000 ;
        RECT 500.100 673.200 501.150 675.000 ;
        RECT 476.550 666.600 478.350 672.600 ;
        RECT 479.850 666.000 481.650 672.600 ;
        RECT 484.350 669.600 486.750 671.700 ;
        RECT 496.350 671.550 498.150 672.300 ;
        RECT 493.200 670.500 498.150 671.550 ;
        RECT 499.350 671.400 501.150 673.200 ;
        RECT 509.550 672.600 510.450 687.300 ;
        RECT 493.200 669.600 494.250 670.500 ;
        RECT 502.050 670.200 504.150 671.700 ;
        RECT 500.250 669.600 504.150 670.200 ;
        RECT 484.950 666.600 486.750 669.600 ;
        RECT 489.450 666.000 491.250 669.600 ;
        RECT 492.450 666.600 494.250 669.600 ;
        RECT 495.750 666.000 497.550 669.600 ;
        RECT 500.250 668.700 503.850 669.600 ;
        RECT 500.250 666.600 502.050 668.700 ;
        RECT 505.050 666.000 506.850 672.600 ;
        RECT 508.050 670.800 510.450 672.600 ;
        RECT 512.550 689.400 514.350 701.400 ;
        RECT 515.550 689.400 517.350 702.000 ;
        RECT 520.350 695.400 522.150 701.400 ;
        RECT 524.850 695.400 526.650 702.000 ;
        RECT 520.350 693.300 522.450 695.400 ;
        RECT 527.850 694.500 529.650 701.400 ;
        RECT 530.850 695.400 532.650 702.000 ;
        RECT 526.950 693.450 533.550 694.500 ;
        RECT 526.950 692.700 528.750 693.450 ;
        RECT 531.750 692.700 533.550 693.450 ;
        RECT 535.650 692.400 537.450 701.400 ;
        RECT 519.450 690.600 522.450 692.400 ;
        RECT 523.350 691.800 525.150 692.400 ;
        RECT 523.350 690.900 529.050 691.800 ;
        RECT 535.650 691.500 537.750 692.400 ;
        RECT 523.350 690.600 525.150 690.900 ;
        RECT 521.250 689.700 522.450 690.600 ;
        RECT 512.550 682.050 513.750 689.400 ;
        RECT 521.250 688.800 526.050 689.700 ;
        RECT 514.650 686.100 516.450 686.550 ;
        RECT 520.350 686.100 522.450 686.700 ;
        RECT 514.650 684.900 522.450 686.100 ;
        RECT 514.650 684.750 516.450 684.900 ;
        RECT 520.350 684.600 522.450 684.900 ;
        RECT 512.550 681.750 517.050 682.050 ;
        RECT 512.550 679.950 518.850 681.750 ;
        RECT 512.550 672.600 513.750 679.950 ;
        RECT 525.150 676.200 526.050 688.800 ;
        RECT 528.150 688.800 529.050 690.900 ;
        RECT 529.950 690.300 537.750 691.500 ;
        RECT 529.950 689.700 531.750 690.300 ;
        RECT 541.050 689.400 542.850 702.000 ;
        RECT 544.050 691.200 545.850 701.400 ;
        RECT 563.100 695.400 564.900 701.400 ;
        RECT 566.100 695.400 567.900 702.000 ;
        RECT 581.100 695.400 582.900 702.000 ;
        RECT 584.100 695.400 585.900 701.400 ;
        RECT 587.100 695.400 588.900 702.000 ;
        RECT 544.050 689.400 546.450 691.200 ;
        RECT 528.150 688.500 536.550 688.800 ;
        RECT 545.550 688.500 546.450 689.400 ;
        RECT 528.150 687.900 546.450 688.500 ;
        RECT 534.750 687.300 546.450 687.900 ;
        RECT 534.750 687.000 536.550 687.300 ;
        RECT 532.800 680.400 534.900 682.050 ;
        RECT 532.800 679.200 540.900 680.400 ;
        RECT 541.950 679.950 544.050 682.050 ;
        RECT 539.100 678.600 540.900 679.200 ;
        RECT 536.100 677.400 537.900 678.000 ;
        RECT 542.250 677.400 544.050 679.950 ;
        RECT 536.100 676.200 544.050 677.400 ;
        RECT 525.150 675.000 537.150 676.200 ;
        RECT 525.150 674.400 526.950 675.000 ;
        RECT 536.100 673.200 537.150 675.000 ;
        RECT 508.050 666.600 509.850 670.800 ;
        RECT 512.550 666.600 514.350 672.600 ;
        RECT 515.850 666.000 517.650 672.600 ;
        RECT 520.350 669.600 522.750 671.700 ;
        RECT 532.350 671.550 534.150 672.300 ;
        RECT 529.200 670.500 534.150 671.550 ;
        RECT 535.350 671.400 537.150 673.200 ;
        RECT 545.550 672.600 546.450 687.300 ;
        RECT 563.700 682.050 564.900 695.400 ;
        RECT 568.950 684.450 571.050 685.050 ;
        RECT 574.950 684.450 577.050 685.050 ;
        RECT 566.100 682.050 567.900 683.850 ;
        RECT 568.950 683.550 577.050 684.450 ;
        RECT 568.950 682.950 571.050 683.550 ;
        RECT 574.950 682.950 577.050 683.550 ;
        RECT 584.700 682.050 585.900 695.400 ;
        RECT 602.100 689.400 603.900 701.400 ;
        RECT 605.100 690.000 606.900 702.000 ;
        RECT 608.100 695.400 609.900 701.400 ;
        RECT 611.100 695.400 612.900 702.000 ;
        RECT 602.700 682.050 603.600 689.400 ;
        RECT 606.000 682.050 607.800 683.850 ;
        RECT 562.950 679.950 565.050 682.050 ;
        RECT 565.950 679.950 568.050 682.050 ;
        RECT 580.950 679.950 583.050 682.050 ;
        RECT 583.950 679.950 586.050 682.050 ;
        RECT 586.950 679.950 589.050 682.050 ;
        RECT 602.100 679.950 604.200 682.050 ;
        RECT 605.400 679.950 607.500 682.050 ;
        RECT 529.200 669.600 530.250 670.500 ;
        RECT 538.050 670.200 540.150 671.700 ;
        RECT 536.250 669.600 540.150 670.200 ;
        RECT 520.950 666.600 522.750 669.600 ;
        RECT 525.450 666.000 527.250 669.600 ;
        RECT 528.450 666.600 530.250 669.600 ;
        RECT 531.750 666.000 533.550 669.600 ;
        RECT 536.250 668.700 539.850 669.600 ;
        RECT 536.250 666.600 538.050 668.700 ;
        RECT 541.050 666.000 542.850 672.600 ;
        RECT 544.050 670.800 546.450 672.600 ;
        RECT 544.050 666.600 545.850 670.800 ;
        RECT 563.700 669.600 564.900 679.950 ;
        RECT 581.100 678.150 582.900 679.950 ;
        RECT 584.700 674.700 585.900 679.950 ;
        RECT 586.950 678.150 588.750 679.950 ;
        RECT 581.700 673.800 585.900 674.700 ;
        RECT 563.100 666.600 564.900 669.600 ;
        RECT 566.100 666.000 567.900 669.600 ;
        RECT 568.950 669.450 571.050 670.050 ;
        RECT 574.950 669.450 577.050 670.050 ;
        RECT 568.950 668.550 577.050 669.450 ;
        RECT 568.950 667.950 571.050 668.550 ;
        RECT 574.950 667.950 577.050 668.550 ;
        RECT 581.700 666.600 583.500 673.800 ;
        RECT 602.700 672.600 603.600 679.950 ;
        RECT 609.000 675.300 609.900 695.400 ;
        RECT 629.400 689.400 631.200 702.000 ;
        RECT 634.500 690.900 636.300 701.400 ;
        RECT 637.500 695.400 639.300 702.000 ;
        RECT 653.100 695.400 654.900 701.400 ;
        RECT 656.100 696.000 657.900 702.000 ;
        RECT 654.000 695.100 654.900 695.400 ;
        RECT 659.100 695.400 660.900 701.400 ;
        RECT 662.100 695.400 663.900 702.000 ;
        RECT 659.100 695.100 660.600 695.400 ;
        RECT 654.000 694.200 660.600 695.100 ;
        RECT 637.200 692.100 639.000 693.900 ;
        RECT 634.500 689.400 636.900 690.900 ;
        RECT 629.100 682.050 630.900 683.850 ;
        RECT 635.700 682.050 636.900 689.400 ;
        RECT 654.000 682.050 654.900 694.200 ;
        RECT 677.100 689.400 678.900 701.400 ;
        RECT 680.100 690.300 681.900 701.400 ;
        RECT 683.100 691.200 684.900 702.000 ;
        RECT 686.100 690.300 687.900 701.400 ;
        RECT 704.100 695.400 705.900 701.400 ;
        RECT 707.100 696.000 708.900 702.000 ;
        RECT 680.100 689.400 687.900 690.300 ;
        RECT 705.000 695.100 705.900 695.400 ;
        RECT 710.100 695.400 711.900 701.400 ;
        RECT 713.100 695.400 714.900 702.000 ;
        RECT 710.100 695.100 711.600 695.400 ;
        RECT 705.000 694.200 711.600 695.100 ;
        RECT 659.100 682.050 660.900 683.850 ;
        RECT 677.400 682.050 678.300 689.400 ;
        RECT 679.950 687.450 682.050 688.050 ;
        RECT 691.950 687.450 694.050 688.050 ;
        RECT 679.950 686.550 694.050 687.450 ;
        RECT 679.950 685.950 682.050 686.550 ;
        RECT 691.950 685.950 694.050 686.550 ;
        RECT 682.950 682.050 684.750 683.850 ;
        RECT 705.000 682.050 705.900 694.200 ;
        RECT 728.100 689.400 729.900 701.400 ;
        RECT 731.100 690.300 732.900 701.400 ;
        RECT 734.100 691.200 735.900 702.000 ;
        RECT 737.100 690.300 738.900 701.400 ;
        RECT 755.100 695.400 756.900 701.400 ;
        RECT 758.100 696.000 759.900 702.000 ;
        RECT 731.100 689.400 738.900 690.300 ;
        RECT 756.000 695.100 756.900 695.400 ;
        RECT 761.100 695.400 762.900 701.400 ;
        RECT 764.100 695.400 765.900 702.000 ;
        RECT 779.700 695.400 781.500 702.000 ;
        RECT 761.100 695.100 762.600 695.400 ;
        RECT 756.000 694.200 762.600 695.100 ;
        RECT 710.100 682.050 711.900 683.850 ;
        RECT 728.400 682.050 729.300 689.400 ;
        RECT 730.950 687.450 733.050 688.050 ;
        RECT 745.950 687.450 748.050 688.050 ;
        RECT 730.950 686.550 748.050 687.450 ;
        RECT 730.950 685.950 733.050 686.550 ;
        RECT 745.950 685.950 748.050 686.550 ;
        RECT 733.950 682.050 735.750 683.850 ;
        RECT 756.000 682.050 756.900 694.200 ;
        RECT 780.000 692.100 781.800 693.900 ;
        RECT 782.700 690.900 784.500 701.400 ;
        RECT 782.100 689.400 784.500 690.900 ;
        RECT 787.800 689.400 789.600 702.000 ;
        RECT 803.100 689.400 804.900 701.400 ;
        RECT 806.100 690.300 807.900 701.400 ;
        RECT 809.100 691.200 810.900 702.000 ;
        RECT 812.100 690.300 813.900 701.400 ;
        RECT 806.100 689.400 813.900 690.300 ;
        RECT 827.100 690.600 828.900 701.400 ;
        RECT 830.100 691.500 831.900 702.000 ;
        RECT 833.100 700.500 840.900 701.400 ;
        RECT 833.100 690.600 834.900 700.500 ;
        RECT 827.100 689.700 834.900 690.600 ;
        RECT 761.100 682.050 762.900 683.850 ;
        RECT 782.100 682.050 783.300 689.400 ;
        RECT 788.100 682.050 789.900 683.850 ;
        RECT 803.400 682.050 804.300 689.400 ;
        RECT 836.100 688.500 837.900 699.600 ;
        RECT 839.100 689.400 840.900 700.500 ;
        RECT 857.100 695.400 858.900 701.400 ;
        RECT 860.100 696.000 861.900 702.000 ;
        RECT 858.000 695.100 858.900 695.400 ;
        RECT 863.100 695.400 864.900 701.400 ;
        RECT 866.100 695.400 867.900 702.000 ;
        RECT 863.100 695.100 864.600 695.400 ;
        RECT 858.000 694.200 864.600 695.100 ;
        RECT 833.100 687.600 837.900 688.500 ;
        RECT 808.950 682.050 810.750 683.850 ;
        RECT 830.250 682.050 832.050 683.850 ;
        RECT 833.100 682.050 834.000 687.600 ;
        RECT 836.100 682.050 837.900 683.850 ;
        RECT 858.000 682.050 858.900 694.200 ;
        RECT 884.100 690.300 885.900 701.400 ;
        RECT 887.100 691.200 888.900 702.000 ;
        RECT 890.100 690.300 891.900 701.400 ;
        RECT 884.100 689.400 891.900 690.300 ;
        RECT 893.100 689.400 894.900 701.400 ;
        RECT 877.950 687.450 880.050 688.050 ;
        RECT 886.950 687.450 889.050 688.050 ;
        RECT 877.950 686.550 889.050 687.450 ;
        RECT 877.950 685.950 880.050 686.550 ;
        RECT 886.950 685.950 889.050 686.550 ;
        RECT 863.100 682.050 864.900 683.850 ;
        RECT 887.250 682.050 889.050 683.850 ;
        RECT 893.700 682.050 894.600 689.400 ;
        RECT 610.800 679.950 612.900 682.050 ;
        RECT 628.950 679.950 631.050 682.050 ;
        RECT 631.950 679.950 634.050 682.050 ;
        RECT 634.950 679.950 637.050 682.050 ;
        RECT 637.950 679.950 640.050 682.050 ;
        RECT 652.950 679.950 655.050 682.050 ;
        RECT 655.950 679.950 658.050 682.050 ;
        RECT 658.950 679.950 661.050 682.050 ;
        RECT 661.950 679.950 664.050 682.050 ;
        RECT 676.950 679.950 679.050 682.050 ;
        RECT 679.950 679.950 682.050 682.050 ;
        RECT 682.950 679.950 685.050 682.050 ;
        RECT 685.950 679.950 688.050 682.050 ;
        RECT 703.950 679.950 706.050 682.050 ;
        RECT 706.950 679.950 709.050 682.050 ;
        RECT 709.950 679.950 712.050 682.050 ;
        RECT 712.950 679.950 715.050 682.050 ;
        RECT 727.950 679.950 730.050 682.050 ;
        RECT 730.950 679.950 733.050 682.050 ;
        RECT 733.950 679.950 736.050 682.050 ;
        RECT 736.950 679.950 739.050 682.050 ;
        RECT 754.950 679.950 757.050 682.050 ;
        RECT 757.950 679.950 760.050 682.050 ;
        RECT 760.950 679.950 763.050 682.050 ;
        RECT 763.950 679.950 766.050 682.050 ;
        RECT 778.950 679.950 781.050 682.050 ;
        RECT 781.950 679.950 784.050 682.050 ;
        RECT 784.950 679.950 787.050 682.050 ;
        RECT 787.950 679.950 790.050 682.050 ;
        RECT 802.950 679.950 805.050 682.050 ;
        RECT 805.950 679.950 808.050 682.050 ;
        RECT 808.950 679.950 811.050 682.050 ;
        RECT 811.950 679.950 814.050 682.050 ;
        RECT 826.950 679.950 829.050 682.050 ;
        RECT 829.950 679.950 832.050 682.050 ;
        RECT 832.950 679.950 835.050 682.050 ;
        RECT 835.950 679.950 838.050 682.050 ;
        RECT 838.950 679.950 841.050 682.050 ;
        RECT 856.950 679.950 859.050 682.050 ;
        RECT 859.950 679.950 862.050 682.050 ;
        RECT 862.950 679.950 865.050 682.050 ;
        RECT 865.950 679.950 868.050 682.050 ;
        RECT 883.950 679.950 886.050 682.050 ;
        RECT 886.950 679.950 889.050 682.050 ;
        RECT 889.950 679.950 892.050 682.050 ;
        RECT 892.950 679.950 895.050 682.050 ;
        RECT 610.950 678.150 612.750 679.950 ;
        RECT 632.100 678.150 633.900 679.950 ;
        RECT 635.700 675.600 636.900 679.950 ;
        RECT 638.100 678.150 639.900 679.950 ;
        RECT 654.000 676.200 654.900 679.950 ;
        RECT 656.100 678.150 657.900 679.950 ;
        RECT 662.100 678.150 663.900 679.950 ;
        RECT 604.500 674.400 612.900 675.300 ;
        RECT 635.700 674.700 639.300 675.600 ;
        RECT 654.000 675.000 657.300 676.200 ;
        RECT 604.500 673.500 606.300 674.400 ;
        RECT 586.800 666.000 588.600 672.600 ;
        RECT 602.700 670.800 605.400 672.600 ;
        RECT 603.600 666.600 605.400 670.800 ;
        RECT 606.600 666.000 608.400 672.600 ;
        RECT 611.100 666.600 612.900 674.400 ;
        RECT 629.100 671.700 636.900 673.050 ;
        RECT 629.100 666.600 630.900 671.700 ;
        RECT 632.100 666.000 633.900 670.800 ;
        RECT 635.100 666.600 636.900 671.700 ;
        RECT 638.100 672.600 639.300 674.700 ;
        RECT 638.100 666.600 639.900 672.600 ;
        RECT 655.500 666.600 657.300 675.000 ;
        RECT 662.100 666.000 663.900 675.600 ;
        RECT 677.400 672.600 678.300 679.950 ;
        RECT 679.950 678.150 681.750 679.950 ;
        RECT 686.100 678.150 687.900 679.950 ;
        RECT 705.000 676.200 705.900 679.950 ;
        RECT 707.100 678.150 708.900 679.950 ;
        RECT 713.100 678.150 714.900 679.950 ;
        RECT 705.000 675.000 708.300 676.200 ;
        RECT 677.400 671.400 682.500 672.600 ;
        RECT 677.700 666.000 679.500 669.600 ;
        RECT 680.700 666.600 682.500 671.400 ;
        RECT 685.200 666.000 687.000 672.600 ;
        RECT 706.500 666.600 708.300 675.000 ;
        RECT 713.100 666.000 714.900 675.600 ;
        RECT 728.400 672.600 729.300 679.950 ;
        RECT 730.950 678.150 732.750 679.950 ;
        RECT 737.100 678.150 738.900 679.950 ;
        RECT 756.000 676.200 756.900 679.950 ;
        RECT 758.100 678.150 759.900 679.950 ;
        RECT 764.100 678.150 765.900 679.950 ;
        RECT 775.950 678.450 778.050 679.050 ;
        RECT 767.550 678.000 778.050 678.450 ;
        RECT 779.100 678.150 780.900 679.950 ;
        RECT 766.950 677.550 778.050 678.000 ;
        RECT 756.000 675.000 759.300 676.200 ;
        RECT 728.400 671.400 733.500 672.600 ;
        RECT 728.700 666.000 730.500 669.600 ;
        RECT 731.700 666.600 733.500 671.400 ;
        RECT 736.200 666.000 738.000 672.600 ;
        RECT 757.500 666.600 759.300 675.000 ;
        RECT 764.100 666.000 765.900 675.600 ;
        RECT 766.950 673.950 769.050 677.550 ;
        RECT 775.950 676.950 778.050 677.550 ;
        RECT 782.100 675.600 783.300 679.950 ;
        RECT 785.100 678.150 786.900 679.950 ;
        RECT 779.700 674.700 783.300 675.600 ;
        RECT 779.700 672.600 780.900 674.700 ;
        RECT 779.100 666.600 780.900 672.600 ;
        RECT 782.100 671.700 789.900 673.050 ;
        RECT 782.100 666.600 783.900 671.700 ;
        RECT 785.100 666.000 786.900 670.800 ;
        RECT 788.100 666.600 789.900 671.700 ;
        RECT 803.400 672.600 804.300 679.950 ;
        RECT 805.950 678.150 807.750 679.950 ;
        RECT 812.100 678.150 813.900 679.950 ;
        RECT 827.250 678.150 829.050 679.950 ;
        RECT 811.950 675.450 814.050 676.050 ;
        RECT 829.950 675.450 832.050 676.050 ;
        RECT 811.950 674.550 832.050 675.450 ;
        RECT 811.950 673.950 814.050 674.550 ;
        RECT 829.950 673.950 832.050 674.550 ;
        RECT 833.100 672.600 834.300 679.950 ;
        RECT 839.100 678.150 840.900 679.950 ;
        RECT 858.000 676.200 858.900 679.950 ;
        RECT 860.100 678.150 861.900 679.950 ;
        RECT 866.100 678.150 867.900 679.950 ;
        RECT 884.100 678.150 885.900 679.950 ;
        RECT 890.250 678.150 892.050 679.950 ;
        RECT 858.000 675.000 861.300 676.200 ;
        RECT 803.400 671.400 808.500 672.600 ;
        RECT 803.700 666.000 805.500 669.600 ;
        RECT 806.700 666.600 808.500 671.400 ;
        RECT 811.200 666.000 813.000 672.600 ;
        RECT 827.700 666.000 829.500 672.600 ;
        RECT 832.200 666.600 834.000 672.600 ;
        RECT 836.700 666.000 838.500 672.600 ;
        RECT 859.500 666.600 861.300 675.000 ;
        RECT 866.100 666.000 867.900 675.600 ;
        RECT 893.700 672.600 894.600 679.950 ;
        RECT 885.000 666.000 886.800 672.600 ;
        RECT 889.500 671.400 894.600 672.600 ;
        RECT 889.500 666.600 891.300 671.400 ;
        RECT 892.500 666.000 894.300 669.600 ;
        RECT 14.100 653.400 15.900 663.000 ;
        RECT 20.700 654.000 22.500 662.400 ;
        RECT 38.100 659.400 39.900 663.000 ;
        RECT 41.100 659.400 42.900 662.400 ;
        RECT 20.700 652.800 24.000 654.000 ;
        RECT 14.100 649.050 15.900 650.850 ;
        RECT 20.100 649.050 21.900 650.850 ;
        RECT 23.100 649.050 24.000 652.800 ;
        RECT 41.100 649.050 42.300 659.400 ;
        RECT 56.100 657.300 57.900 662.400 ;
        RECT 59.100 658.200 60.900 663.000 ;
        RECT 62.100 657.300 63.900 662.400 ;
        RECT 56.100 655.950 63.900 657.300 ;
        RECT 65.100 656.400 66.900 662.400 ;
        RECT 80.100 659.400 81.900 663.000 ;
        RECT 83.100 659.400 84.900 662.400 ;
        RECT 65.100 654.300 66.300 656.400 ;
        RECT 62.700 653.400 66.300 654.300 ;
        RECT 59.100 649.050 60.900 650.850 ;
        RECT 62.700 649.050 63.900 653.400 ;
        RECT 65.100 649.050 66.900 650.850 ;
        RECT 83.100 649.050 84.300 659.400 ;
        RECT 101.100 653.400 102.900 663.000 ;
        RECT 107.700 654.000 109.500 662.400 ;
        RECT 127.500 654.000 129.300 662.400 ;
        RECT 107.700 652.800 111.000 654.000 ;
        RECT 91.950 651.450 94.050 652.050 ;
        RECT 97.950 651.450 100.050 652.050 ;
        RECT 91.950 650.550 100.050 651.450 ;
        RECT 91.950 649.950 94.050 650.550 ;
        RECT 97.950 649.950 100.050 650.550 ;
        RECT 101.100 649.050 102.900 650.850 ;
        RECT 107.100 649.050 108.900 650.850 ;
        RECT 110.100 649.050 111.000 652.800 ;
        RECT 126.000 652.800 129.300 654.000 ;
        RECT 134.100 653.400 135.900 663.000 ;
        RECT 150.000 656.400 151.800 663.000 ;
        RECT 154.500 657.600 156.300 662.400 ;
        RECT 157.500 659.400 159.300 663.000 ;
        RECT 154.500 656.400 159.600 657.600 ;
        RECT 126.000 649.050 126.900 652.800 ;
        RECT 128.100 649.050 129.900 650.850 ;
        RECT 134.100 649.050 135.900 650.850 ;
        RECT 149.100 649.050 150.900 650.850 ;
        RECT 155.250 649.050 157.050 650.850 ;
        RECT 158.700 649.050 159.600 656.400 ;
        RECT 176.100 657.300 177.900 662.400 ;
        RECT 179.100 658.200 180.900 663.000 ;
        RECT 182.100 657.300 183.900 662.400 ;
        RECT 176.100 655.950 183.900 657.300 ;
        RECT 185.100 656.400 186.900 662.400 ;
        RECT 200.100 659.400 201.900 663.000 ;
        RECT 203.100 659.400 204.900 662.400 ;
        RECT 185.100 654.300 186.300 656.400 ;
        RECT 182.700 653.400 186.300 654.300 ;
        RECT 179.100 649.050 180.900 650.850 ;
        RECT 182.700 649.050 183.900 653.400 ;
        RECT 190.950 651.450 193.050 652.050 ;
        RECT 196.950 651.450 199.050 652.050 ;
        RECT 185.100 649.050 186.900 650.850 ;
        RECT 190.950 650.550 199.050 651.450 ;
        RECT 190.950 649.950 193.050 650.550 ;
        RECT 196.950 649.950 199.050 650.550 ;
        RECT 203.100 649.050 204.300 659.400 ;
        RECT 221.100 656.400 222.900 662.400 ;
        RECT 221.700 654.300 222.900 656.400 ;
        RECT 224.100 657.300 225.900 662.400 ;
        RECT 227.100 658.200 228.900 663.000 ;
        RECT 230.100 657.300 231.900 662.400 ;
        RECT 248.100 659.400 249.900 663.000 ;
        RECT 251.100 659.400 252.900 662.400 ;
        RECT 224.100 655.950 231.900 657.300 ;
        RECT 221.700 653.400 225.300 654.300 ;
        RECT 221.100 649.050 222.900 650.850 ;
        RECT 224.100 649.050 225.300 653.400 ;
        RECT 227.100 649.050 228.900 650.850 ;
        RECT 251.100 649.050 252.300 659.400 ;
        RECT 266.100 656.400 267.900 662.400 ;
        RECT 266.700 654.300 267.900 656.400 ;
        RECT 269.100 657.300 270.900 662.400 ;
        RECT 272.100 658.200 273.900 663.000 ;
        RECT 275.100 657.300 276.900 662.400 ;
        RECT 269.100 655.950 276.900 657.300 ;
        RECT 290.400 656.400 292.200 663.000 ;
        RECT 295.500 655.200 297.300 662.400 ;
        RECT 311.400 656.400 313.200 663.000 ;
        RECT 316.500 655.200 318.300 662.400 ;
        RECT 332.400 656.400 334.200 663.000 ;
        RECT 337.500 655.200 339.300 662.400 ;
        RECT 356.100 657.300 357.900 662.400 ;
        RECT 359.100 658.200 360.900 663.000 ;
        RECT 362.100 657.300 363.900 662.400 ;
        RECT 356.100 655.950 363.900 657.300 ;
        RECT 365.100 656.400 366.900 662.400 ;
        RECT 380.100 657.300 381.900 662.400 ;
        RECT 383.100 658.200 384.900 663.000 ;
        RECT 386.100 657.300 387.900 662.400 ;
        RECT 293.100 654.300 297.300 655.200 ;
        RECT 314.100 654.300 318.300 655.200 ;
        RECT 335.100 654.300 339.300 655.200 ;
        RECT 365.100 654.300 366.300 656.400 ;
        RECT 380.100 655.950 387.900 657.300 ;
        RECT 389.100 656.400 390.900 662.400 ;
        RECT 389.100 654.300 390.300 656.400 ;
        RECT 266.700 653.400 270.300 654.300 ;
        RECT 266.100 649.050 267.900 650.850 ;
        RECT 269.100 649.050 270.300 653.400 ;
        RECT 272.100 649.050 273.900 650.850 ;
        RECT 290.250 649.050 292.050 650.850 ;
        RECT 293.100 649.050 294.300 654.300 ;
        RECT 296.100 649.050 297.900 650.850 ;
        RECT 311.250 649.050 313.050 650.850 ;
        RECT 314.100 649.050 315.300 654.300 ;
        RECT 317.100 649.050 318.900 650.850 ;
        RECT 332.250 649.050 334.050 650.850 ;
        RECT 335.100 649.050 336.300 654.300 ;
        RECT 362.700 653.400 366.300 654.300 ;
        RECT 386.700 653.400 390.300 654.300 ;
        RECT 407.100 653.400 408.900 663.000 ;
        RECT 413.700 654.000 415.500 662.400 ;
        RECT 338.100 649.050 339.900 650.850 ;
        RECT 359.100 649.050 360.900 650.850 ;
        RECT 362.700 649.050 363.900 653.400 ;
        RECT 365.100 649.050 366.900 650.850 ;
        RECT 383.100 649.050 384.900 650.850 ;
        RECT 386.700 649.050 387.900 653.400 ;
        RECT 413.700 652.800 417.000 654.000 ;
        RECT 431.100 653.400 432.900 663.000 ;
        RECT 437.700 654.000 439.500 662.400 ;
        RECT 457.500 654.000 459.300 662.400 ;
        RECT 437.700 652.800 441.000 654.000 ;
        RECT 389.100 649.050 390.900 650.850 ;
        RECT 407.100 649.050 408.900 650.850 ;
        RECT 413.100 649.050 414.900 650.850 ;
        RECT 416.100 649.050 417.000 652.800 ;
        RECT 431.100 649.050 432.900 650.850 ;
        RECT 437.100 649.050 438.900 650.850 ;
        RECT 440.100 649.050 441.000 652.800 ;
        RECT 456.000 652.800 459.300 654.000 ;
        RECT 464.100 653.400 465.900 663.000 ;
        RECT 479.700 655.200 481.500 662.400 ;
        RECT 484.800 656.400 486.600 663.000 ;
        RECT 500.100 657.300 501.900 662.400 ;
        RECT 503.100 658.200 504.900 663.000 ;
        RECT 506.100 657.300 507.900 662.400 ;
        RECT 500.100 655.950 507.900 657.300 ;
        RECT 509.100 656.400 510.900 662.400 ;
        RECT 524.400 656.400 526.200 663.000 ;
        RECT 479.700 654.300 483.900 655.200 ;
        RECT 509.100 654.300 510.300 656.400 ;
        RECT 529.500 655.200 531.300 662.400 ;
        RECT 545.100 656.400 546.900 662.400 ;
        RECT 548.400 657.300 550.200 663.000 ;
        RECT 552.900 657.000 554.700 662.400 ;
        RECT 557.100 657.300 558.900 663.000 ;
        RECT 545.100 655.500 549.600 656.400 ;
        RECT 456.000 649.050 456.900 652.800 ;
        RECT 458.100 649.050 459.900 650.850 ;
        RECT 464.100 649.050 465.900 650.850 ;
        RECT 479.100 649.050 480.900 650.850 ;
        RECT 482.700 649.050 483.900 654.300 ;
        RECT 506.700 653.400 510.300 654.300 ;
        RECT 527.100 654.300 531.300 655.200 ;
        RECT 484.950 649.050 486.750 650.850 ;
        RECT 503.100 649.050 504.900 650.850 ;
        RECT 506.700 649.050 507.900 653.400 ;
        RECT 509.100 649.050 510.900 650.850 ;
        RECT 524.250 649.050 526.050 650.850 ;
        RECT 527.100 649.050 528.300 654.300 ;
        RECT 547.500 653.100 549.600 655.500 ;
        RECT 552.900 654.900 553.800 657.000 ;
        RECT 560.100 656.400 561.900 662.400 ;
        RECT 575.100 661.500 582.900 662.400 ;
        RECT 575.100 656.400 576.900 661.500 ;
        RECT 578.100 656.400 579.900 660.600 ;
        RECT 581.100 657.000 582.900 661.500 ;
        RECT 584.100 657.900 585.900 663.000 ;
        RECT 587.100 657.000 588.900 662.400 ;
        RECT 605.100 659.400 606.900 662.400 ;
        RECT 608.100 659.400 609.900 663.000 ;
        RECT 560.400 655.500 561.900 656.400 ;
        RECT 550.800 652.800 553.800 654.900 ;
        RECT 557.400 654.000 561.900 655.500 ;
        RECT 578.700 654.900 579.600 656.400 ;
        RECT 581.100 656.100 588.900 657.000 ;
        RECT 530.100 649.050 531.900 650.850 ;
        RECT 13.950 646.950 16.050 649.050 ;
        RECT 16.950 646.950 19.050 649.050 ;
        RECT 19.950 646.950 22.050 649.050 ;
        RECT 22.950 646.950 25.050 649.050 ;
        RECT 37.950 646.950 40.050 649.050 ;
        RECT 40.950 646.950 43.050 649.050 ;
        RECT 55.950 646.950 58.050 649.050 ;
        RECT 58.950 646.950 61.050 649.050 ;
        RECT 61.950 646.950 64.050 649.050 ;
        RECT 64.950 646.950 67.050 649.050 ;
        RECT 79.950 646.950 82.050 649.050 ;
        RECT 82.950 646.950 85.050 649.050 ;
        RECT 100.950 646.950 103.050 649.050 ;
        RECT 103.950 646.950 106.050 649.050 ;
        RECT 106.950 646.950 109.050 649.050 ;
        RECT 109.950 646.950 112.050 649.050 ;
        RECT 124.950 646.950 127.050 649.050 ;
        RECT 127.950 646.950 130.050 649.050 ;
        RECT 130.950 646.950 133.050 649.050 ;
        RECT 133.950 646.950 136.050 649.050 ;
        RECT 148.950 646.950 151.050 649.050 ;
        RECT 151.950 646.950 154.050 649.050 ;
        RECT 154.950 646.950 157.050 649.050 ;
        RECT 157.950 646.950 160.050 649.050 ;
        RECT 175.950 646.950 178.050 649.050 ;
        RECT 178.950 646.950 181.050 649.050 ;
        RECT 181.950 646.950 184.050 649.050 ;
        RECT 184.950 646.950 187.050 649.050 ;
        RECT 199.950 646.950 202.050 649.050 ;
        RECT 202.950 646.950 205.050 649.050 ;
        RECT 220.950 646.950 223.050 649.050 ;
        RECT 223.950 646.950 226.050 649.050 ;
        RECT 226.950 646.950 229.050 649.050 ;
        RECT 229.950 646.950 232.050 649.050 ;
        RECT 247.950 646.950 250.050 649.050 ;
        RECT 250.950 646.950 253.050 649.050 ;
        RECT 265.950 646.950 268.050 649.050 ;
        RECT 268.950 646.950 271.050 649.050 ;
        RECT 271.950 646.950 274.050 649.050 ;
        RECT 274.950 646.950 277.050 649.050 ;
        RECT 289.950 646.950 292.050 649.050 ;
        RECT 292.950 646.950 295.050 649.050 ;
        RECT 295.950 646.950 298.050 649.050 ;
        RECT 310.950 646.950 313.050 649.050 ;
        RECT 313.950 646.950 316.050 649.050 ;
        RECT 316.950 646.950 319.050 649.050 ;
        RECT 331.950 646.950 334.050 649.050 ;
        RECT 334.950 646.950 337.050 649.050 ;
        RECT 337.950 646.950 340.050 649.050 ;
        RECT 355.950 646.950 358.050 649.050 ;
        RECT 358.950 646.950 361.050 649.050 ;
        RECT 361.950 646.950 364.050 649.050 ;
        RECT 364.950 646.950 367.050 649.050 ;
        RECT 379.950 646.950 382.050 649.050 ;
        RECT 382.950 646.950 385.050 649.050 ;
        RECT 385.950 646.950 388.050 649.050 ;
        RECT 388.950 646.950 391.050 649.050 ;
        RECT 406.950 646.950 409.050 649.050 ;
        RECT 409.950 646.950 412.050 649.050 ;
        RECT 412.950 646.950 415.050 649.050 ;
        RECT 415.950 646.950 418.050 649.050 ;
        RECT 430.950 646.950 433.050 649.050 ;
        RECT 433.950 646.950 436.050 649.050 ;
        RECT 436.950 646.950 439.050 649.050 ;
        RECT 439.950 646.950 442.050 649.050 ;
        RECT 454.950 646.950 457.050 649.050 ;
        RECT 457.950 646.950 460.050 649.050 ;
        RECT 460.950 646.950 463.050 649.050 ;
        RECT 463.950 646.950 466.050 649.050 ;
        RECT 478.950 646.950 481.050 649.050 ;
        RECT 481.950 646.950 484.050 649.050 ;
        RECT 484.950 646.950 487.050 649.050 ;
        RECT 499.950 646.950 502.050 649.050 ;
        RECT 502.950 646.950 505.050 649.050 ;
        RECT 505.950 646.950 508.050 649.050 ;
        RECT 508.950 646.950 511.050 649.050 ;
        RECT 523.950 646.950 526.050 649.050 ;
        RECT 526.950 646.950 529.050 649.050 ;
        RECT 529.950 646.950 532.050 649.050 ;
        RECT 545.100 646.950 547.200 649.050 ;
        RECT 549.900 648.900 552.000 651.000 ;
        RECT 550.200 647.100 552.000 648.900 ;
        RECT 17.100 645.150 18.900 646.950 ;
        RECT 23.100 634.800 24.000 646.950 ;
        RECT 38.100 645.150 39.900 646.950 ;
        RECT 17.400 633.900 24.000 634.800 ;
        RECT 17.400 633.600 18.900 633.900 ;
        RECT 14.100 627.000 15.900 633.600 ;
        RECT 17.100 627.600 18.900 633.600 ;
        RECT 23.100 633.600 24.000 633.900 ;
        RECT 41.100 633.600 42.300 646.950 ;
        RECT 56.100 645.150 57.900 646.950 ;
        RECT 62.700 639.600 63.900 646.950 ;
        RECT 80.100 645.150 81.900 646.950 ;
        RECT 20.100 627.000 21.900 633.000 ;
        RECT 23.100 627.600 24.900 633.600 ;
        RECT 38.100 627.000 39.900 633.600 ;
        RECT 41.100 627.600 42.900 633.600 ;
        RECT 56.400 627.000 58.200 639.600 ;
        RECT 61.500 638.100 63.900 639.600 ;
        RECT 61.500 627.600 63.300 638.100 ;
        RECT 64.200 635.100 66.000 636.900 ;
        RECT 83.100 633.600 84.300 646.950 ;
        RECT 104.100 645.150 105.900 646.950 ;
        RECT 85.950 642.450 88.050 643.050 ;
        RECT 106.950 642.450 109.050 643.050 ;
        RECT 85.950 641.550 109.050 642.450 ;
        RECT 85.950 640.950 88.050 641.550 ;
        RECT 106.950 640.950 109.050 641.550 ;
        RECT 110.100 634.800 111.000 646.950 ;
        RECT 104.400 633.900 111.000 634.800 ;
        RECT 104.400 633.600 105.900 633.900 ;
        RECT 64.500 627.000 66.300 633.600 ;
        RECT 80.100 627.000 81.900 633.600 ;
        RECT 83.100 627.600 84.900 633.600 ;
        RECT 101.100 627.000 102.900 633.600 ;
        RECT 104.100 627.600 105.900 633.600 ;
        RECT 110.100 633.600 111.000 633.900 ;
        RECT 126.000 634.800 126.900 646.950 ;
        RECT 131.100 645.150 132.900 646.950 ;
        RECT 152.250 645.150 154.050 646.950 ;
        RECT 127.950 642.450 130.050 643.050 ;
        RECT 148.950 642.450 151.050 643.050 ;
        RECT 127.950 641.550 151.050 642.450 ;
        RECT 127.950 640.950 130.050 641.550 ;
        RECT 148.950 640.950 151.050 641.550 ;
        RECT 158.700 639.600 159.600 646.950 ;
        RECT 176.100 645.150 177.900 646.950 ;
        RECT 182.700 639.600 183.900 646.950 ;
        RECT 200.100 645.150 201.900 646.950 ;
        RECT 149.100 638.700 156.900 639.600 ;
        RECT 126.000 633.900 132.600 634.800 ;
        RECT 126.000 633.600 126.900 633.900 ;
        RECT 107.100 627.000 108.900 633.000 ;
        RECT 110.100 627.600 111.900 633.600 ;
        RECT 125.100 627.600 126.900 633.600 ;
        RECT 131.100 633.600 132.600 633.900 ;
        RECT 128.100 627.000 129.900 633.000 ;
        RECT 131.100 627.600 132.900 633.600 ;
        RECT 134.100 627.000 135.900 633.600 ;
        RECT 149.100 627.600 150.900 638.700 ;
        RECT 152.100 627.000 153.900 637.800 ;
        RECT 155.100 627.600 156.900 638.700 ;
        RECT 158.100 627.600 159.900 639.600 ;
        RECT 176.400 627.000 178.200 639.600 ;
        RECT 181.500 638.100 183.900 639.600 ;
        RECT 181.500 627.600 183.300 638.100 ;
        RECT 184.200 635.100 186.000 636.900 ;
        RECT 203.100 633.600 204.300 646.950 ;
        RECT 224.100 639.600 225.300 646.950 ;
        RECT 230.100 645.150 231.900 646.950 ;
        RECT 248.100 645.150 249.900 646.950 ;
        RECT 224.100 638.100 226.500 639.600 ;
        RECT 222.000 635.100 223.800 636.900 ;
        RECT 184.500 627.000 186.300 633.600 ;
        RECT 200.100 627.000 201.900 633.600 ;
        RECT 203.100 627.600 204.900 633.600 ;
        RECT 221.700 627.000 223.500 633.600 ;
        RECT 224.700 627.600 226.500 638.100 ;
        RECT 229.800 627.000 231.600 639.600 ;
        RECT 251.100 633.600 252.300 646.950 ;
        RECT 269.100 639.600 270.300 646.950 ;
        RECT 275.100 645.150 276.900 646.950 ;
        RECT 269.100 638.100 271.500 639.600 ;
        RECT 267.000 635.100 268.800 636.900 ;
        RECT 248.100 627.000 249.900 633.600 ;
        RECT 251.100 627.600 252.900 633.600 ;
        RECT 266.700 627.000 268.500 633.600 ;
        RECT 269.700 627.600 271.500 638.100 ;
        RECT 274.800 627.000 276.600 639.600 ;
        RECT 293.100 633.600 294.300 646.950 ;
        RECT 314.100 633.600 315.300 646.950 ;
        RECT 335.100 633.600 336.300 646.950 ;
        RECT 356.100 645.150 357.900 646.950 ;
        RECT 362.700 639.600 363.900 646.950 ;
        RECT 380.100 645.150 381.900 646.950 ;
        RECT 386.700 639.600 387.900 646.950 ;
        RECT 410.100 645.150 411.900 646.950 ;
        RECT 290.100 627.000 291.900 633.600 ;
        RECT 293.100 627.600 294.900 633.600 ;
        RECT 296.100 627.000 297.900 633.600 ;
        RECT 311.100 627.000 312.900 633.600 ;
        RECT 314.100 627.600 315.900 633.600 ;
        RECT 317.100 627.000 318.900 633.600 ;
        RECT 332.100 627.000 333.900 633.600 ;
        RECT 335.100 627.600 336.900 633.600 ;
        RECT 338.100 627.000 339.900 633.600 ;
        RECT 356.400 627.000 358.200 639.600 ;
        RECT 361.500 638.100 363.900 639.600 ;
        RECT 361.500 627.600 363.300 638.100 ;
        RECT 364.200 635.100 366.000 636.900 ;
        RECT 364.500 627.000 366.300 633.600 ;
        RECT 380.400 627.000 382.200 639.600 ;
        RECT 385.500 638.100 387.900 639.600 ;
        RECT 385.500 627.600 387.300 638.100 ;
        RECT 388.200 635.100 390.000 636.900 ;
        RECT 416.100 634.800 417.000 646.950 ;
        RECT 434.100 645.150 435.900 646.950 ;
        RECT 421.950 642.450 424.050 643.050 ;
        RECT 430.950 642.450 433.050 643.050 ;
        RECT 421.950 641.550 433.050 642.450 ;
        RECT 421.950 640.950 424.050 641.550 ;
        RECT 430.950 640.950 433.050 641.550 ;
        RECT 440.100 634.800 441.000 646.950 ;
        RECT 410.400 633.900 417.000 634.800 ;
        RECT 410.400 633.600 411.900 633.900 ;
        RECT 388.500 627.000 390.300 633.600 ;
        RECT 407.100 627.000 408.900 633.600 ;
        RECT 410.100 627.600 411.900 633.600 ;
        RECT 416.100 633.600 417.000 633.900 ;
        RECT 434.400 633.900 441.000 634.800 ;
        RECT 434.400 633.600 435.900 633.900 ;
        RECT 413.100 627.000 414.900 633.000 ;
        RECT 416.100 627.600 417.900 633.600 ;
        RECT 431.100 627.000 432.900 633.600 ;
        RECT 434.100 627.600 435.900 633.600 ;
        RECT 440.100 633.600 441.000 633.900 ;
        RECT 456.000 634.800 456.900 646.950 ;
        RECT 461.100 645.150 462.900 646.950 ;
        RECT 456.000 633.900 462.600 634.800 ;
        RECT 456.000 633.600 456.900 633.900 ;
        RECT 437.100 627.000 438.900 633.000 ;
        RECT 440.100 627.600 441.900 633.600 ;
        RECT 455.100 627.600 456.900 633.600 ;
        RECT 461.100 633.600 462.600 633.900 ;
        RECT 482.700 633.600 483.900 646.950 ;
        RECT 500.100 645.150 501.900 646.950 ;
        RECT 506.700 639.600 507.900 646.950 ;
        RECT 458.100 627.000 459.900 633.000 ;
        RECT 461.100 627.600 462.900 633.600 ;
        RECT 464.100 627.000 465.900 633.600 ;
        RECT 479.100 627.000 480.900 633.600 ;
        RECT 482.100 627.600 483.900 633.600 ;
        RECT 485.100 627.000 486.900 633.600 ;
        RECT 500.400 627.000 502.200 639.600 ;
        RECT 505.500 638.100 507.900 639.600 ;
        RECT 505.500 627.600 507.300 638.100 ;
        RECT 508.200 635.100 510.000 636.900 ;
        RECT 527.100 633.600 528.300 646.950 ;
        RECT 545.400 645.150 547.200 646.950 ;
        RECT 552.900 646.050 553.800 652.800 ;
        RECT 554.700 651.900 556.500 653.700 ;
        RECT 557.400 653.400 559.500 654.000 ;
        RECT 578.700 653.700 583.050 654.900 ;
        RECT 555.000 651.000 557.100 651.900 ;
        RECT 555.000 649.800 561.600 651.000 ;
        RECT 559.800 649.200 561.600 649.800 ;
        RECT 555.000 646.800 557.100 648.900 ;
        RECT 559.800 646.950 561.900 649.200 ;
        RECT 578.250 649.050 580.050 650.850 ;
        RECT 582.000 649.050 583.050 653.700 ;
        RECT 574.950 646.950 577.050 649.050 ;
        RECT 577.950 646.950 580.050 649.050 ;
        RECT 580.950 646.950 583.050 649.050 ;
        RECT 583.950 649.050 585.750 650.850 ;
        RECT 605.700 649.050 606.900 659.400 ;
        RECT 623.400 656.400 625.200 663.000 ;
        RECT 628.500 655.200 630.300 662.400 ;
        RECT 644.400 656.400 646.200 663.000 ;
        RECT 649.500 655.200 651.300 662.400 ;
        RECT 665.100 659.400 666.900 663.000 ;
        RECT 668.100 659.400 669.900 662.400 ;
        RECT 626.100 654.300 630.300 655.200 ;
        RECT 647.100 654.300 651.300 655.200 ;
        RECT 623.250 649.050 625.050 650.850 ;
        RECT 626.100 649.050 627.300 654.300 ;
        RECT 629.100 649.050 630.900 650.850 ;
        RECT 644.250 649.050 646.050 650.850 ;
        RECT 647.100 649.050 648.300 654.300 ;
        RECT 650.100 649.050 651.900 650.850 ;
        RECT 668.100 649.050 669.300 659.400 ;
        RECT 683.100 656.400 684.900 662.400 ;
        RECT 683.700 654.300 684.900 656.400 ;
        RECT 686.100 657.300 687.900 662.400 ;
        RECT 689.100 658.200 690.900 663.000 ;
        RECT 692.100 657.300 693.900 662.400 ;
        RECT 686.100 655.950 693.900 657.300 ;
        RECT 707.100 656.400 708.900 662.400 ;
        RECT 710.100 657.300 711.900 663.000 ;
        RECT 714.600 656.400 716.400 662.400 ;
        RECT 719.100 657.300 720.900 663.000 ;
        RECT 722.100 656.400 723.900 662.400 ;
        RECT 707.700 654.600 708.900 656.400 ;
        RECT 714.900 654.900 716.100 656.400 ;
        RECT 719.100 655.500 723.900 656.400 ;
        RECT 740.100 656.400 741.900 662.400 ;
        RECT 743.100 657.300 744.900 663.000 ;
        RECT 747.300 657.000 749.100 662.400 ;
        RECT 751.800 657.300 753.600 663.000 ;
        RECT 740.100 655.500 741.600 656.400 ;
        RECT 683.700 653.400 687.300 654.300 ;
        RECT 707.700 653.700 714.000 654.600 ;
        RECT 683.100 649.050 684.900 650.850 ;
        RECT 686.100 649.050 687.300 653.400 ;
        RECT 711.900 651.600 714.000 653.700 ;
        RECT 689.100 649.050 690.900 650.850 ;
        RECT 707.400 649.050 709.200 650.850 ;
        RECT 712.200 649.800 714.000 651.600 ;
        RECT 714.900 652.800 717.900 654.900 ;
        RECT 719.100 654.300 721.200 655.500 ;
        RECT 740.100 654.000 744.600 655.500 ;
        RECT 742.500 653.400 744.600 654.000 ;
        RECT 748.200 654.900 749.100 657.000 ;
        RECT 755.100 656.400 756.900 662.400 ;
        RECT 752.400 655.500 756.900 656.400 ;
        RECT 770.100 657.300 771.900 662.400 ;
        RECT 773.100 658.200 774.900 663.000 ;
        RECT 776.100 657.300 777.900 662.400 ;
        RECT 770.100 655.950 777.900 657.300 ;
        RECT 779.100 656.400 780.900 662.400 ;
        RECT 797.400 656.400 799.200 663.000 ;
        RECT 583.950 646.950 586.050 649.050 ;
        RECT 586.950 646.950 589.050 649.050 ;
        RECT 604.950 646.950 607.050 649.050 ;
        RECT 607.950 646.950 610.050 649.050 ;
        RECT 622.950 646.950 625.050 649.050 ;
        RECT 625.950 646.950 628.050 649.050 ;
        RECT 628.950 646.950 631.050 649.050 ;
        RECT 643.950 646.950 646.050 649.050 ;
        RECT 646.950 646.950 649.050 649.050 ;
        RECT 649.950 646.950 652.050 649.050 ;
        RECT 664.950 646.950 667.050 649.050 ;
        RECT 667.950 646.950 670.050 649.050 ;
        RECT 682.950 646.950 685.050 649.050 ;
        RECT 685.950 646.950 688.050 649.050 ;
        RECT 688.950 646.950 691.050 649.050 ;
        RECT 691.950 646.950 694.050 649.050 ;
        RECT 707.100 648.300 709.200 649.050 ;
        RECT 707.100 646.950 714.000 648.300 ;
        RECT 550.800 644.700 553.800 646.050 ;
        RECT 555.300 645.000 557.100 646.800 ;
        RECT 575.250 645.150 577.050 646.950 ;
        RECT 550.800 643.950 552.900 644.700 ;
        RECT 548.100 639.600 550.200 640.500 ;
        RECT 545.100 638.400 550.200 639.600 ;
        RECT 551.100 639.600 552.300 643.950 ;
        RECT 553.800 641.700 555.600 643.500 ;
        RECT 553.800 640.800 559.200 641.700 ;
        RECT 557.100 639.900 559.200 640.800 ;
        RECT 551.100 638.700 554.400 639.600 ;
        RECT 557.100 638.700 561.900 639.900 ;
        RECT 582.000 639.600 583.050 646.950 ;
        RECT 587.100 645.150 588.900 646.950 ;
        RECT 508.500 627.000 510.300 633.600 ;
        RECT 524.100 627.000 525.900 633.600 ;
        RECT 527.100 627.600 528.900 633.600 ;
        RECT 530.100 627.000 531.900 633.600 ;
        RECT 545.100 627.600 546.900 638.400 ;
        RECT 548.100 627.000 550.200 637.500 ;
        RECT 552.600 627.600 554.400 638.700 ;
        RECT 557.100 627.000 558.900 637.500 ;
        RECT 560.100 627.600 561.900 638.700 ;
        RECT 576.600 627.000 578.400 639.600 ;
        RECT 581.100 627.600 584.400 639.600 ;
        RECT 587.100 627.000 588.900 639.600 ;
        RECT 605.700 633.600 606.900 646.950 ;
        RECT 608.100 645.150 609.900 646.950 ;
        RECT 626.100 633.600 627.300 646.950 ;
        RECT 647.100 633.600 648.300 646.950 ;
        RECT 665.100 645.150 666.900 646.950 ;
        RECT 668.100 633.600 669.300 646.950 ;
        RECT 686.100 639.600 687.300 646.950 ;
        RECT 692.100 645.150 693.900 646.950 ;
        RECT 712.200 646.500 714.000 646.950 ;
        RECT 714.900 647.100 716.100 652.800 ;
        RECT 745.500 651.900 747.300 653.700 ;
        RECT 748.200 652.800 751.200 654.900 ;
        RECT 752.400 653.100 754.500 655.500 ;
        RECT 779.100 654.300 780.300 656.400 ;
        RECT 802.500 655.200 804.300 662.400 ;
        RECT 776.700 653.400 780.300 654.300 ;
        RECT 800.100 654.300 804.300 655.200 ;
        RECT 717.000 649.800 719.100 651.900 ;
        RECT 744.900 651.000 747.000 651.900 ;
        RECT 717.300 648.000 719.100 649.800 ;
        RECT 740.400 649.800 747.000 651.000 ;
        RECT 740.400 649.200 742.200 649.800 ;
        RECT 714.900 646.200 717.300 647.100 ;
        RECT 715.800 646.050 717.300 646.200 ;
        RECT 721.800 646.950 723.900 649.050 ;
        RECT 740.100 646.950 742.200 649.200 ;
        RECT 711.000 643.500 714.900 645.300 ;
        RECT 712.800 643.200 714.900 643.500 ;
        RECT 715.800 643.950 717.900 646.050 ;
        RECT 721.800 645.150 723.600 646.950 ;
        RECT 744.900 646.800 747.000 648.900 ;
        RECT 744.900 645.000 746.700 646.800 ;
        RECT 748.200 646.050 749.100 652.800 ;
        RECT 750.000 648.900 752.100 651.000 ;
        RECT 773.100 649.050 774.900 650.850 ;
        RECT 776.700 649.050 777.900 653.400 ;
        RECT 779.100 649.050 780.900 650.850 ;
        RECT 797.250 649.050 799.050 650.850 ;
        RECT 800.100 649.050 801.300 654.300 ;
        RECT 820.500 654.000 822.300 662.400 ;
        RECT 819.000 652.800 822.300 654.000 ;
        RECT 827.100 653.400 828.900 663.000 ;
        RECT 843.000 656.400 844.800 663.000 ;
        RECT 847.500 657.600 849.300 662.400 ;
        RECT 850.500 659.400 852.300 663.000 ;
        RECT 869.100 659.400 870.900 663.000 ;
        RECT 872.100 659.400 873.900 662.400 ;
        RECT 847.500 656.400 852.600 657.600 ;
        RECT 803.100 649.050 804.900 650.850 ;
        RECT 819.000 649.050 819.900 652.800 ;
        RECT 821.100 649.050 822.900 650.850 ;
        RECT 827.100 649.050 828.900 650.850 ;
        RECT 842.100 649.050 843.900 650.850 ;
        RECT 848.250 649.050 850.050 650.850 ;
        RECT 851.700 649.050 852.600 656.400 ;
        RECT 864.000 651.450 868.050 652.050 ;
        RECT 863.550 649.950 868.050 651.450 ;
        RECT 750.000 647.100 751.800 648.900 ;
        RECT 754.800 646.950 756.900 649.050 ;
        RECT 769.950 646.950 772.050 649.050 ;
        RECT 772.950 646.950 775.050 649.050 ;
        RECT 775.950 646.950 778.050 649.050 ;
        RECT 778.950 646.950 781.050 649.050 ;
        RECT 796.950 646.950 799.050 649.050 ;
        RECT 799.950 646.950 802.050 649.050 ;
        RECT 802.950 646.950 805.050 649.050 ;
        RECT 817.950 646.950 820.050 649.050 ;
        RECT 820.950 646.950 823.050 649.050 ;
        RECT 823.950 646.950 826.050 649.050 ;
        RECT 826.950 646.950 829.050 649.050 ;
        RECT 841.950 646.950 844.050 649.050 ;
        RECT 844.950 646.950 847.050 649.050 ;
        RECT 847.950 646.950 850.050 649.050 ;
        RECT 850.950 646.950 853.050 649.050 ;
        RECT 856.950 648.450 859.050 648.900 ;
        RECT 863.550 648.450 864.450 649.950 ;
        RECT 872.100 649.050 873.300 659.400 ;
        RECT 887.100 656.400 888.900 662.400 ;
        RECT 887.700 654.300 888.900 656.400 ;
        RECT 890.100 657.300 891.900 662.400 ;
        RECT 893.100 658.200 894.900 663.000 ;
        RECT 896.100 657.300 897.900 662.400 ;
        RECT 890.100 655.950 897.900 657.300 ;
        RECT 887.700 653.400 891.300 654.300 ;
        RECT 887.100 649.050 888.900 650.850 ;
        RECT 890.100 649.050 891.300 653.400 ;
        RECT 893.100 649.050 894.900 650.850 ;
        RECT 856.950 647.550 864.450 648.450 ;
        RECT 748.200 644.700 751.200 646.050 ;
        RECT 754.800 645.150 756.600 646.950 ;
        RECT 770.100 645.150 771.900 646.950 ;
        RECT 749.100 643.950 751.200 644.700 ;
        RECT 691.950 642.450 694.050 643.050 ;
        RECT 697.950 642.450 700.050 643.050 ;
        RECT 691.950 641.550 700.050 642.450 ;
        RECT 715.800 642.000 716.700 643.950 ;
        RECT 691.950 640.950 694.050 641.550 ;
        RECT 697.950 640.950 700.050 641.550 ;
        RECT 709.500 639.600 711.600 641.700 ;
        RECT 715.200 640.950 716.700 642.000 ;
        RECT 746.400 641.700 748.200 643.500 ;
        RECT 715.200 639.600 716.400 640.950 ;
        RECT 742.800 640.800 748.200 641.700 ;
        RECT 686.100 638.100 688.500 639.600 ;
        RECT 684.000 635.100 685.800 636.900 ;
        RECT 605.100 627.600 606.900 633.600 ;
        RECT 608.100 627.000 609.900 633.600 ;
        RECT 623.100 627.000 624.900 633.600 ;
        RECT 626.100 627.600 627.900 633.600 ;
        RECT 629.100 627.000 630.900 633.600 ;
        RECT 644.100 627.000 645.900 633.600 ;
        RECT 647.100 627.600 648.900 633.600 ;
        RECT 650.100 627.000 651.900 633.600 ;
        RECT 665.100 627.000 666.900 633.600 ;
        RECT 668.100 627.600 669.900 633.600 ;
        RECT 683.700 627.000 685.500 633.600 ;
        RECT 686.700 627.600 688.500 638.100 ;
        RECT 691.800 627.000 693.600 639.600 ;
        RECT 707.100 638.700 711.600 639.600 ;
        RECT 707.100 627.600 708.900 638.700 ;
        RECT 710.100 627.000 711.900 637.500 ;
        RECT 714.600 627.600 716.400 639.600 ;
        RECT 719.100 639.600 721.200 640.500 ;
        RECT 742.800 639.900 744.900 640.800 ;
        RECT 719.100 638.400 723.900 639.600 ;
        RECT 719.100 627.000 720.900 637.500 ;
        RECT 722.100 627.600 723.900 638.400 ;
        RECT 740.100 638.700 744.900 639.900 ;
        RECT 749.700 639.600 750.900 643.950 ;
        RECT 747.600 638.700 750.900 639.600 ;
        RECT 751.800 639.600 753.900 640.500 ;
        RECT 776.700 639.600 777.900 646.950 ;
        RECT 740.100 627.600 741.900 638.700 ;
        RECT 743.100 627.000 744.900 637.500 ;
        RECT 747.600 627.600 749.400 638.700 ;
        RECT 751.800 638.400 756.900 639.600 ;
        RECT 751.800 627.000 753.900 637.500 ;
        RECT 755.100 627.600 756.900 638.400 ;
        RECT 770.400 627.000 772.200 639.600 ;
        RECT 775.500 638.100 777.900 639.600 ;
        RECT 775.500 627.600 777.300 638.100 ;
        RECT 778.200 635.100 780.000 636.900 ;
        RECT 800.100 633.600 801.300 646.950 ;
        RECT 819.000 634.800 819.900 646.950 ;
        RECT 824.100 645.150 825.900 646.950 ;
        RECT 829.950 645.450 832.050 646.050 ;
        RECT 835.950 645.450 838.050 646.050 ;
        RECT 829.950 644.550 838.050 645.450 ;
        RECT 845.250 645.150 847.050 646.950 ;
        RECT 829.950 643.950 832.050 644.550 ;
        RECT 835.950 643.950 838.050 644.550 ;
        RECT 820.950 642.450 823.050 643.050 ;
        RECT 826.950 642.450 829.050 643.050 ;
        RECT 841.950 642.450 844.050 643.050 ;
        RECT 820.950 641.550 844.050 642.450 ;
        RECT 820.950 640.950 823.050 641.550 ;
        RECT 826.950 640.950 829.050 641.550 ;
        RECT 841.950 640.950 844.050 641.550 ;
        RECT 851.700 639.600 852.600 646.950 ;
        RECT 856.950 646.800 859.050 647.550 ;
        RECT 868.950 646.950 871.050 649.050 ;
        RECT 871.950 646.950 874.050 649.050 ;
        RECT 886.950 646.950 889.050 649.050 ;
        RECT 889.950 646.950 892.050 649.050 ;
        RECT 892.950 646.950 895.050 649.050 ;
        RECT 895.950 646.950 898.050 649.050 ;
        RECT 869.100 645.150 870.900 646.950 ;
        RECT 842.100 638.700 849.900 639.600 ;
        RECT 819.000 633.900 825.600 634.800 ;
        RECT 819.000 633.600 819.900 633.900 ;
        RECT 778.500 627.000 780.300 633.600 ;
        RECT 797.100 627.000 798.900 633.600 ;
        RECT 800.100 627.600 801.900 633.600 ;
        RECT 803.100 627.000 804.900 633.600 ;
        RECT 818.100 627.600 819.900 633.600 ;
        RECT 824.100 633.600 825.600 633.900 ;
        RECT 821.100 627.000 822.900 633.000 ;
        RECT 824.100 627.600 825.900 633.600 ;
        RECT 827.100 627.000 828.900 633.600 ;
        RECT 842.100 627.600 843.900 638.700 ;
        RECT 845.100 627.000 846.900 637.800 ;
        RECT 848.100 627.600 849.900 638.700 ;
        RECT 851.100 627.600 852.900 639.600 ;
        RECT 872.100 633.600 873.300 646.950 ;
        RECT 890.100 639.600 891.300 646.950 ;
        RECT 896.100 645.150 897.900 646.950 ;
        RECT 890.100 638.100 892.500 639.600 ;
        RECT 888.000 635.100 889.800 636.900 ;
        RECT 869.100 627.000 870.900 633.600 ;
        RECT 872.100 627.600 873.900 633.600 ;
        RECT 887.700 627.000 889.500 633.600 ;
        RECT 890.700 627.600 892.500 638.100 ;
        RECT 895.800 627.000 897.600 639.600 ;
        RECT 14.100 611.400 15.900 623.400 ;
        RECT 17.100 613.200 18.900 624.000 ;
        RECT 20.100 617.400 21.900 623.400 ;
        RECT 14.100 604.050 15.300 611.400 ;
        RECT 20.700 610.500 21.900 617.400 ;
        RECT 16.200 609.600 21.900 610.500 ;
        RECT 23.550 611.400 25.350 623.400 ;
        RECT 26.550 611.400 28.350 624.000 ;
        RECT 31.350 617.400 33.150 623.400 ;
        RECT 35.850 617.400 37.650 624.000 ;
        RECT 31.350 615.300 33.450 617.400 ;
        RECT 38.850 616.500 40.650 623.400 ;
        RECT 41.850 617.400 43.650 624.000 ;
        RECT 37.950 615.450 44.550 616.500 ;
        RECT 37.950 614.700 39.750 615.450 ;
        RECT 42.750 614.700 44.550 615.450 ;
        RECT 46.650 614.400 48.450 623.400 ;
        RECT 30.450 612.600 33.450 614.400 ;
        RECT 34.350 613.800 36.150 614.400 ;
        RECT 34.350 612.900 40.050 613.800 ;
        RECT 46.650 613.500 48.750 614.400 ;
        RECT 34.350 612.600 36.150 612.900 ;
        RECT 32.250 611.700 33.450 612.600 ;
        RECT 16.200 608.700 18.000 609.600 ;
        RECT 14.100 601.950 16.200 604.050 ;
        RECT 14.100 594.600 15.300 601.950 ;
        RECT 17.100 597.300 18.000 608.700 ;
        RECT 19.800 604.050 21.600 605.850 ;
        RECT 19.500 601.950 21.600 604.050 ;
        RECT 23.550 604.050 24.750 611.400 ;
        RECT 32.250 610.800 37.050 611.700 ;
        RECT 25.650 608.100 27.450 608.550 ;
        RECT 31.350 608.100 33.450 608.700 ;
        RECT 25.650 606.900 33.450 608.100 ;
        RECT 25.650 606.750 27.450 606.900 ;
        RECT 31.350 606.600 33.450 606.900 ;
        RECT 23.550 603.750 28.050 604.050 ;
        RECT 23.550 601.950 29.850 603.750 ;
        RECT 16.200 596.400 18.000 597.300 ;
        RECT 16.200 595.500 21.900 596.400 ;
        RECT 14.100 588.600 15.900 594.600 ;
        RECT 17.100 588.000 18.900 594.600 ;
        RECT 20.700 591.600 21.900 595.500 ;
        RECT 20.100 588.600 21.900 591.600 ;
        RECT 23.550 594.600 24.750 601.950 ;
        RECT 36.150 598.200 37.050 610.800 ;
        RECT 39.150 610.800 40.050 612.900 ;
        RECT 40.950 612.300 48.750 613.500 ;
        RECT 40.950 611.700 42.750 612.300 ;
        RECT 52.050 611.400 53.850 624.000 ;
        RECT 55.050 613.200 56.850 623.400 ;
        RECT 55.050 611.400 57.450 613.200 ;
        RECT 71.100 611.400 72.900 624.000 ;
        RECT 76.200 612.600 78.000 623.400 ;
        RECT 92.100 617.400 93.900 624.000 ;
        RECT 95.100 617.400 96.900 623.400 ;
        RECT 98.100 617.400 99.900 624.000 ;
        RECT 116.100 617.400 117.900 624.000 ;
        RECT 119.100 617.400 120.900 623.400 ;
        RECT 74.400 611.400 78.000 612.600 ;
        RECT 39.150 610.500 47.550 610.800 ;
        RECT 56.550 610.500 57.450 611.400 ;
        RECT 39.150 609.900 57.450 610.500 ;
        RECT 45.750 609.300 57.450 609.900 ;
        RECT 45.750 609.000 47.550 609.300 ;
        RECT 43.800 602.400 45.900 604.050 ;
        RECT 43.800 601.200 51.900 602.400 ;
        RECT 52.950 601.950 55.050 604.050 ;
        RECT 50.100 600.600 51.900 601.200 ;
        RECT 47.100 599.400 48.900 600.000 ;
        RECT 53.250 599.400 55.050 601.950 ;
        RECT 47.100 598.200 55.050 599.400 ;
        RECT 36.150 597.000 48.150 598.200 ;
        RECT 36.150 596.400 37.950 597.000 ;
        RECT 47.100 595.200 48.150 597.000 ;
        RECT 23.550 588.600 25.350 594.600 ;
        RECT 26.850 588.000 28.650 594.600 ;
        RECT 31.350 591.600 33.750 593.700 ;
        RECT 43.350 593.550 45.150 594.300 ;
        RECT 40.200 592.500 45.150 593.550 ;
        RECT 46.350 593.400 48.150 595.200 ;
        RECT 56.550 594.600 57.450 609.300 ;
        RECT 71.250 604.050 73.050 605.850 ;
        RECT 74.400 604.050 75.300 611.400 ;
        RECT 77.100 604.050 78.900 605.850 ;
        RECT 95.100 604.050 96.300 617.400 ;
        RECT 116.100 604.050 117.900 605.850 ;
        RECT 119.100 604.050 120.300 617.400 ;
        RECT 134.100 611.400 135.900 623.400 ;
        RECT 137.100 612.300 138.900 623.400 ;
        RECT 140.100 613.200 141.900 624.000 ;
        RECT 143.100 612.300 144.900 623.400 ;
        RECT 158.100 617.400 159.900 623.400 ;
        RECT 161.100 618.000 162.900 624.000 ;
        RECT 137.100 611.400 144.900 612.300 ;
        RECT 159.000 617.100 159.900 617.400 ;
        RECT 164.100 617.400 165.900 623.400 ;
        RECT 167.100 617.400 168.900 624.000 ;
        RECT 182.100 617.400 183.900 623.400 ;
        RECT 185.100 618.000 186.900 624.000 ;
        RECT 164.100 617.100 165.600 617.400 ;
        RECT 159.000 616.200 165.600 617.100 ;
        RECT 183.000 617.100 183.900 617.400 ;
        RECT 188.100 617.400 189.900 623.400 ;
        RECT 191.100 617.400 192.900 624.000 ;
        RECT 206.100 617.400 207.900 623.400 ;
        RECT 209.100 617.400 210.900 624.000 ;
        RECT 188.100 617.100 189.600 617.400 ;
        RECT 183.000 616.200 189.600 617.100 ;
        RECT 134.400 604.050 135.300 611.400 ;
        RECT 136.950 609.450 139.050 610.050 ;
        RECT 154.950 609.450 157.050 610.050 ;
        RECT 136.950 608.550 157.050 609.450 ;
        RECT 136.950 607.950 139.050 608.550 ;
        RECT 154.950 607.950 157.050 608.550 ;
        RECT 139.950 604.050 141.750 605.850 ;
        RECT 159.000 604.050 159.900 616.200 ;
        RECT 160.950 609.450 163.050 610.050 ;
        RECT 172.950 609.450 175.050 610.050 ;
        RECT 160.950 608.550 175.050 609.450 ;
        RECT 160.950 607.950 163.050 608.550 ;
        RECT 172.950 607.950 175.050 608.550 ;
        RECT 164.100 604.050 165.900 605.850 ;
        RECT 183.000 604.050 183.900 616.200 ;
        RECT 188.100 604.050 189.900 605.850 ;
        RECT 206.700 604.050 207.900 617.400 ;
        RECT 225.000 612.600 226.800 623.400 ;
        RECT 225.000 611.400 228.600 612.600 ;
        RECT 230.100 611.400 231.900 624.000 ;
        RECT 245.400 611.400 247.200 624.000 ;
        RECT 250.500 612.900 252.300 623.400 ;
        RECT 253.500 617.400 255.300 624.000 ;
        RECT 269.100 617.400 270.900 623.400 ;
        RECT 272.100 618.000 273.900 624.000 ;
        RECT 270.000 617.100 270.900 617.400 ;
        RECT 275.100 617.400 276.900 623.400 ;
        RECT 278.100 617.400 279.900 624.000 ;
        RECT 296.100 617.400 297.900 623.400 ;
        RECT 299.100 618.000 300.900 624.000 ;
        RECT 275.100 617.100 276.600 617.400 ;
        RECT 270.000 616.200 276.600 617.100 ;
        RECT 297.000 617.100 297.900 617.400 ;
        RECT 302.100 617.400 303.900 623.400 ;
        RECT 305.100 617.400 306.900 624.000 ;
        RECT 320.100 617.400 321.900 624.000 ;
        RECT 323.100 617.400 324.900 623.400 ;
        RECT 326.100 618.000 327.900 624.000 ;
        RECT 302.100 617.100 303.600 617.400 ;
        RECT 297.000 616.200 303.600 617.100 ;
        RECT 323.400 617.100 324.900 617.400 ;
        RECT 329.100 617.400 330.900 623.400 ;
        RECT 344.100 617.400 345.900 623.400 ;
        RECT 347.100 617.400 348.900 624.000 ;
        RECT 362.100 617.400 363.900 624.000 ;
        RECT 365.100 617.400 366.900 623.400 ;
        RECT 368.100 617.400 369.900 624.000 ;
        RECT 329.100 617.100 330.000 617.400 ;
        RECT 323.400 616.200 330.000 617.100 ;
        RECT 253.200 614.100 255.000 615.900 ;
        RECT 250.500 611.400 252.900 612.900 ;
        RECT 209.100 604.050 210.900 605.850 ;
        RECT 224.100 604.050 225.900 605.850 ;
        RECT 227.700 604.050 228.600 611.400 ;
        RECT 229.950 604.050 231.750 605.850 ;
        RECT 245.100 604.050 246.900 605.850 ;
        RECT 251.700 604.050 252.900 611.400 ;
        RECT 270.000 604.050 270.900 616.200 ;
        RECT 271.950 609.450 274.050 610.050 ;
        RECT 271.950 608.550 282.450 609.450 ;
        RECT 271.950 607.950 274.050 608.550 ;
        RECT 281.550 606.450 282.450 608.550 ;
        RECT 275.100 604.050 276.900 605.850 ;
        RECT 281.550 605.550 285.450 606.450 ;
        RECT 70.950 601.950 73.050 604.050 ;
        RECT 73.950 601.950 76.050 604.050 ;
        RECT 76.950 601.950 79.050 604.050 ;
        RECT 91.950 601.950 94.050 604.050 ;
        RECT 94.950 601.950 97.050 604.050 ;
        RECT 97.950 601.950 100.050 604.050 ;
        RECT 115.950 601.950 118.050 604.050 ;
        RECT 118.950 601.950 121.050 604.050 ;
        RECT 133.950 601.950 136.050 604.050 ;
        RECT 136.950 601.950 139.050 604.050 ;
        RECT 139.950 601.950 142.050 604.050 ;
        RECT 142.950 601.950 145.050 604.050 ;
        RECT 157.950 601.950 160.050 604.050 ;
        RECT 160.950 601.950 163.050 604.050 ;
        RECT 163.950 601.950 166.050 604.050 ;
        RECT 166.950 601.950 169.050 604.050 ;
        RECT 181.950 601.950 184.050 604.050 ;
        RECT 184.950 601.950 187.050 604.050 ;
        RECT 187.950 601.950 190.050 604.050 ;
        RECT 190.950 601.950 193.050 604.050 ;
        RECT 205.950 601.950 208.050 604.050 ;
        RECT 208.950 601.950 211.050 604.050 ;
        RECT 223.950 601.950 226.050 604.050 ;
        RECT 226.950 601.950 229.050 604.050 ;
        RECT 229.950 601.950 232.050 604.050 ;
        RECT 244.950 601.950 247.050 604.050 ;
        RECT 247.950 601.950 250.050 604.050 ;
        RECT 250.950 601.950 253.050 604.050 ;
        RECT 253.950 601.950 256.050 604.050 ;
        RECT 268.950 601.950 271.050 604.050 ;
        RECT 271.950 601.950 274.050 604.050 ;
        RECT 274.950 601.950 277.050 604.050 ;
        RECT 277.950 601.950 280.050 604.050 ;
        RECT 40.200 591.600 41.250 592.500 ;
        RECT 49.050 592.200 51.150 593.700 ;
        RECT 47.250 591.600 51.150 592.200 ;
        RECT 31.950 588.600 33.750 591.600 ;
        RECT 36.450 588.000 38.250 591.600 ;
        RECT 39.450 588.600 41.250 591.600 ;
        RECT 42.750 588.000 44.550 591.600 ;
        RECT 47.250 590.700 50.850 591.600 ;
        RECT 47.250 588.600 49.050 590.700 ;
        RECT 52.050 588.000 53.850 594.600 ;
        RECT 55.050 592.800 57.450 594.600 ;
        RECT 55.050 588.600 56.850 592.800 ;
        RECT 74.400 591.600 75.300 601.950 ;
        RECT 92.250 600.150 94.050 601.950 ;
        RECT 95.100 596.700 96.300 601.950 ;
        RECT 98.100 600.150 99.900 601.950 ;
        RECT 95.100 595.800 99.300 596.700 ;
        RECT 71.100 588.000 72.900 591.600 ;
        RECT 74.100 588.600 75.900 591.600 ;
        RECT 77.100 588.000 78.900 591.600 ;
        RECT 92.400 588.000 94.200 594.600 ;
        RECT 97.500 588.600 99.300 595.800 ;
        RECT 119.100 591.600 120.300 601.950 ;
        RECT 134.400 594.600 135.300 601.950 ;
        RECT 136.950 600.150 138.750 601.950 ;
        RECT 143.100 600.150 144.900 601.950 ;
        RECT 159.000 598.200 159.900 601.950 ;
        RECT 161.100 600.150 162.900 601.950 ;
        RECT 167.100 600.150 168.900 601.950 ;
        RECT 183.000 598.200 183.900 601.950 ;
        RECT 185.100 600.150 186.900 601.950 ;
        RECT 191.100 600.150 192.900 601.950 ;
        RECT 159.000 597.000 162.300 598.200 ;
        RECT 134.400 593.400 139.500 594.600 ;
        RECT 116.100 588.000 117.900 591.600 ;
        RECT 119.100 588.600 120.900 591.600 ;
        RECT 134.700 588.000 136.500 591.600 ;
        RECT 137.700 588.600 139.500 593.400 ;
        RECT 142.200 588.000 144.000 594.600 ;
        RECT 160.500 588.600 162.300 597.000 ;
        RECT 167.100 588.000 168.900 597.600 ;
        RECT 183.000 597.000 186.300 598.200 ;
        RECT 184.500 588.600 186.300 597.000 ;
        RECT 191.100 588.000 192.900 597.600 ;
        RECT 206.700 591.600 207.900 601.950 ;
        RECT 227.700 591.600 228.600 601.950 ;
        RECT 248.100 600.150 249.900 601.950 ;
        RECT 251.700 597.600 252.900 601.950 ;
        RECT 254.100 600.150 255.900 601.950 ;
        RECT 270.000 598.200 270.900 601.950 ;
        RECT 272.100 600.150 273.900 601.950 ;
        RECT 278.100 600.150 279.900 601.950 ;
        RECT 251.700 596.700 255.300 597.600 ;
        RECT 270.000 597.000 273.300 598.200 ;
        RECT 284.550 598.050 285.450 605.550 ;
        RECT 297.000 604.050 297.900 616.200 ;
        RECT 302.100 604.050 303.900 605.850 ;
        RECT 323.100 604.050 324.900 605.850 ;
        RECT 329.100 604.050 330.000 616.200 ;
        RECT 331.950 606.450 336.000 607.050 ;
        RECT 331.950 604.950 336.450 606.450 ;
        RECT 295.950 601.950 298.050 604.050 ;
        RECT 298.950 601.950 301.050 604.050 ;
        RECT 301.950 601.950 304.050 604.050 ;
        RECT 304.950 601.950 307.050 604.050 ;
        RECT 319.950 601.950 322.050 604.050 ;
        RECT 322.950 601.950 325.050 604.050 ;
        RECT 325.950 601.950 328.050 604.050 ;
        RECT 328.950 601.950 331.050 604.050 ;
        RECT 297.000 598.200 297.900 601.950 ;
        RECT 299.100 600.150 300.900 601.950 ;
        RECT 305.100 600.150 306.900 601.950 ;
        RECT 320.100 600.150 321.900 601.950 ;
        RECT 326.100 600.150 327.900 601.950 ;
        RECT 329.100 598.200 330.000 601.950 ;
        RECT 335.550 600.450 336.450 604.950 ;
        RECT 344.700 604.050 345.900 617.400 ;
        RECT 347.100 604.050 348.900 605.850 ;
        RECT 365.700 604.050 366.900 617.400 ;
        RECT 383.400 611.400 385.200 624.000 ;
        RECT 388.500 612.900 390.300 623.400 ;
        RECT 391.500 617.400 393.300 624.000 ;
        RECT 407.100 617.400 408.900 624.000 ;
        RECT 410.100 617.400 411.900 623.400 ;
        RECT 413.100 617.400 414.900 624.000 ;
        RECT 428.100 617.400 429.900 624.000 ;
        RECT 431.100 617.400 432.900 623.400 ;
        RECT 446.100 617.400 447.900 624.000 ;
        RECT 449.100 617.400 450.900 623.400 ;
        RECT 452.100 618.000 453.900 624.000 ;
        RECT 391.200 614.100 393.000 615.900 ;
        RECT 388.500 611.400 390.900 612.900 ;
        RECT 383.100 604.050 384.900 605.850 ;
        RECT 389.700 604.050 390.900 611.400 ;
        RECT 410.100 604.050 411.300 617.400 ;
        RECT 428.100 604.050 429.900 605.850 ;
        RECT 431.100 604.050 432.300 617.400 ;
        RECT 449.400 617.100 450.900 617.400 ;
        RECT 455.100 617.400 456.900 623.400 ;
        RECT 470.100 617.400 471.900 624.000 ;
        RECT 473.100 617.400 474.900 623.400 ;
        RECT 476.100 617.400 477.900 624.000 ;
        RECT 491.100 617.400 492.900 624.000 ;
        RECT 494.100 617.400 495.900 623.400 ;
        RECT 455.100 617.100 456.000 617.400 ;
        RECT 449.400 616.200 456.000 617.100 ;
        RECT 449.100 604.050 450.900 605.850 ;
        RECT 455.100 604.050 456.000 616.200 ;
        RECT 457.950 606.450 460.050 610.050 ;
        RECT 457.950 606.000 462.450 606.450 ;
        RECT 458.550 605.550 462.450 606.000 ;
        RECT 343.950 601.950 346.050 604.050 ;
        RECT 346.950 601.950 349.050 604.050 ;
        RECT 361.950 601.950 364.050 604.050 ;
        RECT 364.950 601.950 367.050 604.050 ;
        RECT 367.950 601.950 370.050 604.050 ;
        RECT 382.950 601.950 385.050 604.050 ;
        RECT 385.950 601.950 388.050 604.050 ;
        RECT 388.950 601.950 391.050 604.050 ;
        RECT 391.950 601.950 394.050 604.050 ;
        RECT 406.950 601.950 409.050 604.050 ;
        RECT 409.950 601.950 412.050 604.050 ;
        RECT 412.950 601.950 415.050 604.050 ;
        RECT 427.950 601.950 430.050 604.050 ;
        RECT 430.950 601.950 433.050 604.050 ;
        RECT 445.950 601.950 448.050 604.050 ;
        RECT 448.950 601.950 451.050 604.050 ;
        RECT 451.950 601.950 454.050 604.050 ;
        RECT 454.950 601.950 457.050 604.050 ;
        RECT 340.950 600.450 343.050 601.050 ;
        RECT 335.550 599.550 343.050 600.450 ;
        RECT 340.950 598.950 343.050 599.550 ;
        RECT 284.550 597.900 288.000 598.050 ;
        RECT 245.100 593.700 252.900 595.050 ;
        RECT 206.100 588.600 207.900 591.600 ;
        RECT 209.100 588.000 210.900 591.600 ;
        RECT 224.100 588.000 225.900 591.600 ;
        RECT 227.100 588.600 228.900 591.600 ;
        RECT 230.100 588.000 231.900 591.600 ;
        RECT 245.100 588.600 246.900 593.700 ;
        RECT 248.100 588.000 249.900 592.800 ;
        RECT 251.100 588.600 252.900 593.700 ;
        RECT 254.100 594.600 255.300 596.700 ;
        RECT 254.100 588.600 255.900 594.600 ;
        RECT 271.500 588.600 273.300 597.000 ;
        RECT 278.100 588.000 279.900 597.600 ;
        RECT 284.550 596.550 289.050 597.900 ;
        RECT 297.000 597.000 300.300 598.200 ;
        RECT 285.000 595.950 289.050 596.550 ;
        RECT 286.950 595.800 289.050 595.950 ;
        RECT 298.500 588.600 300.300 597.000 ;
        RECT 305.100 588.000 306.900 597.600 ;
        RECT 320.100 588.000 321.900 597.600 ;
        RECT 326.700 597.000 330.000 598.200 ;
        RECT 326.700 588.600 328.500 597.000 ;
        RECT 344.700 591.600 345.900 601.950 ;
        RECT 362.100 600.150 363.900 601.950 ;
        RECT 365.700 596.700 366.900 601.950 ;
        RECT 367.950 600.150 369.750 601.950 ;
        RECT 386.100 600.150 387.900 601.950 ;
        RECT 389.700 597.600 390.900 601.950 ;
        RECT 392.100 600.150 393.900 601.950 ;
        RECT 407.250 600.150 409.050 601.950 ;
        RECT 389.700 596.700 393.300 597.600 ;
        RECT 362.700 595.800 366.900 596.700 ;
        RECT 344.100 588.600 345.900 591.600 ;
        RECT 347.100 588.000 348.900 591.600 ;
        RECT 362.700 588.600 364.500 595.800 ;
        RECT 367.800 588.000 369.600 594.600 ;
        RECT 383.100 593.700 390.900 595.050 ;
        RECT 383.100 588.600 384.900 593.700 ;
        RECT 386.100 588.000 387.900 592.800 ;
        RECT 389.100 588.600 390.900 593.700 ;
        RECT 392.100 594.600 393.300 596.700 ;
        RECT 410.100 596.700 411.300 601.950 ;
        RECT 413.100 600.150 414.900 601.950 ;
        RECT 410.100 595.800 414.300 596.700 ;
        RECT 392.100 588.600 393.900 594.600 ;
        RECT 407.400 588.000 409.200 594.600 ;
        RECT 412.500 588.600 414.300 595.800 ;
        RECT 431.100 591.600 432.300 601.950 ;
        RECT 446.100 600.150 447.900 601.950 ;
        RECT 452.100 600.150 453.900 601.950 ;
        RECT 455.100 598.200 456.000 601.950 ;
        RECT 461.550 601.050 462.450 605.550 ;
        RECT 473.100 604.050 474.300 617.400 ;
        RECT 491.100 604.050 492.900 605.850 ;
        RECT 494.100 604.050 495.300 617.400 ;
        RECT 509.100 611.400 510.900 623.400 ;
        RECT 512.100 612.300 513.900 623.400 ;
        RECT 515.100 613.200 516.900 624.000 ;
        RECT 518.100 612.300 519.900 623.400 ;
        RECT 512.100 611.400 519.900 612.300 ;
        RECT 533.400 611.400 535.200 624.000 ;
        RECT 538.500 612.900 540.300 623.400 ;
        RECT 541.500 617.400 543.300 624.000 ;
        RECT 541.200 614.100 543.000 615.900 ;
        RECT 538.500 611.400 540.900 612.900 ;
        RECT 509.400 604.050 510.300 611.400 ;
        RECT 511.950 609.450 514.050 610.050 ;
        RECT 535.950 609.450 538.050 610.200 ;
        RECT 511.950 608.550 538.050 609.450 ;
        RECT 511.950 607.950 514.050 608.550 ;
        RECT 535.950 608.100 538.050 608.550 ;
        RECT 514.950 604.050 516.750 605.850 ;
        RECT 533.100 604.050 534.900 605.850 ;
        RECT 539.700 604.050 540.900 611.400 ;
        RECT 541.950 612.450 544.050 612.900 ;
        RECT 547.950 612.450 550.050 613.050 ;
        RECT 541.950 611.550 550.050 612.450 ;
        RECT 541.950 610.800 544.050 611.550 ;
        RECT 547.950 610.950 550.050 611.550 ;
        RECT 557.100 611.400 558.900 624.000 ;
        RECT 562.200 612.600 564.000 623.400 ;
        RECT 578.100 617.400 579.900 624.000 ;
        RECT 581.100 617.400 582.900 623.400 ;
        RECT 560.400 611.400 564.000 612.600 ;
        RECT 557.250 604.050 559.050 605.850 ;
        RECT 560.400 604.050 561.300 611.400 ;
        RECT 563.100 604.050 564.900 605.850 ;
        RECT 469.950 601.950 472.050 604.050 ;
        RECT 472.950 601.950 475.050 604.050 ;
        RECT 475.950 601.950 478.050 604.050 ;
        RECT 490.950 601.950 493.050 604.050 ;
        RECT 493.950 601.950 496.050 604.050 ;
        RECT 508.950 601.950 511.050 604.050 ;
        RECT 511.950 601.950 514.050 604.050 ;
        RECT 514.950 601.950 517.050 604.050 ;
        RECT 517.950 601.950 520.050 604.050 ;
        RECT 532.950 601.950 535.050 604.050 ;
        RECT 535.950 601.950 538.050 604.050 ;
        RECT 538.950 601.950 541.050 604.050 ;
        RECT 541.950 601.950 544.050 604.050 ;
        RECT 556.950 601.950 559.050 604.050 ;
        RECT 559.950 601.950 562.050 604.050 ;
        RECT 562.950 601.950 565.050 604.050 ;
        RECT 578.100 601.950 580.200 604.050 ;
        RECT 457.950 599.550 462.450 601.050 ;
        RECT 470.250 600.150 472.050 601.950 ;
        RECT 457.950 598.950 462.000 599.550 ;
        RECT 428.100 588.000 429.900 591.600 ;
        RECT 431.100 588.600 432.900 591.600 ;
        RECT 446.100 588.000 447.900 597.600 ;
        RECT 452.700 597.000 456.000 598.200 ;
        RECT 452.700 588.600 454.500 597.000 ;
        RECT 473.100 596.700 474.300 601.950 ;
        RECT 476.100 600.150 477.900 601.950 ;
        RECT 473.100 595.800 477.300 596.700 ;
        RECT 470.400 588.000 472.200 594.600 ;
        RECT 475.500 588.600 477.300 595.800 ;
        RECT 494.100 591.600 495.300 601.950 ;
        RECT 509.400 594.600 510.300 601.950 ;
        RECT 511.950 600.150 513.750 601.950 ;
        RECT 518.100 600.150 519.900 601.950 ;
        RECT 536.100 600.150 537.900 601.950 ;
        RECT 539.700 597.600 540.900 601.950 ;
        RECT 542.100 600.150 543.900 601.950 ;
        RECT 539.700 596.700 543.300 597.600 ;
        RECT 509.400 593.400 514.500 594.600 ;
        RECT 491.100 588.000 492.900 591.600 ;
        RECT 494.100 588.600 495.900 591.600 ;
        RECT 509.700 588.000 511.500 591.600 ;
        RECT 512.700 588.600 514.500 593.400 ;
        RECT 517.200 588.000 519.000 594.600 ;
        RECT 533.100 593.700 540.900 595.050 ;
        RECT 533.100 588.600 534.900 593.700 ;
        RECT 536.100 588.000 537.900 592.800 ;
        RECT 539.100 588.600 540.900 593.700 ;
        RECT 542.100 594.600 543.300 596.700 ;
        RECT 542.100 588.600 543.900 594.600 ;
        RECT 560.400 591.600 561.300 601.950 ;
        RECT 578.250 600.150 580.050 601.950 ;
        RECT 581.100 597.300 582.000 617.400 ;
        RECT 584.100 612.000 585.900 624.000 ;
        RECT 587.100 611.400 588.900 623.400 ;
        RECT 605.100 617.400 606.900 624.000 ;
        RECT 608.100 617.400 609.900 623.400 ;
        RECT 611.100 618.000 612.900 624.000 ;
        RECT 608.400 617.100 609.900 617.400 ;
        RECT 614.100 617.400 615.900 623.400 ;
        RECT 629.100 617.400 630.900 623.400 ;
        RECT 632.100 618.000 633.900 624.000 ;
        RECT 614.100 617.100 615.000 617.400 ;
        RECT 608.400 616.200 615.000 617.100 ;
        RECT 583.200 604.050 585.000 605.850 ;
        RECT 587.400 604.050 588.300 611.400 ;
        RECT 608.100 604.050 609.900 605.850 ;
        RECT 614.100 604.050 615.000 616.200 ;
        RECT 630.000 617.100 630.900 617.400 ;
        RECT 635.100 617.400 636.900 623.400 ;
        RECT 638.100 617.400 639.900 624.000 ;
        RECT 653.100 617.400 654.900 623.400 ;
        RECT 656.100 618.000 657.900 624.000 ;
        RECT 635.100 617.100 636.600 617.400 ;
        RECT 630.000 616.200 636.600 617.100 ;
        RECT 654.000 617.100 654.900 617.400 ;
        RECT 659.100 617.400 660.900 623.400 ;
        RECT 662.100 617.400 663.900 624.000 ;
        RECT 659.100 617.100 660.600 617.400 ;
        RECT 654.000 616.200 660.600 617.100 ;
        RECT 622.950 607.950 625.050 610.050 ;
        RECT 583.500 601.950 585.600 604.050 ;
        RECT 586.800 601.950 588.900 604.050 ;
        RECT 604.950 601.950 607.050 604.050 ;
        RECT 607.950 601.950 610.050 604.050 ;
        RECT 610.950 601.950 613.050 604.050 ;
        RECT 613.950 601.950 616.050 604.050 ;
        RECT 578.100 596.400 586.500 597.300 ;
        RECT 557.100 588.000 558.900 591.600 ;
        RECT 560.100 588.600 561.900 591.600 ;
        RECT 563.100 588.000 564.900 591.600 ;
        RECT 578.100 588.600 579.900 596.400 ;
        RECT 584.700 595.500 586.500 596.400 ;
        RECT 587.400 594.600 588.300 601.950 ;
        RECT 605.100 600.150 606.900 601.950 ;
        RECT 611.100 600.150 612.900 601.950 ;
        RECT 614.100 598.200 615.000 601.950 ;
        RECT 623.550 601.050 624.450 607.950 ;
        RECT 630.000 604.050 630.900 616.200 ;
        RECT 635.100 604.050 636.900 605.850 ;
        RECT 654.000 604.050 654.900 616.200 ;
        RECT 677.100 612.300 678.900 623.400 ;
        RECT 680.100 613.200 681.900 624.000 ;
        RECT 683.100 612.300 684.900 623.400 ;
        RECT 677.100 611.400 684.900 612.300 ;
        RECT 686.100 611.400 687.900 623.400 ;
        RECT 704.100 611.400 705.900 623.400 ;
        RECT 707.100 612.300 708.900 623.400 ;
        RECT 710.100 613.200 711.900 624.000 ;
        RECT 713.100 612.300 714.900 623.400 ;
        RECT 728.100 617.400 729.900 623.400 ;
        RECT 731.100 618.000 732.900 624.000 ;
        RECT 707.100 611.400 714.900 612.300 ;
        RECT 729.000 617.100 729.900 617.400 ;
        RECT 734.100 617.400 735.900 623.400 ;
        RECT 737.100 617.400 738.900 624.000 ;
        RECT 755.100 617.400 756.900 623.400 ;
        RECT 758.100 618.000 759.900 624.000 ;
        RECT 734.100 617.100 735.600 617.400 ;
        RECT 729.000 616.200 735.600 617.100 ;
        RECT 756.000 617.100 756.900 617.400 ;
        RECT 761.100 617.400 762.900 623.400 ;
        RECT 764.100 617.400 765.900 624.000 ;
        RECT 779.700 617.400 781.500 624.000 ;
        RECT 761.100 617.100 762.600 617.400 ;
        RECT 756.000 616.200 762.600 617.100 ;
        RECT 667.950 609.450 670.050 610.050 ;
        RECT 682.950 609.450 685.050 610.050 ;
        RECT 667.950 608.550 685.050 609.450 ;
        RECT 667.950 607.950 670.050 608.550 ;
        RECT 682.950 607.950 685.050 608.550 ;
        RECT 659.100 604.050 660.900 605.850 ;
        RECT 680.250 604.050 682.050 605.850 ;
        RECT 686.700 604.050 687.600 611.400 ;
        RECT 704.400 604.050 705.300 611.400 ;
        RECT 709.950 604.050 711.750 605.850 ;
        RECT 729.000 604.050 729.900 616.200 ;
        RECT 734.100 604.050 735.900 605.850 ;
        RECT 756.000 604.050 756.900 616.200 ;
        RECT 780.000 614.100 781.800 615.900 ;
        RECT 782.700 612.900 784.500 623.400 ;
        RECT 782.100 611.400 784.500 612.900 ;
        RECT 787.800 611.400 789.600 624.000 ;
        RECT 803.700 617.400 805.500 624.000 ;
        RECT 804.000 614.100 805.800 615.900 ;
        RECT 806.700 612.900 808.500 623.400 ;
        RECT 806.100 611.400 808.500 612.900 ;
        RECT 811.800 611.400 813.600 624.000 ;
        RECT 827.100 611.400 828.900 623.400 ;
        RECT 830.100 612.000 831.900 624.000 ;
        RECT 833.100 617.400 834.900 623.400 ;
        RECT 836.100 617.400 837.900 624.000 ;
        RECT 761.100 604.050 762.900 605.850 ;
        RECT 782.100 604.050 783.300 611.400 ;
        RECT 787.950 609.450 790.050 610.050 ;
        RECT 796.950 609.450 799.050 610.050 ;
        RECT 802.950 609.450 805.050 610.050 ;
        RECT 787.950 608.550 805.050 609.450 ;
        RECT 787.950 607.950 790.050 608.550 ;
        RECT 796.950 607.950 799.050 608.550 ;
        RECT 802.950 607.950 805.050 608.550 ;
        RECT 788.100 604.050 789.900 605.850 ;
        RECT 806.100 604.050 807.300 611.400 ;
        RECT 812.100 604.050 813.900 605.850 ;
        RECT 827.700 604.050 828.600 611.400 ;
        RECT 831.000 604.050 832.800 605.850 ;
        RECT 628.950 601.950 631.050 604.050 ;
        RECT 631.950 601.950 634.050 604.050 ;
        RECT 634.950 601.950 637.050 604.050 ;
        RECT 637.950 601.950 640.050 604.050 ;
        RECT 652.950 601.950 655.050 604.050 ;
        RECT 655.950 601.950 658.050 604.050 ;
        RECT 658.950 601.950 661.050 604.050 ;
        RECT 661.950 601.950 664.050 604.050 ;
        RECT 676.950 601.950 679.050 604.050 ;
        RECT 679.950 601.950 682.050 604.050 ;
        RECT 682.950 601.950 685.050 604.050 ;
        RECT 685.950 601.950 688.050 604.050 ;
        RECT 703.950 601.950 706.050 604.050 ;
        RECT 706.950 601.950 709.050 604.050 ;
        RECT 709.950 601.950 712.050 604.050 ;
        RECT 712.950 601.950 715.050 604.050 ;
        RECT 727.950 601.950 730.050 604.050 ;
        RECT 730.950 601.950 733.050 604.050 ;
        RECT 733.950 601.950 736.050 604.050 ;
        RECT 736.950 601.950 739.050 604.050 ;
        RECT 754.950 601.950 757.050 604.050 ;
        RECT 757.950 601.950 760.050 604.050 ;
        RECT 760.950 601.950 763.050 604.050 ;
        RECT 763.950 601.950 766.050 604.050 ;
        RECT 778.950 601.950 781.050 604.050 ;
        RECT 781.950 601.950 784.050 604.050 ;
        RECT 784.950 601.950 787.050 604.050 ;
        RECT 787.950 601.950 790.050 604.050 ;
        RECT 802.950 601.950 805.050 604.050 ;
        RECT 805.950 601.950 808.050 604.050 ;
        RECT 808.950 601.950 811.050 604.050 ;
        RECT 811.950 601.950 814.050 604.050 ;
        RECT 827.100 601.950 829.200 604.050 ;
        RECT 830.400 601.950 832.500 604.050 ;
        RECT 623.550 599.550 628.050 601.050 ;
        RECT 624.000 598.950 628.050 599.550 ;
        RECT 582.600 588.000 584.400 594.600 ;
        RECT 585.600 592.800 588.300 594.600 ;
        RECT 585.600 588.600 587.400 592.800 ;
        RECT 605.100 588.000 606.900 597.600 ;
        RECT 611.700 597.000 615.000 598.200 ;
        RECT 630.000 598.200 630.900 601.950 ;
        RECT 632.100 600.150 633.900 601.950 ;
        RECT 638.100 600.150 639.900 601.950 ;
        RECT 654.000 598.200 654.900 601.950 ;
        RECT 656.100 600.150 657.900 601.950 ;
        RECT 662.100 600.150 663.900 601.950 ;
        RECT 677.100 600.150 678.900 601.950 ;
        RECT 683.250 600.150 685.050 601.950 ;
        RECT 630.000 597.000 633.300 598.200 ;
        RECT 611.700 588.600 613.500 597.000 ;
        RECT 631.500 588.600 633.300 597.000 ;
        RECT 638.100 588.000 639.900 597.600 ;
        RECT 654.000 597.000 657.300 598.200 ;
        RECT 655.500 588.600 657.300 597.000 ;
        RECT 662.100 588.000 663.900 597.600 ;
        RECT 686.700 594.600 687.600 601.950 ;
        RECT 678.000 588.000 679.800 594.600 ;
        RECT 682.500 593.400 687.600 594.600 ;
        RECT 704.400 594.600 705.300 601.950 ;
        RECT 706.950 600.150 708.750 601.950 ;
        RECT 713.100 600.150 714.900 601.950 ;
        RECT 729.000 598.200 729.900 601.950 ;
        RECT 731.100 600.150 732.900 601.950 ;
        RECT 737.100 600.150 738.900 601.950 ;
        RECT 756.000 598.200 756.900 601.950 ;
        RECT 758.100 600.150 759.900 601.950 ;
        RECT 764.100 600.150 765.900 601.950 ;
        RECT 779.100 600.150 780.900 601.950 ;
        RECT 729.000 597.000 732.300 598.200 ;
        RECT 704.400 593.400 709.500 594.600 ;
        RECT 682.500 588.600 684.300 593.400 ;
        RECT 685.500 588.000 687.300 591.600 ;
        RECT 704.700 588.000 706.500 591.600 ;
        RECT 707.700 588.600 709.500 593.400 ;
        RECT 712.200 588.000 714.000 594.600 ;
        RECT 730.500 588.600 732.300 597.000 ;
        RECT 737.100 588.000 738.900 597.600 ;
        RECT 756.000 597.000 759.300 598.200 ;
        RECT 782.100 597.600 783.300 601.950 ;
        RECT 785.100 600.150 786.900 601.950 ;
        RECT 803.100 600.150 804.900 601.950 ;
        RECT 806.100 597.600 807.300 601.950 ;
        RECT 809.100 600.150 810.900 601.950 ;
        RECT 757.500 588.600 759.300 597.000 ;
        RECT 764.100 588.000 765.900 597.600 ;
        RECT 779.700 596.700 783.300 597.600 ;
        RECT 803.700 596.700 807.300 597.600 ;
        RECT 779.700 594.600 780.900 596.700 ;
        RECT 779.100 588.600 780.900 594.600 ;
        RECT 782.100 593.700 789.900 595.050 ;
        RECT 803.700 594.600 804.900 596.700 ;
        RECT 782.100 588.600 783.900 593.700 ;
        RECT 785.100 588.000 786.900 592.800 ;
        RECT 788.100 588.600 789.900 593.700 ;
        RECT 803.100 588.600 804.900 594.600 ;
        RECT 806.100 593.700 813.900 595.050 ;
        RECT 806.100 588.600 807.900 593.700 ;
        RECT 809.100 588.000 810.900 592.800 ;
        RECT 812.100 588.600 813.900 593.700 ;
        RECT 827.700 594.600 828.600 601.950 ;
        RECT 834.000 597.300 834.900 617.400 ;
        RECT 851.100 611.400 852.900 623.400 ;
        RECT 854.100 612.300 855.900 623.400 ;
        RECT 857.100 613.200 858.900 624.000 ;
        RECT 860.100 612.300 861.900 623.400 ;
        RECT 854.100 611.400 861.900 612.300 ;
        RECT 875.400 611.400 877.200 624.000 ;
        RECT 880.500 612.900 882.300 623.400 ;
        RECT 883.500 617.400 885.300 624.000 ;
        RECT 883.200 614.100 885.000 615.900 ;
        RECT 880.500 611.400 882.900 612.900 ;
        RECT 851.400 604.050 852.300 611.400 ;
        RECT 856.950 604.050 858.750 605.850 ;
        RECT 875.100 604.050 876.900 605.850 ;
        RECT 881.700 604.050 882.900 611.400 ;
        RECT 835.800 601.950 837.900 604.050 ;
        RECT 850.950 601.950 853.050 604.050 ;
        RECT 853.950 601.950 856.050 604.050 ;
        RECT 856.950 601.950 859.050 604.050 ;
        RECT 859.950 601.950 862.050 604.050 ;
        RECT 874.950 601.950 877.050 604.050 ;
        RECT 877.950 601.950 880.050 604.050 ;
        RECT 880.950 601.950 883.050 604.050 ;
        RECT 883.950 601.950 886.050 604.050 ;
        RECT 835.950 600.150 837.750 601.950 ;
        RECT 829.500 596.400 837.900 597.300 ;
        RECT 829.500 595.500 831.300 596.400 ;
        RECT 827.700 592.800 830.400 594.600 ;
        RECT 828.600 588.600 830.400 592.800 ;
        RECT 831.600 588.000 833.400 594.600 ;
        RECT 836.100 588.600 837.900 596.400 ;
        RECT 851.400 594.600 852.300 601.950 ;
        RECT 853.950 600.150 855.750 601.950 ;
        RECT 860.100 600.150 861.900 601.950 ;
        RECT 878.100 600.150 879.900 601.950 ;
        RECT 881.700 597.600 882.900 601.950 ;
        RECT 884.100 600.150 885.900 601.950 ;
        RECT 881.700 596.700 885.300 597.600 ;
        RECT 851.400 593.400 856.500 594.600 ;
        RECT 851.700 588.000 853.500 591.600 ;
        RECT 854.700 588.600 856.500 593.400 ;
        RECT 859.200 588.000 861.000 594.600 ;
        RECT 875.100 593.700 882.900 595.050 ;
        RECT 875.100 588.600 876.900 593.700 ;
        RECT 878.100 588.000 879.900 592.800 ;
        RECT 881.100 588.600 882.900 593.700 ;
        RECT 884.100 594.600 885.300 596.700 ;
        RECT 884.100 588.600 885.900 594.600 ;
        RECT 14.100 578.400 15.900 584.400 ;
        RECT 17.100 578.400 18.900 585.000 ;
        RECT 20.100 581.400 21.900 584.400 ;
        RECT 14.100 571.050 15.300 578.400 ;
        RECT 20.700 577.500 21.900 581.400 ;
        RECT 16.200 576.600 21.900 577.500 ;
        RECT 23.550 578.400 25.350 584.400 ;
        RECT 26.850 578.400 28.650 585.000 ;
        RECT 31.950 581.400 33.750 584.400 ;
        RECT 36.450 581.400 38.250 585.000 ;
        RECT 39.450 581.400 41.250 584.400 ;
        RECT 42.750 581.400 44.550 585.000 ;
        RECT 47.250 582.300 49.050 584.400 ;
        RECT 47.250 581.400 50.850 582.300 ;
        RECT 31.350 579.300 33.750 581.400 ;
        RECT 40.200 580.500 41.250 581.400 ;
        RECT 47.250 580.800 51.150 581.400 ;
        RECT 40.200 579.450 45.150 580.500 ;
        RECT 43.350 578.700 45.150 579.450 ;
        RECT 16.200 575.700 18.000 576.600 ;
        RECT 14.100 568.950 16.200 571.050 ;
        RECT 14.100 561.600 15.300 568.950 ;
        RECT 17.100 564.300 18.000 575.700 ;
        RECT 23.550 571.050 24.750 578.400 ;
        RECT 46.350 577.800 48.150 579.600 ;
        RECT 49.050 579.300 51.150 580.800 ;
        RECT 52.050 578.400 53.850 585.000 ;
        RECT 55.050 580.200 56.850 584.400 ;
        RECT 71.100 581.400 72.900 585.000 ;
        RECT 74.100 581.400 75.900 584.400 ;
        RECT 77.100 581.400 78.900 585.000 ;
        RECT 55.050 578.400 57.450 580.200 ;
        RECT 36.150 576.000 37.950 576.600 ;
        RECT 47.100 576.000 48.150 577.800 ;
        RECT 36.150 574.800 48.150 576.000 ;
        RECT 19.500 568.950 21.600 571.050 ;
        RECT 19.800 567.150 21.600 568.950 ;
        RECT 23.550 569.250 29.850 571.050 ;
        RECT 23.550 568.950 28.050 569.250 ;
        RECT 16.200 563.400 18.000 564.300 ;
        RECT 16.200 562.500 21.900 563.400 ;
        RECT 14.100 549.600 15.900 561.600 ;
        RECT 17.100 549.000 18.900 559.800 ;
        RECT 20.700 555.600 21.900 562.500 ;
        RECT 20.100 549.600 21.900 555.600 ;
        RECT 23.550 561.600 24.750 568.950 ;
        RECT 25.650 566.100 27.450 566.250 ;
        RECT 31.350 566.100 33.450 566.400 ;
        RECT 25.650 564.900 33.450 566.100 ;
        RECT 25.650 564.450 27.450 564.900 ;
        RECT 31.350 564.300 33.450 564.900 ;
        RECT 36.150 562.200 37.050 574.800 ;
        RECT 47.100 573.600 55.050 574.800 ;
        RECT 47.100 573.000 48.900 573.600 ;
        RECT 50.100 571.800 51.900 572.400 ;
        RECT 43.800 570.600 51.900 571.800 ;
        RECT 53.250 571.050 55.050 573.600 ;
        RECT 43.800 568.950 45.900 570.600 ;
        RECT 52.950 568.950 55.050 571.050 ;
        RECT 45.750 563.700 47.550 564.000 ;
        RECT 56.550 563.700 57.450 578.400 ;
        RECT 74.400 571.050 75.300 581.400 ;
        RECT 80.550 578.400 82.350 584.400 ;
        RECT 83.850 578.400 85.650 585.000 ;
        RECT 88.950 581.400 90.750 584.400 ;
        RECT 93.450 581.400 95.250 585.000 ;
        RECT 96.450 581.400 98.250 584.400 ;
        RECT 99.750 581.400 101.550 585.000 ;
        RECT 104.250 582.300 106.050 584.400 ;
        RECT 104.250 581.400 107.850 582.300 ;
        RECT 88.350 579.300 90.750 581.400 ;
        RECT 97.200 580.500 98.250 581.400 ;
        RECT 104.250 580.800 108.150 581.400 ;
        RECT 97.200 579.450 102.150 580.500 ;
        RECT 100.350 578.700 102.150 579.450 ;
        RECT 80.550 571.050 81.750 578.400 ;
        RECT 103.350 577.800 105.150 579.600 ;
        RECT 106.050 579.300 108.150 580.800 ;
        RECT 109.050 578.400 110.850 585.000 ;
        RECT 112.050 580.200 113.850 584.400 ;
        RECT 128.100 581.400 129.900 585.000 ;
        RECT 131.100 581.400 132.900 584.400 ;
        RECT 134.100 581.400 135.900 585.000 ;
        RECT 149.100 581.400 150.900 585.000 ;
        RECT 152.100 581.400 153.900 584.400 ;
        RECT 112.050 578.400 114.450 580.200 ;
        RECT 93.150 576.000 94.950 576.600 ;
        RECT 104.100 576.000 105.150 577.800 ;
        RECT 93.150 574.800 105.150 576.000 ;
        RECT 70.950 568.950 73.050 571.050 ;
        RECT 73.950 568.950 76.050 571.050 ;
        RECT 76.950 568.950 79.050 571.050 ;
        RECT 80.550 569.250 86.850 571.050 ;
        RECT 80.550 568.950 85.050 569.250 ;
        RECT 71.250 567.150 73.050 568.950 ;
        RECT 45.750 563.100 57.450 563.700 ;
        RECT 23.550 549.600 25.350 561.600 ;
        RECT 26.550 549.000 28.350 561.600 ;
        RECT 32.250 561.300 37.050 562.200 ;
        RECT 39.150 562.500 57.450 563.100 ;
        RECT 39.150 562.200 47.550 562.500 ;
        RECT 32.250 560.400 33.450 561.300 ;
        RECT 30.450 558.600 33.450 560.400 ;
        RECT 34.350 560.100 36.150 560.400 ;
        RECT 39.150 560.100 40.050 562.200 ;
        RECT 56.550 561.600 57.450 562.500 ;
        RECT 74.400 561.600 75.300 568.950 ;
        RECT 77.100 567.150 78.900 568.950 ;
        RECT 80.550 561.600 81.750 568.950 ;
        RECT 82.650 566.100 84.450 566.250 ;
        RECT 88.350 566.100 90.450 566.400 ;
        RECT 82.650 564.900 90.450 566.100 ;
        RECT 82.650 564.450 84.450 564.900 ;
        RECT 88.350 564.300 90.450 564.900 ;
        RECT 93.150 562.200 94.050 574.800 ;
        RECT 104.100 573.600 112.050 574.800 ;
        RECT 104.100 573.000 105.900 573.600 ;
        RECT 107.100 571.800 108.900 572.400 ;
        RECT 100.800 570.600 108.900 571.800 ;
        RECT 110.250 571.050 112.050 573.600 ;
        RECT 100.800 568.950 102.900 570.600 ;
        RECT 109.950 568.950 112.050 571.050 ;
        RECT 102.750 563.700 104.550 564.000 ;
        RECT 113.550 563.700 114.450 578.400 ;
        RECT 131.400 571.050 132.300 581.400 ;
        RECT 152.100 571.050 153.300 581.400 ;
        RECT 155.550 578.400 157.350 584.400 ;
        RECT 158.850 578.400 160.650 585.000 ;
        RECT 163.950 581.400 165.750 584.400 ;
        RECT 168.450 581.400 170.250 585.000 ;
        RECT 171.450 581.400 173.250 584.400 ;
        RECT 174.750 581.400 176.550 585.000 ;
        RECT 179.250 582.300 181.050 584.400 ;
        RECT 179.250 581.400 182.850 582.300 ;
        RECT 163.350 579.300 165.750 581.400 ;
        RECT 172.200 580.500 173.250 581.400 ;
        RECT 179.250 580.800 183.150 581.400 ;
        RECT 172.200 579.450 177.150 580.500 ;
        RECT 175.350 578.700 177.150 579.450 ;
        RECT 155.550 571.050 156.750 578.400 ;
        RECT 178.350 577.800 180.150 579.600 ;
        RECT 181.050 579.300 183.150 580.800 ;
        RECT 184.050 578.400 185.850 585.000 ;
        RECT 187.050 580.200 188.850 584.400 ;
        RECT 203.100 581.400 204.900 585.000 ;
        RECT 206.100 581.400 207.900 584.400 ;
        RECT 221.100 581.400 222.900 585.000 ;
        RECT 224.100 581.400 225.900 584.400 ;
        RECT 227.100 581.400 228.900 585.000 ;
        RECT 187.050 578.400 189.450 580.200 ;
        RECT 168.150 576.000 169.950 576.600 ;
        RECT 179.100 576.000 180.150 577.800 ;
        RECT 168.150 574.800 180.150 576.000 ;
        RECT 127.950 568.950 130.050 571.050 ;
        RECT 130.950 568.950 133.050 571.050 ;
        RECT 133.950 568.950 136.050 571.050 ;
        RECT 148.950 568.950 151.050 571.050 ;
        RECT 151.950 568.950 154.050 571.050 ;
        RECT 155.550 569.250 161.850 571.050 ;
        RECT 155.550 568.950 160.050 569.250 ;
        RECT 128.250 567.150 130.050 568.950 ;
        RECT 102.750 563.100 114.450 563.700 ;
        RECT 34.350 559.200 40.050 560.100 ;
        RECT 40.950 560.700 42.750 561.300 ;
        RECT 40.950 559.500 48.750 560.700 ;
        RECT 34.350 558.600 36.150 559.200 ;
        RECT 46.650 558.600 48.750 559.500 ;
        RECT 31.350 555.600 33.450 557.700 ;
        RECT 37.950 557.550 39.750 558.300 ;
        RECT 42.750 557.550 44.550 558.300 ;
        RECT 37.950 556.500 44.550 557.550 ;
        RECT 31.350 549.600 33.150 555.600 ;
        RECT 35.850 549.000 37.650 555.600 ;
        RECT 38.850 549.600 40.650 556.500 ;
        RECT 41.850 549.000 43.650 555.600 ;
        RECT 46.650 549.600 48.450 558.600 ;
        RECT 52.050 549.000 53.850 561.600 ;
        RECT 55.050 559.800 57.450 561.600 ;
        RECT 55.050 549.600 56.850 559.800 ;
        RECT 71.100 549.000 72.900 561.600 ;
        RECT 74.400 560.400 78.000 561.600 ;
        RECT 76.200 549.600 78.000 560.400 ;
        RECT 80.550 549.600 82.350 561.600 ;
        RECT 83.550 549.000 85.350 561.600 ;
        RECT 89.250 561.300 94.050 562.200 ;
        RECT 96.150 562.500 114.450 563.100 ;
        RECT 96.150 562.200 104.550 562.500 ;
        RECT 89.250 560.400 90.450 561.300 ;
        RECT 87.450 558.600 90.450 560.400 ;
        RECT 91.350 560.100 93.150 560.400 ;
        RECT 96.150 560.100 97.050 562.200 ;
        RECT 113.550 561.600 114.450 562.500 ;
        RECT 131.400 561.600 132.300 568.950 ;
        RECT 134.100 567.150 135.900 568.950 ;
        RECT 149.100 567.150 150.900 568.950 ;
        RECT 91.350 559.200 97.050 560.100 ;
        RECT 97.950 560.700 99.750 561.300 ;
        RECT 97.950 559.500 105.750 560.700 ;
        RECT 91.350 558.600 93.150 559.200 ;
        RECT 103.650 558.600 105.750 559.500 ;
        RECT 88.350 555.600 90.450 557.700 ;
        RECT 94.950 557.550 96.750 558.300 ;
        RECT 99.750 557.550 101.550 558.300 ;
        RECT 94.950 556.500 101.550 557.550 ;
        RECT 88.350 549.600 90.150 555.600 ;
        RECT 92.850 549.000 94.650 555.600 ;
        RECT 95.850 549.600 97.650 556.500 ;
        RECT 98.850 549.000 100.650 555.600 ;
        RECT 103.650 549.600 105.450 558.600 ;
        RECT 109.050 549.000 110.850 561.600 ;
        RECT 112.050 559.800 114.450 561.600 ;
        RECT 112.050 549.600 113.850 559.800 ;
        RECT 128.100 549.000 129.900 561.600 ;
        RECT 131.400 560.400 135.000 561.600 ;
        RECT 133.200 549.600 135.000 560.400 ;
        RECT 152.100 555.600 153.300 568.950 ;
        RECT 155.550 561.600 156.750 568.950 ;
        RECT 157.650 566.100 159.450 566.250 ;
        RECT 163.350 566.100 165.450 566.400 ;
        RECT 157.650 564.900 165.450 566.100 ;
        RECT 157.650 564.450 159.450 564.900 ;
        RECT 163.350 564.300 165.450 564.900 ;
        RECT 168.150 562.200 169.050 574.800 ;
        RECT 179.100 573.600 187.050 574.800 ;
        RECT 179.100 573.000 180.900 573.600 ;
        RECT 182.100 571.800 183.900 572.400 ;
        RECT 175.800 570.600 183.900 571.800 ;
        RECT 185.250 571.050 187.050 573.600 ;
        RECT 175.800 568.950 177.900 570.600 ;
        RECT 184.950 568.950 187.050 571.050 ;
        RECT 177.750 563.700 179.550 564.000 ;
        RECT 188.550 563.700 189.450 578.400 ;
        RECT 206.100 571.050 207.300 581.400 ;
        RECT 214.950 576.450 217.050 577.050 ;
        RECT 220.950 576.450 223.050 577.050 ;
        RECT 214.950 575.550 223.050 576.450 ;
        RECT 214.950 574.950 217.050 575.550 ;
        RECT 220.950 574.950 223.050 575.550 ;
        RECT 224.400 571.050 225.300 581.400 ;
        RECT 242.700 577.200 244.500 584.400 ;
        RECT 247.800 578.400 249.600 585.000 ;
        RECT 266.100 579.300 267.900 584.400 ;
        RECT 269.100 580.200 270.900 585.000 ;
        RECT 272.100 579.300 273.900 584.400 ;
        RECT 266.100 577.950 273.900 579.300 ;
        RECT 275.100 578.400 276.900 584.400 ;
        RECT 242.700 576.300 246.900 577.200 ;
        RECT 275.100 576.300 276.300 578.400 ;
        RECT 242.100 571.050 243.900 572.850 ;
        RECT 245.700 571.050 246.900 576.300 ;
        RECT 272.700 575.400 276.300 576.300 ;
        RECT 290.100 576.600 291.900 584.400 ;
        RECT 294.600 578.400 296.400 585.000 ;
        RECT 297.600 580.200 299.400 584.400 ;
        RECT 297.600 578.400 300.300 580.200 ;
        RECT 314.400 578.400 316.200 585.000 ;
        RECT 296.700 576.600 298.500 577.500 ;
        RECT 290.100 575.700 298.500 576.600 ;
        RECT 247.950 571.050 249.750 572.850 ;
        RECT 269.100 571.050 270.900 572.850 ;
        RECT 272.700 571.050 273.900 575.400 ;
        RECT 275.100 571.050 276.900 572.850 ;
        RECT 290.250 571.050 292.050 572.850 ;
        RECT 202.950 568.950 205.050 571.050 ;
        RECT 205.950 568.950 208.050 571.050 ;
        RECT 220.950 568.950 223.050 571.050 ;
        RECT 223.950 568.950 226.050 571.050 ;
        RECT 226.950 568.950 229.050 571.050 ;
        RECT 241.950 568.950 244.050 571.050 ;
        RECT 244.950 568.950 247.050 571.050 ;
        RECT 247.950 568.950 250.050 571.050 ;
        RECT 265.950 568.950 268.050 571.050 ;
        RECT 268.950 568.950 271.050 571.050 ;
        RECT 271.950 568.950 274.050 571.050 ;
        RECT 274.950 568.950 277.050 571.050 ;
        RECT 290.100 568.950 292.200 571.050 ;
        RECT 203.100 567.150 204.900 568.950 ;
        RECT 177.750 563.100 189.450 563.700 ;
        RECT 149.100 549.000 150.900 555.600 ;
        RECT 152.100 549.600 153.900 555.600 ;
        RECT 155.550 549.600 157.350 561.600 ;
        RECT 158.550 549.000 160.350 561.600 ;
        RECT 164.250 561.300 169.050 562.200 ;
        RECT 171.150 562.500 189.450 563.100 ;
        RECT 171.150 562.200 179.550 562.500 ;
        RECT 164.250 560.400 165.450 561.300 ;
        RECT 162.450 558.600 165.450 560.400 ;
        RECT 166.350 560.100 168.150 560.400 ;
        RECT 171.150 560.100 172.050 562.200 ;
        RECT 188.550 561.600 189.450 562.500 ;
        RECT 166.350 559.200 172.050 560.100 ;
        RECT 172.950 560.700 174.750 561.300 ;
        RECT 172.950 559.500 180.750 560.700 ;
        RECT 166.350 558.600 168.150 559.200 ;
        RECT 178.650 558.600 180.750 559.500 ;
        RECT 163.350 555.600 165.450 557.700 ;
        RECT 169.950 557.550 171.750 558.300 ;
        RECT 174.750 557.550 176.550 558.300 ;
        RECT 169.950 556.500 176.550 557.550 ;
        RECT 163.350 549.600 165.150 555.600 ;
        RECT 167.850 549.000 169.650 555.600 ;
        RECT 170.850 549.600 172.650 556.500 ;
        RECT 173.850 549.000 175.650 555.600 ;
        RECT 178.650 549.600 180.450 558.600 ;
        RECT 184.050 549.000 185.850 561.600 ;
        RECT 187.050 559.800 189.450 561.600 ;
        RECT 187.050 549.600 188.850 559.800 ;
        RECT 206.100 555.600 207.300 568.950 ;
        RECT 221.250 567.150 223.050 568.950 ;
        RECT 224.400 561.600 225.300 568.950 ;
        RECT 227.100 567.150 228.900 568.950 ;
        RECT 203.100 549.000 204.900 555.600 ;
        RECT 206.100 549.600 207.900 555.600 ;
        RECT 221.100 549.000 222.900 561.600 ;
        RECT 224.400 560.400 228.000 561.600 ;
        RECT 226.200 549.600 228.000 560.400 ;
        RECT 245.700 555.600 246.900 568.950 ;
        RECT 266.100 567.150 267.900 568.950 ;
        RECT 272.700 561.600 273.900 568.950 ;
        RECT 242.100 549.000 243.900 555.600 ;
        RECT 245.100 549.600 246.900 555.600 ;
        RECT 248.100 549.000 249.900 555.600 ;
        RECT 266.400 549.000 268.200 561.600 ;
        RECT 271.500 560.100 273.900 561.600 ;
        RECT 271.500 549.600 273.300 560.100 ;
        RECT 274.200 557.100 276.000 558.900 ;
        RECT 293.100 555.600 294.000 575.700 ;
        RECT 299.400 571.050 300.300 578.400 ;
        RECT 319.500 577.200 321.300 584.400 ;
        RECT 317.100 576.300 321.300 577.200 ;
        RECT 314.250 571.050 316.050 572.850 ;
        RECT 317.100 571.050 318.300 576.300 ;
        RECT 335.100 575.400 336.900 585.000 ;
        RECT 341.700 576.000 343.500 584.400 ;
        RECT 362.400 578.400 364.200 585.000 ;
        RECT 367.500 577.200 369.300 584.400 ;
        RECT 383.100 578.400 384.900 584.400 ;
        RECT 365.100 576.300 369.300 577.200 ;
        RECT 383.700 576.300 384.900 578.400 ;
        RECT 386.100 579.300 387.900 584.400 ;
        RECT 389.100 580.200 390.900 585.000 ;
        RECT 392.100 579.300 393.900 584.400 ;
        RECT 407.100 581.400 408.900 585.000 ;
        RECT 410.100 581.400 411.900 584.400 ;
        RECT 386.100 577.950 393.900 579.300 ;
        RECT 341.700 574.800 345.000 576.000 ;
        RECT 320.100 571.050 321.900 572.850 ;
        RECT 335.100 571.050 336.900 572.850 ;
        RECT 341.100 571.050 342.900 572.850 ;
        RECT 344.100 571.050 345.000 574.800 ;
        RECT 362.250 571.050 364.050 572.850 ;
        RECT 365.100 571.050 366.300 576.300 ;
        RECT 383.700 575.400 387.300 576.300 ;
        RECT 368.100 571.050 369.900 572.850 ;
        RECT 383.100 571.050 384.900 572.850 ;
        RECT 386.100 571.050 387.300 575.400 ;
        RECT 389.100 571.050 390.900 572.850 ;
        RECT 410.100 571.050 411.300 581.400 ;
        RECT 425.100 576.600 426.900 584.400 ;
        RECT 429.600 578.400 431.400 585.000 ;
        RECT 432.600 580.200 434.400 584.400 ;
        RECT 432.600 578.400 435.300 580.200 ;
        RECT 452.400 578.400 454.200 585.000 ;
        RECT 431.700 576.600 433.500 577.500 ;
        RECT 425.100 575.700 433.500 576.600 ;
        RECT 425.250 571.050 427.050 572.850 ;
        RECT 295.500 568.950 297.600 571.050 ;
        RECT 298.800 568.950 300.900 571.050 ;
        RECT 313.950 568.950 316.050 571.050 ;
        RECT 316.950 568.950 319.050 571.050 ;
        RECT 319.950 568.950 322.050 571.050 ;
        RECT 334.950 568.950 337.050 571.050 ;
        RECT 337.950 568.950 340.050 571.050 ;
        RECT 340.950 568.950 343.050 571.050 ;
        RECT 343.950 568.950 346.050 571.050 ;
        RECT 361.950 568.950 364.050 571.050 ;
        RECT 364.950 568.950 367.050 571.050 ;
        RECT 367.950 568.950 370.050 571.050 ;
        RECT 382.950 568.950 385.050 571.050 ;
        RECT 385.950 568.950 388.050 571.050 ;
        RECT 388.950 568.950 391.050 571.050 ;
        RECT 391.950 568.950 394.050 571.050 ;
        RECT 406.950 568.950 409.050 571.050 ;
        RECT 409.950 568.950 412.050 571.050 ;
        RECT 425.100 568.950 427.200 571.050 ;
        RECT 295.200 567.150 297.000 568.950 ;
        RECT 299.400 561.600 300.300 568.950 ;
        RECT 274.500 549.000 276.300 555.600 ;
        RECT 290.100 549.000 291.900 555.600 ;
        RECT 293.100 549.600 294.900 555.600 ;
        RECT 296.100 549.000 297.900 561.000 ;
        RECT 299.100 549.600 300.900 561.600 ;
        RECT 317.100 555.600 318.300 568.950 ;
        RECT 338.100 567.150 339.900 568.950 ;
        RECT 344.100 556.800 345.000 568.950 ;
        RECT 338.400 555.900 345.000 556.800 ;
        RECT 338.400 555.600 339.900 555.900 ;
        RECT 314.100 549.000 315.900 555.600 ;
        RECT 317.100 549.600 318.900 555.600 ;
        RECT 320.100 549.000 321.900 555.600 ;
        RECT 335.100 549.000 336.900 555.600 ;
        RECT 338.100 549.600 339.900 555.600 ;
        RECT 344.100 555.600 345.000 555.900 ;
        RECT 365.100 555.600 366.300 568.950 ;
        RECT 386.100 561.600 387.300 568.950 ;
        RECT 392.100 567.150 393.900 568.950 ;
        RECT 407.100 567.150 408.900 568.950 ;
        RECT 386.100 560.100 388.500 561.600 ;
        RECT 384.000 557.100 385.800 558.900 ;
        RECT 341.100 549.000 342.900 555.000 ;
        RECT 344.100 549.600 345.900 555.600 ;
        RECT 362.100 549.000 363.900 555.600 ;
        RECT 365.100 549.600 366.900 555.600 ;
        RECT 368.100 549.000 369.900 555.600 ;
        RECT 383.700 549.000 385.500 555.600 ;
        RECT 386.700 549.600 388.500 560.100 ;
        RECT 391.800 549.000 393.600 561.600 ;
        RECT 410.100 555.600 411.300 568.950 ;
        RECT 428.100 555.600 429.000 575.700 ;
        RECT 434.400 571.050 435.300 578.400 ;
        RECT 457.500 577.200 459.300 584.400 ;
        RECT 473.100 578.400 474.900 584.400 ;
        RECT 476.100 578.400 477.900 585.000 ;
        RECT 455.100 576.300 459.300 577.200 ;
        RECT 452.250 571.050 454.050 572.850 ;
        RECT 455.100 571.050 456.300 576.300 ;
        RECT 458.100 571.050 459.900 572.850 ;
        RECT 473.700 571.050 474.900 578.400 ;
        RECT 491.100 576.600 492.900 584.400 ;
        RECT 495.600 578.400 497.400 585.000 ;
        RECT 498.600 580.200 500.400 584.400 ;
        RECT 515.100 581.400 516.900 585.000 ;
        RECT 518.100 581.400 519.900 584.400 ;
        RECT 498.600 578.400 501.300 580.200 ;
        RECT 497.700 576.600 499.500 577.500 ;
        RECT 491.100 575.700 499.500 576.600 ;
        RECT 476.100 571.050 477.900 572.850 ;
        RECT 491.250 571.050 493.050 572.850 ;
        RECT 430.500 568.950 432.600 571.050 ;
        RECT 433.800 568.950 435.900 571.050 ;
        RECT 451.950 568.950 454.050 571.050 ;
        RECT 454.950 568.950 457.050 571.050 ;
        RECT 457.950 568.950 460.050 571.050 ;
        RECT 472.950 568.950 475.050 571.050 ;
        RECT 475.950 568.950 478.050 571.050 ;
        RECT 491.100 568.950 493.200 571.050 ;
        RECT 430.200 567.150 432.000 568.950 ;
        RECT 434.400 561.600 435.300 568.950 ;
        RECT 407.100 549.000 408.900 555.600 ;
        RECT 410.100 549.600 411.900 555.600 ;
        RECT 425.100 549.000 426.900 555.600 ;
        RECT 428.100 549.600 429.900 555.600 ;
        RECT 431.100 549.000 432.900 561.000 ;
        RECT 434.100 549.600 435.900 561.600 ;
        RECT 455.100 555.600 456.300 568.950 ;
        RECT 473.700 561.600 474.900 568.950 ;
        RECT 452.100 549.000 453.900 555.600 ;
        RECT 455.100 549.600 456.900 555.600 ;
        RECT 458.100 549.000 459.900 555.600 ;
        RECT 473.100 549.600 474.900 561.600 ;
        RECT 476.100 549.000 477.900 561.600 ;
        RECT 494.100 555.600 495.000 575.700 ;
        RECT 500.400 571.050 501.300 578.400 ;
        RECT 518.100 571.050 519.300 581.400 ;
        RECT 533.100 579.300 534.900 584.400 ;
        RECT 536.100 580.200 537.900 585.000 ;
        RECT 539.100 579.300 540.900 584.400 ;
        RECT 533.100 577.950 540.900 579.300 ;
        RECT 542.100 578.400 543.900 584.400 ;
        RECT 557.100 579.300 558.900 584.400 ;
        RECT 560.100 580.200 561.900 585.000 ;
        RECT 563.100 579.300 564.900 584.400 ;
        RECT 542.100 576.300 543.300 578.400 ;
        RECT 557.100 577.950 564.900 579.300 ;
        RECT 566.100 578.400 567.900 584.400 ;
        RECT 566.100 576.300 567.300 578.400 ;
        RECT 539.700 575.400 543.300 576.300 ;
        RECT 563.700 575.400 567.300 576.300 ;
        RECT 581.100 575.400 582.900 585.000 ;
        RECT 587.700 576.000 589.500 584.400 ;
        RECT 605.100 579.300 606.900 584.400 ;
        RECT 608.100 580.200 609.900 585.000 ;
        RECT 611.100 579.300 612.900 584.400 ;
        RECT 605.100 577.950 612.900 579.300 ;
        RECT 614.100 578.400 615.900 584.400 ;
        RECT 614.100 576.300 615.300 578.400 ;
        RECT 629.700 577.200 631.500 584.400 ;
        RECT 634.800 578.400 636.600 585.000 ;
        RECT 652.500 578.400 654.300 585.000 ;
        RECT 657.000 578.400 658.800 584.400 ;
        RECT 661.500 578.400 663.300 585.000 ;
        RECT 680.400 578.400 682.200 585.000 ;
        RECT 629.700 576.300 633.900 577.200 ;
        RECT 536.100 571.050 537.900 572.850 ;
        RECT 539.700 571.050 540.900 575.400 ;
        RECT 542.100 571.050 543.900 572.850 ;
        RECT 560.100 571.050 561.900 572.850 ;
        RECT 563.700 571.050 564.900 575.400 ;
        RECT 587.700 574.800 591.000 576.000 ;
        RECT 568.950 573.450 571.050 574.050 ;
        RECT 574.950 573.450 577.050 573.900 ;
        RECT 566.100 571.050 567.900 572.850 ;
        RECT 568.950 572.550 577.050 573.450 ;
        RECT 568.950 571.950 571.050 572.550 ;
        RECT 574.950 571.800 577.050 572.550 ;
        RECT 581.100 571.050 582.900 572.850 ;
        RECT 587.100 571.050 588.900 572.850 ;
        RECT 590.100 571.050 591.000 574.800 ;
        RECT 611.700 575.400 615.300 576.300 ;
        RECT 608.100 571.050 609.900 572.850 ;
        RECT 611.700 571.050 612.900 575.400 ;
        RECT 614.100 571.050 615.900 572.850 ;
        RECT 629.100 571.050 630.900 572.850 ;
        RECT 632.700 571.050 633.900 576.300 ;
        RECT 634.950 571.050 636.750 572.850 ;
        RECT 650.100 571.050 651.900 572.850 ;
        RECT 656.700 571.050 657.900 578.400 ;
        RECT 685.500 577.200 687.300 584.400 ;
        RECT 705.000 578.400 706.800 585.000 ;
        RECT 709.500 579.600 711.300 584.400 ;
        RECT 712.500 581.400 714.300 585.000 ;
        RECT 728.100 581.400 729.900 584.400 ;
        RECT 731.100 581.400 732.900 585.000 ;
        RECT 709.500 578.400 714.600 579.600 ;
        RECT 683.100 576.300 687.300 577.200 ;
        RECT 661.950 571.050 663.750 572.850 ;
        RECT 680.250 571.050 682.050 572.850 ;
        RECT 683.100 571.050 684.300 576.300 ;
        RECT 686.100 571.050 687.900 572.850 ;
        RECT 704.100 571.050 705.900 572.850 ;
        RECT 710.250 571.050 712.050 572.850 ;
        RECT 713.700 571.050 714.600 578.400 ;
        RECT 728.700 571.050 729.900 581.400 ;
        RECT 746.100 579.300 747.900 584.400 ;
        RECT 749.100 580.200 750.900 585.000 ;
        RECT 752.100 579.300 753.900 584.400 ;
        RECT 746.100 577.950 753.900 579.300 ;
        RECT 755.100 578.400 756.900 584.400 ;
        RECT 770.700 581.400 772.500 585.000 ;
        RECT 773.700 579.600 775.500 584.400 ;
        RECT 770.400 578.400 775.500 579.600 ;
        RECT 778.200 578.400 780.000 585.000 ;
        RECT 755.100 576.300 756.300 578.400 ;
        RECT 752.700 575.400 756.300 576.300 ;
        RECT 749.100 571.050 750.900 572.850 ;
        RECT 752.700 571.050 753.900 575.400 ;
        RECT 755.100 571.050 756.900 572.850 ;
        RECT 770.400 571.050 771.300 578.400 ;
        RECT 772.950 576.450 775.050 577.050 ;
        RECT 790.950 576.450 793.050 577.050 ;
        RECT 772.950 575.550 793.050 576.450 ;
        RECT 796.500 576.000 798.300 584.400 ;
        RECT 772.950 574.950 775.050 575.550 ;
        RECT 790.950 574.950 793.050 575.550 ;
        RECT 795.000 574.800 798.300 576.000 ;
        RECT 803.100 575.400 804.900 585.000 ;
        RECT 818.100 575.400 819.900 585.000 ;
        RECT 824.700 576.000 826.500 584.400 ;
        RECT 847.500 576.000 849.300 584.400 ;
        RECT 824.700 574.800 828.000 576.000 ;
        RECT 772.950 571.050 774.750 572.850 ;
        RECT 779.100 571.050 780.900 572.850 ;
        RECT 795.000 571.050 795.900 574.800 ;
        RECT 797.100 571.050 798.900 572.850 ;
        RECT 803.100 571.050 804.900 572.850 ;
        RECT 818.100 571.050 819.900 572.850 ;
        RECT 824.100 571.050 825.900 572.850 ;
        RECT 827.100 571.050 828.000 574.800 ;
        RECT 846.000 574.800 849.300 576.000 ;
        RECT 854.100 575.400 855.900 585.000 ;
        RECT 869.100 578.400 870.900 584.400 ;
        RECT 869.700 576.300 870.900 578.400 ;
        RECT 872.100 579.300 873.900 584.400 ;
        RECT 875.100 580.200 876.900 585.000 ;
        RECT 878.100 579.300 879.900 584.400 ;
        RECT 872.100 577.950 879.900 579.300 ;
        RECT 869.700 575.400 873.300 576.300 ;
        RECT 840.000 573.450 844.050 574.050 ;
        RECT 839.550 571.950 844.050 573.450 ;
        RECT 496.500 568.950 498.600 571.050 ;
        RECT 499.800 568.950 501.900 571.050 ;
        RECT 514.950 568.950 517.050 571.050 ;
        RECT 517.950 568.950 520.050 571.050 ;
        RECT 532.950 568.950 535.050 571.050 ;
        RECT 535.950 568.950 538.050 571.050 ;
        RECT 538.950 568.950 541.050 571.050 ;
        RECT 541.950 568.950 544.050 571.050 ;
        RECT 556.950 568.950 559.050 571.050 ;
        RECT 559.950 568.950 562.050 571.050 ;
        RECT 562.950 568.950 565.050 571.050 ;
        RECT 565.950 568.950 568.050 571.050 ;
        RECT 580.950 568.950 583.050 571.050 ;
        RECT 583.950 568.950 586.050 571.050 ;
        RECT 586.950 568.950 589.050 571.050 ;
        RECT 589.950 568.950 592.050 571.050 ;
        RECT 604.950 568.950 607.050 571.050 ;
        RECT 607.950 568.950 610.050 571.050 ;
        RECT 610.950 568.950 613.050 571.050 ;
        RECT 613.950 568.950 616.050 571.050 ;
        RECT 628.950 568.950 631.050 571.050 ;
        RECT 631.950 568.950 634.050 571.050 ;
        RECT 634.950 568.950 637.050 571.050 ;
        RECT 649.950 568.950 652.050 571.050 ;
        RECT 652.950 568.950 655.050 571.050 ;
        RECT 655.950 568.950 658.050 571.050 ;
        RECT 658.950 568.950 661.050 571.050 ;
        RECT 661.950 568.950 664.050 571.050 ;
        RECT 679.950 568.950 682.050 571.050 ;
        RECT 682.950 568.950 685.050 571.050 ;
        RECT 685.950 568.950 688.050 571.050 ;
        RECT 703.950 568.950 706.050 571.050 ;
        RECT 706.950 568.950 709.050 571.050 ;
        RECT 709.950 568.950 712.050 571.050 ;
        RECT 712.950 568.950 715.050 571.050 ;
        RECT 727.950 568.950 730.050 571.050 ;
        RECT 730.950 568.950 733.050 571.050 ;
        RECT 745.950 568.950 748.050 571.050 ;
        RECT 748.950 568.950 751.050 571.050 ;
        RECT 751.950 568.950 754.050 571.050 ;
        RECT 754.950 568.950 757.050 571.050 ;
        RECT 769.950 568.950 772.050 571.050 ;
        RECT 772.950 568.950 775.050 571.050 ;
        RECT 775.950 568.950 778.050 571.050 ;
        RECT 778.950 568.950 781.050 571.050 ;
        RECT 793.950 568.950 796.050 571.050 ;
        RECT 796.950 568.950 799.050 571.050 ;
        RECT 799.950 568.950 802.050 571.050 ;
        RECT 802.950 568.950 805.050 571.050 ;
        RECT 817.950 568.950 820.050 571.050 ;
        RECT 820.950 568.950 823.050 571.050 ;
        RECT 823.950 568.950 826.050 571.050 ;
        RECT 826.950 568.950 829.050 571.050 ;
        RECT 496.200 567.150 498.000 568.950 ;
        RECT 500.400 561.600 501.300 568.950 ;
        RECT 515.100 567.150 516.900 568.950 ;
        RECT 491.100 549.000 492.900 555.600 ;
        RECT 494.100 549.600 495.900 555.600 ;
        RECT 497.100 549.000 498.900 561.000 ;
        RECT 500.100 549.600 501.900 561.600 ;
        RECT 518.100 555.600 519.300 568.950 ;
        RECT 533.100 567.150 534.900 568.950 ;
        RECT 539.700 561.600 540.900 568.950 ;
        RECT 557.100 567.150 558.900 568.950 ;
        RECT 563.700 561.600 564.900 568.950 ;
        RECT 584.100 567.150 585.900 568.950 ;
        RECT 574.950 564.450 577.050 565.050 ;
        RECT 586.950 564.450 589.050 565.050 ;
        RECT 574.950 563.550 589.050 564.450 ;
        RECT 574.950 562.950 577.050 563.550 ;
        RECT 586.950 562.950 589.050 563.550 ;
        RECT 515.100 549.000 516.900 555.600 ;
        RECT 518.100 549.600 519.900 555.600 ;
        RECT 533.400 549.000 535.200 561.600 ;
        RECT 538.500 560.100 540.900 561.600 ;
        RECT 538.500 549.600 540.300 560.100 ;
        RECT 541.200 557.100 543.000 558.900 ;
        RECT 541.500 549.000 543.300 555.600 ;
        RECT 557.400 549.000 559.200 561.600 ;
        RECT 562.500 560.100 564.900 561.600 ;
        RECT 562.500 549.600 564.300 560.100 ;
        RECT 565.200 557.100 567.000 558.900 ;
        RECT 590.100 556.800 591.000 568.950 ;
        RECT 605.100 567.150 606.900 568.950 ;
        RECT 595.950 564.450 598.050 565.050 ;
        RECT 607.950 564.450 610.050 565.050 ;
        RECT 595.950 563.550 610.050 564.450 ;
        RECT 595.950 562.950 598.050 563.550 ;
        RECT 607.950 562.950 610.050 563.550 ;
        RECT 611.700 561.600 612.900 568.950 ;
        RECT 584.400 555.900 591.000 556.800 ;
        RECT 584.400 555.600 585.900 555.900 ;
        RECT 565.500 549.000 567.300 555.600 ;
        RECT 581.100 549.000 582.900 555.600 ;
        RECT 584.100 549.600 585.900 555.600 ;
        RECT 590.100 555.600 591.000 555.900 ;
        RECT 587.100 549.000 588.900 555.000 ;
        RECT 590.100 549.600 591.900 555.600 ;
        RECT 605.400 549.000 607.200 561.600 ;
        RECT 610.500 560.100 612.900 561.600 ;
        RECT 610.500 549.600 612.300 560.100 ;
        RECT 613.200 557.100 615.000 558.900 ;
        RECT 632.700 555.600 633.900 568.950 ;
        RECT 653.100 567.150 654.900 568.950 ;
        RECT 657.000 563.400 657.900 568.950 ;
        RECT 658.950 567.150 660.750 568.950 ;
        RECT 653.100 562.500 657.900 563.400 ;
        RECT 613.500 549.000 615.300 555.600 ;
        RECT 629.100 549.000 630.900 555.600 ;
        RECT 632.100 549.600 633.900 555.600 ;
        RECT 635.100 549.000 636.900 555.600 ;
        RECT 650.100 550.500 651.900 561.600 ;
        RECT 653.100 551.400 654.900 562.500 ;
        RECT 656.100 560.400 663.900 561.300 ;
        RECT 656.100 550.500 657.900 560.400 ;
        RECT 650.100 549.600 657.900 550.500 ;
        RECT 659.100 549.000 660.900 559.500 ;
        RECT 662.100 549.600 663.900 560.400 ;
        RECT 683.100 555.600 684.300 568.950 ;
        RECT 707.250 567.150 709.050 568.950 ;
        RECT 713.700 561.600 714.600 568.950 ;
        RECT 704.100 560.700 711.900 561.600 ;
        RECT 680.100 549.000 681.900 555.600 ;
        RECT 683.100 549.600 684.900 555.600 ;
        RECT 686.100 549.000 687.900 555.600 ;
        RECT 704.100 549.600 705.900 560.700 ;
        RECT 707.100 549.000 708.900 559.800 ;
        RECT 710.100 549.600 711.900 560.700 ;
        RECT 713.100 549.600 714.900 561.600 ;
        RECT 728.700 555.600 729.900 568.950 ;
        RECT 731.100 567.150 732.900 568.950 ;
        RECT 746.100 567.150 747.900 568.950 ;
        RECT 752.700 561.600 753.900 568.950 ;
        RECT 770.400 561.600 771.300 568.950 ;
        RECT 775.950 567.150 777.750 568.950 ;
        RECT 728.100 549.600 729.900 555.600 ;
        RECT 731.100 549.000 732.900 555.600 ;
        RECT 746.400 549.000 748.200 561.600 ;
        RECT 751.500 560.100 753.900 561.600 ;
        RECT 751.500 549.600 753.300 560.100 ;
        RECT 754.200 557.100 756.000 558.900 ;
        RECT 754.500 549.000 756.300 555.600 ;
        RECT 770.100 549.600 771.900 561.600 ;
        RECT 773.100 560.700 780.900 561.600 ;
        RECT 773.100 549.600 774.900 560.700 ;
        RECT 776.100 549.000 777.900 559.800 ;
        RECT 779.100 549.600 780.900 560.700 ;
        RECT 795.000 556.800 795.900 568.950 ;
        RECT 800.100 567.150 801.900 568.950 ;
        RECT 821.100 567.150 822.900 568.950 ;
        RECT 811.950 564.450 814.050 565.050 ;
        RECT 823.950 564.450 826.050 564.750 ;
        RECT 811.950 563.550 826.050 564.450 ;
        RECT 811.950 562.950 814.050 563.550 ;
        RECT 823.950 562.650 826.050 563.550 ;
        RECT 827.100 556.800 828.000 568.950 ;
        RECT 839.550 568.050 840.450 571.950 ;
        RECT 846.000 571.050 846.900 574.800 ;
        RECT 859.950 573.450 862.050 574.050 ;
        RECT 865.950 573.450 868.050 574.050 ;
        RECT 848.100 571.050 849.900 572.850 ;
        RECT 854.100 571.050 855.900 572.850 ;
        RECT 859.950 572.550 868.050 573.450 ;
        RECT 859.950 571.950 862.050 572.550 ;
        RECT 865.950 571.950 868.050 572.550 ;
        RECT 869.100 571.050 870.900 572.850 ;
        RECT 872.100 571.050 873.300 575.400 ;
        RECT 875.100 571.050 876.900 572.850 ;
        RECT 844.950 568.950 847.050 571.050 ;
        RECT 847.950 568.950 850.050 571.050 ;
        RECT 850.950 568.950 853.050 571.050 ;
        RECT 853.950 568.950 856.050 571.050 ;
        RECT 868.950 568.950 871.050 571.050 ;
        RECT 871.950 568.950 874.050 571.050 ;
        RECT 874.950 568.950 877.050 571.050 ;
        RECT 877.950 568.950 880.050 571.050 ;
        RECT 839.550 566.550 844.050 568.050 ;
        RECT 840.000 565.950 844.050 566.550 ;
        RECT 795.000 555.900 801.600 556.800 ;
        RECT 795.000 555.600 795.900 555.900 ;
        RECT 794.100 549.600 795.900 555.600 ;
        RECT 800.100 555.600 801.600 555.900 ;
        RECT 821.400 555.900 828.000 556.800 ;
        RECT 821.400 555.600 822.900 555.900 ;
        RECT 797.100 549.000 798.900 555.000 ;
        RECT 800.100 549.600 801.900 555.600 ;
        RECT 803.100 549.000 804.900 555.600 ;
        RECT 818.100 549.000 819.900 555.600 ;
        RECT 821.100 549.600 822.900 555.600 ;
        RECT 827.100 555.600 828.000 555.900 ;
        RECT 846.000 556.800 846.900 568.950 ;
        RECT 851.100 567.150 852.900 568.950 ;
        RECT 872.100 561.600 873.300 568.950 ;
        RECT 878.100 567.150 879.900 568.950 ;
        RECT 872.100 560.100 874.500 561.600 ;
        RECT 870.000 557.100 871.800 558.900 ;
        RECT 846.000 555.900 852.600 556.800 ;
        RECT 846.000 555.600 846.900 555.900 ;
        RECT 824.100 549.000 825.900 555.000 ;
        RECT 827.100 549.600 828.900 555.600 ;
        RECT 845.100 549.600 846.900 555.600 ;
        RECT 851.100 555.600 852.600 555.900 ;
        RECT 848.100 549.000 849.900 555.000 ;
        RECT 851.100 549.600 852.900 555.600 ;
        RECT 854.100 549.000 855.900 555.600 ;
        RECT 869.700 549.000 871.500 555.600 ;
        RECT 872.700 549.600 874.500 560.100 ;
        RECT 877.800 549.000 879.600 561.600 ;
        RECT 14.100 533.400 15.900 545.400 ;
        RECT 17.100 535.200 18.900 546.000 ;
        RECT 20.100 539.400 21.900 545.400 ;
        RECT 14.100 526.050 15.300 533.400 ;
        RECT 20.700 532.500 21.900 539.400 ;
        RECT 16.200 531.600 21.900 532.500 ;
        RECT 23.550 533.400 25.350 545.400 ;
        RECT 26.550 533.400 28.350 546.000 ;
        RECT 31.350 539.400 33.150 545.400 ;
        RECT 35.850 539.400 37.650 546.000 ;
        RECT 31.350 537.300 33.450 539.400 ;
        RECT 38.850 538.500 40.650 545.400 ;
        RECT 41.850 539.400 43.650 546.000 ;
        RECT 37.950 537.450 44.550 538.500 ;
        RECT 37.950 536.700 39.750 537.450 ;
        RECT 42.750 536.700 44.550 537.450 ;
        RECT 46.650 536.400 48.450 545.400 ;
        RECT 30.450 534.600 33.450 536.400 ;
        RECT 34.350 535.800 36.150 536.400 ;
        RECT 34.350 534.900 40.050 535.800 ;
        RECT 46.650 535.500 48.750 536.400 ;
        RECT 34.350 534.600 36.150 534.900 ;
        RECT 32.250 533.700 33.450 534.600 ;
        RECT 16.200 530.700 18.000 531.600 ;
        RECT 14.100 523.950 16.200 526.050 ;
        RECT 14.100 516.600 15.300 523.950 ;
        RECT 17.100 519.300 18.000 530.700 ;
        RECT 19.800 526.050 21.600 527.850 ;
        RECT 19.500 523.950 21.600 526.050 ;
        RECT 23.550 526.050 24.750 533.400 ;
        RECT 32.250 532.800 37.050 533.700 ;
        RECT 25.650 530.100 27.450 530.550 ;
        RECT 31.350 530.100 33.450 530.700 ;
        RECT 25.650 528.900 33.450 530.100 ;
        RECT 25.650 528.750 27.450 528.900 ;
        RECT 31.350 528.600 33.450 528.900 ;
        RECT 23.550 525.750 28.050 526.050 ;
        RECT 23.550 523.950 29.850 525.750 ;
        RECT 16.200 518.400 18.000 519.300 ;
        RECT 16.200 517.500 21.900 518.400 ;
        RECT 14.100 510.600 15.900 516.600 ;
        RECT 17.100 510.000 18.900 516.600 ;
        RECT 20.700 513.600 21.900 517.500 ;
        RECT 20.100 510.600 21.900 513.600 ;
        RECT 23.550 516.600 24.750 523.950 ;
        RECT 36.150 520.200 37.050 532.800 ;
        RECT 39.150 532.800 40.050 534.900 ;
        RECT 40.950 534.300 48.750 535.500 ;
        RECT 40.950 533.700 42.750 534.300 ;
        RECT 52.050 533.400 53.850 546.000 ;
        RECT 55.050 535.200 56.850 545.400 ;
        RECT 55.050 533.400 57.450 535.200 ;
        RECT 39.150 532.500 47.550 532.800 ;
        RECT 56.550 532.500 57.450 533.400 ;
        RECT 39.150 531.900 57.450 532.500 ;
        RECT 45.750 531.300 57.450 531.900 ;
        RECT 45.750 531.000 47.550 531.300 ;
        RECT 43.800 524.400 45.900 526.050 ;
        RECT 43.800 523.200 51.900 524.400 ;
        RECT 52.950 523.950 55.050 526.050 ;
        RECT 50.100 522.600 51.900 523.200 ;
        RECT 47.100 521.400 48.900 522.000 ;
        RECT 53.250 521.400 55.050 523.950 ;
        RECT 47.100 520.200 55.050 521.400 ;
        RECT 36.150 519.000 48.150 520.200 ;
        RECT 36.150 518.400 37.950 519.000 ;
        RECT 47.100 517.200 48.150 519.000 ;
        RECT 23.550 510.600 25.350 516.600 ;
        RECT 26.850 510.000 28.650 516.600 ;
        RECT 31.350 513.600 33.750 515.700 ;
        RECT 43.350 515.550 45.150 516.300 ;
        RECT 40.200 514.500 45.150 515.550 ;
        RECT 46.350 515.400 48.150 517.200 ;
        RECT 56.550 516.600 57.450 531.300 ;
        RECT 40.200 513.600 41.250 514.500 ;
        RECT 49.050 514.200 51.150 515.700 ;
        RECT 47.250 513.600 51.150 514.200 ;
        RECT 31.950 510.600 33.750 513.600 ;
        RECT 36.450 510.000 38.250 513.600 ;
        RECT 39.450 510.600 41.250 513.600 ;
        RECT 42.750 510.000 44.550 513.600 ;
        RECT 47.250 512.700 50.850 513.600 ;
        RECT 47.250 510.600 49.050 512.700 ;
        RECT 52.050 510.000 53.850 516.600 ;
        RECT 55.050 514.800 57.450 516.600 ;
        RECT 59.550 533.400 61.350 545.400 ;
        RECT 62.550 533.400 64.350 546.000 ;
        RECT 67.350 539.400 69.150 545.400 ;
        RECT 71.850 539.400 73.650 546.000 ;
        RECT 67.350 537.300 69.450 539.400 ;
        RECT 74.850 538.500 76.650 545.400 ;
        RECT 77.850 539.400 79.650 546.000 ;
        RECT 73.950 537.450 80.550 538.500 ;
        RECT 73.950 536.700 75.750 537.450 ;
        RECT 78.750 536.700 80.550 537.450 ;
        RECT 82.650 536.400 84.450 545.400 ;
        RECT 66.450 534.600 69.450 536.400 ;
        RECT 70.350 535.800 72.150 536.400 ;
        RECT 70.350 534.900 76.050 535.800 ;
        RECT 82.650 535.500 84.750 536.400 ;
        RECT 70.350 534.600 72.150 534.900 ;
        RECT 68.250 533.700 69.450 534.600 ;
        RECT 59.550 526.050 60.750 533.400 ;
        RECT 68.250 532.800 73.050 533.700 ;
        RECT 61.650 530.100 63.450 530.550 ;
        RECT 67.350 530.100 69.450 530.700 ;
        RECT 61.650 528.900 69.450 530.100 ;
        RECT 61.650 528.750 63.450 528.900 ;
        RECT 67.350 528.600 69.450 528.900 ;
        RECT 59.550 525.750 64.050 526.050 ;
        RECT 59.550 523.950 65.850 525.750 ;
        RECT 59.550 516.600 60.750 523.950 ;
        RECT 72.150 520.200 73.050 532.800 ;
        RECT 75.150 532.800 76.050 534.900 ;
        RECT 76.950 534.300 84.750 535.500 ;
        RECT 76.950 533.700 78.750 534.300 ;
        RECT 88.050 533.400 89.850 546.000 ;
        RECT 91.050 535.200 92.850 545.400 ;
        RECT 91.050 533.400 93.450 535.200 ;
        RECT 110.100 533.400 111.900 546.000 ;
        RECT 115.200 534.600 117.000 545.400 ;
        RECT 113.400 533.400 117.000 534.600 ;
        RECT 131.100 533.400 132.900 545.400 ;
        RECT 134.100 534.300 135.900 545.400 ;
        RECT 137.100 535.200 138.900 546.000 ;
        RECT 140.100 534.300 141.900 545.400 ;
        RECT 155.100 539.400 156.900 546.000 ;
        RECT 158.100 539.400 159.900 545.400 ;
        RECT 161.100 540.000 162.900 546.000 ;
        RECT 158.400 539.100 159.900 539.400 ;
        RECT 164.100 539.400 165.900 545.400 ;
        RECT 179.100 539.400 180.900 545.400 ;
        RECT 182.100 539.400 183.900 546.000 ;
        RECT 164.100 539.100 165.000 539.400 ;
        RECT 158.400 538.200 165.000 539.100 ;
        RECT 134.100 533.400 141.900 534.300 ;
        RECT 75.150 532.500 83.550 532.800 ;
        RECT 92.550 532.500 93.450 533.400 ;
        RECT 75.150 531.900 93.450 532.500 ;
        RECT 81.750 531.300 93.450 531.900 ;
        RECT 81.750 531.000 83.550 531.300 ;
        RECT 79.800 524.400 81.900 526.050 ;
        RECT 79.800 523.200 87.900 524.400 ;
        RECT 88.950 523.950 91.050 526.050 ;
        RECT 86.100 522.600 87.900 523.200 ;
        RECT 83.100 521.400 84.900 522.000 ;
        RECT 89.250 521.400 91.050 523.950 ;
        RECT 83.100 520.200 91.050 521.400 ;
        RECT 72.150 519.000 84.150 520.200 ;
        RECT 72.150 518.400 73.950 519.000 ;
        RECT 83.100 517.200 84.150 519.000 ;
        RECT 55.050 510.600 56.850 514.800 ;
        RECT 59.550 510.600 61.350 516.600 ;
        RECT 62.850 510.000 64.650 516.600 ;
        RECT 67.350 513.600 69.750 515.700 ;
        RECT 79.350 515.550 81.150 516.300 ;
        RECT 76.200 514.500 81.150 515.550 ;
        RECT 82.350 515.400 84.150 517.200 ;
        RECT 92.550 516.600 93.450 531.300 ;
        RECT 110.250 526.050 112.050 527.850 ;
        RECT 113.400 526.050 114.300 533.400 ;
        RECT 116.100 526.050 117.900 527.850 ;
        RECT 131.400 526.050 132.300 533.400 ;
        RECT 136.950 526.050 138.750 527.850 ;
        RECT 158.100 526.050 159.900 527.850 ;
        RECT 164.100 526.050 165.000 538.200 ;
        RECT 179.700 526.050 180.900 539.400 ;
        RECT 197.100 533.400 198.900 546.000 ;
        RECT 200.100 532.500 201.900 545.400 ;
        RECT 203.100 533.400 204.900 546.000 ;
        RECT 206.100 532.500 207.900 545.400 ;
        RECT 209.100 533.400 210.900 546.000 ;
        RECT 212.100 532.500 213.900 545.400 ;
        RECT 215.100 533.400 216.900 546.000 ;
        RECT 218.100 532.500 219.900 545.400 ;
        RECT 221.100 533.400 222.900 546.000 ;
        RECT 236.100 539.400 237.900 545.400 ;
        RECT 199.050 531.300 201.900 532.500 ;
        RECT 204.000 531.300 207.900 532.500 ;
        RECT 210.000 531.300 213.900 532.500 ;
        RECT 216.000 531.300 219.900 532.500 ;
        RECT 236.100 532.500 237.300 539.400 ;
        RECT 239.100 535.200 240.900 546.000 ;
        RECT 242.100 533.400 243.900 545.400 ;
        RECT 257.100 539.400 258.900 546.000 ;
        RECT 260.100 539.400 261.900 545.400 ;
        RECT 236.100 531.600 241.800 532.500 ;
        RECT 182.100 526.050 183.900 527.850 ;
        RECT 199.050 526.050 200.100 531.300 ;
        RECT 109.950 523.950 112.050 526.050 ;
        RECT 112.950 523.950 115.050 526.050 ;
        RECT 115.950 523.950 118.050 526.050 ;
        RECT 130.950 523.950 133.050 526.050 ;
        RECT 133.950 523.950 136.050 526.050 ;
        RECT 136.950 523.950 139.050 526.050 ;
        RECT 139.950 523.950 142.050 526.050 ;
        RECT 154.950 523.950 157.050 526.050 ;
        RECT 157.950 523.950 160.050 526.050 ;
        RECT 160.950 523.950 163.050 526.050 ;
        RECT 163.950 523.950 166.050 526.050 ;
        RECT 178.950 523.950 181.050 526.050 ;
        RECT 181.950 523.950 184.050 526.050 ;
        RECT 199.050 523.950 202.200 526.050 ;
        RECT 76.200 513.600 77.250 514.500 ;
        RECT 85.050 514.200 87.150 515.700 ;
        RECT 83.250 513.600 87.150 514.200 ;
        RECT 67.950 510.600 69.750 513.600 ;
        RECT 72.450 510.000 74.250 513.600 ;
        RECT 75.450 510.600 77.250 513.600 ;
        RECT 78.750 510.000 80.550 513.600 ;
        RECT 83.250 512.700 86.850 513.600 ;
        RECT 83.250 510.600 85.050 512.700 ;
        RECT 88.050 510.000 89.850 516.600 ;
        RECT 91.050 514.800 93.450 516.600 ;
        RECT 91.050 510.600 92.850 514.800 ;
        RECT 113.400 513.600 114.300 523.950 ;
        RECT 131.400 516.600 132.300 523.950 ;
        RECT 133.950 522.150 135.750 523.950 ;
        RECT 140.100 522.150 141.900 523.950 ;
        RECT 155.100 522.150 156.900 523.950 ;
        RECT 161.100 522.150 162.900 523.950 ;
        RECT 164.100 520.200 165.000 523.950 ;
        RECT 131.400 515.400 136.500 516.600 ;
        RECT 110.100 510.000 111.900 513.600 ;
        RECT 113.100 510.600 114.900 513.600 ;
        RECT 116.100 510.000 117.900 513.600 ;
        RECT 131.700 510.000 133.500 513.600 ;
        RECT 134.700 510.600 136.500 515.400 ;
        RECT 139.200 510.000 141.000 516.600 ;
        RECT 155.100 510.000 156.900 519.600 ;
        RECT 161.700 519.000 165.000 520.200 ;
        RECT 161.700 510.600 163.500 519.000 ;
        RECT 179.700 513.600 180.900 523.950 ;
        RECT 199.050 518.700 200.100 523.950 ;
        RECT 201.000 520.800 202.800 521.400 ;
        RECT 204.000 520.800 205.200 531.300 ;
        RECT 201.000 519.600 205.200 520.800 ;
        RECT 207.000 520.800 208.800 521.400 ;
        RECT 210.000 520.800 211.200 531.300 ;
        RECT 207.000 519.600 211.200 520.800 ;
        RECT 213.000 520.800 214.800 521.400 ;
        RECT 216.000 520.800 217.200 531.300 ;
        RECT 240.000 530.700 241.800 531.600 ;
        RECT 236.400 526.050 238.200 527.850 ;
        RECT 218.100 523.950 220.200 526.050 ;
        RECT 236.400 523.950 238.500 526.050 ;
        RECT 218.400 522.150 220.200 523.950 ;
        RECT 213.000 519.600 217.200 520.800 ;
        RECT 204.000 518.700 205.200 519.600 ;
        RECT 210.000 518.700 211.200 519.600 ;
        RECT 216.000 518.700 217.200 519.600 ;
        RECT 240.000 519.300 240.900 530.700 ;
        RECT 242.700 526.050 243.900 533.400 ;
        RECT 257.100 526.050 258.900 527.850 ;
        RECT 260.100 526.050 261.300 539.400 ;
        RECT 275.100 533.400 276.900 546.000 ;
        RECT 280.200 534.600 282.000 545.400 ;
        RECT 278.400 533.400 282.000 534.600 ;
        RECT 296.100 534.300 297.900 545.400 ;
        RECT 299.100 535.200 300.900 546.000 ;
        RECT 302.100 534.300 303.900 545.400 ;
        RECT 296.100 533.400 303.900 534.300 ;
        RECT 305.100 533.400 306.900 545.400 ;
        RECT 323.100 539.400 324.900 546.000 ;
        RECT 326.100 539.400 327.900 545.400 ;
        RECT 329.100 539.400 330.900 546.000 ;
        RECT 344.100 539.400 345.900 546.000 ;
        RECT 347.100 539.400 348.900 545.400 ;
        RECT 350.100 539.400 351.900 546.000 ;
        RECT 365.100 539.400 366.900 546.000 ;
        RECT 368.100 539.400 369.900 545.400 ;
        RECT 371.100 540.000 372.900 546.000 ;
        RECT 275.250 526.050 277.050 527.850 ;
        RECT 278.400 526.050 279.300 533.400 ;
        RECT 281.100 526.050 282.900 527.850 ;
        RECT 299.250 526.050 301.050 527.850 ;
        RECT 305.700 526.050 306.600 533.400 ;
        RECT 326.700 526.050 327.900 539.400 ;
        RECT 347.700 526.050 348.900 539.400 ;
        RECT 368.400 539.100 369.900 539.400 ;
        RECT 374.100 539.400 375.900 545.400 ;
        RECT 374.100 539.100 375.000 539.400 ;
        RECT 368.400 538.200 375.000 539.100 ;
        RECT 368.100 526.050 369.900 527.850 ;
        RECT 374.100 526.050 375.000 538.200 ;
        RECT 389.100 534.300 390.900 545.400 ;
        RECT 392.100 535.200 393.900 546.000 ;
        RECT 395.100 534.300 396.900 545.400 ;
        RECT 389.100 533.400 396.900 534.300 ;
        RECT 398.100 533.400 399.900 545.400 ;
        RECT 413.400 533.400 415.200 546.000 ;
        RECT 418.500 534.900 420.300 545.400 ;
        RECT 421.500 539.400 423.300 546.000 ;
        RECT 421.200 536.100 423.000 537.900 ;
        RECT 418.500 533.400 420.900 534.900 ;
        RECT 437.400 533.400 439.200 546.000 ;
        RECT 442.500 534.900 444.300 545.400 ;
        RECT 445.500 539.400 447.300 546.000 ;
        RECT 464.100 539.400 465.900 546.000 ;
        RECT 467.100 539.400 468.900 545.400 ;
        RECT 470.100 540.000 471.900 546.000 ;
        RECT 467.400 539.100 468.900 539.400 ;
        RECT 473.100 539.400 474.900 545.400 ;
        RECT 488.100 539.400 489.900 546.000 ;
        RECT 491.100 539.400 492.900 545.400 ;
        RECT 494.100 540.000 495.900 546.000 ;
        RECT 473.100 539.100 474.000 539.400 ;
        RECT 467.400 538.200 474.000 539.100 ;
        RECT 491.400 539.100 492.900 539.400 ;
        RECT 497.100 539.400 498.900 545.400 ;
        RECT 512.100 539.400 513.900 546.000 ;
        RECT 515.100 539.400 516.900 545.400 ;
        RECT 518.100 540.000 519.900 546.000 ;
        RECT 497.100 539.100 498.000 539.400 ;
        RECT 491.400 538.200 498.000 539.100 ;
        RECT 515.400 539.100 516.900 539.400 ;
        RECT 521.100 539.400 522.900 545.400 ;
        RECT 536.100 539.400 537.900 546.000 ;
        RECT 539.100 539.400 540.900 545.400 ;
        RECT 554.100 539.400 555.900 546.000 ;
        RECT 557.100 539.400 558.900 545.400 ;
        RECT 560.100 540.000 561.900 546.000 ;
        RECT 521.100 539.100 522.000 539.400 ;
        RECT 515.400 538.200 522.000 539.100 ;
        RECT 445.200 536.100 447.000 537.900 ;
        RECT 442.500 533.400 444.900 534.900 ;
        RECT 392.250 526.050 394.050 527.850 ;
        RECT 398.700 526.050 399.600 533.400 ;
        RECT 413.100 526.050 414.900 527.850 ;
        RECT 419.700 526.050 420.900 533.400 ;
        RECT 437.100 526.050 438.900 527.850 ;
        RECT 443.700 526.050 444.900 533.400 ;
        RECT 448.950 531.450 451.050 532.050 ;
        RECT 469.950 531.450 472.050 532.200 ;
        RECT 448.950 530.550 472.050 531.450 ;
        RECT 448.950 529.950 451.050 530.550 ;
        RECT 469.950 530.100 472.050 530.550 ;
        RECT 467.100 526.050 468.900 527.850 ;
        RECT 473.100 526.050 474.000 538.200 ;
        RECT 475.950 531.450 478.050 532.050 ;
        RECT 493.950 531.450 496.050 532.050 ;
        RECT 475.950 530.550 496.050 531.450 ;
        RECT 475.950 529.950 478.050 530.550 ;
        RECT 493.950 529.950 496.050 530.550 ;
        RECT 491.100 526.050 492.900 527.850 ;
        RECT 497.100 526.050 498.000 538.200 ;
        RECT 515.100 526.050 516.900 527.850 ;
        RECT 521.100 526.050 522.000 538.200 ;
        RECT 531.000 528.450 535.050 529.050 ;
        RECT 530.550 526.950 535.050 528.450 ;
        RECT 241.800 523.950 243.900 526.050 ;
        RECT 256.950 523.950 259.050 526.050 ;
        RECT 259.950 523.950 262.050 526.050 ;
        RECT 274.950 523.950 277.050 526.050 ;
        RECT 277.950 523.950 280.050 526.050 ;
        RECT 280.950 523.950 283.050 526.050 ;
        RECT 295.950 523.950 298.050 526.050 ;
        RECT 298.950 523.950 301.050 526.050 ;
        RECT 301.950 523.950 304.050 526.050 ;
        RECT 304.950 523.950 307.050 526.050 ;
        RECT 322.950 523.950 325.050 526.050 ;
        RECT 325.950 523.950 328.050 526.050 ;
        RECT 328.950 523.950 331.050 526.050 ;
        RECT 343.950 523.950 346.050 526.050 ;
        RECT 346.950 523.950 349.050 526.050 ;
        RECT 349.950 523.950 352.050 526.050 ;
        RECT 364.950 523.950 367.050 526.050 ;
        RECT 367.950 523.950 370.050 526.050 ;
        RECT 370.950 523.950 373.050 526.050 ;
        RECT 373.950 523.950 376.050 526.050 ;
        RECT 388.950 523.950 391.050 526.050 ;
        RECT 391.950 523.950 394.050 526.050 ;
        RECT 394.950 523.950 397.050 526.050 ;
        RECT 397.950 523.950 400.050 526.050 ;
        RECT 412.950 523.950 415.050 526.050 ;
        RECT 415.950 523.950 418.050 526.050 ;
        RECT 418.950 523.950 421.050 526.050 ;
        RECT 421.950 523.950 424.050 526.050 ;
        RECT 436.950 523.950 439.050 526.050 ;
        RECT 439.950 523.950 442.050 526.050 ;
        RECT 442.950 523.950 445.050 526.050 ;
        RECT 445.950 523.950 448.050 526.050 ;
        RECT 463.950 523.950 466.050 526.050 ;
        RECT 466.950 523.950 469.050 526.050 ;
        RECT 469.950 523.950 472.050 526.050 ;
        RECT 472.950 523.950 475.050 526.050 ;
        RECT 487.950 523.950 490.050 526.050 ;
        RECT 490.950 523.950 493.050 526.050 ;
        RECT 493.950 523.950 496.050 526.050 ;
        RECT 496.950 523.950 499.050 526.050 ;
        RECT 511.950 523.950 514.050 526.050 ;
        RECT 514.950 523.950 517.050 526.050 ;
        RECT 517.950 523.950 520.050 526.050 ;
        RECT 520.950 523.950 523.050 526.050 ;
        RECT 199.050 517.500 201.900 518.700 ;
        RECT 204.000 517.500 207.900 518.700 ;
        RECT 210.000 517.500 213.900 518.700 ;
        RECT 216.000 517.500 219.900 518.700 ;
        RECT 240.000 518.400 241.800 519.300 ;
        RECT 179.100 510.600 180.900 513.600 ;
        RECT 182.100 510.000 183.900 513.600 ;
        RECT 197.100 510.000 198.900 516.600 ;
        RECT 200.100 510.600 201.900 517.500 ;
        RECT 203.100 510.000 204.900 516.600 ;
        RECT 206.100 510.600 207.900 517.500 ;
        RECT 209.100 510.000 210.900 516.600 ;
        RECT 212.100 510.600 213.900 517.500 ;
        RECT 215.100 510.000 216.900 516.600 ;
        RECT 218.100 510.600 219.900 517.500 ;
        RECT 236.100 517.500 241.800 518.400 ;
        RECT 221.100 510.000 222.900 516.600 ;
        RECT 236.100 513.600 237.300 517.500 ;
        RECT 242.700 516.600 243.900 523.950 ;
        RECT 236.100 510.600 237.900 513.600 ;
        RECT 239.100 510.000 240.900 516.600 ;
        RECT 242.100 510.600 243.900 516.600 ;
        RECT 260.100 513.600 261.300 523.950 ;
        RECT 278.400 513.600 279.300 523.950 ;
        RECT 296.100 522.150 297.900 523.950 ;
        RECT 302.250 522.150 304.050 523.950 ;
        RECT 305.700 516.600 306.600 523.950 ;
        RECT 323.100 522.150 324.900 523.950 ;
        RECT 326.700 518.700 327.900 523.950 ;
        RECT 328.950 522.150 330.750 523.950 ;
        RECT 344.100 522.150 345.900 523.950 ;
        RECT 347.700 518.700 348.900 523.950 ;
        RECT 349.950 522.150 351.750 523.950 ;
        RECT 365.100 522.150 366.900 523.950 ;
        RECT 371.100 522.150 372.900 523.950 ;
        RECT 374.100 520.200 375.000 523.950 ;
        RECT 389.100 522.150 390.900 523.950 ;
        RECT 395.250 522.150 397.050 523.950 ;
        RECT 257.100 510.000 258.900 513.600 ;
        RECT 260.100 510.600 261.900 513.600 ;
        RECT 275.100 510.000 276.900 513.600 ;
        RECT 278.100 510.600 279.900 513.600 ;
        RECT 281.100 510.000 282.900 513.600 ;
        RECT 297.000 510.000 298.800 516.600 ;
        RECT 301.500 515.400 306.600 516.600 ;
        RECT 323.700 517.800 327.900 518.700 ;
        RECT 344.700 517.800 348.900 518.700 ;
        RECT 301.500 510.600 303.300 515.400 ;
        RECT 304.500 510.000 306.300 513.600 ;
        RECT 323.700 510.600 325.500 517.800 ;
        RECT 328.800 510.000 330.600 516.600 ;
        RECT 344.700 510.600 346.500 517.800 ;
        RECT 349.800 510.000 351.600 516.600 ;
        RECT 365.100 510.000 366.900 519.600 ;
        RECT 371.700 519.000 375.000 520.200 ;
        RECT 371.700 510.600 373.500 519.000 ;
        RECT 398.700 516.600 399.600 523.950 ;
        RECT 416.100 522.150 417.900 523.950 ;
        RECT 419.700 519.600 420.900 523.950 ;
        RECT 422.100 522.150 423.900 523.950 ;
        RECT 440.100 522.150 441.900 523.950 ;
        RECT 443.700 519.600 444.900 523.950 ;
        RECT 446.100 522.150 447.900 523.950 ;
        RECT 464.100 522.150 465.900 523.950 ;
        RECT 470.100 522.150 471.900 523.950 ;
        RECT 473.100 520.200 474.000 523.950 ;
        RECT 488.100 522.150 489.900 523.950 ;
        RECT 494.100 522.150 495.900 523.950 ;
        RECT 497.100 520.200 498.000 523.950 ;
        RECT 512.100 522.150 513.900 523.950 ;
        RECT 518.100 522.150 519.900 523.950 ;
        RECT 521.100 520.200 522.000 523.950 ;
        RECT 530.550 523.050 531.450 526.950 ;
        RECT 536.100 526.050 537.900 527.850 ;
        RECT 539.100 526.050 540.300 539.400 ;
        RECT 557.400 539.100 558.900 539.400 ;
        RECT 563.100 539.400 564.900 545.400 ;
        RECT 578.100 539.400 579.900 546.000 ;
        RECT 581.100 539.400 582.900 545.400 ;
        RECT 584.100 539.400 585.900 546.000 ;
        RECT 599.100 539.400 600.900 546.000 ;
        RECT 602.100 539.400 603.900 545.400 ;
        RECT 605.100 539.400 606.900 546.000 ;
        RECT 623.700 539.400 625.500 546.000 ;
        RECT 563.100 539.100 564.000 539.400 ;
        RECT 557.400 538.200 564.000 539.100 ;
        RECT 541.950 531.450 544.050 532.050 ;
        RECT 559.950 531.450 562.050 532.050 ;
        RECT 541.950 530.550 562.050 531.450 ;
        RECT 541.950 529.950 544.050 530.550 ;
        RECT 559.950 529.950 562.050 530.550 ;
        RECT 544.950 528.450 547.050 529.050 ;
        RECT 550.950 528.450 553.050 529.050 ;
        RECT 544.950 527.550 553.050 528.450 ;
        RECT 544.950 526.950 547.050 527.550 ;
        RECT 550.950 526.950 553.050 527.550 ;
        RECT 557.100 526.050 558.900 527.850 ;
        RECT 563.100 526.050 564.000 538.200 ;
        RECT 581.100 526.050 582.300 539.400 ;
        RECT 602.100 526.050 603.300 539.400 ;
        RECT 624.000 536.100 625.800 537.900 ;
        RECT 626.700 534.900 628.500 545.400 ;
        RECT 626.100 533.400 628.500 534.900 ;
        RECT 631.800 533.400 633.600 546.000 ;
        RECT 647.100 539.400 648.900 546.000 ;
        RECT 650.100 539.400 651.900 545.400 ;
        RECT 653.100 539.400 654.900 546.000 ;
        RECT 668.100 539.400 669.900 546.000 ;
        RECT 671.100 539.400 672.900 545.400 ;
        RECT 674.100 539.400 675.900 546.000 ;
        RECT 689.100 539.400 690.900 546.000 ;
        RECT 692.100 539.400 693.900 545.400 ;
        RECT 626.100 526.050 627.300 533.400 ;
        RECT 632.100 526.050 633.900 527.850 ;
        RECT 650.100 526.050 651.300 539.400 ;
        RECT 671.700 526.050 672.900 539.400 ;
        RECT 535.950 523.950 538.050 526.050 ;
        RECT 538.950 523.950 541.050 526.050 ;
        RECT 553.950 523.950 556.050 526.050 ;
        RECT 556.950 523.950 559.050 526.050 ;
        RECT 559.950 523.950 562.050 526.050 ;
        RECT 562.950 523.950 565.050 526.050 ;
        RECT 577.950 523.950 580.050 526.050 ;
        RECT 580.950 523.950 583.050 526.050 ;
        RECT 583.950 523.950 586.050 526.050 ;
        RECT 598.950 523.950 601.050 526.050 ;
        RECT 601.950 523.950 604.050 526.050 ;
        RECT 604.950 523.950 607.050 526.050 ;
        RECT 622.950 523.950 625.050 526.050 ;
        RECT 625.950 523.950 628.050 526.050 ;
        RECT 628.950 523.950 631.050 526.050 ;
        RECT 631.950 523.950 634.050 526.050 ;
        RECT 646.950 523.950 649.050 526.050 ;
        RECT 649.950 523.950 652.050 526.050 ;
        RECT 652.950 523.950 655.050 526.050 ;
        RECT 667.950 523.950 670.050 526.050 ;
        RECT 670.950 523.950 673.050 526.050 ;
        RECT 673.950 523.950 676.050 526.050 ;
        RECT 689.100 523.950 691.200 526.050 ;
        RECT 530.550 521.550 535.050 523.050 ;
        RECT 531.000 520.950 535.050 521.550 ;
        RECT 419.700 518.700 423.300 519.600 ;
        RECT 443.700 518.700 447.300 519.600 ;
        RECT 390.000 510.000 391.800 516.600 ;
        RECT 394.500 515.400 399.600 516.600 ;
        RECT 413.100 515.700 420.900 517.050 ;
        RECT 394.500 510.600 396.300 515.400 ;
        RECT 397.500 510.000 399.300 513.600 ;
        RECT 413.100 510.600 414.900 515.700 ;
        RECT 416.100 510.000 417.900 514.800 ;
        RECT 419.100 510.600 420.900 515.700 ;
        RECT 422.100 516.600 423.300 518.700 ;
        RECT 422.100 510.600 423.900 516.600 ;
        RECT 437.100 515.700 444.900 517.050 ;
        RECT 437.100 510.600 438.900 515.700 ;
        RECT 440.100 510.000 441.900 514.800 ;
        RECT 443.100 510.600 444.900 515.700 ;
        RECT 446.100 516.600 447.300 518.700 ;
        RECT 446.100 510.600 447.900 516.600 ;
        RECT 464.100 510.000 465.900 519.600 ;
        RECT 470.700 519.000 474.000 520.200 ;
        RECT 470.700 510.600 472.500 519.000 ;
        RECT 488.100 510.000 489.900 519.600 ;
        RECT 494.700 519.000 498.000 520.200 ;
        RECT 494.700 510.600 496.500 519.000 ;
        RECT 512.100 510.000 513.900 519.600 ;
        RECT 518.700 519.000 522.000 520.200 ;
        RECT 523.950 519.450 526.050 520.050 ;
        RECT 529.950 519.450 532.050 520.050 ;
        RECT 518.700 510.600 520.500 519.000 ;
        RECT 523.950 518.550 532.050 519.450 ;
        RECT 523.950 517.950 526.050 518.550 ;
        RECT 529.950 517.950 532.050 518.550 ;
        RECT 539.100 513.600 540.300 523.950 ;
        RECT 554.100 522.150 555.900 523.950 ;
        RECT 560.100 522.150 561.900 523.950 ;
        RECT 563.100 520.200 564.000 523.950 ;
        RECT 578.250 522.150 580.050 523.950 ;
        RECT 536.100 510.000 537.900 513.600 ;
        RECT 539.100 510.600 540.900 513.600 ;
        RECT 541.950 513.450 544.050 514.050 ;
        RECT 550.950 513.450 553.050 513.900 ;
        RECT 541.950 512.550 553.050 513.450 ;
        RECT 541.950 511.950 544.050 512.550 ;
        RECT 550.950 511.800 553.050 512.550 ;
        RECT 554.100 510.000 555.900 519.600 ;
        RECT 560.700 519.000 564.000 520.200 ;
        RECT 560.700 510.600 562.500 519.000 ;
        RECT 581.100 518.700 582.300 523.950 ;
        RECT 584.100 522.150 585.900 523.950 ;
        RECT 599.250 522.150 601.050 523.950 ;
        RECT 602.100 518.700 603.300 523.950 ;
        RECT 605.100 522.150 606.900 523.950 ;
        RECT 623.100 522.150 624.900 523.950 ;
        RECT 626.100 519.600 627.300 523.950 ;
        RECT 629.100 522.150 630.900 523.950 ;
        RECT 647.250 522.150 649.050 523.950 ;
        RECT 623.700 518.700 627.300 519.600 ;
        RECT 650.100 518.700 651.300 523.950 ;
        RECT 653.100 522.150 654.900 523.950 ;
        RECT 668.100 522.150 669.900 523.950 ;
        RECT 671.700 518.700 672.900 523.950 ;
        RECT 673.950 522.150 675.750 523.950 ;
        RECT 689.250 522.150 691.050 523.950 ;
        RECT 692.100 519.300 693.000 539.400 ;
        RECT 695.100 534.000 696.900 546.000 ;
        RECT 698.100 533.400 699.900 545.400 ;
        RECT 713.400 533.400 715.200 546.000 ;
        RECT 718.500 534.900 720.300 545.400 ;
        RECT 721.500 539.400 723.300 546.000 ;
        RECT 740.100 539.400 741.900 546.000 ;
        RECT 743.100 539.400 744.900 545.400 ;
        RECT 746.100 540.000 747.900 546.000 ;
        RECT 743.400 539.100 744.900 539.400 ;
        RECT 749.100 539.400 750.900 545.400 ;
        RECT 749.100 539.100 750.000 539.400 ;
        RECT 743.400 538.200 750.000 539.100 ;
        RECT 721.200 536.100 723.000 537.900 ;
        RECT 718.500 533.400 720.900 534.900 ;
        RECT 694.200 526.050 696.000 527.850 ;
        RECT 698.400 526.050 699.300 533.400 ;
        RECT 713.100 526.050 714.900 527.850 ;
        RECT 719.700 526.050 720.900 533.400 ;
        RECT 743.100 526.050 744.900 527.850 ;
        RECT 749.100 526.050 750.000 538.200 ;
        RECT 767.100 534.300 768.900 545.400 ;
        RECT 770.100 535.200 771.900 546.000 ;
        RECT 773.100 534.300 774.900 545.400 ;
        RECT 767.100 533.400 774.900 534.300 ;
        RECT 776.100 533.400 777.900 545.400 ;
        RECT 791.100 533.400 792.900 545.400 ;
        RECT 794.100 534.300 795.900 545.400 ;
        RECT 797.100 535.200 798.900 546.000 ;
        RECT 800.100 534.300 801.900 545.400 ;
        RECT 815.100 539.400 816.900 545.400 ;
        RECT 818.100 540.000 819.900 546.000 ;
        RECT 794.100 533.400 801.900 534.300 ;
        RECT 816.000 539.100 816.900 539.400 ;
        RECT 821.100 539.400 822.900 545.400 ;
        RECT 824.100 539.400 825.900 546.000 ;
        RECT 839.100 539.400 840.900 545.400 ;
        RECT 842.100 540.000 843.900 546.000 ;
        RECT 821.100 539.100 822.600 539.400 ;
        RECT 816.000 538.200 822.600 539.100 ;
        RECT 840.000 539.100 840.900 539.400 ;
        RECT 845.100 539.400 846.900 545.400 ;
        RECT 848.100 539.400 849.900 546.000 ;
        RECT 845.100 539.100 846.600 539.400 ;
        RECT 840.000 538.200 846.600 539.100 ;
        RECT 754.950 528.450 757.050 529.050 ;
        RECT 763.950 528.450 766.050 529.050 ;
        RECT 754.950 527.550 766.050 528.450 ;
        RECT 754.950 526.950 757.050 527.550 ;
        RECT 763.950 526.950 766.050 527.550 ;
        RECT 770.250 526.050 772.050 527.850 ;
        RECT 776.700 526.050 777.600 533.400 ;
        RECT 778.950 528.450 781.050 529.050 ;
        RECT 784.950 528.450 787.050 528.900 ;
        RECT 778.950 527.550 787.050 528.450 ;
        RECT 778.950 526.950 781.050 527.550 ;
        RECT 784.950 526.800 787.050 527.550 ;
        RECT 791.400 526.050 792.300 533.400 ;
        RECT 796.950 526.050 798.750 527.850 ;
        RECT 816.000 526.050 816.900 538.200 ;
        RECT 834.000 528.450 838.050 529.050 ;
        RECT 821.100 526.050 822.900 527.850 ;
        RECT 833.550 526.950 838.050 528.450 ;
        RECT 694.500 523.950 696.600 526.050 ;
        RECT 697.800 523.950 699.900 526.050 ;
        RECT 712.950 523.950 715.050 526.050 ;
        RECT 715.950 523.950 718.050 526.050 ;
        RECT 718.950 523.950 721.050 526.050 ;
        RECT 721.950 523.950 724.050 526.050 ;
        RECT 739.950 523.950 742.050 526.050 ;
        RECT 742.950 523.950 745.050 526.050 ;
        RECT 745.950 523.950 748.050 526.050 ;
        RECT 748.950 523.950 751.050 526.050 ;
        RECT 766.950 523.950 769.050 526.050 ;
        RECT 769.950 523.950 772.050 526.050 ;
        RECT 772.950 523.950 775.050 526.050 ;
        RECT 775.950 523.950 778.050 526.050 ;
        RECT 790.950 523.950 793.050 526.050 ;
        RECT 793.950 523.950 796.050 526.050 ;
        RECT 796.950 523.950 799.050 526.050 ;
        RECT 799.950 523.950 802.050 526.050 ;
        RECT 814.950 523.950 817.050 526.050 ;
        RECT 817.950 523.950 820.050 526.050 ;
        RECT 820.950 523.950 823.050 526.050 ;
        RECT 823.950 523.950 826.050 526.050 ;
        RECT 581.100 517.800 585.300 518.700 ;
        RECT 602.100 517.800 606.300 518.700 ;
        RECT 578.400 510.000 580.200 516.600 ;
        RECT 583.500 510.600 585.300 517.800 ;
        RECT 599.400 510.000 601.200 516.600 ;
        RECT 604.500 510.600 606.300 517.800 ;
        RECT 623.700 516.600 624.900 518.700 ;
        RECT 650.100 517.800 654.300 518.700 ;
        RECT 623.100 510.600 624.900 516.600 ;
        RECT 626.100 515.700 633.900 517.050 ;
        RECT 626.100 510.600 627.900 515.700 ;
        RECT 629.100 510.000 630.900 514.800 ;
        RECT 632.100 510.600 633.900 515.700 ;
        RECT 647.400 510.000 649.200 516.600 ;
        RECT 652.500 510.600 654.300 517.800 ;
        RECT 668.700 517.800 672.900 518.700 ;
        RECT 689.100 518.400 697.500 519.300 ;
        RECT 668.700 510.600 670.500 517.800 ;
        RECT 673.800 510.000 675.600 516.600 ;
        RECT 689.100 510.600 690.900 518.400 ;
        RECT 695.700 517.500 697.500 518.400 ;
        RECT 698.400 516.600 699.300 523.950 ;
        RECT 716.100 522.150 717.900 523.950 ;
        RECT 719.700 519.600 720.900 523.950 ;
        RECT 722.100 522.150 723.900 523.950 ;
        RECT 740.100 522.150 741.900 523.950 ;
        RECT 746.100 522.150 747.900 523.950 ;
        RECT 749.100 520.200 750.000 523.950 ;
        RECT 767.100 522.150 768.900 523.950 ;
        RECT 773.250 522.150 775.050 523.950 ;
        RECT 719.700 518.700 723.300 519.600 ;
        RECT 693.600 510.000 695.400 516.600 ;
        RECT 696.600 514.800 699.300 516.600 ;
        RECT 713.100 515.700 720.900 517.050 ;
        RECT 696.600 510.600 698.400 514.800 ;
        RECT 713.100 510.600 714.900 515.700 ;
        RECT 716.100 510.000 717.900 514.800 ;
        RECT 719.100 510.600 720.900 515.700 ;
        RECT 722.100 516.600 723.300 518.700 ;
        RECT 722.100 510.600 723.900 516.600 ;
        RECT 740.100 510.000 741.900 519.600 ;
        RECT 746.700 519.000 750.000 520.200 ;
        RECT 746.700 510.600 748.500 519.000 ;
        RECT 776.700 516.600 777.600 523.950 ;
        RECT 768.000 510.000 769.800 516.600 ;
        RECT 772.500 515.400 777.600 516.600 ;
        RECT 791.400 516.600 792.300 523.950 ;
        RECT 793.950 522.150 795.750 523.950 ;
        RECT 800.100 522.150 801.900 523.950 ;
        RECT 816.000 520.200 816.900 523.950 ;
        RECT 818.100 522.150 819.900 523.950 ;
        RECT 824.100 522.150 825.900 523.950 ;
        RECT 833.550 523.050 834.450 526.950 ;
        RECT 840.000 526.050 840.900 538.200 ;
        RECT 863.100 534.300 864.900 545.400 ;
        RECT 866.100 535.200 867.900 546.000 ;
        RECT 869.100 534.300 870.900 545.400 ;
        RECT 863.100 533.400 870.900 534.300 ;
        RECT 872.100 533.400 873.900 545.400 ;
        RECT 887.700 539.400 889.500 546.000 ;
        RECT 888.000 536.100 889.800 537.900 ;
        RECT 890.700 534.900 892.500 545.400 ;
        RECT 890.100 533.400 892.500 534.900 ;
        RECT 895.800 533.400 897.600 546.000 ;
        RECT 847.950 531.450 850.050 532.050 ;
        RECT 853.950 531.450 856.050 532.050 ;
        RECT 868.950 531.450 871.050 532.050 ;
        RECT 847.950 530.550 871.050 531.450 ;
        RECT 847.950 529.950 850.050 530.550 ;
        RECT 853.950 529.950 856.050 530.550 ;
        RECT 868.950 529.950 871.050 530.550 ;
        RECT 845.100 526.050 846.900 527.850 ;
        RECT 866.250 526.050 868.050 527.850 ;
        RECT 872.700 526.050 873.600 533.400 ;
        RECT 882.000 528.450 886.050 529.050 ;
        RECT 881.550 526.950 886.050 528.450 ;
        RECT 838.950 523.950 841.050 526.050 ;
        RECT 841.950 523.950 844.050 526.050 ;
        RECT 844.950 523.950 847.050 526.050 ;
        RECT 847.950 523.950 850.050 526.050 ;
        RECT 862.950 523.950 865.050 526.050 ;
        RECT 865.950 523.950 868.050 526.050 ;
        RECT 868.950 523.950 871.050 526.050 ;
        RECT 871.950 523.950 874.050 526.050 ;
        RECT 833.550 521.550 838.050 523.050 ;
        RECT 834.000 520.950 838.050 521.550 ;
        RECT 840.000 520.200 840.900 523.950 ;
        RECT 842.100 522.150 843.900 523.950 ;
        RECT 848.100 522.150 849.900 523.950 ;
        RECT 863.100 522.150 864.900 523.950 ;
        RECT 869.250 522.150 871.050 523.950 ;
        RECT 816.000 519.000 819.300 520.200 ;
        RECT 791.400 515.400 796.500 516.600 ;
        RECT 772.500 510.600 774.300 515.400 ;
        RECT 775.500 510.000 777.300 513.600 ;
        RECT 791.700 510.000 793.500 513.600 ;
        RECT 794.700 510.600 796.500 515.400 ;
        RECT 799.200 510.000 801.000 516.600 ;
        RECT 817.500 510.600 819.300 519.000 ;
        RECT 824.100 510.000 825.900 519.600 ;
        RECT 840.000 519.000 843.300 520.200 ;
        RECT 841.500 510.600 843.300 519.000 ;
        RECT 848.100 510.000 849.900 519.600 ;
        RECT 850.950 519.450 853.050 520.050 ;
        RECT 865.950 519.450 868.050 520.050 ;
        RECT 850.950 518.550 868.050 519.450 ;
        RECT 850.950 517.950 853.050 518.550 ;
        RECT 865.950 517.950 868.050 518.550 ;
        RECT 872.700 516.600 873.600 523.950 ;
        RECT 874.950 522.450 877.050 523.050 ;
        RECT 881.550 522.450 882.450 526.950 ;
        RECT 890.100 526.050 891.300 533.400 ;
        RECT 896.100 526.050 897.900 527.850 ;
        RECT 886.950 523.950 889.050 526.050 ;
        RECT 889.950 523.950 892.050 526.050 ;
        RECT 892.950 523.950 895.050 526.050 ;
        RECT 895.950 523.950 898.050 526.050 ;
        RECT 874.950 521.550 882.450 522.450 ;
        RECT 887.100 522.150 888.900 523.950 ;
        RECT 874.950 520.950 877.050 521.550 ;
        RECT 890.100 519.600 891.300 523.950 ;
        RECT 893.100 522.150 894.900 523.950 ;
        RECT 887.700 518.700 891.300 519.600 ;
        RECT 887.700 516.600 888.900 518.700 ;
        RECT 864.000 510.000 865.800 516.600 ;
        RECT 868.500 515.400 873.600 516.600 ;
        RECT 868.500 510.600 870.300 515.400 ;
        RECT 871.500 510.000 873.300 513.600 ;
        RECT 887.100 510.600 888.900 516.600 ;
        RECT 890.100 515.700 897.900 517.050 ;
        RECT 890.100 510.600 891.900 515.700 ;
        RECT 893.100 510.000 894.900 514.800 ;
        RECT 896.100 510.600 897.900 515.700 ;
        RECT 14.100 500.400 15.900 506.400 ;
        RECT 17.100 500.400 18.900 507.000 ;
        RECT 20.100 503.400 21.900 506.400 ;
        RECT 14.100 493.050 15.300 500.400 ;
        RECT 20.700 499.500 21.900 503.400 ;
        RECT 16.200 498.600 21.900 499.500 ;
        RECT 23.550 500.400 25.350 506.400 ;
        RECT 26.850 500.400 28.650 507.000 ;
        RECT 31.950 503.400 33.750 506.400 ;
        RECT 36.450 503.400 38.250 507.000 ;
        RECT 39.450 503.400 41.250 506.400 ;
        RECT 42.750 503.400 44.550 507.000 ;
        RECT 47.250 504.300 49.050 506.400 ;
        RECT 47.250 503.400 50.850 504.300 ;
        RECT 31.350 501.300 33.750 503.400 ;
        RECT 40.200 502.500 41.250 503.400 ;
        RECT 47.250 502.800 51.150 503.400 ;
        RECT 40.200 501.450 45.150 502.500 ;
        RECT 43.350 500.700 45.150 501.450 ;
        RECT 16.200 497.700 18.000 498.600 ;
        RECT 14.100 490.950 16.200 493.050 ;
        RECT 14.100 483.600 15.300 490.950 ;
        RECT 17.100 486.300 18.000 497.700 ;
        RECT 23.550 493.050 24.750 500.400 ;
        RECT 46.350 499.800 48.150 501.600 ;
        RECT 49.050 501.300 51.150 502.800 ;
        RECT 52.050 500.400 53.850 507.000 ;
        RECT 55.050 502.200 56.850 506.400 ;
        RECT 55.050 500.400 57.450 502.200 ;
        RECT 36.150 498.000 37.950 498.600 ;
        RECT 47.100 498.000 48.150 499.800 ;
        RECT 36.150 496.800 48.150 498.000 ;
        RECT 19.500 490.950 21.600 493.050 ;
        RECT 19.800 489.150 21.600 490.950 ;
        RECT 23.550 491.250 29.850 493.050 ;
        RECT 23.550 490.950 28.050 491.250 ;
        RECT 16.200 485.400 18.000 486.300 ;
        RECT 16.200 484.500 21.900 485.400 ;
        RECT 14.100 471.600 15.900 483.600 ;
        RECT 17.100 471.000 18.900 481.800 ;
        RECT 20.700 477.600 21.900 484.500 ;
        RECT 20.100 471.600 21.900 477.600 ;
        RECT 23.550 483.600 24.750 490.950 ;
        RECT 25.650 488.100 27.450 488.250 ;
        RECT 31.350 488.100 33.450 488.400 ;
        RECT 25.650 486.900 33.450 488.100 ;
        RECT 25.650 486.450 27.450 486.900 ;
        RECT 31.350 486.300 33.450 486.900 ;
        RECT 36.150 484.200 37.050 496.800 ;
        RECT 47.100 495.600 55.050 496.800 ;
        RECT 47.100 495.000 48.900 495.600 ;
        RECT 50.100 493.800 51.900 494.400 ;
        RECT 43.800 492.600 51.900 493.800 ;
        RECT 53.250 493.050 55.050 495.600 ;
        RECT 43.800 490.950 45.900 492.600 ;
        RECT 52.950 490.950 55.050 493.050 ;
        RECT 45.750 485.700 47.550 486.000 ;
        RECT 56.550 485.700 57.450 500.400 ;
        RECT 76.500 498.000 78.300 506.400 ;
        RECT 75.000 496.800 78.300 498.000 ;
        RECT 83.100 497.400 84.900 507.000 ;
        RECT 99.000 500.400 100.800 507.000 ;
        RECT 103.500 501.600 105.300 506.400 ;
        RECT 106.500 503.400 108.300 507.000 ;
        RECT 122.100 503.400 123.900 507.000 ;
        RECT 125.100 503.400 126.900 506.400 ;
        RECT 103.500 500.400 108.600 501.600 ;
        RECT 75.000 493.050 75.900 496.800 ;
        RECT 77.100 493.050 78.900 494.850 ;
        RECT 83.100 493.050 84.900 494.850 ;
        RECT 98.100 493.050 99.900 494.850 ;
        RECT 104.250 493.050 106.050 494.850 ;
        RECT 107.700 493.050 108.600 500.400 ;
        RECT 125.100 493.050 126.300 503.400 ;
        RECT 142.500 498.000 144.300 506.400 ;
        RECT 141.000 496.800 144.300 498.000 ;
        RECT 149.100 497.400 150.900 507.000 ;
        RECT 167.100 500.400 168.900 507.000 ;
        RECT 170.100 499.500 171.900 506.400 ;
        RECT 173.100 500.400 174.900 507.000 ;
        RECT 176.100 499.500 177.900 506.400 ;
        RECT 179.100 500.400 180.900 507.000 ;
        RECT 182.100 499.500 183.900 506.400 ;
        RECT 185.100 500.400 186.900 507.000 ;
        RECT 188.100 499.500 189.900 506.400 ;
        RECT 191.100 500.400 192.900 507.000 ;
        RECT 169.050 498.300 171.900 499.500 ;
        RECT 174.000 498.300 177.900 499.500 ;
        RECT 180.000 498.300 183.900 499.500 ;
        RECT 186.000 498.300 189.900 499.500 ;
        RECT 209.100 498.600 210.900 506.400 ;
        RECT 213.600 500.400 215.400 507.000 ;
        RECT 216.600 502.200 218.400 506.400 ;
        RECT 216.600 500.400 219.300 502.200 ;
        RECT 215.700 498.600 217.500 499.500 ;
        RECT 141.000 493.050 141.900 496.800 ;
        RECT 143.100 493.050 144.900 494.850 ;
        RECT 149.100 493.050 150.900 494.850 ;
        RECT 169.050 493.050 170.100 498.300 ;
        RECT 174.000 497.400 175.200 498.300 ;
        RECT 180.000 497.400 181.200 498.300 ;
        RECT 186.000 497.400 187.200 498.300 ;
        RECT 209.100 497.700 217.500 498.600 ;
        RECT 171.000 496.200 175.200 497.400 ;
        RECT 171.000 495.600 172.800 496.200 ;
        RECT 73.950 490.950 76.050 493.050 ;
        RECT 76.950 490.950 79.050 493.050 ;
        RECT 79.950 490.950 82.050 493.050 ;
        RECT 82.950 490.950 85.050 493.050 ;
        RECT 97.950 490.950 100.050 493.050 ;
        RECT 100.950 490.950 103.050 493.050 ;
        RECT 103.950 490.950 106.050 493.050 ;
        RECT 106.950 490.950 109.050 493.050 ;
        RECT 121.950 490.950 124.050 493.050 ;
        RECT 124.950 490.950 127.050 493.050 ;
        RECT 139.950 490.950 142.050 493.050 ;
        RECT 142.950 490.950 145.050 493.050 ;
        RECT 145.950 490.950 148.050 493.050 ;
        RECT 148.950 490.950 151.050 493.050 ;
        RECT 169.050 490.950 172.200 493.050 ;
        RECT 45.750 485.100 57.450 485.700 ;
        RECT 23.550 471.600 25.350 483.600 ;
        RECT 26.550 471.000 28.350 483.600 ;
        RECT 32.250 483.300 37.050 484.200 ;
        RECT 39.150 484.500 57.450 485.100 ;
        RECT 39.150 484.200 47.550 484.500 ;
        RECT 32.250 482.400 33.450 483.300 ;
        RECT 30.450 480.600 33.450 482.400 ;
        RECT 34.350 482.100 36.150 482.400 ;
        RECT 39.150 482.100 40.050 484.200 ;
        RECT 56.550 483.600 57.450 484.500 ;
        RECT 34.350 481.200 40.050 482.100 ;
        RECT 40.950 482.700 42.750 483.300 ;
        RECT 40.950 481.500 48.750 482.700 ;
        RECT 34.350 480.600 36.150 481.200 ;
        RECT 46.650 480.600 48.750 481.500 ;
        RECT 31.350 477.600 33.450 479.700 ;
        RECT 37.950 479.550 39.750 480.300 ;
        RECT 42.750 479.550 44.550 480.300 ;
        RECT 37.950 478.500 44.550 479.550 ;
        RECT 31.350 471.600 33.150 477.600 ;
        RECT 35.850 471.000 37.650 477.600 ;
        RECT 38.850 471.600 40.650 478.500 ;
        RECT 41.850 471.000 43.650 477.600 ;
        RECT 46.650 471.600 48.450 480.600 ;
        RECT 52.050 471.000 53.850 483.600 ;
        RECT 55.050 481.800 57.450 483.600 ;
        RECT 55.050 471.600 56.850 481.800 ;
        RECT 75.000 478.800 75.900 490.950 ;
        RECT 80.100 489.150 81.900 490.950 ;
        RECT 101.250 489.150 103.050 490.950 ;
        RECT 107.700 483.600 108.600 490.950 ;
        RECT 122.100 489.150 123.900 490.950 ;
        RECT 98.100 482.700 105.900 483.600 ;
        RECT 75.000 477.900 81.600 478.800 ;
        RECT 75.000 477.600 75.900 477.900 ;
        RECT 74.100 471.600 75.900 477.600 ;
        RECT 80.100 477.600 81.600 477.900 ;
        RECT 77.100 471.000 78.900 477.000 ;
        RECT 80.100 471.600 81.900 477.600 ;
        RECT 83.100 471.000 84.900 477.600 ;
        RECT 98.100 471.600 99.900 482.700 ;
        RECT 101.100 471.000 102.900 481.800 ;
        RECT 104.100 471.600 105.900 482.700 ;
        RECT 107.100 471.600 108.900 483.600 ;
        RECT 125.100 477.600 126.300 490.950 ;
        RECT 141.000 478.800 141.900 490.950 ;
        RECT 146.100 489.150 147.900 490.950 ;
        RECT 169.050 485.700 170.100 490.950 ;
        RECT 174.000 485.700 175.200 496.200 ;
        RECT 177.000 496.200 181.200 497.400 ;
        RECT 177.000 495.600 178.800 496.200 ;
        RECT 180.000 485.700 181.200 496.200 ;
        RECT 183.000 496.200 187.200 497.400 ;
        RECT 183.000 495.600 184.800 496.200 ;
        RECT 186.000 485.700 187.200 496.200 ;
        RECT 188.400 493.050 190.200 494.850 ;
        RECT 209.250 493.050 211.050 494.850 ;
        RECT 188.100 490.950 190.200 493.050 ;
        RECT 209.100 490.950 211.200 493.050 ;
        RECT 169.050 484.500 171.900 485.700 ;
        RECT 174.000 484.500 177.900 485.700 ;
        RECT 180.000 484.500 183.900 485.700 ;
        RECT 186.000 484.500 189.900 485.700 ;
        RECT 141.000 477.900 147.600 478.800 ;
        RECT 141.000 477.600 141.900 477.900 ;
        RECT 122.100 471.000 123.900 477.600 ;
        RECT 125.100 471.600 126.900 477.600 ;
        RECT 140.100 471.600 141.900 477.600 ;
        RECT 146.100 477.600 147.600 477.900 ;
        RECT 143.100 471.000 144.900 477.000 ;
        RECT 146.100 471.600 147.900 477.600 ;
        RECT 149.100 471.000 150.900 477.600 ;
        RECT 167.100 471.000 168.900 483.600 ;
        RECT 170.100 471.600 171.900 484.500 ;
        RECT 173.100 471.000 174.900 483.600 ;
        RECT 176.100 471.600 177.900 484.500 ;
        RECT 179.100 471.000 180.900 483.600 ;
        RECT 182.100 471.600 183.900 484.500 ;
        RECT 185.100 471.000 186.900 483.600 ;
        RECT 188.100 471.600 189.900 484.500 ;
        RECT 191.100 471.000 192.900 483.600 ;
        RECT 212.100 477.600 213.000 497.700 ;
        RECT 218.400 493.050 219.300 500.400 ;
        RECT 233.700 499.200 235.500 506.400 ;
        RECT 238.800 500.400 240.600 507.000 ;
        RECT 254.100 503.400 255.900 506.400 ;
        RECT 254.100 499.500 255.300 503.400 ;
        RECT 257.100 500.400 258.900 507.000 ;
        RECT 260.100 500.400 261.900 506.400 ;
        RECT 233.700 498.300 237.900 499.200 ;
        RECT 254.100 498.600 259.800 499.500 ;
        RECT 233.100 493.050 234.900 494.850 ;
        RECT 236.700 493.050 237.900 498.300 ;
        RECT 258.000 497.700 259.800 498.600 ;
        RECT 238.950 493.050 240.750 494.850 ;
        RECT 214.500 490.950 216.600 493.050 ;
        RECT 217.800 490.950 219.900 493.050 ;
        RECT 232.950 490.950 235.050 493.050 ;
        RECT 235.950 490.950 238.050 493.050 ;
        RECT 238.950 490.950 241.050 493.050 ;
        RECT 254.400 490.950 256.500 493.050 ;
        RECT 214.200 489.150 216.000 490.950 ;
        RECT 218.400 483.600 219.300 490.950 ;
        RECT 209.100 471.000 210.900 477.600 ;
        RECT 212.100 471.600 213.900 477.600 ;
        RECT 215.100 471.000 216.900 483.000 ;
        RECT 218.100 471.600 219.900 483.600 ;
        RECT 236.700 477.600 237.900 490.950 ;
        RECT 254.400 489.150 256.200 490.950 ;
        RECT 258.000 486.300 258.900 497.700 ;
        RECT 260.700 493.050 261.900 500.400 ;
        RECT 275.100 501.300 276.900 506.400 ;
        RECT 278.100 502.200 279.900 507.000 ;
        RECT 281.100 501.300 282.900 506.400 ;
        RECT 275.100 499.950 282.900 501.300 ;
        RECT 284.100 500.400 285.900 506.400 ;
        RECT 299.400 500.400 301.200 507.000 ;
        RECT 284.100 498.300 285.300 500.400 ;
        RECT 304.500 499.200 306.300 506.400 ;
        RECT 320.100 500.400 321.900 507.000 ;
        RECT 323.100 500.400 324.900 506.400 ;
        RECT 281.700 497.400 285.300 498.300 ;
        RECT 302.100 498.300 306.300 499.200 ;
        RECT 278.100 493.050 279.900 494.850 ;
        RECT 281.700 493.050 282.900 497.400 ;
        RECT 284.100 493.050 285.900 494.850 ;
        RECT 299.250 493.050 301.050 494.850 ;
        RECT 302.100 493.050 303.300 498.300 ;
        RECT 305.100 493.050 306.900 494.850 ;
        RECT 320.100 493.050 321.900 494.850 ;
        RECT 323.100 493.050 324.300 500.400 ;
        RECT 338.700 499.200 340.500 506.400 ;
        RECT 343.800 500.400 345.600 507.000 ;
        RECT 359.400 500.400 361.200 507.000 ;
        RECT 364.500 499.200 366.300 506.400 ;
        RECT 383.700 500.400 385.500 507.000 ;
        RECT 388.200 500.400 390.000 506.400 ;
        RECT 392.700 500.400 394.500 507.000 ;
        RECT 410.100 503.400 411.900 507.000 ;
        RECT 413.100 503.400 414.900 506.400 ;
        RECT 338.700 498.300 342.900 499.200 ;
        RECT 338.100 493.050 339.900 494.850 ;
        RECT 341.700 493.050 342.900 498.300 ;
        RECT 362.100 498.300 366.300 499.200 ;
        RECT 343.950 493.050 345.750 494.850 ;
        RECT 359.250 493.050 361.050 494.850 ;
        RECT 362.100 493.050 363.300 498.300 ;
        RECT 367.950 495.450 370.050 496.050 ;
        RECT 376.950 495.450 379.050 496.050 ;
        RECT 365.100 493.050 366.900 494.850 ;
        RECT 367.950 494.550 379.050 495.450 ;
        RECT 367.950 493.950 370.050 494.550 ;
        RECT 376.950 493.950 379.050 494.550 ;
        RECT 383.250 493.050 385.050 494.850 ;
        RECT 389.100 493.050 390.300 500.400 ;
        RECT 395.100 493.050 396.900 494.850 ;
        RECT 413.100 493.050 414.300 503.400 ;
        RECT 428.100 497.400 429.900 507.000 ;
        RECT 434.700 498.000 436.500 506.400 ;
        RECT 455.100 501.300 456.900 506.400 ;
        RECT 458.100 502.200 459.900 507.000 ;
        RECT 461.100 501.300 462.900 506.400 ;
        RECT 455.100 499.950 462.900 501.300 ;
        RECT 464.100 500.400 465.900 506.400 ;
        RECT 464.100 498.300 465.300 500.400 ;
        RECT 434.700 496.800 438.000 498.000 ;
        RECT 428.100 493.050 429.900 494.850 ;
        RECT 434.100 493.050 435.900 494.850 ;
        RECT 437.100 493.050 438.000 496.800 ;
        RECT 461.700 497.400 465.300 498.300 ;
        RECT 482.100 498.600 483.900 506.400 ;
        RECT 486.600 500.400 488.400 507.000 ;
        RECT 489.600 502.200 491.400 506.400 ;
        RECT 489.600 500.400 492.300 502.200 ;
        RECT 488.700 498.600 490.500 499.500 ;
        RECT 482.100 497.700 490.500 498.600 ;
        RECT 458.100 493.050 459.900 494.850 ;
        RECT 461.700 493.050 462.900 497.400 ;
        RECT 464.100 493.050 465.900 494.850 ;
        RECT 482.250 493.050 484.050 494.850 ;
        RECT 259.800 490.950 261.900 493.050 ;
        RECT 274.950 490.950 277.050 493.050 ;
        RECT 277.950 490.950 280.050 493.050 ;
        RECT 280.950 490.950 283.050 493.050 ;
        RECT 283.950 490.950 286.050 493.050 ;
        RECT 298.950 490.950 301.050 493.050 ;
        RECT 301.950 490.950 304.050 493.050 ;
        RECT 304.950 490.950 307.050 493.050 ;
        RECT 319.950 490.950 322.050 493.050 ;
        RECT 322.950 490.950 325.050 493.050 ;
        RECT 337.950 490.950 340.050 493.050 ;
        RECT 340.950 490.950 343.050 493.050 ;
        RECT 343.950 490.950 346.050 493.050 ;
        RECT 358.950 490.950 361.050 493.050 ;
        RECT 361.950 490.950 364.050 493.050 ;
        RECT 364.950 490.950 367.050 493.050 ;
        RECT 382.950 490.950 385.050 493.050 ;
        RECT 385.950 490.950 388.050 493.050 ;
        RECT 388.950 490.950 391.050 493.050 ;
        RECT 391.950 490.950 394.050 493.050 ;
        RECT 394.950 490.950 397.050 493.050 ;
        RECT 409.950 490.950 412.050 493.050 ;
        RECT 412.950 490.950 415.050 493.050 ;
        RECT 427.950 490.950 430.050 493.050 ;
        RECT 430.950 490.950 433.050 493.050 ;
        RECT 433.950 490.950 436.050 493.050 ;
        RECT 436.950 490.950 439.050 493.050 ;
        RECT 454.950 490.950 457.050 493.050 ;
        RECT 457.950 490.950 460.050 493.050 ;
        RECT 460.950 490.950 463.050 493.050 ;
        RECT 463.950 490.950 466.050 493.050 ;
        RECT 482.100 490.950 484.200 493.050 ;
        RECT 258.000 485.400 259.800 486.300 ;
        RECT 254.100 484.500 259.800 485.400 ;
        RECT 254.100 477.600 255.300 484.500 ;
        RECT 260.700 483.600 261.900 490.950 ;
        RECT 275.100 489.150 276.900 490.950 ;
        RECT 281.700 483.600 282.900 490.950 ;
        RECT 233.100 471.000 234.900 477.600 ;
        RECT 236.100 471.600 237.900 477.600 ;
        RECT 239.100 471.000 240.900 477.600 ;
        RECT 254.100 471.600 255.900 477.600 ;
        RECT 257.100 471.000 258.900 481.800 ;
        RECT 260.100 471.600 261.900 483.600 ;
        RECT 275.400 471.000 277.200 483.600 ;
        RECT 280.500 482.100 282.900 483.600 ;
        RECT 280.500 471.600 282.300 482.100 ;
        RECT 283.200 479.100 285.000 480.900 ;
        RECT 302.100 477.600 303.300 490.950 ;
        RECT 323.100 483.600 324.300 490.950 ;
        RECT 283.500 471.000 285.300 477.600 ;
        RECT 299.100 471.000 300.900 477.600 ;
        RECT 302.100 471.600 303.900 477.600 ;
        RECT 305.100 471.000 306.900 477.600 ;
        RECT 320.100 471.000 321.900 483.600 ;
        RECT 323.100 471.600 324.900 483.600 ;
        RECT 341.700 477.600 342.900 490.950 ;
        RECT 362.100 477.600 363.300 490.950 ;
        RECT 386.250 489.150 388.050 490.950 ;
        RECT 389.100 485.400 390.000 490.950 ;
        RECT 392.100 489.150 393.900 490.950 ;
        RECT 410.100 489.150 411.900 490.950 ;
        RECT 389.100 484.500 393.900 485.400 ;
        RECT 383.100 482.400 390.900 483.300 ;
        RECT 338.100 471.000 339.900 477.600 ;
        RECT 341.100 471.600 342.900 477.600 ;
        RECT 344.100 471.000 345.900 477.600 ;
        RECT 359.100 471.000 360.900 477.600 ;
        RECT 362.100 471.600 363.900 477.600 ;
        RECT 365.100 471.000 366.900 477.600 ;
        RECT 383.100 471.600 384.900 482.400 ;
        RECT 386.100 471.000 387.900 481.500 ;
        RECT 389.100 472.500 390.900 482.400 ;
        RECT 392.100 473.400 393.900 484.500 ;
        RECT 395.100 472.500 396.900 483.600 ;
        RECT 413.100 477.600 414.300 490.950 ;
        RECT 431.100 489.150 432.900 490.950 ;
        RECT 437.100 478.800 438.000 490.950 ;
        RECT 455.100 489.150 456.900 490.950 ;
        RECT 461.700 483.600 462.900 490.950 ;
        RECT 431.400 477.900 438.000 478.800 ;
        RECT 431.400 477.600 432.900 477.900 ;
        RECT 389.100 471.600 396.900 472.500 ;
        RECT 410.100 471.000 411.900 477.600 ;
        RECT 413.100 471.600 414.900 477.600 ;
        RECT 428.100 471.000 429.900 477.600 ;
        RECT 431.100 471.600 432.900 477.600 ;
        RECT 437.100 477.600 438.000 477.900 ;
        RECT 434.100 471.000 435.900 477.000 ;
        RECT 437.100 471.600 438.900 477.600 ;
        RECT 455.400 471.000 457.200 483.600 ;
        RECT 460.500 482.100 462.900 483.600 ;
        RECT 460.500 471.600 462.300 482.100 ;
        RECT 463.200 479.100 465.000 480.900 ;
        RECT 485.100 477.600 486.000 497.700 ;
        RECT 491.400 493.050 492.300 500.400 ;
        RECT 509.100 498.600 510.900 506.400 ;
        RECT 513.600 500.400 515.400 507.000 ;
        RECT 516.600 502.200 518.400 506.400 ;
        RECT 516.600 500.400 519.300 502.200 ;
        RECT 533.700 500.400 535.500 507.000 ;
        RECT 538.200 500.400 540.000 506.400 ;
        RECT 542.700 500.400 544.500 507.000 ;
        RECT 560.100 501.300 561.900 506.400 ;
        RECT 563.100 502.200 564.900 507.000 ;
        RECT 566.100 501.300 567.900 506.400 ;
        RECT 515.700 498.600 517.500 499.500 ;
        RECT 509.100 497.700 517.500 498.600 ;
        RECT 509.250 493.050 511.050 494.850 ;
        RECT 487.500 490.950 489.600 493.050 ;
        RECT 490.800 490.950 492.900 493.050 ;
        RECT 509.100 490.950 511.200 493.050 ;
        RECT 487.200 489.150 489.000 490.950 ;
        RECT 491.400 483.600 492.300 490.950 ;
        RECT 463.500 471.000 465.300 477.600 ;
        RECT 482.100 471.000 483.900 477.600 ;
        RECT 485.100 471.600 486.900 477.600 ;
        RECT 488.100 471.000 489.900 483.000 ;
        RECT 491.100 471.600 492.900 483.600 ;
        RECT 512.100 477.600 513.000 497.700 ;
        RECT 518.400 493.050 519.300 500.400 ;
        RECT 528.000 495.450 532.050 496.050 ;
        RECT 527.550 493.950 532.050 495.450 ;
        RECT 514.500 490.950 516.600 493.050 ;
        RECT 517.800 490.950 519.900 493.050 ;
        RECT 514.200 489.150 516.000 490.950 ;
        RECT 518.400 483.600 519.300 490.950 ;
        RECT 527.550 490.050 528.450 493.950 ;
        RECT 533.250 493.050 535.050 494.850 ;
        RECT 539.100 493.050 540.300 500.400 ;
        RECT 560.100 499.950 567.900 501.300 ;
        RECT 569.100 500.400 570.900 506.400 ;
        RECT 584.100 503.400 585.900 507.000 ;
        RECT 587.100 503.400 588.900 506.400 ;
        RECT 569.100 498.300 570.300 500.400 ;
        RECT 566.700 497.400 570.300 498.300 ;
        RECT 545.100 493.050 546.900 494.850 ;
        RECT 563.100 493.050 564.900 494.850 ;
        RECT 566.700 493.050 567.900 497.400 ;
        RECT 569.100 493.050 570.900 494.850 ;
        RECT 587.100 493.050 588.300 503.400 ;
        RECT 605.100 497.400 606.900 507.000 ;
        RECT 611.700 498.000 613.500 506.400 ;
        RECT 611.700 496.800 615.000 498.000 ;
        RECT 629.100 497.400 630.900 507.000 ;
        RECT 635.700 498.000 637.500 506.400 ;
        RECT 653.400 500.400 655.200 507.000 ;
        RECT 658.500 499.200 660.300 506.400 ;
        RECT 675.600 502.200 677.400 506.400 ;
        RECT 656.100 498.300 660.300 499.200 ;
        RECT 674.700 500.400 677.400 502.200 ;
        RECT 678.600 500.400 680.400 507.000 ;
        RECT 635.700 496.800 639.000 498.000 ;
        RECT 605.100 493.050 606.900 494.850 ;
        RECT 611.100 493.050 612.900 494.850 ;
        RECT 614.100 493.050 615.000 496.800 ;
        RECT 629.100 493.050 630.900 494.850 ;
        RECT 635.100 493.050 636.900 494.850 ;
        RECT 638.100 493.050 639.000 496.800 ;
        RECT 648.000 495.450 652.050 496.050 ;
        RECT 647.550 493.950 652.050 495.450 ;
        RECT 532.950 490.950 535.050 493.050 ;
        RECT 535.950 490.950 538.050 493.050 ;
        RECT 538.950 490.950 541.050 493.050 ;
        RECT 541.950 490.950 544.050 493.050 ;
        RECT 544.950 490.950 547.050 493.050 ;
        RECT 559.950 490.950 562.050 493.050 ;
        RECT 562.950 490.950 565.050 493.050 ;
        RECT 565.950 490.950 568.050 493.050 ;
        RECT 568.950 490.950 571.050 493.050 ;
        RECT 583.950 490.950 586.050 493.050 ;
        RECT 586.950 490.950 589.050 493.050 ;
        RECT 604.950 490.950 607.050 493.050 ;
        RECT 607.950 490.950 610.050 493.050 ;
        RECT 610.950 490.950 613.050 493.050 ;
        RECT 613.950 490.950 616.050 493.050 ;
        RECT 628.950 490.950 631.050 493.050 ;
        RECT 631.950 490.950 634.050 493.050 ;
        RECT 634.950 490.950 637.050 493.050 ;
        RECT 637.950 490.950 640.050 493.050 ;
        RECT 527.550 488.550 532.050 490.050 ;
        RECT 536.250 489.150 538.050 490.950 ;
        RECT 528.000 487.950 532.050 488.550 ;
        RECT 539.100 485.400 540.000 490.950 ;
        RECT 542.100 489.150 543.900 490.950 ;
        RECT 560.100 489.150 561.900 490.950 ;
        RECT 547.950 486.450 550.050 487.050 ;
        RECT 559.950 486.450 562.050 487.050 ;
        RECT 547.950 485.550 562.050 486.450 ;
        RECT 539.100 484.500 543.900 485.400 ;
        RECT 547.950 484.950 550.050 485.550 ;
        RECT 559.950 484.950 562.050 485.550 ;
        RECT 509.100 471.000 510.900 477.600 ;
        RECT 512.100 471.600 513.900 477.600 ;
        RECT 515.100 471.000 516.900 483.000 ;
        RECT 518.100 471.600 519.900 483.600 ;
        RECT 533.100 482.400 540.900 483.300 ;
        RECT 533.100 471.600 534.900 482.400 ;
        RECT 536.100 471.000 537.900 481.500 ;
        RECT 539.100 472.500 540.900 482.400 ;
        RECT 542.100 473.400 543.900 484.500 ;
        RECT 566.700 483.600 567.900 490.950 ;
        RECT 584.100 489.150 585.900 490.950 ;
        RECT 545.100 472.500 546.900 483.600 ;
        RECT 539.100 471.600 546.900 472.500 ;
        RECT 560.400 471.000 562.200 483.600 ;
        RECT 565.500 482.100 567.900 483.600 ;
        RECT 565.500 471.600 567.300 482.100 ;
        RECT 568.200 479.100 570.000 480.900 ;
        RECT 587.100 477.600 588.300 490.950 ;
        RECT 608.100 489.150 609.900 490.950 ;
        RECT 598.950 486.450 601.050 487.050 ;
        RECT 604.950 486.450 607.050 487.050 ;
        RECT 598.950 485.550 607.050 486.450 ;
        RECT 598.950 484.950 601.050 485.550 ;
        RECT 604.950 484.950 607.050 485.550 ;
        RECT 614.100 478.800 615.000 490.950 ;
        RECT 632.100 489.150 633.900 490.950 ;
        RECT 638.100 478.800 639.000 490.950 ;
        RECT 647.550 490.050 648.450 493.950 ;
        RECT 653.250 493.050 655.050 494.850 ;
        RECT 656.100 493.050 657.300 498.300 ;
        RECT 659.100 493.050 660.900 494.850 ;
        RECT 674.700 493.050 675.600 500.400 ;
        RECT 676.500 498.600 678.300 499.500 ;
        RECT 683.100 498.600 684.900 506.400 ;
        RECT 698.700 503.400 700.500 507.000 ;
        RECT 701.700 501.600 703.500 506.400 ;
        RECT 676.500 497.700 684.900 498.600 ;
        RECT 698.400 500.400 703.500 501.600 ;
        RECT 706.200 500.400 708.000 507.000 ;
        RECT 725.100 503.400 726.900 506.400 ;
        RECT 728.100 503.400 729.900 507.000 ;
        RECT 652.950 490.950 655.050 493.050 ;
        RECT 655.950 490.950 658.050 493.050 ;
        RECT 658.950 490.950 661.050 493.050 ;
        RECT 674.100 490.950 676.200 493.050 ;
        RECT 677.400 490.950 679.500 493.050 ;
        RECT 647.550 488.550 652.050 490.050 ;
        RECT 648.000 487.950 652.050 488.550 ;
        RECT 608.400 477.900 615.000 478.800 ;
        RECT 608.400 477.600 609.900 477.900 ;
        RECT 568.500 471.000 570.300 477.600 ;
        RECT 584.100 471.000 585.900 477.600 ;
        RECT 587.100 471.600 588.900 477.600 ;
        RECT 605.100 471.000 606.900 477.600 ;
        RECT 608.100 471.600 609.900 477.600 ;
        RECT 614.100 477.600 615.000 477.900 ;
        RECT 632.400 477.900 639.000 478.800 ;
        RECT 632.400 477.600 633.900 477.900 ;
        RECT 611.100 471.000 612.900 477.000 ;
        RECT 614.100 471.600 615.900 477.600 ;
        RECT 629.100 471.000 630.900 477.600 ;
        RECT 632.100 471.600 633.900 477.600 ;
        RECT 638.100 477.600 639.000 477.900 ;
        RECT 656.100 477.600 657.300 490.950 ;
        RECT 674.700 483.600 675.600 490.950 ;
        RECT 678.000 489.150 679.800 490.950 ;
        RECT 635.100 471.000 636.900 477.000 ;
        RECT 638.100 471.600 639.900 477.600 ;
        RECT 653.100 471.000 654.900 477.600 ;
        RECT 656.100 471.600 657.900 477.600 ;
        RECT 659.100 471.000 660.900 477.600 ;
        RECT 674.100 471.600 675.900 483.600 ;
        RECT 677.100 471.000 678.900 483.000 ;
        RECT 681.000 477.600 681.900 497.700 ;
        RECT 688.950 495.450 691.050 496.050 ;
        RECT 694.950 495.450 697.050 496.050 ;
        RECT 682.950 493.050 684.750 494.850 ;
        RECT 688.950 494.550 697.050 495.450 ;
        RECT 688.950 493.950 691.050 494.550 ;
        RECT 694.950 493.950 697.050 494.550 ;
        RECT 698.400 493.050 699.300 500.400 ;
        RECT 700.950 498.450 703.050 499.050 ;
        RECT 721.950 498.450 724.050 499.050 ;
        RECT 700.950 497.550 724.050 498.450 ;
        RECT 700.950 496.950 703.050 497.550 ;
        RECT 721.950 496.950 724.050 497.550 ;
        RECT 700.950 493.050 702.750 494.850 ;
        RECT 707.100 493.050 708.900 494.850 ;
        RECT 725.700 493.050 726.900 503.400 ;
        RECT 744.600 502.200 746.400 506.400 ;
        RECT 743.700 500.400 746.400 502.200 ;
        RECT 747.600 500.400 749.400 507.000 ;
        RECT 743.700 493.050 744.600 500.400 ;
        RECT 745.500 498.600 747.300 499.500 ;
        RECT 752.100 498.600 753.900 506.400 ;
        RECT 745.500 497.700 753.900 498.600 ;
        RECT 682.800 490.950 684.900 493.050 ;
        RECT 697.950 490.950 700.050 493.050 ;
        RECT 700.950 490.950 703.050 493.050 ;
        RECT 703.950 490.950 706.050 493.050 ;
        RECT 706.950 490.950 709.050 493.050 ;
        RECT 724.950 490.950 727.050 493.050 ;
        RECT 727.950 490.950 730.050 493.050 ;
        RECT 743.100 490.950 745.200 493.050 ;
        RECT 746.400 490.950 748.500 493.050 ;
        RECT 688.950 483.450 691.050 484.050 ;
        RECT 694.950 483.450 697.050 484.050 ;
        RECT 698.400 483.600 699.300 490.950 ;
        RECT 703.950 489.150 705.750 490.950 ;
        RECT 700.950 486.450 703.050 487.050 ;
        RECT 721.950 486.450 724.050 487.050 ;
        RECT 700.950 485.550 724.050 486.450 ;
        RECT 700.950 484.950 703.050 485.550 ;
        RECT 721.950 484.950 724.050 485.550 ;
        RECT 688.950 482.550 697.050 483.450 ;
        RECT 688.950 481.950 691.050 482.550 ;
        RECT 694.950 481.950 697.050 482.550 ;
        RECT 680.100 471.600 681.900 477.600 ;
        RECT 683.100 471.000 684.900 477.600 ;
        RECT 698.100 471.600 699.900 483.600 ;
        RECT 701.100 482.700 708.900 483.600 ;
        RECT 701.100 471.600 702.900 482.700 ;
        RECT 704.100 471.000 705.900 481.800 ;
        RECT 707.100 471.600 708.900 482.700 ;
        RECT 725.700 477.600 726.900 490.950 ;
        RECT 728.100 489.150 729.900 490.950 ;
        RECT 743.700 483.600 744.600 490.950 ;
        RECT 747.000 489.150 748.800 490.950 ;
        RECT 725.100 471.600 726.900 477.600 ;
        RECT 728.100 471.000 729.900 477.600 ;
        RECT 743.100 471.600 744.900 483.600 ;
        RECT 746.100 471.000 747.900 483.000 ;
        RECT 750.000 477.600 750.900 497.700 ;
        RECT 767.100 497.400 768.900 507.000 ;
        RECT 773.700 498.000 775.500 506.400 ;
        RECT 794.400 500.400 796.200 507.000 ;
        RECT 799.500 499.200 801.300 506.400 ;
        RECT 815.700 500.400 817.500 507.000 ;
        RECT 820.200 500.400 822.000 506.400 ;
        RECT 824.700 500.400 826.500 507.000 ;
        RECT 797.100 498.300 801.300 499.200 ;
        RECT 773.700 496.800 777.000 498.000 ;
        RECT 751.950 493.050 753.750 494.850 ;
        RECT 767.100 493.050 768.900 494.850 ;
        RECT 773.100 493.050 774.900 494.850 ;
        RECT 776.100 493.050 777.000 496.800 ;
        RECT 794.250 493.050 796.050 494.850 ;
        RECT 797.100 493.050 798.300 498.300 ;
        RECT 800.100 493.050 801.900 494.850 ;
        RECT 815.250 493.050 817.050 494.850 ;
        RECT 821.100 493.050 822.300 500.400 ;
        RECT 842.100 497.400 843.900 507.000 ;
        RECT 848.700 498.000 850.500 506.400 ;
        RECT 866.100 503.400 867.900 507.000 ;
        RECT 869.100 503.400 870.900 506.400 ;
        RECT 848.700 496.800 852.000 498.000 ;
        RECT 827.100 493.050 828.900 494.850 ;
        RECT 842.100 493.050 843.900 494.850 ;
        RECT 848.100 493.050 849.900 494.850 ;
        RECT 851.100 493.050 852.000 496.800 ;
        RECT 869.100 493.050 870.300 503.400 ;
        RECT 884.100 500.400 885.900 506.400 ;
        RECT 884.700 498.300 885.900 500.400 ;
        RECT 887.100 501.300 888.900 506.400 ;
        RECT 890.100 502.200 891.900 507.000 ;
        RECT 893.100 501.300 894.900 506.400 ;
        RECT 887.100 499.950 894.900 501.300 ;
        RECT 884.700 497.400 888.300 498.300 ;
        RECT 884.100 493.050 885.900 494.850 ;
        RECT 887.100 493.050 888.300 497.400 ;
        RECT 890.100 493.050 891.900 494.850 ;
        RECT 751.800 490.950 753.900 493.050 ;
        RECT 766.950 490.950 769.050 493.050 ;
        RECT 769.950 490.950 772.050 493.050 ;
        RECT 772.950 490.950 775.050 493.050 ;
        RECT 775.950 490.950 778.050 493.050 ;
        RECT 793.950 490.950 796.050 493.050 ;
        RECT 796.950 490.950 799.050 493.050 ;
        RECT 799.950 490.950 802.050 493.050 ;
        RECT 814.950 490.950 817.050 493.050 ;
        RECT 817.950 490.950 820.050 493.050 ;
        RECT 820.950 490.950 823.050 493.050 ;
        RECT 823.950 490.950 826.050 493.050 ;
        RECT 826.950 490.950 829.050 493.050 ;
        RECT 841.950 490.950 844.050 493.050 ;
        RECT 844.950 490.950 847.050 493.050 ;
        RECT 847.950 490.950 850.050 493.050 ;
        RECT 850.950 490.950 853.050 493.050 ;
        RECT 865.950 490.950 868.050 493.050 ;
        RECT 868.950 490.950 871.050 493.050 ;
        RECT 883.950 490.950 886.050 493.050 ;
        RECT 886.950 490.950 889.050 493.050 ;
        RECT 889.950 490.950 892.050 493.050 ;
        RECT 892.950 490.950 895.050 493.050 ;
        RECT 770.100 489.150 771.900 490.950 ;
        RECT 776.100 478.800 777.000 490.950 ;
        RECT 770.400 477.900 777.000 478.800 ;
        RECT 770.400 477.600 771.900 477.900 ;
        RECT 749.100 471.600 750.900 477.600 ;
        RECT 752.100 471.000 753.900 477.600 ;
        RECT 767.100 471.000 768.900 477.600 ;
        RECT 770.100 471.600 771.900 477.600 ;
        RECT 776.100 477.600 777.000 477.900 ;
        RECT 797.100 477.600 798.300 490.950 ;
        RECT 818.250 489.150 820.050 490.950 ;
        RECT 799.950 486.450 802.050 487.050 ;
        RECT 808.950 486.450 811.050 487.050 ;
        RECT 799.950 485.550 811.050 486.450 ;
        RECT 799.950 484.950 802.050 485.550 ;
        RECT 808.950 484.950 811.050 485.550 ;
        RECT 821.100 485.400 822.000 490.950 ;
        RECT 824.100 489.150 825.900 490.950 ;
        RECT 845.100 489.150 846.900 490.950 ;
        RECT 821.100 484.500 825.900 485.400 ;
        RECT 815.100 482.400 822.900 483.300 ;
        RECT 773.100 471.000 774.900 477.000 ;
        RECT 776.100 471.600 777.900 477.600 ;
        RECT 794.100 471.000 795.900 477.600 ;
        RECT 797.100 471.600 798.900 477.600 ;
        RECT 800.100 471.000 801.900 477.600 ;
        RECT 815.100 471.600 816.900 482.400 ;
        RECT 818.100 471.000 819.900 481.500 ;
        RECT 821.100 472.500 822.900 482.400 ;
        RECT 824.100 473.400 825.900 484.500 ;
        RECT 827.100 472.500 828.900 483.600 ;
        RECT 851.100 478.800 852.000 490.950 ;
        RECT 866.100 489.150 867.900 490.950 ;
        RECT 845.400 477.900 852.000 478.800 ;
        RECT 845.400 477.600 846.900 477.900 ;
        RECT 821.100 471.600 828.900 472.500 ;
        RECT 842.100 471.000 843.900 477.600 ;
        RECT 845.100 471.600 846.900 477.600 ;
        RECT 851.100 477.600 852.000 477.900 ;
        RECT 869.100 477.600 870.300 490.950 ;
        RECT 887.100 483.600 888.300 490.950 ;
        RECT 893.100 489.150 894.900 490.950 ;
        RECT 887.100 482.100 889.500 483.600 ;
        RECT 885.000 479.100 886.800 480.900 ;
        RECT 848.100 471.000 849.900 477.000 ;
        RECT 851.100 471.600 852.900 477.600 ;
        RECT 866.100 471.000 867.900 477.600 ;
        RECT 869.100 471.600 870.900 477.600 ;
        RECT 884.700 471.000 886.500 477.600 ;
        RECT 887.700 471.600 889.500 482.100 ;
        RECT 892.800 471.000 894.600 483.600 ;
        RECT 17.100 455.400 18.900 467.400 ;
        RECT 20.100 457.200 21.900 468.000 ;
        RECT 23.100 461.400 24.900 467.400 ;
        RECT 17.100 448.050 18.300 455.400 ;
        RECT 23.700 454.500 24.900 461.400 ;
        RECT 19.200 453.600 24.900 454.500 ;
        RECT 26.550 455.400 28.350 467.400 ;
        RECT 29.550 455.400 31.350 468.000 ;
        RECT 34.350 461.400 36.150 467.400 ;
        RECT 38.850 461.400 40.650 468.000 ;
        RECT 34.350 459.300 36.450 461.400 ;
        RECT 41.850 460.500 43.650 467.400 ;
        RECT 44.850 461.400 46.650 468.000 ;
        RECT 40.950 459.450 47.550 460.500 ;
        RECT 40.950 458.700 42.750 459.450 ;
        RECT 45.750 458.700 47.550 459.450 ;
        RECT 49.650 458.400 51.450 467.400 ;
        RECT 33.450 456.600 36.450 458.400 ;
        RECT 37.350 457.800 39.150 458.400 ;
        RECT 37.350 456.900 43.050 457.800 ;
        RECT 49.650 457.500 51.750 458.400 ;
        RECT 37.350 456.600 39.150 456.900 ;
        RECT 35.250 455.700 36.450 456.600 ;
        RECT 19.200 452.700 21.000 453.600 ;
        RECT 17.100 445.950 19.200 448.050 ;
        RECT 17.100 438.600 18.300 445.950 ;
        RECT 20.100 441.300 21.000 452.700 ;
        RECT 22.800 448.050 24.600 449.850 ;
        RECT 22.500 445.950 24.600 448.050 ;
        RECT 26.550 448.050 27.750 455.400 ;
        RECT 35.250 454.800 40.050 455.700 ;
        RECT 28.650 452.100 30.450 452.550 ;
        RECT 34.350 452.100 36.450 452.700 ;
        RECT 28.650 450.900 36.450 452.100 ;
        RECT 28.650 450.750 30.450 450.900 ;
        RECT 34.350 450.600 36.450 450.900 ;
        RECT 26.550 447.750 31.050 448.050 ;
        RECT 26.550 445.950 32.850 447.750 ;
        RECT 19.200 440.400 21.000 441.300 ;
        RECT 19.200 439.500 24.900 440.400 ;
        RECT 17.100 432.600 18.900 438.600 ;
        RECT 20.100 432.000 21.900 438.600 ;
        RECT 23.700 435.600 24.900 439.500 ;
        RECT 23.100 432.600 24.900 435.600 ;
        RECT 26.550 438.600 27.750 445.950 ;
        RECT 39.150 442.200 40.050 454.800 ;
        RECT 42.150 454.800 43.050 456.900 ;
        RECT 43.950 456.300 51.750 457.500 ;
        RECT 43.950 455.700 45.750 456.300 ;
        RECT 55.050 455.400 56.850 468.000 ;
        RECT 58.050 457.200 59.850 467.400 ;
        RECT 58.050 455.400 60.450 457.200 ;
        RECT 42.150 454.500 50.550 454.800 ;
        RECT 59.550 454.500 60.450 455.400 ;
        RECT 42.150 453.900 60.450 454.500 ;
        RECT 48.750 453.300 60.450 453.900 ;
        RECT 48.750 453.000 50.550 453.300 ;
        RECT 46.800 446.400 48.900 448.050 ;
        RECT 46.800 445.200 54.900 446.400 ;
        RECT 55.950 445.950 58.050 448.050 ;
        RECT 53.100 444.600 54.900 445.200 ;
        RECT 50.100 443.400 51.900 444.000 ;
        RECT 56.250 443.400 58.050 445.950 ;
        RECT 50.100 442.200 58.050 443.400 ;
        RECT 39.150 441.000 51.150 442.200 ;
        RECT 39.150 440.400 40.950 441.000 ;
        RECT 50.100 439.200 51.150 441.000 ;
        RECT 26.550 432.600 28.350 438.600 ;
        RECT 29.850 432.000 31.650 438.600 ;
        RECT 34.350 435.600 36.750 437.700 ;
        RECT 46.350 437.550 48.150 438.300 ;
        RECT 43.200 436.500 48.150 437.550 ;
        RECT 49.350 437.400 51.150 439.200 ;
        RECT 59.550 438.600 60.450 453.300 ;
        RECT 43.200 435.600 44.250 436.500 ;
        RECT 52.050 436.200 54.150 437.700 ;
        RECT 50.250 435.600 54.150 436.200 ;
        RECT 34.950 432.600 36.750 435.600 ;
        RECT 39.450 432.000 41.250 435.600 ;
        RECT 42.450 432.600 44.250 435.600 ;
        RECT 45.750 432.000 47.550 435.600 ;
        RECT 50.250 434.700 53.850 435.600 ;
        RECT 50.250 432.600 52.050 434.700 ;
        RECT 55.050 432.000 56.850 438.600 ;
        RECT 58.050 436.800 60.450 438.600 ;
        RECT 62.550 455.400 64.350 467.400 ;
        RECT 65.550 455.400 67.350 468.000 ;
        RECT 70.350 461.400 72.150 467.400 ;
        RECT 74.850 461.400 76.650 468.000 ;
        RECT 70.350 459.300 72.450 461.400 ;
        RECT 77.850 460.500 79.650 467.400 ;
        RECT 80.850 461.400 82.650 468.000 ;
        RECT 76.950 459.450 83.550 460.500 ;
        RECT 76.950 458.700 78.750 459.450 ;
        RECT 81.750 458.700 83.550 459.450 ;
        RECT 85.650 458.400 87.450 467.400 ;
        RECT 69.450 456.600 72.450 458.400 ;
        RECT 73.350 457.800 75.150 458.400 ;
        RECT 73.350 456.900 79.050 457.800 ;
        RECT 85.650 457.500 87.750 458.400 ;
        RECT 73.350 456.600 75.150 456.900 ;
        RECT 71.250 455.700 72.450 456.600 ;
        RECT 62.550 448.050 63.750 455.400 ;
        RECT 71.250 454.800 76.050 455.700 ;
        RECT 64.650 452.100 66.450 452.550 ;
        RECT 70.350 452.100 72.450 452.700 ;
        RECT 64.650 450.900 72.450 452.100 ;
        RECT 64.650 450.750 66.450 450.900 ;
        RECT 70.350 450.600 72.450 450.900 ;
        RECT 62.550 447.750 67.050 448.050 ;
        RECT 62.550 445.950 68.850 447.750 ;
        RECT 62.550 438.600 63.750 445.950 ;
        RECT 75.150 442.200 76.050 454.800 ;
        RECT 78.150 454.800 79.050 456.900 ;
        RECT 79.950 456.300 87.750 457.500 ;
        RECT 79.950 455.700 81.750 456.300 ;
        RECT 91.050 455.400 92.850 468.000 ;
        RECT 94.050 457.200 95.850 467.400 ;
        RECT 113.100 461.400 114.900 468.000 ;
        RECT 116.100 461.400 117.900 467.400 ;
        RECT 94.050 455.400 96.450 457.200 ;
        RECT 78.150 454.500 86.550 454.800 ;
        RECT 95.550 454.500 96.450 455.400 ;
        RECT 78.150 453.900 96.450 454.500 ;
        RECT 84.750 453.300 96.450 453.900 ;
        RECT 84.750 453.000 86.550 453.300 ;
        RECT 82.800 446.400 84.900 448.050 ;
        RECT 82.800 445.200 90.900 446.400 ;
        RECT 91.950 445.950 94.050 448.050 ;
        RECT 89.100 444.600 90.900 445.200 ;
        RECT 86.100 443.400 87.900 444.000 ;
        RECT 92.250 443.400 94.050 445.950 ;
        RECT 86.100 442.200 94.050 443.400 ;
        RECT 75.150 441.000 87.150 442.200 ;
        RECT 75.150 440.400 76.950 441.000 ;
        RECT 86.100 439.200 87.150 441.000 ;
        RECT 58.050 432.600 59.850 436.800 ;
        RECT 62.550 432.600 64.350 438.600 ;
        RECT 65.850 432.000 67.650 438.600 ;
        RECT 70.350 435.600 72.750 437.700 ;
        RECT 82.350 437.550 84.150 438.300 ;
        RECT 79.200 436.500 84.150 437.550 ;
        RECT 85.350 437.400 87.150 439.200 ;
        RECT 95.550 438.600 96.450 453.300 ;
        RECT 113.100 448.050 114.900 449.850 ;
        RECT 116.100 448.050 117.300 461.400 ;
        RECT 131.400 455.400 133.200 468.000 ;
        RECT 136.500 456.900 138.300 467.400 ;
        RECT 139.500 461.400 141.300 468.000 ;
        RECT 155.700 461.400 157.500 468.000 ;
        RECT 139.200 458.100 141.000 459.900 ;
        RECT 156.000 458.100 157.800 459.900 ;
        RECT 158.700 456.900 160.500 467.400 ;
        RECT 136.500 455.400 138.900 456.900 ;
        RECT 131.100 448.050 132.900 449.850 ;
        RECT 137.700 448.050 138.900 455.400 ;
        RECT 158.100 455.400 160.500 456.900 ;
        RECT 163.800 455.400 165.600 468.000 ;
        RECT 179.100 461.400 180.900 468.000 ;
        RECT 182.100 461.400 183.900 467.400 ;
        RECT 185.100 461.400 186.900 468.000 ;
        RECT 200.100 461.400 201.900 468.000 ;
        RECT 203.100 461.400 204.900 467.400 ;
        RECT 158.100 448.050 159.300 455.400 ;
        RECT 164.100 448.050 165.900 449.850 ;
        RECT 182.700 448.050 183.900 461.400 ;
        RECT 200.100 448.050 201.900 449.850 ;
        RECT 203.100 448.050 204.300 461.400 ;
        RECT 218.100 456.600 219.900 467.400 ;
        RECT 221.100 457.500 222.900 468.000 ;
        RECT 224.100 466.500 231.900 467.400 ;
        RECT 224.100 456.600 225.900 466.500 ;
        RECT 218.100 455.700 225.900 456.600 ;
        RECT 227.100 454.500 228.900 465.600 ;
        RECT 230.100 455.400 231.900 466.500 ;
        RECT 245.100 455.400 246.900 467.400 ;
        RECT 248.100 455.400 249.900 468.000 ;
        RECT 263.100 461.400 264.900 468.000 ;
        RECT 266.100 461.400 267.900 467.400 ;
        RECT 269.100 461.400 270.900 468.000 ;
        RECT 224.100 453.600 228.900 454.500 ;
        RECT 221.250 448.050 223.050 449.850 ;
        RECT 224.100 448.050 225.000 453.600 ;
        RECT 227.100 448.050 228.900 449.850 ;
        RECT 245.700 448.050 246.900 455.400 ;
        RECT 266.700 448.050 267.900 461.400 ;
        RECT 287.100 455.400 288.900 467.400 ;
        RECT 290.100 456.000 291.900 468.000 ;
        RECT 293.100 461.400 294.900 467.400 ;
        RECT 296.100 461.400 297.900 468.000 ;
        RECT 314.100 461.400 315.900 468.000 ;
        RECT 317.100 461.400 318.900 467.400 ;
        RECT 320.100 461.400 321.900 468.000 ;
        RECT 335.100 461.400 336.900 468.000 ;
        RECT 338.100 461.400 339.900 467.400 ;
        RECT 341.100 461.400 342.900 468.000 ;
        RECT 356.700 461.400 358.500 468.000 ;
        RECT 268.950 453.450 271.050 454.050 ;
        RECT 280.950 453.450 283.050 454.050 ;
        RECT 268.950 452.550 283.050 453.450 ;
        RECT 268.950 451.950 271.050 452.550 ;
        RECT 280.950 451.950 283.050 452.550 ;
        RECT 287.700 448.050 288.600 455.400 ;
        RECT 291.000 448.050 292.800 449.850 ;
        RECT 112.950 445.950 115.050 448.050 ;
        RECT 115.950 445.950 118.050 448.050 ;
        RECT 130.950 445.950 133.050 448.050 ;
        RECT 133.950 445.950 136.050 448.050 ;
        RECT 136.950 445.950 139.050 448.050 ;
        RECT 139.950 445.950 142.050 448.050 ;
        RECT 154.950 445.950 157.050 448.050 ;
        RECT 157.950 445.950 160.050 448.050 ;
        RECT 160.950 445.950 163.050 448.050 ;
        RECT 163.950 445.950 166.050 448.050 ;
        RECT 178.950 445.950 181.050 448.050 ;
        RECT 181.950 445.950 184.050 448.050 ;
        RECT 184.950 445.950 187.050 448.050 ;
        RECT 199.950 445.950 202.050 448.050 ;
        RECT 202.950 445.950 205.050 448.050 ;
        RECT 217.950 445.950 220.050 448.050 ;
        RECT 220.950 445.950 223.050 448.050 ;
        RECT 223.950 445.950 226.050 448.050 ;
        RECT 226.950 445.950 229.050 448.050 ;
        RECT 229.950 445.950 232.050 448.050 ;
        RECT 244.950 445.950 247.050 448.050 ;
        RECT 247.950 445.950 250.050 448.050 ;
        RECT 262.950 445.950 265.050 448.050 ;
        RECT 265.950 445.950 268.050 448.050 ;
        RECT 268.950 445.950 271.050 448.050 ;
        RECT 287.100 445.950 289.200 448.050 ;
        RECT 290.400 445.950 292.500 448.050 ;
        RECT 79.200 435.600 80.250 436.500 ;
        RECT 88.050 436.200 90.150 437.700 ;
        RECT 86.250 435.600 90.150 436.200 ;
        RECT 70.950 432.600 72.750 435.600 ;
        RECT 75.450 432.000 77.250 435.600 ;
        RECT 78.450 432.600 80.250 435.600 ;
        RECT 81.750 432.000 83.550 435.600 ;
        RECT 86.250 434.700 89.850 435.600 ;
        RECT 86.250 432.600 88.050 434.700 ;
        RECT 91.050 432.000 92.850 438.600 ;
        RECT 94.050 436.800 96.450 438.600 ;
        RECT 94.050 432.600 95.850 436.800 ;
        RECT 116.100 435.600 117.300 445.950 ;
        RECT 134.100 444.150 135.900 445.950 ;
        RECT 137.700 441.600 138.900 445.950 ;
        RECT 140.100 444.150 141.900 445.950 ;
        RECT 142.950 444.450 145.050 445.050 ;
        RECT 148.950 444.450 151.050 445.050 ;
        RECT 142.950 443.550 151.050 444.450 ;
        RECT 155.100 444.150 156.900 445.950 ;
        RECT 142.950 442.950 145.050 443.550 ;
        RECT 148.950 442.950 151.050 443.550 ;
        RECT 158.100 441.600 159.300 445.950 ;
        RECT 161.100 444.150 162.900 445.950 ;
        RECT 179.100 444.150 180.900 445.950 ;
        RECT 137.700 440.700 141.300 441.600 ;
        RECT 131.100 437.700 138.900 439.050 ;
        RECT 113.100 432.000 114.900 435.600 ;
        RECT 116.100 432.600 117.900 435.600 ;
        RECT 131.100 432.600 132.900 437.700 ;
        RECT 134.100 432.000 135.900 436.800 ;
        RECT 137.100 432.600 138.900 437.700 ;
        RECT 140.100 438.600 141.300 440.700 ;
        RECT 155.700 440.700 159.300 441.600 ;
        RECT 182.700 440.700 183.900 445.950 ;
        RECT 184.950 444.150 186.750 445.950 ;
        RECT 155.700 438.600 156.900 440.700 ;
        RECT 179.700 439.800 183.900 440.700 ;
        RECT 140.100 432.600 141.900 438.600 ;
        RECT 155.100 432.600 156.900 438.600 ;
        RECT 158.100 437.700 165.900 439.050 ;
        RECT 158.100 432.600 159.900 437.700 ;
        RECT 161.100 432.000 162.900 436.800 ;
        RECT 164.100 432.600 165.900 437.700 ;
        RECT 179.700 432.600 181.500 439.800 ;
        RECT 184.800 432.000 186.600 438.600 ;
        RECT 203.100 435.600 204.300 445.950 ;
        RECT 218.250 444.150 220.050 445.950 ;
        RECT 224.100 438.600 225.300 445.950 ;
        RECT 230.100 444.150 231.900 445.950 ;
        RECT 245.700 438.600 246.900 445.950 ;
        RECT 248.100 444.150 249.900 445.950 ;
        RECT 263.100 444.150 264.900 445.950 ;
        RECT 266.700 440.700 267.900 445.950 ;
        RECT 268.950 444.150 270.750 445.950 ;
        RECT 263.700 439.800 267.900 440.700 ;
        RECT 200.100 432.000 201.900 435.600 ;
        RECT 203.100 432.600 204.900 435.600 ;
        RECT 218.700 432.000 220.500 438.600 ;
        RECT 223.200 432.600 225.000 438.600 ;
        RECT 227.700 432.000 229.500 438.600 ;
        RECT 245.100 432.600 246.900 438.600 ;
        RECT 248.100 432.000 249.900 438.600 ;
        RECT 263.700 432.600 265.500 439.800 ;
        RECT 287.700 438.600 288.600 445.950 ;
        RECT 294.000 441.300 294.900 461.400 ;
        RECT 317.100 448.050 318.300 461.400 ;
        RECT 338.100 448.050 339.300 461.400 ;
        RECT 357.000 458.100 358.800 459.900 ;
        RECT 359.700 456.900 361.500 467.400 ;
        RECT 359.100 455.400 361.500 456.900 ;
        RECT 364.800 455.400 366.600 468.000 ;
        RECT 380.100 456.300 381.900 467.400 ;
        RECT 383.100 457.200 384.900 468.000 ;
        RECT 386.100 456.300 387.900 467.400 ;
        RECT 380.100 455.400 387.900 456.300 ;
        RECT 389.100 455.400 390.900 467.400 ;
        RECT 404.100 461.400 405.900 468.000 ;
        RECT 407.100 461.400 408.900 467.400 ;
        RECT 410.100 462.000 411.900 468.000 ;
        RECT 407.400 461.100 408.900 461.400 ;
        RECT 413.100 461.400 414.900 467.400 ;
        RECT 413.100 461.100 414.000 461.400 ;
        RECT 407.400 460.200 414.000 461.100 ;
        RECT 400.950 456.450 403.050 457.050 ;
        RECT 406.950 456.450 409.050 457.050 ;
        RECT 400.950 455.550 409.050 456.450 ;
        RECT 359.100 448.050 360.300 455.400 ;
        RECT 370.950 453.450 373.050 454.050 ;
        RECT 385.950 453.450 388.050 454.050 ;
        RECT 370.950 452.550 388.050 453.450 ;
        RECT 370.950 451.950 373.050 452.550 ;
        RECT 385.950 451.950 388.050 452.550 ;
        RECT 365.100 448.050 366.900 449.850 ;
        RECT 383.250 448.050 385.050 449.850 ;
        RECT 389.700 448.050 390.600 455.400 ;
        RECT 400.950 454.950 403.050 455.550 ;
        RECT 406.950 454.950 409.050 455.550 ;
        RECT 409.950 453.450 412.050 453.900 ;
        RECT 401.550 452.550 412.050 453.450 ;
        RECT 401.550 450.450 402.450 452.550 ;
        RECT 409.950 451.800 412.050 452.550 ;
        RECT 398.550 449.550 402.450 450.450 ;
        RECT 295.800 445.950 297.900 448.050 ;
        RECT 313.950 445.950 316.050 448.050 ;
        RECT 316.950 445.950 319.050 448.050 ;
        RECT 319.950 445.950 322.050 448.050 ;
        RECT 334.950 445.950 337.050 448.050 ;
        RECT 337.950 445.950 340.050 448.050 ;
        RECT 340.950 445.950 343.050 448.050 ;
        RECT 355.950 445.950 358.050 448.050 ;
        RECT 358.950 445.950 361.050 448.050 ;
        RECT 361.950 445.950 364.050 448.050 ;
        RECT 364.950 445.950 367.050 448.050 ;
        RECT 379.950 445.950 382.050 448.050 ;
        RECT 382.950 445.950 385.050 448.050 ;
        RECT 385.950 445.950 388.050 448.050 ;
        RECT 388.950 445.950 391.050 448.050 ;
        RECT 295.950 444.150 297.750 445.950 ;
        RECT 314.250 444.150 316.050 445.950 ;
        RECT 289.500 440.400 297.900 441.300 ;
        RECT 289.500 439.500 291.300 440.400 ;
        RECT 268.800 432.000 270.600 438.600 ;
        RECT 287.700 436.800 290.400 438.600 ;
        RECT 288.600 432.600 290.400 436.800 ;
        RECT 291.600 432.000 293.400 438.600 ;
        RECT 296.100 432.600 297.900 440.400 ;
        RECT 317.100 440.700 318.300 445.950 ;
        RECT 320.100 444.150 321.900 445.950 ;
        RECT 335.250 444.150 337.050 445.950 ;
        RECT 338.100 440.700 339.300 445.950 ;
        RECT 341.100 444.150 342.900 445.950 ;
        RECT 356.100 444.150 357.900 445.950 ;
        RECT 359.100 441.600 360.300 445.950 ;
        RECT 362.100 444.150 363.900 445.950 ;
        RECT 380.100 444.150 381.900 445.950 ;
        RECT 386.250 444.150 388.050 445.950 ;
        RECT 356.700 440.700 360.300 441.600 ;
        RECT 317.100 439.800 321.300 440.700 ;
        RECT 338.100 439.800 342.300 440.700 ;
        RECT 314.400 432.000 316.200 438.600 ;
        RECT 319.500 432.600 321.300 439.800 ;
        RECT 335.400 432.000 337.200 438.600 ;
        RECT 340.500 432.600 342.300 439.800 ;
        RECT 356.700 438.600 357.900 440.700 ;
        RECT 356.100 432.600 357.900 438.600 ;
        RECT 359.100 437.700 366.900 439.050 ;
        RECT 389.700 438.600 390.600 445.950 ;
        RECT 398.550 445.050 399.450 449.550 ;
        RECT 407.100 448.050 408.900 449.850 ;
        RECT 413.100 448.050 414.000 460.200 ;
        RECT 428.400 455.400 430.200 468.000 ;
        RECT 433.500 456.900 435.300 467.400 ;
        RECT 436.500 461.400 438.300 468.000 ;
        RECT 436.200 458.100 438.000 459.900 ;
        RECT 433.500 455.400 435.900 456.900 ;
        RECT 452.400 455.400 454.200 468.000 ;
        RECT 457.500 456.900 459.300 467.400 ;
        RECT 460.500 461.400 462.300 468.000 ;
        RECT 476.100 461.400 477.900 468.000 ;
        RECT 479.100 461.400 480.900 467.400 ;
        RECT 482.100 462.000 483.900 468.000 ;
        RECT 479.400 461.100 480.900 461.400 ;
        RECT 485.100 461.400 486.900 467.400 ;
        RECT 500.100 461.400 501.900 468.000 ;
        RECT 503.100 461.400 504.900 467.400 ;
        RECT 506.100 462.000 507.900 468.000 ;
        RECT 485.100 461.100 486.000 461.400 ;
        RECT 479.400 460.200 486.000 461.100 ;
        RECT 503.400 461.100 504.900 461.400 ;
        RECT 509.100 461.400 510.900 467.400 ;
        RECT 524.100 461.400 525.900 468.000 ;
        RECT 527.100 461.400 528.900 467.400 ;
        RECT 509.100 461.100 510.000 461.400 ;
        RECT 503.400 460.200 510.000 461.100 ;
        RECT 460.200 458.100 462.000 459.900 ;
        RECT 457.500 455.400 459.900 456.900 ;
        RECT 428.100 448.050 429.900 449.850 ;
        RECT 434.700 448.050 435.900 455.400 ;
        RECT 452.100 448.050 453.900 449.850 ;
        RECT 458.700 448.050 459.900 455.400 ;
        RECT 466.950 453.450 469.050 454.050 ;
        RECT 481.950 453.450 484.050 454.200 ;
        RECT 466.950 452.550 484.050 453.450 ;
        RECT 466.950 451.950 469.050 452.550 ;
        RECT 481.950 452.100 484.050 452.550 ;
        RECT 479.100 448.050 480.900 449.850 ;
        RECT 485.100 448.050 486.000 460.200 ;
        RECT 487.950 453.450 490.050 454.050 ;
        RECT 505.950 453.450 508.050 454.050 ;
        RECT 487.950 452.550 508.050 453.450 ;
        RECT 487.950 451.950 490.050 452.550 ;
        RECT 505.950 451.950 508.050 452.550 ;
        RECT 503.100 448.050 504.900 449.850 ;
        RECT 509.100 448.050 510.000 460.200 ;
        RECT 524.100 448.050 525.900 449.850 ;
        RECT 527.100 448.050 528.300 461.400 ;
        RECT 542.400 455.400 544.200 468.000 ;
        RECT 547.500 456.900 549.300 467.400 ;
        RECT 550.500 461.400 552.300 468.000 ;
        RECT 566.100 461.400 567.900 468.000 ;
        RECT 569.100 461.400 570.900 467.400 ;
        RECT 572.100 461.400 573.900 468.000 ;
        RECT 550.200 458.100 552.000 459.900 ;
        RECT 547.500 455.400 549.900 456.900 ;
        RECT 542.100 448.050 543.900 449.850 ;
        RECT 548.700 448.050 549.900 455.400 ;
        RECT 561.000 450.450 565.050 451.050 ;
        RECT 560.550 448.950 565.050 450.450 ;
        RECT 403.950 445.950 406.050 448.050 ;
        RECT 406.950 445.950 409.050 448.050 ;
        RECT 409.950 445.950 412.050 448.050 ;
        RECT 412.950 445.950 415.050 448.050 ;
        RECT 427.950 445.950 430.050 448.050 ;
        RECT 430.950 445.950 433.050 448.050 ;
        RECT 433.950 445.950 436.050 448.050 ;
        RECT 436.950 445.950 439.050 448.050 ;
        RECT 451.950 445.950 454.050 448.050 ;
        RECT 454.950 445.950 457.050 448.050 ;
        RECT 457.950 445.950 460.050 448.050 ;
        RECT 460.950 445.950 463.050 448.050 ;
        RECT 475.950 445.950 478.050 448.050 ;
        RECT 478.950 445.950 481.050 448.050 ;
        RECT 481.950 445.950 484.050 448.050 ;
        RECT 484.950 445.950 487.050 448.050 ;
        RECT 499.950 445.950 502.050 448.050 ;
        RECT 502.950 445.950 505.050 448.050 ;
        RECT 505.950 445.950 508.050 448.050 ;
        RECT 508.950 445.950 511.050 448.050 ;
        RECT 523.950 445.950 526.050 448.050 ;
        RECT 526.950 445.950 529.050 448.050 ;
        RECT 541.950 445.950 544.050 448.050 ;
        RECT 544.950 445.950 547.050 448.050 ;
        RECT 547.950 445.950 550.050 448.050 ;
        RECT 550.950 445.950 553.050 448.050 ;
        RECT 398.550 443.550 403.050 445.050 ;
        RECT 404.100 444.150 405.900 445.950 ;
        RECT 410.100 444.150 411.900 445.950 ;
        RECT 399.000 442.950 403.050 443.550 ;
        RECT 413.100 442.200 414.000 445.950 ;
        RECT 431.100 444.150 432.900 445.950 ;
        RECT 359.100 432.600 360.900 437.700 ;
        RECT 362.100 432.000 363.900 436.800 ;
        RECT 365.100 432.600 366.900 437.700 ;
        RECT 381.000 432.000 382.800 438.600 ;
        RECT 385.500 437.400 390.600 438.600 ;
        RECT 385.500 432.600 387.300 437.400 ;
        RECT 388.500 432.000 390.300 435.600 ;
        RECT 404.100 432.000 405.900 441.600 ;
        RECT 410.700 441.000 414.000 442.200 ;
        RECT 434.700 441.600 435.900 445.950 ;
        RECT 437.100 444.150 438.900 445.950 ;
        RECT 455.100 444.150 456.900 445.950 ;
        RECT 458.700 441.600 459.900 445.950 ;
        RECT 461.100 444.150 462.900 445.950 ;
        RECT 476.100 444.150 477.900 445.950 ;
        RECT 482.100 444.150 483.900 445.950 ;
        RECT 485.100 442.200 486.000 445.950 ;
        RECT 500.100 444.150 501.900 445.950 ;
        RECT 506.100 444.150 507.900 445.950 ;
        RECT 509.100 442.200 510.000 445.950 ;
        RECT 410.700 432.600 412.500 441.000 ;
        RECT 434.700 440.700 438.300 441.600 ;
        RECT 458.700 440.700 462.300 441.600 ;
        RECT 428.100 437.700 435.900 439.050 ;
        RECT 428.100 432.600 429.900 437.700 ;
        RECT 431.100 432.000 432.900 436.800 ;
        RECT 434.100 432.600 435.900 437.700 ;
        RECT 437.100 438.600 438.300 440.700 ;
        RECT 437.100 432.600 438.900 438.600 ;
        RECT 452.100 437.700 459.900 439.050 ;
        RECT 452.100 432.600 453.900 437.700 ;
        RECT 455.100 432.000 456.900 436.800 ;
        RECT 458.100 432.600 459.900 437.700 ;
        RECT 461.100 438.600 462.300 440.700 ;
        RECT 461.100 432.600 462.900 438.600 ;
        RECT 476.100 432.000 477.900 441.600 ;
        RECT 482.700 441.000 486.000 442.200 ;
        RECT 482.700 432.600 484.500 441.000 ;
        RECT 500.100 432.000 501.900 441.600 ;
        RECT 506.700 441.000 510.000 442.200 ;
        RECT 506.700 432.600 508.500 441.000 ;
        RECT 527.100 435.600 528.300 445.950 ;
        RECT 545.100 444.150 546.900 445.950 ;
        RECT 548.700 441.600 549.900 445.950 ;
        RECT 551.100 444.150 552.900 445.950 ;
        RECT 553.950 444.450 556.050 445.050 ;
        RECT 560.550 444.450 561.450 448.950 ;
        RECT 569.700 448.050 570.900 461.400 ;
        RECT 590.400 455.400 592.200 468.000 ;
        RECT 595.500 456.900 597.300 467.400 ;
        RECT 598.500 461.400 600.300 468.000 ;
        RECT 617.100 461.400 618.900 467.400 ;
        RECT 620.100 462.000 621.900 468.000 ;
        RECT 618.000 461.100 618.900 461.400 ;
        RECT 623.100 461.400 624.900 467.400 ;
        RECT 626.100 461.400 627.900 468.000 ;
        RECT 623.100 461.100 624.600 461.400 ;
        RECT 618.000 460.200 624.600 461.100 ;
        RECT 598.200 458.100 600.000 459.900 ;
        RECT 595.500 455.400 597.900 456.900 ;
        RECT 590.100 448.050 591.900 449.850 ;
        RECT 596.700 448.050 597.900 455.400 ;
        RECT 618.000 448.050 618.900 460.200 ;
        RECT 644.100 455.400 645.900 467.400 ;
        RECT 647.100 456.300 648.900 467.400 ;
        RECT 650.100 457.200 651.900 468.000 ;
        RECT 653.100 456.300 654.900 467.400 ;
        RECT 668.100 461.400 669.900 467.400 ;
        RECT 671.100 462.000 672.900 468.000 ;
        RECT 647.100 455.400 654.900 456.300 ;
        RECT 669.000 461.100 669.900 461.400 ;
        RECT 674.100 461.400 675.900 467.400 ;
        RECT 677.100 461.400 678.900 468.000 ;
        RECT 692.100 461.400 693.900 467.400 ;
        RECT 695.100 462.000 696.900 468.000 ;
        RECT 674.100 461.100 675.600 461.400 ;
        RECT 669.000 460.200 675.600 461.100 ;
        RECT 693.000 461.100 693.900 461.400 ;
        RECT 698.100 461.400 699.900 467.400 ;
        RECT 701.100 461.400 702.900 468.000 ;
        RECT 716.100 461.400 717.900 467.400 ;
        RECT 719.100 462.000 720.900 468.000 ;
        RECT 698.100 461.100 699.600 461.400 ;
        RECT 693.000 460.200 699.600 461.100 ;
        RECT 717.000 461.100 717.900 461.400 ;
        RECT 722.100 461.400 723.900 467.400 ;
        RECT 725.100 461.400 726.900 468.000 ;
        RECT 722.100 461.100 723.600 461.400 ;
        RECT 717.000 460.200 723.600 461.100 ;
        RECT 623.100 448.050 624.900 449.850 ;
        RECT 644.400 448.050 645.300 455.400 ;
        RECT 652.950 453.450 655.050 454.050 ;
        RECT 664.950 453.450 667.050 454.050 ;
        RECT 652.950 452.550 667.050 453.450 ;
        RECT 652.950 451.950 655.050 452.550 ;
        RECT 664.950 451.950 667.050 452.550 ;
        RECT 649.950 448.050 651.750 449.850 ;
        RECT 669.000 448.050 669.900 460.200 ;
        RECT 670.950 453.450 673.050 454.050 ;
        RECT 670.950 452.550 681.450 453.450 ;
        RECT 670.950 451.950 673.050 452.550 ;
        RECT 680.550 450.450 681.450 452.550 ;
        RECT 674.100 448.050 675.900 449.850 ;
        RECT 680.550 449.550 684.450 450.450 ;
        RECT 565.950 445.950 568.050 448.050 ;
        RECT 568.950 445.950 571.050 448.050 ;
        RECT 571.950 445.950 574.050 448.050 ;
        RECT 589.950 445.950 592.050 448.050 ;
        RECT 592.950 445.950 595.050 448.050 ;
        RECT 595.950 445.950 598.050 448.050 ;
        RECT 598.950 445.950 601.050 448.050 ;
        RECT 616.950 445.950 619.050 448.050 ;
        RECT 619.950 445.950 622.050 448.050 ;
        RECT 622.950 445.950 625.050 448.050 ;
        RECT 625.950 445.950 628.050 448.050 ;
        RECT 643.950 445.950 646.050 448.050 ;
        RECT 646.950 445.950 649.050 448.050 ;
        RECT 649.950 445.950 652.050 448.050 ;
        RECT 652.950 445.950 655.050 448.050 ;
        RECT 667.950 445.950 670.050 448.050 ;
        RECT 670.950 445.950 673.050 448.050 ;
        RECT 673.950 445.950 676.050 448.050 ;
        RECT 676.950 445.950 679.050 448.050 ;
        RECT 553.950 443.550 561.450 444.450 ;
        RECT 566.100 444.150 567.900 445.950 ;
        RECT 553.950 442.950 556.050 443.550 ;
        RECT 548.700 440.700 552.300 441.600 ;
        RECT 569.700 440.700 570.900 445.950 ;
        RECT 571.950 444.150 573.750 445.950 ;
        RECT 593.100 444.150 594.900 445.950 ;
        RECT 596.700 441.600 597.900 445.950 ;
        RECT 599.100 444.150 600.900 445.950 ;
        RECT 618.000 442.200 618.900 445.950 ;
        RECT 620.100 444.150 621.900 445.950 ;
        RECT 626.100 444.150 627.900 445.950 ;
        RECT 596.700 440.700 600.300 441.600 ;
        RECT 618.000 441.000 621.300 442.200 ;
        RECT 542.100 437.700 549.900 439.050 ;
        RECT 524.100 432.000 525.900 435.600 ;
        RECT 527.100 432.600 528.900 435.600 ;
        RECT 542.100 432.600 543.900 437.700 ;
        RECT 545.100 432.000 546.900 436.800 ;
        RECT 548.100 432.600 549.900 437.700 ;
        RECT 551.100 438.600 552.300 440.700 ;
        RECT 566.700 439.800 570.900 440.700 ;
        RECT 551.100 432.600 552.900 438.600 ;
        RECT 566.700 432.600 568.500 439.800 ;
        RECT 571.800 432.000 573.600 438.600 ;
        RECT 590.100 437.700 597.900 439.050 ;
        RECT 590.100 432.600 591.900 437.700 ;
        RECT 593.100 432.000 594.900 436.800 ;
        RECT 596.100 432.600 597.900 437.700 ;
        RECT 599.100 438.600 600.300 440.700 ;
        RECT 599.100 432.600 600.900 438.600 ;
        RECT 619.500 432.600 621.300 441.000 ;
        RECT 626.100 432.000 627.900 441.600 ;
        RECT 644.400 438.600 645.300 445.950 ;
        RECT 646.950 444.150 648.750 445.950 ;
        RECT 653.100 444.150 654.900 445.950 ;
        RECT 669.000 442.200 669.900 445.950 ;
        RECT 671.100 444.150 672.900 445.950 ;
        RECT 677.100 444.150 678.900 445.950 ;
        RECT 683.550 444.450 684.450 449.550 ;
        RECT 693.000 448.050 693.900 460.200 ;
        RECT 698.100 448.050 699.900 449.850 ;
        RECT 717.000 448.050 717.900 460.200 ;
        RECT 740.100 455.400 741.900 467.400 ;
        RECT 743.100 456.300 744.900 467.400 ;
        RECT 746.100 457.200 747.900 468.000 ;
        RECT 749.100 456.300 750.900 467.400 ;
        RECT 764.100 461.400 765.900 467.400 ;
        RECT 767.100 461.400 768.900 468.000 ;
        RECT 782.700 461.400 784.500 468.000 ;
        RECT 743.100 455.400 750.900 456.300 ;
        RECT 724.950 453.450 727.050 454.050 ;
        RECT 733.950 453.450 736.050 454.050 ;
        RECT 724.950 452.550 736.050 453.450 ;
        RECT 724.950 451.950 727.050 452.550 ;
        RECT 733.950 451.950 736.050 452.550 ;
        RECT 722.100 448.050 723.900 449.850 ;
        RECT 740.400 448.050 741.300 455.400 ;
        RECT 745.950 448.050 747.750 449.850 ;
        RECT 764.700 448.050 765.900 461.400 ;
        RECT 783.000 458.100 784.800 459.900 ;
        RECT 785.700 456.900 787.500 467.400 ;
        RECT 785.100 455.400 787.500 456.900 ;
        RECT 790.800 455.400 792.600 468.000 ;
        RECT 809.100 455.400 810.900 467.400 ;
        RECT 812.100 456.300 813.900 467.400 ;
        RECT 815.100 457.200 816.900 468.000 ;
        RECT 818.100 456.300 819.900 467.400 ;
        RECT 833.100 461.400 834.900 467.400 ;
        RECT 836.100 462.000 837.900 468.000 ;
        RECT 812.100 455.400 819.900 456.300 ;
        RECT 834.000 461.100 834.900 461.400 ;
        RECT 839.100 461.400 840.900 467.400 ;
        RECT 842.100 461.400 843.900 468.000 ;
        RECT 857.100 461.400 858.900 467.400 ;
        RECT 860.100 462.000 861.900 468.000 ;
        RECT 839.100 461.100 840.600 461.400 ;
        RECT 834.000 460.200 840.600 461.100 ;
        RECT 858.000 461.100 858.900 461.400 ;
        RECT 863.100 461.400 864.900 467.400 ;
        RECT 866.100 461.400 867.900 468.000 ;
        RECT 863.100 461.100 864.600 461.400 ;
        RECT 858.000 460.200 864.600 461.100 ;
        RECT 767.100 448.050 768.900 449.850 ;
        RECT 785.100 448.050 786.300 455.400 ;
        RECT 791.100 448.050 792.900 449.850 ;
        RECT 809.400 448.050 810.300 455.400 ;
        RECT 814.950 448.050 816.750 449.850 ;
        RECT 834.000 448.050 834.900 460.200 ;
        RECT 835.950 453.450 838.050 454.050 ;
        RECT 850.950 453.450 853.050 454.050 ;
        RECT 835.950 452.550 853.050 453.450 ;
        RECT 835.950 451.950 838.050 452.550 ;
        RECT 850.950 451.950 853.050 452.550 ;
        RECT 839.100 448.050 840.900 449.850 ;
        RECT 858.000 448.050 858.900 460.200 ;
        RECT 884.100 456.300 885.900 467.400 ;
        RECT 887.100 457.200 888.900 468.000 ;
        RECT 890.100 456.300 891.900 467.400 ;
        RECT 884.100 455.400 891.900 456.300 ;
        RECT 893.100 455.400 894.900 467.400 ;
        RECT 865.950 453.450 868.050 454.050 ;
        RECT 889.950 453.450 892.050 454.050 ;
        RECT 865.950 452.550 892.050 453.450 ;
        RECT 865.950 451.950 868.050 452.550 ;
        RECT 889.950 451.950 892.050 452.550 ;
        RECT 863.100 448.050 864.900 449.850 ;
        RECT 887.250 448.050 889.050 449.850 ;
        RECT 893.700 448.050 894.600 455.400 ;
        RECT 691.950 445.950 694.050 448.050 ;
        RECT 694.950 445.950 697.050 448.050 ;
        RECT 697.950 445.950 700.050 448.050 ;
        RECT 700.950 445.950 703.050 448.050 ;
        RECT 715.950 445.950 718.050 448.050 ;
        RECT 718.950 445.950 721.050 448.050 ;
        RECT 721.950 445.950 724.050 448.050 ;
        RECT 724.950 445.950 727.050 448.050 ;
        RECT 739.950 445.950 742.050 448.050 ;
        RECT 742.950 445.950 745.050 448.050 ;
        RECT 745.950 445.950 748.050 448.050 ;
        RECT 748.950 445.950 751.050 448.050 ;
        RECT 763.950 445.950 766.050 448.050 ;
        RECT 766.950 445.950 769.050 448.050 ;
        RECT 781.950 445.950 784.050 448.050 ;
        RECT 784.950 445.950 787.050 448.050 ;
        RECT 787.950 445.950 790.050 448.050 ;
        RECT 790.950 445.950 793.050 448.050 ;
        RECT 808.950 445.950 811.050 448.050 ;
        RECT 811.950 445.950 814.050 448.050 ;
        RECT 814.950 445.950 817.050 448.050 ;
        RECT 817.950 445.950 820.050 448.050 ;
        RECT 832.950 445.950 835.050 448.050 ;
        RECT 835.950 445.950 838.050 448.050 ;
        RECT 838.950 445.950 841.050 448.050 ;
        RECT 841.950 445.950 844.050 448.050 ;
        RECT 856.950 445.950 859.050 448.050 ;
        RECT 859.950 445.950 862.050 448.050 ;
        RECT 862.950 445.950 865.050 448.050 ;
        RECT 865.950 445.950 868.050 448.050 ;
        RECT 688.950 444.450 691.050 445.050 ;
        RECT 683.550 443.550 691.050 444.450 ;
        RECT 688.950 442.950 691.050 443.550 ;
        RECT 693.000 442.200 693.900 445.950 ;
        RECT 695.100 444.150 696.900 445.950 ;
        RECT 701.100 444.150 702.900 445.950 ;
        RECT 717.000 442.200 717.900 445.950 ;
        RECT 719.100 444.150 720.900 445.950 ;
        RECT 725.100 444.150 726.900 445.950 ;
        RECT 669.000 441.000 672.300 442.200 ;
        RECT 644.400 437.400 649.500 438.600 ;
        RECT 644.700 432.000 646.500 435.600 ;
        RECT 647.700 432.600 649.500 437.400 ;
        RECT 652.200 432.000 654.000 438.600 ;
        RECT 670.500 432.600 672.300 441.000 ;
        RECT 677.100 432.000 678.900 441.600 ;
        RECT 693.000 441.000 696.300 442.200 ;
        RECT 694.500 432.600 696.300 441.000 ;
        RECT 701.100 432.000 702.900 441.600 ;
        RECT 717.000 441.000 720.300 442.200 ;
        RECT 718.500 432.600 720.300 441.000 ;
        RECT 725.100 432.000 726.900 441.600 ;
        RECT 740.400 438.600 741.300 445.950 ;
        RECT 742.950 444.150 744.750 445.950 ;
        RECT 749.100 444.150 750.900 445.950 ;
        RECT 740.400 437.400 745.500 438.600 ;
        RECT 740.700 432.000 742.500 435.600 ;
        RECT 743.700 432.600 745.500 437.400 ;
        RECT 748.200 432.000 750.000 438.600 ;
        RECT 764.700 435.600 765.900 445.950 ;
        RECT 782.100 444.150 783.900 445.950 ;
        RECT 785.100 441.600 786.300 445.950 ;
        RECT 788.100 444.150 789.900 445.950 ;
        RECT 782.700 440.700 786.300 441.600 ;
        RECT 782.700 438.600 783.900 440.700 ;
        RECT 764.100 432.600 765.900 435.600 ;
        RECT 767.100 432.000 768.900 435.600 ;
        RECT 782.100 432.600 783.900 438.600 ;
        RECT 785.100 437.700 792.900 439.050 ;
        RECT 785.100 432.600 786.900 437.700 ;
        RECT 788.100 432.000 789.900 436.800 ;
        RECT 791.100 432.600 792.900 437.700 ;
        RECT 809.400 438.600 810.300 445.950 ;
        RECT 811.950 444.150 813.750 445.950 ;
        RECT 818.100 444.150 819.900 445.950 ;
        RECT 834.000 442.200 834.900 445.950 ;
        RECT 836.100 444.150 837.900 445.950 ;
        RECT 842.100 444.150 843.900 445.950 ;
        RECT 858.000 442.200 858.900 445.950 ;
        RECT 860.100 444.150 861.900 445.950 ;
        RECT 866.100 444.150 867.900 445.950 ;
        RECT 877.950 444.450 880.050 448.050 ;
        RECT 883.950 445.950 886.050 448.050 ;
        RECT 886.950 445.950 889.050 448.050 ;
        RECT 889.950 445.950 892.050 448.050 ;
        RECT 892.950 445.950 895.050 448.050 ;
        RECT 877.950 444.000 882.450 444.450 ;
        RECT 884.100 444.150 885.900 445.950 ;
        RECT 890.250 444.150 892.050 445.950 ;
        RECT 878.550 443.550 882.450 444.000 ;
        RECT 834.000 441.000 837.300 442.200 ;
        RECT 809.400 437.400 814.500 438.600 ;
        RECT 809.700 432.000 811.500 435.600 ;
        RECT 812.700 432.600 814.500 437.400 ;
        RECT 817.200 432.000 819.000 438.600 ;
        RECT 835.500 432.600 837.300 441.000 ;
        RECT 842.100 432.000 843.900 441.600 ;
        RECT 858.000 441.000 861.300 442.200 ;
        RECT 859.500 432.600 861.300 441.000 ;
        RECT 866.100 432.000 867.900 441.600 ;
        RECT 881.550 441.450 882.450 443.550 ;
        RECT 889.950 441.450 892.050 442.050 ;
        RECT 881.550 440.550 892.050 441.450 ;
        RECT 889.950 439.950 892.050 440.550 ;
        RECT 893.700 438.600 894.600 445.950 ;
        RECT 885.000 432.000 886.800 438.600 ;
        RECT 889.500 437.400 894.600 438.600 ;
        RECT 889.500 432.600 891.300 437.400 ;
        RECT 892.500 432.000 894.300 435.600 ;
        RECT 14.100 422.400 15.900 428.400 ;
        RECT 17.100 422.400 18.900 429.000 ;
        RECT 20.100 425.400 21.900 428.400 ;
        RECT 14.100 415.050 15.300 422.400 ;
        RECT 20.700 421.500 21.900 425.400 ;
        RECT 16.200 420.600 21.900 421.500 ;
        RECT 35.100 422.400 36.900 428.400 ;
        RECT 38.100 422.400 39.900 429.000 ;
        RECT 41.100 425.400 42.900 428.400 ;
        RECT 16.200 419.700 18.000 420.600 ;
        RECT 14.100 412.950 16.200 415.050 ;
        RECT 14.100 405.600 15.300 412.950 ;
        RECT 17.100 408.300 18.000 419.700 ;
        RECT 35.100 415.050 36.300 422.400 ;
        RECT 41.700 421.500 42.900 425.400 ;
        RECT 37.200 420.600 42.900 421.500 ;
        RECT 56.100 422.400 57.900 428.400 ;
        RECT 59.100 422.400 60.900 429.000 ;
        RECT 62.100 425.400 63.900 428.400 ;
        RECT 37.200 419.700 39.000 420.600 ;
        RECT 19.500 412.950 21.600 415.050 ;
        RECT 19.800 411.150 21.600 412.950 ;
        RECT 35.100 412.950 37.200 415.050 ;
        RECT 16.200 407.400 18.000 408.300 ;
        RECT 16.200 406.500 21.900 407.400 ;
        RECT 14.100 393.600 15.900 405.600 ;
        RECT 17.100 393.000 18.900 403.800 ;
        RECT 20.700 399.600 21.900 406.500 ;
        RECT 20.100 393.600 21.900 399.600 ;
        RECT 35.100 405.600 36.300 412.950 ;
        RECT 38.100 408.300 39.000 419.700 ;
        RECT 56.100 415.050 57.300 422.400 ;
        RECT 62.700 421.500 63.900 425.400 ;
        RECT 58.200 420.600 63.900 421.500 ;
        RECT 65.550 422.400 67.350 428.400 ;
        RECT 68.850 422.400 70.650 429.000 ;
        RECT 73.950 425.400 75.750 428.400 ;
        RECT 78.450 425.400 80.250 429.000 ;
        RECT 81.450 425.400 83.250 428.400 ;
        RECT 84.750 425.400 86.550 429.000 ;
        RECT 89.250 426.300 91.050 428.400 ;
        RECT 89.250 425.400 92.850 426.300 ;
        RECT 73.350 423.300 75.750 425.400 ;
        RECT 82.200 424.500 83.250 425.400 ;
        RECT 89.250 424.800 93.150 425.400 ;
        RECT 82.200 423.450 87.150 424.500 ;
        RECT 85.350 422.700 87.150 423.450 ;
        RECT 58.200 419.700 60.000 420.600 ;
        RECT 40.500 412.950 42.600 415.050 ;
        RECT 40.800 411.150 42.600 412.950 ;
        RECT 56.100 412.950 58.200 415.050 ;
        RECT 37.200 407.400 39.000 408.300 ;
        RECT 37.200 406.500 42.900 407.400 ;
        RECT 35.100 393.600 36.900 405.600 ;
        RECT 38.100 393.000 39.900 403.800 ;
        RECT 41.700 399.600 42.900 406.500 ;
        RECT 41.100 393.600 42.900 399.600 ;
        RECT 56.100 405.600 57.300 412.950 ;
        RECT 59.100 408.300 60.000 419.700 ;
        RECT 65.550 415.050 66.750 422.400 ;
        RECT 88.350 421.800 90.150 423.600 ;
        RECT 91.050 423.300 93.150 424.800 ;
        RECT 94.050 422.400 95.850 429.000 ;
        RECT 97.050 424.200 98.850 428.400 ;
        RECT 97.050 422.400 99.450 424.200 ;
        RECT 78.150 420.000 79.950 420.600 ;
        RECT 89.100 420.000 90.150 421.800 ;
        RECT 78.150 418.800 90.150 420.000 ;
        RECT 61.500 412.950 63.600 415.050 ;
        RECT 61.800 411.150 63.600 412.950 ;
        RECT 65.550 413.250 71.850 415.050 ;
        RECT 65.550 412.950 70.050 413.250 ;
        RECT 58.200 407.400 60.000 408.300 ;
        RECT 58.200 406.500 63.900 407.400 ;
        RECT 56.100 393.600 57.900 405.600 ;
        RECT 59.100 393.000 60.900 403.800 ;
        RECT 62.700 399.600 63.900 406.500 ;
        RECT 62.100 393.600 63.900 399.600 ;
        RECT 65.550 405.600 66.750 412.950 ;
        RECT 67.650 410.100 69.450 410.250 ;
        RECT 73.350 410.100 75.450 410.400 ;
        RECT 67.650 408.900 75.450 410.100 ;
        RECT 67.650 408.450 69.450 408.900 ;
        RECT 73.350 408.300 75.450 408.900 ;
        RECT 78.150 406.200 79.050 418.800 ;
        RECT 89.100 417.600 97.050 418.800 ;
        RECT 89.100 417.000 90.900 417.600 ;
        RECT 92.100 415.800 93.900 416.400 ;
        RECT 85.800 414.600 93.900 415.800 ;
        RECT 95.250 415.050 97.050 417.600 ;
        RECT 85.800 412.950 87.900 414.600 ;
        RECT 94.950 412.950 97.050 415.050 ;
        RECT 87.750 407.700 89.550 408.000 ;
        RECT 98.550 407.700 99.450 422.400 ;
        RECT 87.750 407.100 99.450 407.700 ;
        RECT 65.550 393.600 67.350 405.600 ;
        RECT 68.550 393.000 70.350 405.600 ;
        RECT 74.250 405.300 79.050 406.200 ;
        RECT 81.150 406.500 99.450 407.100 ;
        RECT 81.150 406.200 89.550 406.500 ;
        RECT 74.250 404.400 75.450 405.300 ;
        RECT 72.450 402.600 75.450 404.400 ;
        RECT 76.350 404.100 78.150 404.400 ;
        RECT 81.150 404.100 82.050 406.200 ;
        RECT 98.550 405.600 99.450 406.500 ;
        RECT 76.350 403.200 82.050 404.100 ;
        RECT 82.950 404.700 84.750 405.300 ;
        RECT 82.950 403.500 90.750 404.700 ;
        RECT 76.350 402.600 78.150 403.200 ;
        RECT 88.650 402.600 90.750 403.500 ;
        RECT 73.350 399.600 75.450 401.700 ;
        RECT 79.950 401.550 81.750 402.300 ;
        RECT 84.750 401.550 86.550 402.300 ;
        RECT 79.950 400.500 86.550 401.550 ;
        RECT 73.350 393.600 75.150 399.600 ;
        RECT 77.850 393.000 79.650 399.600 ;
        RECT 80.850 393.600 82.650 400.500 ;
        RECT 83.850 393.000 85.650 399.600 ;
        RECT 88.650 393.600 90.450 402.600 ;
        RECT 94.050 393.000 95.850 405.600 ;
        RECT 97.050 403.800 99.450 405.600 ;
        RECT 101.550 422.400 103.350 428.400 ;
        RECT 104.850 422.400 106.650 429.000 ;
        RECT 109.950 425.400 111.750 428.400 ;
        RECT 114.450 425.400 116.250 429.000 ;
        RECT 117.450 425.400 119.250 428.400 ;
        RECT 120.750 425.400 122.550 429.000 ;
        RECT 125.250 426.300 127.050 428.400 ;
        RECT 125.250 425.400 128.850 426.300 ;
        RECT 109.350 423.300 111.750 425.400 ;
        RECT 118.200 424.500 119.250 425.400 ;
        RECT 125.250 424.800 129.150 425.400 ;
        RECT 118.200 423.450 123.150 424.500 ;
        RECT 121.350 422.700 123.150 423.450 ;
        RECT 101.550 415.050 102.750 422.400 ;
        RECT 124.350 421.800 126.150 423.600 ;
        RECT 127.050 423.300 129.150 424.800 ;
        RECT 130.050 422.400 131.850 429.000 ;
        RECT 133.050 424.200 134.850 428.400 ;
        RECT 149.100 425.400 150.900 429.000 ;
        RECT 152.100 425.400 153.900 428.400 ;
        RECT 133.050 422.400 135.450 424.200 ;
        RECT 114.150 420.000 115.950 420.600 ;
        RECT 125.100 420.000 126.150 421.800 ;
        RECT 114.150 418.800 126.150 420.000 ;
        RECT 101.550 413.250 107.850 415.050 ;
        RECT 101.550 412.950 106.050 413.250 ;
        RECT 101.550 405.600 102.750 412.950 ;
        RECT 103.650 410.100 105.450 410.250 ;
        RECT 109.350 410.100 111.450 410.400 ;
        RECT 103.650 408.900 111.450 410.100 ;
        RECT 103.650 408.450 105.450 408.900 ;
        RECT 109.350 408.300 111.450 408.900 ;
        RECT 114.150 406.200 115.050 418.800 ;
        RECT 125.100 417.600 133.050 418.800 ;
        RECT 125.100 417.000 126.900 417.600 ;
        RECT 128.100 415.800 129.900 416.400 ;
        RECT 121.800 414.600 129.900 415.800 ;
        RECT 131.250 415.050 133.050 417.600 ;
        RECT 121.800 412.950 123.900 414.600 ;
        RECT 130.950 412.950 133.050 415.050 ;
        RECT 123.750 407.700 125.550 408.000 ;
        RECT 134.550 407.700 135.450 422.400 ;
        RECT 152.100 415.050 153.300 425.400 ;
        RECT 167.100 422.400 168.900 429.000 ;
        RECT 170.100 421.500 171.900 428.400 ;
        RECT 173.100 422.400 174.900 429.000 ;
        RECT 176.100 421.500 177.900 428.400 ;
        RECT 179.100 422.400 180.900 429.000 ;
        RECT 182.100 421.500 183.900 428.400 ;
        RECT 185.100 422.400 186.900 429.000 ;
        RECT 188.100 421.500 189.900 428.400 ;
        RECT 191.100 422.400 192.900 429.000 ;
        RECT 206.100 425.400 207.900 428.400 ;
        RECT 209.100 425.400 210.900 429.000 ;
        RECT 169.050 420.300 171.900 421.500 ;
        RECT 174.000 420.300 177.900 421.500 ;
        RECT 180.000 420.300 183.900 421.500 ;
        RECT 186.000 420.300 189.900 421.500 ;
        RECT 169.050 415.050 170.100 420.300 ;
        RECT 174.000 419.400 175.200 420.300 ;
        RECT 180.000 419.400 181.200 420.300 ;
        RECT 186.000 419.400 187.200 420.300 ;
        RECT 171.000 418.200 175.200 419.400 ;
        RECT 171.000 417.600 172.800 418.200 ;
        RECT 148.950 412.950 151.050 415.050 ;
        RECT 151.950 412.950 154.050 415.050 ;
        RECT 169.050 412.950 172.200 415.050 ;
        RECT 149.100 411.150 150.900 412.950 ;
        RECT 123.750 407.100 135.450 407.700 ;
        RECT 97.050 393.600 98.850 403.800 ;
        RECT 101.550 393.600 103.350 405.600 ;
        RECT 104.550 393.000 106.350 405.600 ;
        RECT 110.250 405.300 115.050 406.200 ;
        RECT 117.150 406.500 135.450 407.100 ;
        RECT 117.150 406.200 125.550 406.500 ;
        RECT 110.250 404.400 111.450 405.300 ;
        RECT 108.450 402.600 111.450 404.400 ;
        RECT 112.350 404.100 114.150 404.400 ;
        RECT 117.150 404.100 118.050 406.200 ;
        RECT 134.550 405.600 135.450 406.500 ;
        RECT 112.350 403.200 118.050 404.100 ;
        RECT 118.950 404.700 120.750 405.300 ;
        RECT 118.950 403.500 126.750 404.700 ;
        RECT 112.350 402.600 114.150 403.200 ;
        RECT 124.650 402.600 126.750 403.500 ;
        RECT 109.350 399.600 111.450 401.700 ;
        RECT 115.950 401.550 117.750 402.300 ;
        RECT 120.750 401.550 122.550 402.300 ;
        RECT 115.950 400.500 122.550 401.550 ;
        RECT 109.350 393.600 111.150 399.600 ;
        RECT 113.850 393.000 115.650 399.600 ;
        RECT 116.850 393.600 118.650 400.500 ;
        RECT 119.850 393.000 121.650 399.600 ;
        RECT 124.650 393.600 126.450 402.600 ;
        RECT 130.050 393.000 131.850 405.600 ;
        RECT 133.050 403.800 135.450 405.600 ;
        RECT 133.050 393.600 134.850 403.800 ;
        RECT 152.100 399.600 153.300 412.950 ;
        RECT 169.050 407.700 170.100 412.950 ;
        RECT 174.000 407.700 175.200 418.200 ;
        RECT 177.000 418.200 181.200 419.400 ;
        RECT 177.000 417.600 178.800 418.200 ;
        RECT 180.000 407.700 181.200 418.200 ;
        RECT 183.000 418.200 187.200 419.400 ;
        RECT 183.000 417.600 184.800 418.200 ;
        RECT 186.000 407.700 187.200 418.200 ;
        RECT 188.400 415.050 190.200 416.850 ;
        RECT 206.700 415.050 207.900 425.400 ;
        RECT 224.100 422.400 225.900 429.000 ;
        RECT 227.100 421.500 228.900 428.400 ;
        RECT 230.100 422.400 231.900 429.000 ;
        RECT 233.100 421.500 234.900 428.400 ;
        RECT 236.100 422.400 237.900 429.000 ;
        RECT 239.100 421.500 240.900 428.400 ;
        RECT 242.100 422.400 243.900 429.000 ;
        RECT 245.100 421.500 246.900 428.400 ;
        RECT 248.100 422.400 249.900 429.000 ;
        RECT 263.100 423.300 264.900 428.400 ;
        RECT 266.100 424.200 267.900 429.000 ;
        RECT 269.100 423.300 270.900 428.400 ;
        RECT 263.100 421.950 270.900 423.300 ;
        RECT 272.100 422.400 273.900 428.400 ;
        RECT 287.100 423.300 288.900 428.400 ;
        RECT 290.100 424.200 291.900 429.000 ;
        RECT 293.100 423.300 294.900 428.400 ;
        RECT 227.100 420.300 231.000 421.500 ;
        RECT 233.100 420.300 237.000 421.500 ;
        RECT 239.100 420.300 243.000 421.500 ;
        RECT 245.100 420.300 247.950 421.500 ;
        RECT 272.100 420.300 273.300 422.400 ;
        RECT 287.100 421.950 294.900 423.300 ;
        RECT 296.100 422.400 297.900 428.400 ;
        RECT 296.100 420.300 297.300 422.400 ;
        RECT 229.800 419.400 231.000 420.300 ;
        RECT 235.800 419.400 237.000 420.300 ;
        RECT 241.800 419.400 243.000 420.300 ;
        RECT 229.800 418.200 234.000 419.400 ;
        RECT 226.800 415.050 228.600 416.850 ;
        RECT 188.100 412.950 190.200 415.050 ;
        RECT 205.950 412.950 208.050 415.050 ;
        RECT 208.950 412.950 211.050 415.050 ;
        RECT 226.800 412.950 228.900 415.050 ;
        RECT 169.050 406.500 171.900 407.700 ;
        RECT 174.000 406.500 177.900 407.700 ;
        RECT 180.000 406.500 183.900 407.700 ;
        RECT 186.000 406.500 189.900 407.700 ;
        RECT 149.100 393.000 150.900 399.600 ;
        RECT 152.100 393.600 153.900 399.600 ;
        RECT 167.100 393.000 168.900 405.600 ;
        RECT 170.100 393.600 171.900 406.500 ;
        RECT 173.100 393.000 174.900 405.600 ;
        RECT 176.100 393.600 177.900 406.500 ;
        RECT 179.100 393.000 180.900 405.600 ;
        RECT 182.100 393.600 183.900 406.500 ;
        RECT 185.100 393.000 186.900 405.600 ;
        RECT 188.100 393.600 189.900 406.500 ;
        RECT 191.100 393.000 192.900 405.600 ;
        RECT 206.700 399.600 207.900 412.950 ;
        RECT 209.100 411.150 210.900 412.950 ;
        RECT 229.800 407.700 231.000 418.200 ;
        RECT 232.200 417.600 234.000 418.200 ;
        RECT 235.800 418.200 240.000 419.400 ;
        RECT 235.800 407.700 237.000 418.200 ;
        RECT 238.200 417.600 240.000 418.200 ;
        RECT 241.800 418.200 246.000 419.400 ;
        RECT 241.800 407.700 243.000 418.200 ;
        RECT 244.200 417.600 246.000 418.200 ;
        RECT 246.900 415.050 247.950 420.300 ;
        RECT 269.700 419.400 273.300 420.300 ;
        RECT 293.700 419.400 297.300 420.300 ;
        RECT 314.100 420.600 315.900 428.400 ;
        RECT 318.600 422.400 320.400 429.000 ;
        RECT 321.600 424.200 323.400 428.400 ;
        RECT 321.600 422.400 324.300 424.200 ;
        RECT 320.700 420.600 322.500 421.500 ;
        RECT 314.100 419.700 322.500 420.600 ;
        RECT 266.100 415.050 267.900 416.850 ;
        RECT 269.700 415.050 270.900 419.400 ;
        RECT 272.100 415.050 273.900 416.850 ;
        RECT 290.100 415.050 291.900 416.850 ;
        RECT 293.700 415.050 294.900 419.400 ;
        RECT 296.100 415.050 297.900 416.850 ;
        RECT 314.250 415.050 316.050 416.850 ;
        RECT 244.800 412.950 247.950 415.050 ;
        RECT 262.950 412.950 265.050 415.050 ;
        RECT 265.950 412.950 268.050 415.050 ;
        RECT 268.950 412.950 271.050 415.050 ;
        RECT 271.950 412.950 274.050 415.050 ;
        RECT 286.950 412.950 289.050 415.050 ;
        RECT 289.950 412.950 292.050 415.050 ;
        RECT 292.950 412.950 295.050 415.050 ;
        RECT 295.950 412.950 298.050 415.050 ;
        RECT 314.100 412.950 316.200 415.050 ;
        RECT 246.900 407.700 247.950 412.950 ;
        RECT 263.100 411.150 264.900 412.950 ;
        RECT 227.100 406.500 231.000 407.700 ;
        RECT 233.100 406.500 237.000 407.700 ;
        RECT 239.100 406.500 243.000 407.700 ;
        RECT 245.100 406.500 247.950 407.700 ;
        RECT 206.100 393.600 207.900 399.600 ;
        RECT 209.100 393.000 210.900 399.600 ;
        RECT 224.100 393.000 225.900 405.600 ;
        RECT 227.100 393.600 228.900 406.500 ;
        RECT 230.100 393.000 231.900 405.600 ;
        RECT 233.100 393.600 234.900 406.500 ;
        RECT 236.100 393.000 237.900 405.600 ;
        RECT 239.100 393.600 240.900 406.500 ;
        RECT 242.100 393.000 243.900 405.600 ;
        RECT 245.100 393.600 246.900 406.500 ;
        RECT 269.700 405.600 270.900 412.950 ;
        RECT 287.100 411.150 288.900 412.950 ;
        RECT 271.950 408.450 274.050 409.050 ;
        RECT 277.950 408.450 280.050 409.050 ;
        RECT 271.950 407.550 280.050 408.450 ;
        RECT 271.950 406.950 274.050 407.550 ;
        RECT 277.950 406.950 280.050 407.550 ;
        RECT 293.700 405.600 294.900 412.950 ;
        RECT 248.100 393.000 249.900 405.600 ;
        RECT 263.400 393.000 265.200 405.600 ;
        RECT 268.500 404.100 270.900 405.600 ;
        RECT 268.500 393.600 270.300 404.100 ;
        RECT 271.200 401.100 273.000 402.900 ;
        RECT 271.500 393.000 273.300 399.600 ;
        RECT 287.400 393.000 289.200 405.600 ;
        RECT 292.500 404.100 294.900 405.600 ;
        RECT 292.500 393.600 294.300 404.100 ;
        RECT 295.200 401.100 297.000 402.900 ;
        RECT 317.100 399.600 318.000 419.700 ;
        RECT 323.400 415.050 324.300 422.400 ;
        RECT 338.100 420.600 339.900 428.400 ;
        RECT 342.600 422.400 344.400 429.000 ;
        RECT 345.600 424.200 347.400 428.400 ;
        RECT 345.600 422.400 348.300 424.200 ;
        RECT 362.400 422.400 364.200 429.000 ;
        RECT 344.700 420.600 346.500 421.500 ;
        RECT 338.100 419.700 346.500 420.600 ;
        RECT 338.250 415.050 340.050 416.850 ;
        RECT 319.500 412.950 321.600 415.050 ;
        RECT 322.800 412.950 324.900 415.050 ;
        RECT 338.100 412.950 340.200 415.050 ;
        RECT 319.200 411.150 321.000 412.950 ;
        RECT 323.400 405.600 324.300 412.950 ;
        RECT 295.500 393.000 297.300 399.600 ;
        RECT 314.100 393.000 315.900 399.600 ;
        RECT 317.100 393.600 318.900 399.600 ;
        RECT 320.100 393.000 321.900 405.000 ;
        RECT 323.100 393.600 324.900 405.600 ;
        RECT 341.100 399.600 342.000 419.700 ;
        RECT 347.400 415.050 348.300 422.400 ;
        RECT 367.500 421.200 369.300 428.400 ;
        RECT 383.100 425.400 384.900 429.000 ;
        RECT 386.100 425.400 387.900 428.400 ;
        RECT 365.100 420.300 369.300 421.200 ;
        RECT 362.250 415.050 364.050 416.850 ;
        RECT 365.100 415.050 366.300 420.300 ;
        RECT 368.100 415.050 369.900 416.850 ;
        RECT 386.100 415.050 387.300 425.400 ;
        RECT 402.000 422.400 403.800 429.000 ;
        RECT 406.500 423.600 408.300 428.400 ;
        RECT 409.500 425.400 411.300 429.000 ;
        RECT 406.500 422.400 411.600 423.600 ;
        RECT 401.100 415.050 402.900 416.850 ;
        RECT 407.250 415.050 409.050 416.850 ;
        RECT 410.700 415.050 411.600 422.400 ;
        RECT 428.100 419.400 429.900 429.000 ;
        RECT 434.700 420.000 436.500 428.400 ;
        RECT 454.500 420.000 456.300 428.400 ;
        RECT 434.700 418.800 438.000 420.000 ;
        RECT 428.100 415.050 429.900 416.850 ;
        RECT 434.100 415.050 435.900 416.850 ;
        RECT 437.100 415.050 438.000 418.800 ;
        RECT 453.000 418.800 456.300 420.000 ;
        RECT 461.100 419.400 462.900 429.000 ;
        RECT 476.100 419.400 477.900 429.000 ;
        RECT 482.700 420.000 484.500 428.400 ;
        RECT 500.400 422.400 502.200 429.000 ;
        RECT 505.500 421.200 507.300 428.400 ;
        RECT 503.100 420.300 507.300 421.200 ;
        RECT 509.550 422.400 511.350 428.400 ;
        RECT 512.850 422.400 514.650 429.000 ;
        RECT 517.950 425.400 519.750 428.400 ;
        RECT 522.450 425.400 524.250 429.000 ;
        RECT 525.450 425.400 527.250 428.400 ;
        RECT 528.750 425.400 530.550 429.000 ;
        RECT 533.250 426.300 535.050 428.400 ;
        RECT 533.250 425.400 536.850 426.300 ;
        RECT 517.350 423.300 519.750 425.400 ;
        RECT 526.200 424.500 527.250 425.400 ;
        RECT 533.250 424.800 537.150 425.400 ;
        RECT 526.200 423.450 531.150 424.500 ;
        RECT 529.350 422.700 531.150 423.450 ;
        RECT 482.700 418.800 486.000 420.000 ;
        RECT 453.000 415.050 453.900 418.800 ;
        RECT 455.100 415.050 456.900 416.850 ;
        RECT 461.100 415.050 462.900 416.850 ;
        RECT 476.100 415.050 477.900 416.850 ;
        RECT 482.100 415.050 483.900 416.850 ;
        RECT 485.100 415.050 486.000 418.800 ;
        RECT 500.250 415.050 502.050 416.850 ;
        RECT 503.100 415.050 504.300 420.300 ;
        RECT 506.100 415.050 507.900 416.850 ;
        RECT 509.550 415.050 510.750 422.400 ;
        RECT 532.350 421.800 534.150 423.600 ;
        RECT 535.050 423.300 537.150 424.800 ;
        RECT 538.050 422.400 539.850 429.000 ;
        RECT 541.050 424.200 542.850 428.400 ;
        RECT 541.050 422.400 543.450 424.200 ;
        RECT 522.150 420.000 523.950 420.600 ;
        RECT 533.100 420.000 534.150 421.800 ;
        RECT 522.150 418.800 534.150 420.000 ;
        RECT 343.500 412.950 345.600 415.050 ;
        RECT 346.800 412.950 348.900 415.050 ;
        RECT 361.950 412.950 364.050 415.050 ;
        RECT 364.950 412.950 367.050 415.050 ;
        RECT 367.950 412.950 370.050 415.050 ;
        RECT 382.950 412.950 385.050 415.050 ;
        RECT 385.950 412.950 388.050 415.050 ;
        RECT 400.950 412.950 403.050 415.050 ;
        RECT 403.950 412.950 406.050 415.050 ;
        RECT 406.950 412.950 409.050 415.050 ;
        RECT 409.950 412.950 412.050 415.050 ;
        RECT 427.950 412.950 430.050 415.050 ;
        RECT 430.950 412.950 433.050 415.050 ;
        RECT 433.950 412.950 436.050 415.050 ;
        RECT 436.950 412.950 439.050 415.050 ;
        RECT 451.950 412.950 454.050 415.050 ;
        RECT 454.950 412.950 457.050 415.050 ;
        RECT 457.950 412.950 460.050 415.050 ;
        RECT 460.950 412.950 463.050 415.050 ;
        RECT 475.950 412.950 478.050 415.050 ;
        RECT 478.950 412.950 481.050 415.050 ;
        RECT 481.950 412.950 484.050 415.050 ;
        RECT 484.950 412.950 487.050 415.050 ;
        RECT 499.950 412.950 502.050 415.050 ;
        RECT 502.950 412.950 505.050 415.050 ;
        RECT 505.950 412.950 508.050 415.050 ;
        RECT 509.550 413.250 515.850 415.050 ;
        RECT 509.550 412.950 514.050 413.250 ;
        RECT 343.200 411.150 345.000 412.950 ;
        RECT 347.400 405.600 348.300 412.950 ;
        RECT 338.100 393.000 339.900 399.600 ;
        RECT 341.100 393.600 342.900 399.600 ;
        RECT 344.100 393.000 345.900 405.000 ;
        RECT 347.100 393.600 348.900 405.600 ;
        RECT 365.100 399.600 366.300 412.950 ;
        RECT 383.100 411.150 384.900 412.950 ;
        RECT 386.100 399.600 387.300 412.950 ;
        RECT 404.250 411.150 406.050 412.950 ;
        RECT 388.950 408.450 391.050 409.050 ;
        RECT 406.950 408.450 409.050 409.050 ;
        RECT 388.950 407.550 409.050 408.450 ;
        RECT 388.950 406.950 391.050 407.550 ;
        RECT 406.950 406.950 409.050 407.550 ;
        RECT 410.700 405.600 411.600 412.950 ;
        RECT 431.100 411.150 432.900 412.950 ;
        RECT 401.100 404.700 408.900 405.600 ;
        RECT 362.100 393.000 363.900 399.600 ;
        RECT 365.100 393.600 366.900 399.600 ;
        RECT 368.100 393.000 369.900 399.600 ;
        RECT 383.100 393.000 384.900 399.600 ;
        RECT 386.100 393.600 387.900 399.600 ;
        RECT 401.100 393.600 402.900 404.700 ;
        RECT 404.100 393.000 405.900 403.800 ;
        RECT 407.100 393.600 408.900 404.700 ;
        RECT 410.100 393.600 411.900 405.600 ;
        RECT 437.100 400.800 438.000 412.950 ;
        RECT 431.400 399.900 438.000 400.800 ;
        RECT 431.400 399.600 432.900 399.900 ;
        RECT 428.100 393.000 429.900 399.600 ;
        RECT 431.100 393.600 432.900 399.600 ;
        RECT 437.100 399.600 438.000 399.900 ;
        RECT 453.000 400.800 453.900 412.950 ;
        RECT 458.100 411.150 459.900 412.950 ;
        RECT 479.100 411.150 480.900 412.950 ;
        RECT 485.100 400.800 486.000 412.950 ;
        RECT 453.000 399.900 459.600 400.800 ;
        RECT 453.000 399.600 453.900 399.900 ;
        RECT 434.100 393.000 435.900 399.000 ;
        RECT 437.100 393.600 438.900 399.600 ;
        RECT 439.950 396.450 442.050 397.050 ;
        RECT 448.950 396.450 451.050 397.050 ;
        RECT 439.950 395.550 451.050 396.450 ;
        RECT 439.950 394.950 442.050 395.550 ;
        RECT 448.950 394.950 451.050 395.550 ;
        RECT 452.100 393.600 453.900 399.600 ;
        RECT 458.100 399.600 459.600 399.900 ;
        RECT 479.400 399.900 486.000 400.800 ;
        RECT 479.400 399.600 480.900 399.900 ;
        RECT 455.100 393.000 456.900 399.000 ;
        RECT 458.100 393.600 459.900 399.600 ;
        RECT 461.100 393.000 462.900 399.600 ;
        RECT 476.100 393.000 477.900 399.600 ;
        RECT 479.100 393.600 480.900 399.600 ;
        RECT 485.100 399.600 486.000 399.900 ;
        RECT 503.100 399.600 504.300 412.950 ;
        RECT 509.550 405.600 510.750 412.950 ;
        RECT 511.650 410.100 513.450 410.250 ;
        RECT 517.350 410.100 519.450 410.400 ;
        RECT 511.650 408.900 519.450 410.100 ;
        RECT 511.650 408.450 513.450 408.900 ;
        RECT 517.350 408.300 519.450 408.900 ;
        RECT 522.150 406.200 523.050 418.800 ;
        RECT 533.100 417.600 541.050 418.800 ;
        RECT 533.100 417.000 534.900 417.600 ;
        RECT 536.100 415.800 537.900 416.400 ;
        RECT 529.800 414.600 537.900 415.800 ;
        RECT 539.250 415.050 541.050 417.600 ;
        RECT 529.800 412.950 531.900 414.600 ;
        RECT 538.950 412.950 541.050 415.050 ;
        RECT 531.750 407.700 533.550 408.000 ;
        RECT 542.550 407.700 543.450 422.400 ;
        RECT 557.700 421.200 559.500 428.400 ;
        RECT 562.800 422.400 564.600 429.000 ;
        RECT 557.700 420.300 561.900 421.200 ;
        RECT 557.100 415.050 558.900 416.850 ;
        RECT 560.700 415.050 561.900 420.300 ;
        RECT 562.950 420.450 565.050 421.050 ;
        RECT 574.950 420.450 577.050 421.050 ;
        RECT 562.950 419.550 577.050 420.450 ;
        RECT 581.100 420.600 582.900 428.400 ;
        RECT 585.600 422.400 587.400 429.000 ;
        RECT 588.600 424.200 590.400 428.400 ;
        RECT 605.700 425.400 607.500 429.000 ;
        RECT 588.600 422.400 591.300 424.200 ;
        RECT 608.700 423.600 610.500 428.400 ;
        RECT 587.700 420.600 589.500 421.500 ;
        RECT 581.100 419.700 589.500 420.600 ;
        RECT 562.950 418.950 565.050 419.550 ;
        RECT 574.950 418.950 577.050 419.550 ;
        RECT 562.950 415.050 564.750 416.850 ;
        RECT 581.250 415.050 583.050 416.850 ;
        RECT 556.950 412.950 559.050 415.050 ;
        RECT 559.950 412.950 562.050 415.050 ;
        RECT 562.950 412.950 565.050 415.050 ;
        RECT 581.100 412.950 583.200 415.050 ;
        RECT 531.750 407.100 543.450 407.700 ;
        RECT 482.100 393.000 483.900 399.000 ;
        RECT 485.100 393.600 486.900 399.600 ;
        RECT 500.100 393.000 501.900 399.600 ;
        RECT 503.100 393.600 504.900 399.600 ;
        RECT 506.100 393.000 507.900 399.600 ;
        RECT 509.550 393.600 511.350 405.600 ;
        RECT 512.550 393.000 514.350 405.600 ;
        RECT 518.250 405.300 523.050 406.200 ;
        RECT 525.150 406.500 543.450 407.100 ;
        RECT 525.150 406.200 533.550 406.500 ;
        RECT 518.250 404.400 519.450 405.300 ;
        RECT 516.450 402.600 519.450 404.400 ;
        RECT 520.350 404.100 522.150 404.400 ;
        RECT 525.150 404.100 526.050 406.200 ;
        RECT 542.550 405.600 543.450 406.500 ;
        RECT 520.350 403.200 526.050 404.100 ;
        RECT 526.950 404.700 528.750 405.300 ;
        RECT 526.950 403.500 534.750 404.700 ;
        RECT 520.350 402.600 522.150 403.200 ;
        RECT 532.650 402.600 534.750 403.500 ;
        RECT 517.350 399.600 519.450 401.700 ;
        RECT 523.950 401.550 525.750 402.300 ;
        RECT 528.750 401.550 530.550 402.300 ;
        RECT 523.950 400.500 530.550 401.550 ;
        RECT 517.350 393.600 519.150 399.600 ;
        RECT 521.850 393.000 523.650 399.600 ;
        RECT 524.850 393.600 526.650 400.500 ;
        RECT 527.850 393.000 529.650 399.600 ;
        RECT 532.650 393.600 534.450 402.600 ;
        RECT 538.050 393.000 539.850 405.600 ;
        RECT 541.050 403.800 543.450 405.600 ;
        RECT 541.050 393.600 542.850 403.800 ;
        RECT 560.700 399.600 561.900 412.950 ;
        RECT 562.950 408.450 565.050 409.050 ;
        RECT 577.950 408.450 580.050 409.050 ;
        RECT 562.950 407.550 580.050 408.450 ;
        RECT 562.950 406.950 565.050 407.550 ;
        RECT 577.950 406.950 580.050 407.550 ;
        RECT 584.100 399.600 585.000 419.700 ;
        RECT 590.400 415.050 591.300 422.400 ;
        RECT 605.400 422.400 610.500 423.600 ;
        RECT 613.200 422.400 615.000 429.000 ;
        RECT 605.400 415.050 606.300 422.400 ;
        RECT 631.500 420.000 633.300 428.400 ;
        RECT 630.000 418.800 633.300 420.000 ;
        RECT 638.100 419.400 639.900 429.000 ;
        RECT 653.100 425.400 654.900 429.000 ;
        RECT 656.100 425.400 657.900 428.400 ;
        RECT 607.950 415.050 609.750 416.850 ;
        RECT 614.100 415.050 615.900 416.850 ;
        RECT 630.000 415.050 630.900 418.800 ;
        RECT 632.100 415.050 633.900 416.850 ;
        RECT 638.100 415.050 639.900 416.850 ;
        RECT 656.100 415.050 657.300 425.400 ;
        RECT 671.100 422.400 672.900 428.400 ;
        RECT 671.700 420.300 672.900 422.400 ;
        RECT 674.100 423.300 675.900 428.400 ;
        RECT 677.100 424.200 678.900 429.000 ;
        RECT 680.100 423.300 681.900 428.400 ;
        RECT 674.100 421.950 681.900 423.300 ;
        RECT 695.100 423.300 696.900 428.400 ;
        RECT 698.100 424.200 699.900 429.000 ;
        RECT 701.100 423.300 702.900 428.400 ;
        RECT 695.100 421.950 702.900 423.300 ;
        RECT 704.100 422.400 705.900 428.400 ;
        RECT 719.700 425.400 721.500 429.000 ;
        RECT 722.700 423.600 724.500 428.400 ;
        RECT 719.400 422.400 724.500 423.600 ;
        RECT 727.200 422.400 729.000 429.000 ;
        RECT 743.700 425.400 745.500 429.000 ;
        RECT 746.700 423.600 748.500 428.400 ;
        RECT 743.400 422.400 748.500 423.600 ;
        RECT 751.200 422.400 753.000 429.000 ;
        RECT 682.950 420.450 685.050 421.050 ;
        RECT 688.950 420.450 691.050 421.050 ;
        RECT 671.700 419.400 675.300 420.300 ;
        RECT 671.100 415.050 672.900 416.850 ;
        RECT 674.100 415.050 675.300 419.400 ;
        RECT 682.950 419.550 691.050 420.450 ;
        RECT 704.100 420.300 705.300 422.400 ;
        RECT 682.950 418.950 685.050 419.550 ;
        RECT 688.950 418.950 691.050 419.550 ;
        RECT 701.700 419.400 705.300 420.300 ;
        RECT 677.100 415.050 678.900 416.850 ;
        RECT 698.100 415.050 699.900 416.850 ;
        RECT 701.700 415.050 702.900 419.400 ;
        RECT 706.950 417.450 709.050 421.050 ;
        RECT 706.950 417.000 711.450 417.450 ;
        RECT 704.100 415.050 705.900 416.850 ;
        RECT 707.550 416.550 711.450 417.000 ;
        RECT 586.500 412.950 588.600 415.050 ;
        RECT 589.800 412.950 591.900 415.050 ;
        RECT 604.950 412.950 607.050 415.050 ;
        RECT 607.950 412.950 610.050 415.050 ;
        RECT 610.950 412.950 613.050 415.050 ;
        RECT 613.950 412.950 616.050 415.050 ;
        RECT 628.950 412.950 631.050 415.050 ;
        RECT 631.950 412.950 634.050 415.050 ;
        RECT 634.950 412.950 637.050 415.050 ;
        RECT 637.950 412.950 640.050 415.050 ;
        RECT 652.950 412.950 655.050 415.050 ;
        RECT 655.950 412.950 658.050 415.050 ;
        RECT 670.950 412.950 673.050 415.050 ;
        RECT 673.950 412.950 676.050 415.050 ;
        RECT 676.950 412.950 679.050 415.050 ;
        RECT 679.950 412.950 682.050 415.050 ;
        RECT 694.950 412.950 697.050 415.050 ;
        RECT 697.950 412.950 700.050 415.050 ;
        RECT 700.950 412.950 703.050 415.050 ;
        RECT 703.950 412.950 706.050 415.050 ;
        RECT 586.200 411.150 588.000 412.950 ;
        RECT 590.400 405.600 591.300 412.950 ;
        RECT 605.400 405.600 606.300 412.950 ;
        RECT 610.950 411.150 612.750 412.950 ;
        RECT 557.100 393.000 558.900 399.600 ;
        RECT 560.100 393.600 561.900 399.600 ;
        RECT 563.100 393.000 564.900 399.600 ;
        RECT 581.100 393.000 582.900 399.600 ;
        RECT 584.100 393.600 585.900 399.600 ;
        RECT 587.100 393.000 588.900 405.000 ;
        RECT 590.100 393.600 591.900 405.600 ;
        RECT 605.100 393.600 606.900 405.600 ;
        RECT 608.100 404.700 615.900 405.600 ;
        RECT 608.100 393.600 609.900 404.700 ;
        RECT 611.100 393.000 612.900 403.800 ;
        RECT 614.100 393.600 615.900 404.700 ;
        RECT 630.000 400.800 630.900 412.950 ;
        RECT 635.100 411.150 636.900 412.950 ;
        RECT 653.100 411.150 654.900 412.950 ;
        RECT 630.000 399.900 636.600 400.800 ;
        RECT 630.000 399.600 630.900 399.900 ;
        RECT 629.100 393.600 630.900 399.600 ;
        RECT 635.100 399.600 636.600 399.900 ;
        RECT 656.100 399.600 657.300 412.950 ;
        RECT 674.100 405.600 675.300 412.950 ;
        RECT 680.100 411.150 681.900 412.950 ;
        RECT 695.100 411.150 696.900 412.950 ;
        RECT 676.950 408.450 679.050 409.050 ;
        RECT 697.950 408.450 700.050 409.050 ;
        RECT 676.950 407.550 700.050 408.450 ;
        RECT 676.950 406.950 679.050 407.550 ;
        RECT 697.950 406.950 700.050 407.550 ;
        RECT 701.700 405.600 702.900 412.950 ;
        RECT 710.550 412.050 711.450 416.550 ;
        RECT 719.400 415.050 720.300 422.400 ;
        RECT 721.950 415.050 723.750 416.850 ;
        RECT 728.100 415.050 729.900 416.850 ;
        RECT 743.400 415.050 744.300 422.400 ;
        RECT 767.100 419.400 768.900 429.000 ;
        RECT 773.700 420.000 775.500 428.400 ;
        RECT 791.100 425.400 792.900 428.400 ;
        RECT 794.100 425.400 795.900 429.000 ;
        RECT 773.700 418.800 777.000 420.000 ;
        RECT 745.950 415.050 747.750 416.850 ;
        RECT 752.100 415.050 753.900 416.850 ;
        RECT 767.100 415.050 768.900 416.850 ;
        RECT 773.100 415.050 774.900 416.850 ;
        RECT 776.100 415.050 777.000 418.800 ;
        RECT 791.700 415.050 792.900 425.400 ;
        RECT 811.500 420.000 813.300 428.400 ;
        RECT 810.000 418.800 813.300 420.000 ;
        RECT 818.100 419.400 819.900 429.000 ;
        RECT 834.000 422.400 835.800 429.000 ;
        RECT 838.500 423.600 840.300 428.400 ;
        RECT 841.500 425.400 843.300 429.000 ;
        RECT 838.500 422.400 843.600 423.600 ;
        RECT 810.000 415.050 810.900 418.800 ;
        RECT 812.100 415.050 813.900 416.850 ;
        RECT 818.100 415.050 819.900 416.850 ;
        RECT 833.100 415.050 834.900 416.850 ;
        RECT 839.250 415.050 841.050 416.850 ;
        RECT 842.700 415.050 843.600 422.400 ;
        RECT 857.100 419.400 858.900 429.000 ;
        RECT 863.700 420.000 865.500 428.400 ;
        RECT 881.100 425.400 882.900 429.000 ;
        RECT 884.100 425.400 885.900 428.400 ;
        RECT 863.700 418.800 867.000 420.000 ;
        RECT 857.100 415.050 858.900 416.850 ;
        RECT 863.100 415.050 864.900 416.850 ;
        RECT 866.100 415.050 867.000 418.800 ;
        RECT 884.100 415.050 885.300 425.400 ;
        RECT 718.950 412.950 721.050 415.050 ;
        RECT 721.950 412.950 724.050 415.050 ;
        RECT 724.950 412.950 727.050 415.050 ;
        RECT 727.950 412.950 730.050 415.050 ;
        RECT 742.950 412.950 745.050 415.050 ;
        RECT 745.950 412.950 748.050 415.050 ;
        RECT 748.950 412.950 751.050 415.050 ;
        RECT 751.950 412.950 754.050 415.050 ;
        RECT 766.950 412.950 769.050 415.050 ;
        RECT 769.950 412.950 772.050 415.050 ;
        RECT 772.950 412.950 775.050 415.050 ;
        RECT 775.950 412.950 778.050 415.050 ;
        RECT 790.950 412.950 793.050 415.050 ;
        RECT 793.950 412.950 796.050 415.050 ;
        RECT 808.950 412.950 811.050 415.050 ;
        RECT 811.950 412.950 814.050 415.050 ;
        RECT 814.950 412.950 817.050 415.050 ;
        RECT 817.950 412.950 820.050 415.050 ;
        RECT 832.950 412.950 835.050 415.050 ;
        RECT 835.950 412.950 838.050 415.050 ;
        RECT 838.950 412.950 841.050 415.050 ;
        RECT 841.950 412.950 844.050 415.050 ;
        RECT 856.950 412.950 859.050 415.050 ;
        RECT 859.950 412.950 862.050 415.050 ;
        RECT 862.950 412.950 865.050 415.050 ;
        RECT 865.950 412.950 868.050 415.050 ;
        RECT 880.950 412.950 883.050 415.050 ;
        RECT 883.950 412.950 886.050 415.050 ;
        RECT 706.950 410.550 711.450 412.050 ;
        RECT 706.950 409.950 711.000 410.550 ;
        RECT 719.400 405.600 720.300 412.950 ;
        RECT 724.950 411.150 726.750 412.950 ;
        RECT 743.400 405.600 744.300 412.950 ;
        RECT 748.950 411.150 750.750 412.950 ;
        RECT 770.100 411.150 771.900 412.950 ;
        RECT 745.950 408.450 748.050 409.050 ;
        RECT 766.950 408.450 769.050 409.050 ;
        RECT 745.950 407.550 769.050 408.450 ;
        RECT 745.950 406.950 748.050 407.550 ;
        RECT 766.950 406.950 769.050 407.550 ;
        RECT 674.100 404.100 676.500 405.600 ;
        RECT 672.000 401.100 673.800 402.900 ;
        RECT 632.100 393.000 633.900 399.000 ;
        RECT 635.100 393.600 636.900 399.600 ;
        RECT 638.100 393.000 639.900 399.600 ;
        RECT 653.100 393.000 654.900 399.600 ;
        RECT 656.100 393.600 657.900 399.600 ;
        RECT 671.700 393.000 673.500 399.600 ;
        RECT 674.700 393.600 676.500 404.100 ;
        RECT 679.800 393.000 681.600 405.600 ;
        RECT 695.400 393.000 697.200 405.600 ;
        RECT 700.500 404.100 702.900 405.600 ;
        RECT 700.500 393.600 702.300 404.100 ;
        RECT 703.200 401.100 705.000 402.900 ;
        RECT 703.500 393.000 705.300 399.600 ;
        RECT 719.100 393.600 720.900 405.600 ;
        RECT 722.100 404.700 729.900 405.600 ;
        RECT 722.100 393.600 723.900 404.700 ;
        RECT 725.100 393.000 726.900 403.800 ;
        RECT 728.100 393.600 729.900 404.700 ;
        RECT 743.100 393.600 744.900 405.600 ;
        RECT 746.100 404.700 753.900 405.600 ;
        RECT 746.100 393.600 747.900 404.700 ;
        RECT 749.100 393.000 750.900 403.800 ;
        RECT 752.100 393.600 753.900 404.700 ;
        RECT 776.100 400.800 777.000 412.950 ;
        RECT 770.400 399.900 777.000 400.800 ;
        RECT 770.400 399.600 771.900 399.900 ;
        RECT 767.100 393.000 768.900 399.600 ;
        RECT 770.100 393.600 771.900 399.600 ;
        RECT 776.100 399.600 777.000 399.900 ;
        RECT 791.700 399.600 792.900 412.950 ;
        RECT 794.100 411.150 795.900 412.950 ;
        RECT 810.000 400.800 810.900 412.950 ;
        RECT 815.100 411.150 816.900 412.950 ;
        RECT 836.250 411.150 838.050 412.950 ;
        RECT 842.700 405.600 843.600 412.950 ;
        RECT 860.100 411.150 861.900 412.950 ;
        RECT 833.100 404.700 840.900 405.600 ;
        RECT 810.000 399.900 816.600 400.800 ;
        RECT 810.000 399.600 810.900 399.900 ;
        RECT 773.100 393.000 774.900 399.000 ;
        RECT 776.100 393.600 777.900 399.600 ;
        RECT 791.100 393.600 792.900 399.600 ;
        RECT 794.100 393.000 795.900 399.600 ;
        RECT 809.100 393.600 810.900 399.600 ;
        RECT 815.100 399.600 816.600 399.900 ;
        RECT 812.100 393.000 813.900 399.000 ;
        RECT 815.100 393.600 816.900 399.600 ;
        RECT 818.100 393.000 819.900 399.600 ;
        RECT 833.100 393.600 834.900 404.700 ;
        RECT 836.100 393.000 837.900 403.800 ;
        RECT 839.100 393.600 840.900 404.700 ;
        RECT 842.100 393.600 843.900 405.600 ;
        RECT 850.950 405.450 853.050 405.900 ;
        RECT 862.950 405.450 865.050 406.050 ;
        RECT 850.950 404.550 865.050 405.450 ;
        RECT 850.950 403.800 853.050 404.550 ;
        RECT 862.950 403.950 865.050 404.550 ;
        RECT 866.100 400.800 867.000 412.950 ;
        RECT 881.100 411.150 882.900 412.950 ;
        RECT 860.400 399.900 867.000 400.800 ;
        RECT 860.400 399.600 861.900 399.900 ;
        RECT 857.100 393.000 858.900 399.600 ;
        RECT 860.100 393.600 861.900 399.600 ;
        RECT 866.100 399.600 867.000 399.900 ;
        RECT 884.100 399.600 885.300 412.950 ;
        RECT 863.100 393.000 864.900 399.000 ;
        RECT 866.100 393.600 867.900 399.600 ;
        RECT 881.100 393.000 882.900 399.600 ;
        RECT 884.100 393.600 885.900 399.600 ;
        RECT 14.100 377.400 15.900 389.400 ;
        RECT 17.100 379.200 18.900 390.000 ;
        RECT 20.100 383.400 21.900 389.400 ;
        RECT 14.100 370.050 15.300 377.400 ;
        RECT 20.700 376.500 21.900 383.400 ;
        RECT 16.200 375.600 21.900 376.500 ;
        RECT 23.550 377.400 25.350 389.400 ;
        RECT 26.550 377.400 28.350 390.000 ;
        RECT 31.350 383.400 33.150 389.400 ;
        RECT 35.850 383.400 37.650 390.000 ;
        RECT 31.350 381.300 33.450 383.400 ;
        RECT 38.850 382.500 40.650 389.400 ;
        RECT 41.850 383.400 43.650 390.000 ;
        RECT 37.950 381.450 44.550 382.500 ;
        RECT 37.950 380.700 39.750 381.450 ;
        RECT 42.750 380.700 44.550 381.450 ;
        RECT 46.650 380.400 48.450 389.400 ;
        RECT 30.450 378.600 33.450 380.400 ;
        RECT 34.350 379.800 36.150 380.400 ;
        RECT 34.350 378.900 40.050 379.800 ;
        RECT 46.650 379.500 48.750 380.400 ;
        RECT 34.350 378.600 36.150 378.900 ;
        RECT 32.250 377.700 33.450 378.600 ;
        RECT 16.200 374.700 18.000 375.600 ;
        RECT 14.100 367.950 16.200 370.050 ;
        RECT 14.100 360.600 15.300 367.950 ;
        RECT 17.100 363.300 18.000 374.700 ;
        RECT 19.800 370.050 21.600 371.850 ;
        RECT 19.500 367.950 21.600 370.050 ;
        RECT 23.550 370.050 24.750 377.400 ;
        RECT 32.250 376.800 37.050 377.700 ;
        RECT 25.650 374.100 27.450 374.550 ;
        RECT 31.350 374.100 33.450 374.700 ;
        RECT 25.650 372.900 33.450 374.100 ;
        RECT 25.650 372.750 27.450 372.900 ;
        RECT 31.350 372.600 33.450 372.900 ;
        RECT 23.550 369.750 28.050 370.050 ;
        RECT 23.550 367.950 29.850 369.750 ;
        RECT 16.200 362.400 18.000 363.300 ;
        RECT 16.200 361.500 21.900 362.400 ;
        RECT 14.100 354.600 15.900 360.600 ;
        RECT 17.100 354.000 18.900 360.600 ;
        RECT 20.700 357.600 21.900 361.500 ;
        RECT 20.100 354.600 21.900 357.600 ;
        RECT 23.550 360.600 24.750 367.950 ;
        RECT 36.150 364.200 37.050 376.800 ;
        RECT 39.150 376.800 40.050 378.900 ;
        RECT 40.950 378.300 48.750 379.500 ;
        RECT 40.950 377.700 42.750 378.300 ;
        RECT 52.050 377.400 53.850 390.000 ;
        RECT 55.050 379.200 56.850 389.400 ;
        RECT 55.050 377.400 57.450 379.200 ;
        RECT 39.150 376.500 47.550 376.800 ;
        RECT 56.550 376.500 57.450 377.400 ;
        RECT 39.150 375.900 57.450 376.500 ;
        RECT 45.750 375.300 57.450 375.900 ;
        RECT 45.750 375.000 47.550 375.300 ;
        RECT 43.800 368.400 45.900 370.050 ;
        RECT 43.800 367.200 51.900 368.400 ;
        RECT 52.950 367.950 55.050 370.050 ;
        RECT 50.100 366.600 51.900 367.200 ;
        RECT 47.100 365.400 48.900 366.000 ;
        RECT 53.250 365.400 55.050 367.950 ;
        RECT 47.100 364.200 55.050 365.400 ;
        RECT 36.150 363.000 48.150 364.200 ;
        RECT 36.150 362.400 37.950 363.000 ;
        RECT 47.100 361.200 48.150 363.000 ;
        RECT 23.550 354.600 25.350 360.600 ;
        RECT 26.850 354.000 28.650 360.600 ;
        RECT 31.350 357.600 33.750 359.700 ;
        RECT 43.350 359.550 45.150 360.300 ;
        RECT 40.200 358.500 45.150 359.550 ;
        RECT 46.350 359.400 48.150 361.200 ;
        RECT 56.550 360.600 57.450 375.300 ;
        RECT 40.200 357.600 41.250 358.500 ;
        RECT 49.050 358.200 51.150 359.700 ;
        RECT 47.250 357.600 51.150 358.200 ;
        RECT 31.950 354.600 33.750 357.600 ;
        RECT 36.450 354.000 38.250 357.600 ;
        RECT 39.450 354.600 41.250 357.600 ;
        RECT 42.750 354.000 44.550 357.600 ;
        RECT 47.250 356.700 50.850 357.600 ;
        RECT 47.250 354.600 49.050 356.700 ;
        RECT 52.050 354.000 53.850 360.600 ;
        RECT 55.050 358.800 57.450 360.600 ;
        RECT 59.550 377.400 61.350 389.400 ;
        RECT 62.550 377.400 64.350 390.000 ;
        RECT 67.350 383.400 69.150 389.400 ;
        RECT 71.850 383.400 73.650 390.000 ;
        RECT 67.350 381.300 69.450 383.400 ;
        RECT 74.850 382.500 76.650 389.400 ;
        RECT 77.850 383.400 79.650 390.000 ;
        RECT 73.950 381.450 80.550 382.500 ;
        RECT 73.950 380.700 75.750 381.450 ;
        RECT 78.750 380.700 80.550 381.450 ;
        RECT 82.650 380.400 84.450 389.400 ;
        RECT 66.450 378.600 69.450 380.400 ;
        RECT 70.350 379.800 72.150 380.400 ;
        RECT 70.350 378.900 76.050 379.800 ;
        RECT 82.650 379.500 84.750 380.400 ;
        RECT 70.350 378.600 72.150 378.900 ;
        RECT 68.250 377.700 69.450 378.600 ;
        RECT 59.550 370.050 60.750 377.400 ;
        RECT 68.250 376.800 73.050 377.700 ;
        RECT 61.650 374.100 63.450 374.550 ;
        RECT 67.350 374.100 69.450 374.700 ;
        RECT 61.650 372.900 69.450 374.100 ;
        RECT 61.650 372.750 63.450 372.900 ;
        RECT 67.350 372.600 69.450 372.900 ;
        RECT 59.550 369.750 64.050 370.050 ;
        RECT 59.550 367.950 65.850 369.750 ;
        RECT 59.550 360.600 60.750 367.950 ;
        RECT 72.150 364.200 73.050 376.800 ;
        RECT 75.150 376.800 76.050 378.900 ;
        RECT 76.950 378.300 84.750 379.500 ;
        RECT 76.950 377.700 78.750 378.300 ;
        RECT 88.050 377.400 89.850 390.000 ;
        RECT 91.050 379.200 92.850 389.400 ;
        RECT 107.100 383.400 108.900 390.000 ;
        RECT 110.100 383.400 111.900 389.400 ;
        RECT 113.100 383.400 114.900 390.000 ;
        RECT 91.050 377.400 93.450 379.200 ;
        RECT 75.150 376.500 83.550 376.800 ;
        RECT 92.550 376.500 93.450 377.400 ;
        RECT 75.150 375.900 93.450 376.500 ;
        RECT 81.750 375.300 93.450 375.900 ;
        RECT 81.750 375.000 83.550 375.300 ;
        RECT 79.800 368.400 81.900 370.050 ;
        RECT 79.800 367.200 87.900 368.400 ;
        RECT 88.950 367.950 91.050 370.050 ;
        RECT 86.100 366.600 87.900 367.200 ;
        RECT 83.100 365.400 84.900 366.000 ;
        RECT 89.250 365.400 91.050 367.950 ;
        RECT 83.100 364.200 91.050 365.400 ;
        RECT 72.150 363.000 84.150 364.200 ;
        RECT 72.150 362.400 73.950 363.000 ;
        RECT 83.100 361.200 84.150 363.000 ;
        RECT 55.050 354.600 56.850 358.800 ;
        RECT 59.550 354.600 61.350 360.600 ;
        RECT 62.850 354.000 64.650 360.600 ;
        RECT 67.350 357.600 69.750 359.700 ;
        RECT 79.350 359.550 81.150 360.300 ;
        RECT 76.200 358.500 81.150 359.550 ;
        RECT 82.350 359.400 84.150 361.200 ;
        RECT 92.550 360.600 93.450 375.300 ;
        RECT 110.100 370.050 111.300 383.400 ;
        RECT 128.100 377.400 129.900 390.000 ;
        RECT 132.600 377.400 135.900 389.400 ;
        RECT 138.600 377.400 140.400 390.000 ;
        RECT 155.100 383.400 156.900 390.000 ;
        RECT 158.100 383.400 159.900 389.400 ;
        RECT 161.100 383.400 162.900 390.000 ;
        RECT 176.100 383.400 177.900 390.000 ;
        RECT 179.100 383.400 180.900 389.400 ;
        RECT 128.100 370.050 129.900 371.850 ;
        RECT 133.950 370.050 135.000 377.400 ;
        RECT 139.950 370.050 141.750 371.850 ;
        RECT 158.100 370.050 159.300 383.400 ;
        RECT 176.100 370.050 177.900 371.850 ;
        RECT 179.100 370.050 180.300 383.400 ;
        RECT 194.400 377.400 196.200 390.000 ;
        RECT 199.500 378.900 201.300 389.400 ;
        RECT 202.500 383.400 204.300 390.000 ;
        RECT 218.100 383.400 219.900 390.000 ;
        RECT 221.100 383.400 222.900 389.400 ;
        RECT 224.100 383.400 225.900 390.000 ;
        RECT 239.100 383.400 240.900 390.000 ;
        RECT 242.100 383.400 243.900 389.400 ;
        RECT 245.100 383.400 246.900 390.000 ;
        RECT 260.100 388.500 267.900 389.400 ;
        RECT 202.200 380.100 204.000 381.900 ;
        RECT 199.500 377.400 201.900 378.900 ;
        RECT 194.100 370.050 195.900 371.850 ;
        RECT 200.700 370.050 201.900 377.400 ;
        RECT 221.100 370.050 222.300 383.400 ;
        RECT 242.100 370.050 243.300 383.400 ;
        RECT 260.100 377.400 261.900 388.500 ;
        RECT 263.100 376.500 264.900 387.600 ;
        RECT 266.100 378.600 267.900 388.500 ;
        RECT 269.100 379.500 270.900 390.000 ;
        RECT 272.100 378.600 273.900 389.400 ;
        RECT 287.100 383.400 288.900 390.000 ;
        RECT 290.100 383.400 291.900 389.400 ;
        RECT 266.100 377.700 273.900 378.600 ;
        RECT 263.100 375.600 267.900 376.500 ;
        RECT 263.100 370.050 264.900 371.850 ;
        RECT 267.000 370.050 267.900 375.600 ;
        RECT 268.950 370.050 270.750 371.850 ;
        RECT 106.950 367.950 109.050 370.050 ;
        RECT 109.950 367.950 112.050 370.050 ;
        RECT 112.950 367.950 115.050 370.050 ;
        RECT 127.950 367.950 130.050 370.050 ;
        RECT 130.950 367.950 133.050 370.050 ;
        RECT 107.250 366.150 109.050 367.950 ;
        RECT 110.100 362.700 111.300 367.950 ;
        RECT 113.100 366.150 114.900 367.950 ;
        RECT 131.250 366.150 133.050 367.950 ;
        RECT 133.950 367.950 136.050 370.050 ;
        RECT 136.950 367.950 139.050 370.050 ;
        RECT 139.950 367.950 142.050 370.050 ;
        RECT 154.950 367.950 157.050 370.050 ;
        RECT 157.950 367.950 160.050 370.050 ;
        RECT 160.950 367.950 163.050 370.050 ;
        RECT 175.950 367.950 178.050 370.050 ;
        RECT 178.950 367.950 181.050 370.050 ;
        RECT 193.950 367.950 196.050 370.050 ;
        RECT 196.950 367.950 199.050 370.050 ;
        RECT 199.950 367.950 202.050 370.050 ;
        RECT 202.950 367.950 205.050 370.050 ;
        RECT 217.950 367.950 220.050 370.050 ;
        RECT 220.950 367.950 223.050 370.050 ;
        RECT 223.950 367.950 226.050 370.050 ;
        RECT 238.950 367.950 241.050 370.050 ;
        RECT 241.950 367.950 244.050 370.050 ;
        RECT 244.950 367.950 247.050 370.050 ;
        RECT 259.950 367.950 262.050 370.050 ;
        RECT 262.950 367.950 265.050 370.050 ;
        RECT 265.950 367.950 268.050 370.050 ;
        RECT 268.950 367.950 271.050 370.050 ;
        RECT 271.950 367.950 274.050 370.050 ;
        RECT 287.100 367.950 289.200 370.050 ;
        RECT 133.950 363.300 135.000 367.950 ;
        RECT 136.950 366.150 138.750 367.950 ;
        RECT 155.250 366.150 157.050 367.950 ;
        RECT 110.100 361.800 114.300 362.700 ;
        RECT 133.950 362.100 138.300 363.300 ;
        RECT 76.200 357.600 77.250 358.500 ;
        RECT 85.050 358.200 87.150 359.700 ;
        RECT 83.250 357.600 87.150 358.200 ;
        RECT 67.950 354.600 69.750 357.600 ;
        RECT 72.450 354.000 74.250 357.600 ;
        RECT 75.450 354.600 77.250 357.600 ;
        RECT 78.750 354.000 80.550 357.600 ;
        RECT 83.250 356.700 86.850 357.600 ;
        RECT 83.250 354.600 85.050 356.700 ;
        RECT 88.050 354.000 89.850 360.600 ;
        RECT 91.050 358.800 93.450 360.600 ;
        RECT 91.050 354.600 92.850 358.800 ;
        RECT 107.400 354.000 109.200 360.600 ;
        RECT 112.500 354.600 114.300 361.800 ;
        RECT 128.100 360.000 135.900 360.900 ;
        RECT 137.400 360.600 138.300 362.100 ;
        RECT 158.100 362.700 159.300 367.950 ;
        RECT 161.100 366.150 162.900 367.950 ;
        RECT 158.100 361.800 162.300 362.700 ;
        RECT 128.100 354.600 129.900 360.000 ;
        RECT 131.100 354.000 132.900 359.100 ;
        RECT 134.100 355.500 135.900 360.000 ;
        RECT 137.100 356.400 138.900 360.600 ;
        RECT 140.100 355.500 141.900 360.600 ;
        RECT 134.100 354.600 141.900 355.500 ;
        RECT 155.400 354.000 157.200 360.600 ;
        RECT 160.500 354.600 162.300 361.800 ;
        RECT 179.100 357.600 180.300 367.950 ;
        RECT 197.100 366.150 198.900 367.950 ;
        RECT 200.700 363.600 201.900 367.950 ;
        RECT 203.100 366.150 204.900 367.950 ;
        RECT 218.250 366.150 220.050 367.950 ;
        RECT 200.700 362.700 204.300 363.600 ;
        RECT 194.100 359.700 201.900 361.050 ;
        RECT 176.100 354.000 177.900 357.600 ;
        RECT 179.100 354.600 180.900 357.600 ;
        RECT 194.100 354.600 195.900 359.700 ;
        RECT 197.100 354.000 198.900 358.800 ;
        RECT 200.100 354.600 201.900 359.700 ;
        RECT 203.100 360.600 204.300 362.700 ;
        RECT 221.100 362.700 222.300 367.950 ;
        RECT 224.100 366.150 225.900 367.950 ;
        RECT 239.250 366.150 241.050 367.950 ;
        RECT 242.100 362.700 243.300 367.950 ;
        RECT 245.100 366.150 246.900 367.950 ;
        RECT 260.100 366.150 261.900 367.950 ;
        RECT 221.100 361.800 225.300 362.700 ;
        RECT 242.100 361.800 246.300 362.700 ;
        RECT 203.100 354.600 204.900 360.600 ;
        RECT 218.400 354.000 220.200 360.600 ;
        RECT 223.500 354.600 225.300 361.800 ;
        RECT 239.400 354.000 241.200 360.600 ;
        RECT 244.500 354.600 246.300 361.800 ;
        RECT 266.700 360.600 267.900 367.950 ;
        RECT 271.950 366.150 273.750 367.950 ;
        RECT 287.250 366.150 289.050 367.950 ;
        RECT 290.100 363.300 291.000 383.400 ;
        RECT 293.100 378.000 294.900 390.000 ;
        RECT 296.100 377.400 297.900 389.400 ;
        RECT 311.100 383.400 312.900 390.000 ;
        RECT 314.100 383.400 315.900 389.400 ;
        RECT 317.100 383.400 318.900 390.000 ;
        RECT 332.100 383.400 333.900 390.000 ;
        RECT 335.100 383.400 336.900 389.400 ;
        RECT 338.100 383.400 339.900 390.000 ;
        RECT 353.100 383.400 354.900 390.000 ;
        RECT 356.100 383.400 357.900 389.400 ;
        RECT 359.100 383.400 360.900 390.000 ;
        RECT 292.200 370.050 294.000 371.850 ;
        RECT 296.400 370.050 297.300 377.400 ;
        RECT 304.950 375.450 307.050 376.050 ;
        RECT 310.950 375.450 313.050 376.050 ;
        RECT 304.950 374.550 313.050 375.450 ;
        RECT 304.950 373.950 307.050 374.550 ;
        RECT 310.950 373.950 313.050 374.550 ;
        RECT 314.100 370.050 315.300 383.400 ;
        RECT 335.700 370.050 336.900 383.400 ;
        RECT 356.700 370.050 357.900 383.400 ;
        RECT 374.100 377.400 375.900 389.400 ;
        RECT 377.100 378.000 378.900 390.000 ;
        RECT 380.100 383.400 381.900 389.400 ;
        RECT 383.100 383.400 384.900 390.000 ;
        RECT 398.100 383.400 399.900 390.000 ;
        RECT 401.100 383.400 402.900 389.400 ;
        RECT 404.100 383.400 405.900 390.000 ;
        RECT 374.700 370.050 375.600 377.400 ;
        RECT 378.000 370.050 379.800 371.850 ;
        RECT 292.500 367.950 294.600 370.050 ;
        RECT 295.800 367.950 297.900 370.050 ;
        RECT 310.950 367.950 313.050 370.050 ;
        RECT 313.950 367.950 316.050 370.050 ;
        RECT 316.950 367.950 319.050 370.050 ;
        RECT 331.950 367.950 334.050 370.050 ;
        RECT 334.950 367.950 337.050 370.050 ;
        RECT 337.950 367.950 340.050 370.050 ;
        RECT 352.950 367.950 355.050 370.050 ;
        RECT 355.950 367.950 358.050 370.050 ;
        RECT 358.950 367.950 361.050 370.050 ;
        RECT 374.100 367.950 376.200 370.050 ;
        RECT 377.400 367.950 379.500 370.050 ;
        RECT 287.100 362.400 295.500 363.300 ;
        RECT 262.500 354.000 264.300 360.600 ;
        RECT 267.000 354.600 268.800 360.600 ;
        RECT 271.500 354.000 273.300 360.600 ;
        RECT 287.100 354.600 288.900 362.400 ;
        RECT 293.700 361.500 295.500 362.400 ;
        RECT 296.400 360.600 297.300 367.950 ;
        RECT 311.250 366.150 313.050 367.950 ;
        RECT 314.100 362.700 315.300 367.950 ;
        RECT 317.100 366.150 318.900 367.950 ;
        RECT 332.100 366.150 333.900 367.950 ;
        RECT 335.700 362.700 336.900 367.950 ;
        RECT 337.950 366.150 339.750 367.950 ;
        RECT 353.100 366.150 354.900 367.950 ;
        RECT 356.700 362.700 357.900 367.950 ;
        RECT 358.950 366.150 360.750 367.950 ;
        RECT 314.100 361.800 318.300 362.700 ;
        RECT 291.600 354.000 293.400 360.600 ;
        RECT 294.600 358.800 297.300 360.600 ;
        RECT 294.600 354.600 296.400 358.800 ;
        RECT 311.400 354.000 313.200 360.600 ;
        RECT 316.500 354.600 318.300 361.800 ;
        RECT 332.700 361.800 336.900 362.700 ;
        RECT 353.700 361.800 357.900 362.700 ;
        RECT 332.700 354.600 334.500 361.800 ;
        RECT 337.800 354.000 339.600 360.600 ;
        RECT 353.700 354.600 355.500 361.800 ;
        RECT 374.700 360.600 375.600 367.950 ;
        RECT 381.000 363.300 381.900 383.400 ;
        RECT 401.700 370.050 402.900 383.400 ;
        RECT 419.100 377.400 420.900 389.400 ;
        RECT 422.100 379.200 423.900 390.000 ;
        RECT 425.100 383.400 426.900 389.400 ;
        RECT 419.100 370.050 420.300 377.400 ;
        RECT 425.700 376.500 426.900 383.400 ;
        RECT 440.400 377.400 442.200 390.000 ;
        RECT 445.500 378.900 447.300 389.400 ;
        RECT 448.500 383.400 450.300 390.000 ;
        RECT 464.100 383.400 465.900 390.000 ;
        RECT 467.100 383.400 468.900 389.400 ;
        RECT 448.200 380.100 450.000 381.900 ;
        RECT 445.500 377.400 447.900 378.900 ;
        RECT 421.200 375.600 426.900 376.500 ;
        RECT 421.200 374.700 423.000 375.600 ;
        RECT 382.800 367.950 384.900 370.050 ;
        RECT 397.950 367.950 400.050 370.050 ;
        RECT 400.950 367.950 403.050 370.050 ;
        RECT 403.950 367.950 406.050 370.050 ;
        RECT 419.100 367.950 421.200 370.050 ;
        RECT 382.950 366.150 384.750 367.950 ;
        RECT 398.100 366.150 399.900 367.950 ;
        RECT 376.500 362.400 384.900 363.300 ;
        RECT 401.700 362.700 402.900 367.950 ;
        RECT 403.950 366.150 405.750 367.950 ;
        RECT 376.500 361.500 378.300 362.400 ;
        RECT 358.800 354.000 360.600 360.600 ;
        RECT 374.700 358.800 377.400 360.600 ;
        RECT 375.600 354.600 377.400 358.800 ;
        RECT 378.600 354.000 380.400 360.600 ;
        RECT 383.100 354.600 384.900 362.400 ;
        RECT 398.700 361.800 402.900 362.700 ;
        RECT 398.700 354.600 400.500 361.800 ;
        RECT 419.100 360.600 420.300 367.950 ;
        RECT 422.100 363.300 423.000 374.700 ;
        RECT 424.800 370.050 426.600 371.850 ;
        RECT 440.100 370.050 441.900 371.850 ;
        RECT 446.700 370.050 447.900 377.400 ;
        RECT 448.950 375.450 451.050 376.050 ;
        RECT 463.950 375.450 466.050 376.050 ;
        RECT 448.950 374.550 466.050 375.450 ;
        RECT 448.950 373.950 451.050 374.550 ;
        RECT 463.950 373.950 466.050 374.550 ;
        RECT 424.500 367.950 426.600 370.050 ;
        RECT 439.950 367.950 442.050 370.050 ;
        RECT 442.950 367.950 445.050 370.050 ;
        RECT 445.950 367.950 448.050 370.050 ;
        RECT 448.950 367.950 451.050 370.050 ;
        RECT 464.100 367.950 466.200 370.050 ;
        RECT 443.100 366.150 444.900 367.950 ;
        RECT 421.200 362.400 423.000 363.300 ;
        RECT 446.700 363.600 447.900 367.950 ;
        RECT 449.100 366.150 450.900 367.950 ;
        RECT 464.250 366.150 466.050 367.950 ;
        RECT 446.700 362.700 450.300 363.600 ;
        RECT 467.100 363.300 468.000 383.400 ;
        RECT 470.100 378.000 471.900 390.000 ;
        RECT 473.100 377.400 474.900 389.400 ;
        RECT 488.100 378.600 489.900 389.400 ;
        RECT 491.100 379.500 493.200 390.000 ;
        RECT 488.100 377.400 493.200 378.600 ;
        RECT 495.600 378.300 497.400 389.400 ;
        RECT 500.100 379.500 501.900 390.000 ;
        RECT 503.100 378.300 504.900 389.400 ;
        RECT 518.100 383.400 519.900 390.000 ;
        RECT 521.100 383.400 522.900 389.400 ;
        RECT 524.100 384.000 525.900 390.000 ;
        RECT 521.400 383.100 522.900 383.400 ;
        RECT 527.100 383.400 528.900 389.400 ;
        RECT 527.100 383.100 528.000 383.400 ;
        RECT 521.400 382.200 528.000 383.100 ;
        RECT 469.200 370.050 471.000 371.850 ;
        RECT 473.400 370.050 474.300 377.400 ;
        RECT 491.100 376.500 493.200 377.400 ;
        RECT 494.100 377.400 497.400 378.300 ;
        RECT 494.100 373.050 495.300 377.400 ;
        RECT 500.100 377.100 504.900 378.300 ;
        RECT 500.100 376.200 502.200 377.100 ;
        RECT 496.800 375.300 502.200 376.200 ;
        RECT 505.950 375.450 508.050 376.050 ;
        RECT 520.950 375.450 523.050 376.050 ;
        RECT 496.800 373.500 498.600 375.300 ;
        RECT 505.950 374.550 523.050 375.450 ;
        RECT 505.950 373.950 508.050 374.550 ;
        RECT 520.950 373.950 523.050 374.550 ;
        RECT 493.800 372.300 495.900 373.050 ;
        RECT 488.400 370.050 490.200 371.850 ;
        RECT 493.800 370.950 496.800 372.300 ;
        RECT 469.500 367.950 471.600 370.050 ;
        RECT 472.800 367.950 474.900 370.050 ;
        RECT 488.100 367.950 490.200 370.050 ;
        RECT 493.200 368.100 495.000 369.900 ;
        RECT 421.200 361.500 426.900 362.400 ;
        RECT 403.800 354.000 405.600 360.600 ;
        RECT 419.100 354.600 420.900 360.600 ;
        RECT 422.100 354.000 423.900 360.600 ;
        RECT 425.700 357.600 426.900 361.500 ;
        RECT 425.100 354.600 426.900 357.600 ;
        RECT 440.100 359.700 447.900 361.050 ;
        RECT 440.100 354.600 441.900 359.700 ;
        RECT 443.100 354.000 444.900 358.800 ;
        RECT 446.100 354.600 447.900 359.700 ;
        RECT 449.100 360.600 450.300 362.700 ;
        RECT 464.100 362.400 472.500 363.300 ;
        RECT 449.100 354.600 450.900 360.600 ;
        RECT 464.100 354.600 465.900 362.400 ;
        RECT 470.700 361.500 472.500 362.400 ;
        RECT 473.400 360.600 474.300 367.950 ;
        RECT 492.900 366.000 495.000 368.100 ;
        RECT 495.900 364.200 496.800 370.950 ;
        RECT 498.300 370.200 500.100 372.000 ;
        RECT 498.000 368.100 500.100 370.200 ;
        RECT 521.100 370.050 522.900 371.850 ;
        RECT 527.100 370.050 528.000 382.200 ;
        RECT 542.100 378.600 543.900 389.400 ;
        RECT 545.100 379.500 547.200 390.000 ;
        RECT 542.100 377.400 547.200 378.600 ;
        RECT 549.600 378.300 551.400 389.400 ;
        RECT 554.100 379.500 555.900 390.000 ;
        RECT 557.100 378.300 558.900 389.400 ;
        RECT 572.100 383.400 573.900 390.000 ;
        RECT 575.100 383.400 576.900 389.400 ;
        RECT 545.100 376.500 547.200 377.400 ;
        RECT 548.100 377.400 551.400 378.300 ;
        RECT 548.100 373.050 549.300 377.400 ;
        RECT 554.100 377.100 558.900 378.300 ;
        RECT 554.100 376.200 556.200 377.100 ;
        RECT 550.800 375.300 556.200 376.200 ;
        RECT 550.800 373.500 552.600 375.300 ;
        RECT 547.800 372.300 549.900 373.050 ;
        RECT 542.400 370.050 544.200 371.850 ;
        RECT 547.800 370.950 550.800 372.300 ;
        RECT 502.800 367.800 504.900 370.050 ;
        RECT 517.950 367.950 520.050 370.050 ;
        RECT 520.950 367.950 523.050 370.050 ;
        RECT 523.950 367.950 526.050 370.050 ;
        RECT 526.950 367.950 529.050 370.050 ;
        RECT 542.100 367.950 544.200 370.050 ;
        RECT 547.200 368.100 549.000 369.900 ;
        RECT 502.800 367.200 504.600 367.800 ;
        RECT 498.000 366.000 504.600 367.200 ;
        RECT 518.100 366.150 519.900 367.950 ;
        RECT 524.100 366.150 525.900 367.950 ;
        RECT 498.000 365.100 500.100 366.000 ;
        RECT 490.500 361.500 492.600 363.900 ;
        RECT 493.800 362.100 496.800 364.200 ;
        RECT 497.700 363.300 499.500 365.100 ;
        RECT 527.100 364.200 528.000 367.950 ;
        RECT 546.900 366.000 549.000 368.100 ;
        RECT 549.900 364.200 550.800 370.950 ;
        RECT 552.300 370.200 554.100 372.000 ;
        RECT 552.000 368.100 554.100 370.200 ;
        RECT 572.100 370.050 573.900 371.850 ;
        RECT 575.100 370.050 576.300 383.400 ;
        RECT 593.400 377.400 595.200 390.000 ;
        RECT 598.500 378.900 600.300 389.400 ;
        RECT 601.500 383.400 603.300 390.000 ;
        RECT 617.100 383.400 618.900 390.000 ;
        RECT 620.100 383.400 621.900 389.400 ;
        RECT 623.100 383.400 624.900 390.000 ;
        RECT 638.100 383.400 639.900 390.000 ;
        RECT 641.100 383.400 642.900 389.400 ;
        RECT 601.200 380.100 603.000 381.900 ;
        RECT 598.500 377.400 600.900 378.900 ;
        RECT 577.950 375.450 580.050 376.050 ;
        RECT 595.950 375.450 598.050 375.900 ;
        RECT 577.950 374.550 598.050 375.450 ;
        RECT 577.950 373.950 580.050 374.550 ;
        RECT 595.950 373.800 598.050 374.550 ;
        RECT 593.100 370.050 594.900 371.850 ;
        RECT 599.700 370.050 600.900 377.400 ;
        RECT 620.100 370.050 621.300 383.400 ;
        RECT 638.100 370.050 639.900 371.850 ;
        RECT 641.100 370.050 642.300 383.400 ;
        RECT 656.100 378.300 657.900 389.400 ;
        RECT 659.100 379.200 660.900 390.000 ;
        RECT 662.100 378.300 663.900 389.400 ;
        RECT 656.100 377.400 663.900 378.300 ;
        RECT 665.100 377.400 666.900 389.400 ;
        RECT 680.400 377.400 682.200 390.000 ;
        RECT 685.500 378.900 687.300 389.400 ;
        RECT 688.500 383.400 690.300 390.000 ;
        RECT 688.200 380.100 690.000 381.900 ;
        RECT 685.500 377.400 687.900 378.900 ;
        RECT 704.100 377.400 705.900 389.400 ;
        RECT 707.100 378.300 708.900 389.400 ;
        RECT 710.100 379.200 711.900 390.000 ;
        RECT 713.100 378.300 714.900 389.400 ;
        RECT 728.100 383.400 729.900 389.400 ;
        RECT 731.100 384.000 732.900 390.000 ;
        RECT 707.100 377.400 714.900 378.300 ;
        RECT 729.000 383.100 729.900 383.400 ;
        RECT 734.100 383.400 735.900 389.400 ;
        RECT 737.100 383.400 738.900 390.000 ;
        RECT 752.100 383.400 753.900 389.400 ;
        RECT 755.100 384.000 756.900 390.000 ;
        RECT 734.100 383.100 735.600 383.400 ;
        RECT 729.000 382.200 735.600 383.100 ;
        RECT 753.000 383.100 753.900 383.400 ;
        RECT 758.100 383.400 759.900 389.400 ;
        RECT 761.100 383.400 762.900 390.000 ;
        RECT 758.100 383.100 759.600 383.400 ;
        RECT 753.000 382.200 759.600 383.100 ;
        RECT 659.250 370.050 661.050 371.850 ;
        RECT 665.700 370.050 666.600 377.400 ;
        RECT 680.100 370.050 681.900 371.850 ;
        RECT 686.700 370.050 687.900 377.400 ;
        RECT 704.400 370.050 705.300 377.400 ;
        RECT 709.950 370.050 711.750 371.850 ;
        RECT 729.000 370.050 729.900 382.200 ;
        RECT 734.100 370.050 735.900 371.850 ;
        RECT 753.000 370.050 753.900 382.200 ;
        RECT 776.100 378.300 777.900 389.400 ;
        RECT 779.100 379.200 780.900 390.000 ;
        RECT 782.100 378.300 783.900 389.400 ;
        RECT 776.100 377.400 783.900 378.300 ;
        RECT 785.100 377.400 786.900 389.400 ;
        RECT 803.400 377.400 805.200 390.000 ;
        RECT 808.500 378.900 810.300 389.400 ;
        RECT 811.500 383.400 813.300 390.000 ;
        RECT 827.100 383.400 828.900 390.000 ;
        RECT 830.100 383.400 831.900 389.400 ;
        RECT 833.100 383.400 834.900 390.000 ;
        RECT 851.100 383.400 852.900 389.400 ;
        RECT 854.100 383.400 855.900 390.000 ;
        RECT 872.100 383.400 873.900 390.000 ;
        RECT 875.100 383.400 876.900 389.400 ;
        RECT 878.100 383.400 879.900 390.000 ;
        RECT 811.200 380.100 813.000 381.900 ;
        RECT 808.500 377.400 810.900 378.900 ;
        RECT 758.100 370.050 759.900 371.850 ;
        RECT 779.250 370.050 781.050 371.850 ;
        RECT 785.700 370.050 786.600 377.400 ;
        RECT 803.100 370.050 804.900 371.850 ;
        RECT 809.700 370.050 810.900 377.400 ;
        RECT 830.700 370.050 831.900 383.400 ;
        RECT 851.700 370.050 852.900 383.400 ;
        RECT 854.100 370.050 855.900 371.850 ;
        RECT 875.100 370.050 876.300 383.400 ;
        RECT 556.800 367.800 558.900 370.050 ;
        RECT 571.950 367.950 574.050 370.050 ;
        RECT 574.950 367.950 577.050 370.050 ;
        RECT 592.950 367.950 595.050 370.050 ;
        RECT 595.950 367.950 598.050 370.050 ;
        RECT 598.950 367.950 601.050 370.050 ;
        RECT 601.950 367.950 604.050 370.050 ;
        RECT 616.950 367.950 619.050 370.050 ;
        RECT 619.950 367.950 622.050 370.050 ;
        RECT 622.950 367.950 625.050 370.050 ;
        RECT 637.950 367.950 640.050 370.050 ;
        RECT 640.950 367.950 643.050 370.050 ;
        RECT 655.950 367.950 658.050 370.050 ;
        RECT 658.950 367.950 661.050 370.050 ;
        RECT 661.950 367.950 664.050 370.050 ;
        RECT 664.950 367.950 667.050 370.050 ;
        RECT 679.950 367.950 682.050 370.050 ;
        RECT 682.950 367.950 685.050 370.050 ;
        RECT 685.950 367.950 688.050 370.050 ;
        RECT 688.950 367.950 691.050 370.050 ;
        RECT 703.950 367.950 706.050 370.050 ;
        RECT 706.950 367.950 709.050 370.050 ;
        RECT 709.950 367.950 712.050 370.050 ;
        RECT 712.950 367.950 715.050 370.050 ;
        RECT 727.950 367.950 730.050 370.050 ;
        RECT 730.950 367.950 733.050 370.050 ;
        RECT 733.950 367.950 736.050 370.050 ;
        RECT 736.950 367.950 739.050 370.050 ;
        RECT 751.950 367.950 754.050 370.050 ;
        RECT 754.950 367.950 757.050 370.050 ;
        RECT 757.950 367.950 760.050 370.050 ;
        RECT 760.950 367.950 763.050 370.050 ;
        RECT 775.950 367.950 778.050 370.050 ;
        RECT 778.950 367.950 781.050 370.050 ;
        RECT 781.950 367.950 784.050 370.050 ;
        RECT 784.950 367.950 787.050 370.050 ;
        RECT 802.950 367.950 805.050 370.050 ;
        RECT 805.950 367.950 808.050 370.050 ;
        RECT 808.950 367.950 811.050 370.050 ;
        RECT 811.950 367.950 814.050 370.050 ;
        RECT 826.950 367.950 829.050 370.050 ;
        RECT 829.950 367.950 832.050 370.050 ;
        RECT 832.950 367.950 835.050 370.050 ;
        RECT 850.950 367.950 853.050 370.050 ;
        RECT 853.950 367.950 856.050 370.050 ;
        RECT 871.950 367.950 874.050 370.050 ;
        RECT 874.950 367.950 877.050 370.050 ;
        RECT 877.950 367.950 880.050 370.050 ;
        RECT 556.800 367.200 558.600 367.800 ;
        RECT 552.000 366.000 558.600 367.200 ;
        RECT 552.000 365.100 554.100 366.000 ;
        RECT 468.600 354.000 470.400 360.600 ;
        RECT 471.600 358.800 474.300 360.600 ;
        RECT 488.100 360.600 492.600 361.500 ;
        RECT 471.600 354.600 473.400 358.800 ;
        RECT 488.100 354.600 489.900 360.600 ;
        RECT 495.900 360.000 496.800 362.100 ;
        RECT 500.400 363.000 502.500 363.600 ;
        RECT 500.400 361.500 504.900 363.000 ;
        RECT 503.400 360.600 504.900 361.500 ;
        RECT 491.400 354.000 493.200 359.700 ;
        RECT 495.900 354.600 497.700 360.000 ;
        RECT 500.100 354.000 501.900 359.700 ;
        RECT 503.100 354.600 504.900 360.600 ;
        RECT 518.100 354.000 519.900 363.600 ;
        RECT 524.700 363.000 528.000 364.200 ;
        RECT 524.700 354.600 526.500 363.000 ;
        RECT 544.500 361.500 546.600 363.900 ;
        RECT 547.800 362.100 550.800 364.200 ;
        RECT 551.700 363.300 553.500 365.100 ;
        RECT 542.100 360.600 546.600 361.500 ;
        RECT 542.100 354.600 543.900 360.600 ;
        RECT 549.900 360.000 550.800 362.100 ;
        RECT 554.400 363.000 556.500 363.600 ;
        RECT 554.400 361.500 558.900 363.000 ;
        RECT 557.400 360.600 558.900 361.500 ;
        RECT 545.400 354.000 547.200 359.700 ;
        RECT 549.900 354.600 551.700 360.000 ;
        RECT 554.100 354.000 555.900 359.700 ;
        RECT 557.100 354.600 558.900 360.600 ;
        RECT 575.100 357.600 576.300 367.950 ;
        RECT 583.950 366.450 586.050 367.050 ;
        RECT 589.950 366.450 592.050 367.050 ;
        RECT 583.950 365.550 592.050 366.450 ;
        RECT 596.100 366.150 597.900 367.950 ;
        RECT 583.950 364.950 586.050 365.550 ;
        RECT 589.950 364.950 592.050 365.550 ;
        RECT 599.700 363.600 600.900 367.950 ;
        RECT 602.100 366.150 603.900 367.950 ;
        RECT 617.250 366.150 619.050 367.950 ;
        RECT 599.700 362.700 603.300 363.600 ;
        RECT 593.100 359.700 600.900 361.050 ;
        RECT 572.100 354.000 573.900 357.600 ;
        RECT 575.100 354.600 576.900 357.600 ;
        RECT 593.100 354.600 594.900 359.700 ;
        RECT 596.100 354.000 597.900 358.800 ;
        RECT 599.100 354.600 600.900 359.700 ;
        RECT 602.100 360.600 603.300 362.700 ;
        RECT 620.100 362.700 621.300 367.950 ;
        RECT 623.100 366.150 624.900 367.950 ;
        RECT 620.100 361.800 624.300 362.700 ;
        RECT 602.100 354.600 603.900 360.600 ;
        RECT 617.400 354.000 619.200 360.600 ;
        RECT 622.500 354.600 624.300 361.800 ;
        RECT 641.100 357.600 642.300 367.950 ;
        RECT 656.100 366.150 657.900 367.950 ;
        RECT 662.250 366.150 664.050 367.950 ;
        RECT 665.700 360.600 666.600 367.950 ;
        RECT 683.100 366.150 684.900 367.950 ;
        RECT 686.700 363.600 687.900 367.950 ;
        RECT 689.100 366.150 690.900 367.950 ;
        RECT 686.700 362.700 690.300 363.600 ;
        RECT 638.100 354.000 639.900 357.600 ;
        RECT 641.100 354.600 642.900 357.600 ;
        RECT 657.000 354.000 658.800 360.600 ;
        RECT 661.500 359.400 666.600 360.600 ;
        RECT 680.100 359.700 687.900 361.050 ;
        RECT 661.500 354.600 663.300 359.400 ;
        RECT 664.500 354.000 666.300 357.600 ;
        RECT 680.100 354.600 681.900 359.700 ;
        RECT 683.100 354.000 684.900 358.800 ;
        RECT 686.100 354.600 687.900 359.700 ;
        RECT 689.100 360.600 690.300 362.700 ;
        RECT 704.400 360.600 705.300 367.950 ;
        RECT 706.950 366.150 708.750 367.950 ;
        RECT 713.100 366.150 714.900 367.950 ;
        RECT 729.000 364.200 729.900 367.950 ;
        RECT 731.100 366.150 732.900 367.950 ;
        RECT 737.100 366.150 738.900 367.950 ;
        RECT 753.000 364.200 753.900 367.950 ;
        RECT 755.100 366.150 756.900 367.950 ;
        RECT 761.100 366.150 762.900 367.950 ;
        RECT 776.100 366.150 777.900 367.950 ;
        RECT 782.250 366.150 784.050 367.950 ;
        RECT 729.000 363.000 732.300 364.200 ;
        RECT 689.100 354.600 690.900 360.600 ;
        RECT 704.400 359.400 709.500 360.600 ;
        RECT 704.700 354.000 706.500 357.600 ;
        RECT 707.700 354.600 709.500 359.400 ;
        RECT 712.200 354.000 714.000 360.600 ;
        RECT 730.500 354.600 732.300 363.000 ;
        RECT 737.100 354.000 738.900 363.600 ;
        RECT 753.000 363.000 756.300 364.200 ;
        RECT 754.500 354.600 756.300 363.000 ;
        RECT 761.100 354.000 762.900 363.600 ;
        RECT 769.950 363.450 772.050 364.050 ;
        RECT 778.950 363.450 781.050 363.750 ;
        RECT 769.950 362.550 781.050 363.450 ;
        RECT 769.950 361.950 772.050 362.550 ;
        RECT 778.950 361.650 781.050 362.550 ;
        RECT 785.700 360.600 786.600 367.950 ;
        RECT 806.100 366.150 807.900 367.950 ;
        RECT 809.700 363.600 810.900 367.950 ;
        RECT 812.100 366.150 813.900 367.950 ;
        RECT 827.100 366.150 828.900 367.950 ;
        RECT 809.700 362.700 813.300 363.600 ;
        RECT 830.700 362.700 831.900 367.950 ;
        RECT 832.950 366.150 834.750 367.950 ;
        RECT 777.000 354.000 778.800 360.600 ;
        RECT 781.500 359.400 786.600 360.600 ;
        RECT 803.100 359.700 810.900 361.050 ;
        RECT 781.500 354.600 783.300 359.400 ;
        RECT 784.500 354.000 786.300 357.600 ;
        RECT 803.100 354.600 804.900 359.700 ;
        RECT 806.100 354.000 807.900 358.800 ;
        RECT 809.100 354.600 810.900 359.700 ;
        RECT 812.100 360.600 813.300 362.700 ;
        RECT 827.700 361.800 831.900 362.700 ;
        RECT 812.100 354.600 813.900 360.600 ;
        RECT 827.700 354.600 829.500 361.800 ;
        RECT 832.800 354.000 834.600 360.600 ;
        RECT 838.950 357.450 841.050 358.050 ;
        RECT 847.950 357.450 850.050 358.050 ;
        RECT 851.700 357.600 852.900 367.950 ;
        RECT 872.250 366.150 874.050 367.950 ;
        RECT 875.100 362.700 876.300 367.950 ;
        RECT 878.100 366.150 879.900 367.950 ;
        RECT 875.100 361.800 879.300 362.700 ;
        RECT 838.950 356.550 850.050 357.450 ;
        RECT 838.950 355.950 841.050 356.550 ;
        RECT 847.950 355.950 850.050 356.550 ;
        RECT 851.100 354.600 852.900 357.600 ;
        RECT 854.100 354.000 855.900 357.600 ;
        RECT 872.400 354.000 874.200 360.600 ;
        RECT 877.500 354.600 879.300 361.800 ;
        RECT 17.100 344.400 18.900 350.400 ;
        RECT 20.100 344.400 21.900 351.000 ;
        RECT 23.100 347.400 24.900 350.400 ;
        RECT 17.100 337.050 18.300 344.400 ;
        RECT 23.700 343.500 24.900 347.400 ;
        RECT 19.200 342.600 24.900 343.500 ;
        RECT 38.100 344.400 39.900 350.400 ;
        RECT 41.100 344.400 42.900 351.000 ;
        RECT 44.100 347.400 45.900 350.400 ;
        RECT 19.200 341.700 21.000 342.600 ;
        RECT 17.100 334.950 19.200 337.050 ;
        RECT 17.100 327.600 18.300 334.950 ;
        RECT 20.100 330.300 21.000 341.700 ;
        RECT 38.100 337.050 39.300 344.400 ;
        RECT 44.700 343.500 45.900 347.400 ;
        RECT 40.200 342.600 45.900 343.500 ;
        RECT 47.550 344.400 49.350 350.400 ;
        RECT 50.850 344.400 52.650 351.000 ;
        RECT 55.950 347.400 57.750 350.400 ;
        RECT 60.450 347.400 62.250 351.000 ;
        RECT 63.450 347.400 65.250 350.400 ;
        RECT 66.750 347.400 68.550 351.000 ;
        RECT 71.250 348.300 73.050 350.400 ;
        RECT 71.250 347.400 74.850 348.300 ;
        RECT 55.350 345.300 57.750 347.400 ;
        RECT 64.200 346.500 65.250 347.400 ;
        RECT 71.250 346.800 75.150 347.400 ;
        RECT 64.200 345.450 69.150 346.500 ;
        RECT 67.350 344.700 69.150 345.450 ;
        RECT 40.200 341.700 42.000 342.600 ;
        RECT 22.500 334.950 24.600 337.050 ;
        RECT 22.800 333.150 24.600 334.950 ;
        RECT 38.100 334.950 40.200 337.050 ;
        RECT 19.200 329.400 21.000 330.300 ;
        RECT 19.200 328.500 24.900 329.400 ;
        RECT 17.100 315.600 18.900 327.600 ;
        RECT 20.100 315.000 21.900 325.800 ;
        RECT 23.700 321.600 24.900 328.500 ;
        RECT 23.100 315.600 24.900 321.600 ;
        RECT 38.100 327.600 39.300 334.950 ;
        RECT 41.100 330.300 42.000 341.700 ;
        RECT 47.550 337.050 48.750 344.400 ;
        RECT 70.350 343.800 72.150 345.600 ;
        RECT 73.050 345.300 75.150 346.800 ;
        RECT 76.050 344.400 77.850 351.000 ;
        RECT 79.050 346.200 80.850 350.400 ;
        RECT 95.100 347.400 96.900 350.400 ;
        RECT 98.100 347.400 99.900 351.000 ;
        RECT 79.050 344.400 81.450 346.200 ;
        RECT 60.150 342.000 61.950 342.600 ;
        RECT 71.100 342.000 72.150 343.800 ;
        RECT 60.150 340.800 72.150 342.000 ;
        RECT 43.500 334.950 45.600 337.050 ;
        RECT 43.800 333.150 45.600 334.950 ;
        RECT 47.550 335.250 53.850 337.050 ;
        RECT 47.550 334.950 52.050 335.250 ;
        RECT 40.200 329.400 42.000 330.300 ;
        RECT 40.200 328.500 45.900 329.400 ;
        RECT 38.100 315.600 39.900 327.600 ;
        RECT 41.100 315.000 42.900 325.800 ;
        RECT 44.700 321.600 45.900 328.500 ;
        RECT 44.100 315.600 45.900 321.600 ;
        RECT 47.550 327.600 48.750 334.950 ;
        RECT 49.650 332.100 51.450 332.250 ;
        RECT 55.350 332.100 57.450 332.400 ;
        RECT 49.650 330.900 57.450 332.100 ;
        RECT 49.650 330.450 51.450 330.900 ;
        RECT 55.350 330.300 57.450 330.900 ;
        RECT 60.150 328.200 61.050 340.800 ;
        RECT 71.100 339.600 79.050 340.800 ;
        RECT 71.100 339.000 72.900 339.600 ;
        RECT 74.100 337.800 75.900 338.400 ;
        RECT 67.800 336.600 75.900 337.800 ;
        RECT 77.250 337.050 79.050 339.600 ;
        RECT 67.800 334.950 69.900 336.600 ;
        RECT 76.950 334.950 79.050 337.050 ;
        RECT 69.750 329.700 71.550 330.000 ;
        RECT 80.550 329.700 81.450 344.400 ;
        RECT 95.700 337.050 96.900 347.400 ;
        RECT 101.550 344.400 103.350 350.400 ;
        RECT 104.850 344.400 106.650 351.000 ;
        RECT 109.950 347.400 111.750 350.400 ;
        RECT 114.450 347.400 116.250 351.000 ;
        RECT 117.450 347.400 119.250 350.400 ;
        RECT 120.750 347.400 122.550 351.000 ;
        RECT 125.250 348.300 127.050 350.400 ;
        RECT 125.250 347.400 128.850 348.300 ;
        RECT 109.350 345.300 111.750 347.400 ;
        RECT 118.200 346.500 119.250 347.400 ;
        RECT 125.250 346.800 129.150 347.400 ;
        RECT 118.200 345.450 123.150 346.500 ;
        RECT 121.350 344.700 123.150 345.450 ;
        RECT 101.550 337.050 102.750 344.400 ;
        RECT 124.350 343.800 126.150 345.600 ;
        RECT 127.050 345.300 129.150 346.800 ;
        RECT 130.050 344.400 131.850 351.000 ;
        RECT 152.100 350.400 153.300 351.000 ;
        RECT 133.050 346.200 134.850 350.400 ;
        RECT 152.100 347.400 153.900 350.400 ;
        RECT 155.100 347.400 156.900 350.400 ;
        RECT 133.050 344.400 135.450 346.200 ;
        RECT 114.150 342.000 115.950 342.600 ;
        RECT 125.100 342.000 126.150 343.800 ;
        RECT 114.150 340.800 126.150 342.000 ;
        RECT 94.950 334.950 97.050 337.050 ;
        RECT 97.950 334.950 100.050 337.050 ;
        RECT 101.550 335.250 107.850 337.050 ;
        RECT 101.550 334.950 106.050 335.250 ;
        RECT 69.750 329.100 81.450 329.700 ;
        RECT 47.550 315.600 49.350 327.600 ;
        RECT 50.550 315.000 52.350 327.600 ;
        RECT 56.250 327.300 61.050 328.200 ;
        RECT 63.150 328.500 81.450 329.100 ;
        RECT 63.150 328.200 71.550 328.500 ;
        RECT 56.250 326.400 57.450 327.300 ;
        RECT 54.450 324.600 57.450 326.400 ;
        RECT 58.350 326.100 60.150 326.400 ;
        RECT 63.150 326.100 64.050 328.200 ;
        RECT 80.550 327.600 81.450 328.500 ;
        RECT 58.350 325.200 64.050 326.100 ;
        RECT 64.950 326.700 66.750 327.300 ;
        RECT 64.950 325.500 72.750 326.700 ;
        RECT 58.350 324.600 60.150 325.200 ;
        RECT 70.650 324.600 72.750 325.500 ;
        RECT 55.350 321.600 57.450 323.700 ;
        RECT 61.950 323.550 63.750 324.300 ;
        RECT 66.750 323.550 68.550 324.300 ;
        RECT 61.950 322.500 68.550 323.550 ;
        RECT 55.350 315.600 57.150 321.600 ;
        RECT 59.850 315.000 61.650 321.600 ;
        RECT 62.850 315.600 64.650 322.500 ;
        RECT 65.850 315.000 67.650 321.600 ;
        RECT 70.650 315.600 72.450 324.600 ;
        RECT 76.050 315.000 77.850 327.600 ;
        RECT 79.050 325.800 81.450 327.600 ;
        RECT 79.050 315.600 80.850 325.800 ;
        RECT 95.700 321.600 96.900 334.950 ;
        RECT 98.100 333.150 99.900 334.950 ;
        RECT 101.550 327.600 102.750 334.950 ;
        RECT 103.650 332.100 105.450 332.250 ;
        RECT 109.350 332.100 111.450 332.400 ;
        RECT 103.650 330.900 111.450 332.100 ;
        RECT 103.650 330.450 105.450 330.900 ;
        RECT 109.350 330.300 111.450 330.900 ;
        RECT 114.150 328.200 115.050 340.800 ;
        RECT 125.100 339.600 133.050 340.800 ;
        RECT 125.100 339.000 126.900 339.600 ;
        RECT 128.100 337.800 129.900 338.400 ;
        RECT 121.800 336.600 129.900 337.800 ;
        RECT 131.250 337.050 133.050 339.600 ;
        RECT 121.800 334.950 123.900 336.600 ;
        RECT 130.950 334.950 133.050 337.050 ;
        RECT 123.750 329.700 125.550 330.000 ;
        RECT 134.550 329.700 135.450 344.400 ;
        RECT 155.400 343.200 156.300 347.400 ;
        RECT 158.100 345.000 159.900 351.000 ;
        RECT 161.100 344.400 162.900 350.400 ;
        RECT 155.400 342.300 160.800 343.200 ;
        RECT 158.700 341.400 160.800 342.300 ;
        RECT 152.400 337.050 154.200 338.850 ;
        RECT 152.100 334.950 154.200 337.050 ;
        RECT 155.400 334.950 157.500 337.050 ;
        RECT 156.000 333.150 157.800 334.950 ;
        RECT 158.700 330.900 159.600 341.400 ;
        RECT 162.000 337.050 162.900 344.400 ;
        RECT 176.100 345.300 177.900 350.400 ;
        RECT 179.100 346.200 180.900 351.000 ;
        RECT 182.100 345.300 183.900 350.400 ;
        RECT 176.100 343.950 183.900 345.300 ;
        RECT 185.100 344.400 186.900 350.400 ;
        RECT 203.100 344.400 204.900 350.400 ;
        RECT 185.100 342.300 186.300 344.400 ;
        RECT 182.700 341.400 186.300 342.300 ;
        RECT 203.700 342.300 204.900 344.400 ;
        RECT 206.100 345.300 207.900 350.400 ;
        RECT 209.100 346.200 210.900 351.000 ;
        RECT 212.100 345.300 213.900 350.400 ;
        RECT 206.100 343.950 213.900 345.300 ;
        RECT 230.700 343.200 232.500 350.400 ;
        RECT 235.800 344.400 237.600 351.000 ;
        RECT 254.400 344.400 256.200 351.000 ;
        RECT 259.500 343.200 261.300 350.400 ;
        RECT 275.100 347.400 276.900 351.000 ;
        RECT 278.100 347.400 279.900 350.400 ;
        RECT 281.100 347.400 282.900 351.000 ;
        RECT 230.700 342.300 234.900 343.200 ;
        RECT 203.700 341.400 207.300 342.300 ;
        RECT 179.100 337.050 180.900 338.850 ;
        RECT 182.700 337.050 183.900 341.400 ;
        RECT 185.100 337.050 186.900 338.850 ;
        RECT 203.100 337.050 204.900 338.850 ;
        RECT 206.100 337.050 207.300 341.400 ;
        RECT 209.100 337.050 210.900 338.850 ;
        RECT 230.100 337.050 231.900 338.850 ;
        RECT 233.700 337.050 234.900 342.300 ;
        RECT 257.100 342.300 261.300 343.200 ;
        RECT 235.950 337.050 237.750 338.850 ;
        RECT 254.250 337.050 256.050 338.850 ;
        RECT 257.100 337.050 258.300 342.300 ;
        RECT 260.100 337.050 261.900 338.850 ;
        RECT 278.700 337.050 279.600 347.400 ;
        RECT 296.700 343.200 298.500 350.400 ;
        RECT 301.800 344.400 303.600 351.000 ;
        RECT 317.700 344.400 319.500 351.000 ;
        RECT 322.200 344.400 324.000 350.400 ;
        RECT 326.700 344.400 328.500 351.000 ;
        RECT 347.100 347.400 348.900 351.000 ;
        RECT 350.100 347.400 351.900 350.400 ;
        RECT 367.800 347.400 369.900 351.000 ;
        RECT 371.100 347.400 372.900 350.400 ;
        RECT 374.100 347.400 375.900 351.000 ;
        RECT 377.100 347.400 379.800 350.400 ;
        RECT 296.700 342.300 300.900 343.200 ;
        RECT 283.950 339.450 286.050 340.050 ;
        RECT 289.950 339.450 292.050 340.050 ;
        RECT 283.950 338.550 292.050 339.450 ;
        RECT 283.950 337.950 286.050 338.550 ;
        RECT 289.950 337.950 292.050 338.550 ;
        RECT 296.100 337.050 297.900 338.850 ;
        RECT 299.700 337.050 300.900 342.300 ;
        RECT 301.950 337.050 303.750 338.850 ;
        RECT 317.250 337.050 319.050 338.850 ;
        RECT 323.100 337.050 324.300 344.400 ;
        RECT 329.100 337.050 330.900 338.850 ;
        RECT 350.100 337.050 351.300 347.400 ;
        RECT 371.700 346.500 372.600 347.400 ;
        RECT 378.900 346.500 379.800 347.400 ;
        RECT 371.700 345.600 384.300 346.500 ;
        RECT 373.950 337.050 375.750 338.850 ;
        RECT 383.100 337.050 384.300 345.600 ;
        RECT 388.950 345.450 391.050 346.050 ;
        RECT 394.950 345.450 397.050 346.050 ;
        RECT 388.950 344.550 397.050 345.450 ;
        RECT 388.950 343.950 391.050 344.550 ;
        RECT 394.950 343.950 397.050 344.550 ;
        RECT 401.100 345.300 402.900 350.400 ;
        RECT 404.100 346.200 405.900 351.000 ;
        RECT 407.100 345.300 408.900 350.400 ;
        RECT 401.100 343.950 408.900 345.300 ;
        RECT 410.100 344.400 411.900 350.400 ;
        RECT 426.000 344.400 427.800 351.000 ;
        RECT 430.500 345.600 432.300 350.400 ;
        RECT 433.500 347.400 435.300 351.000 ;
        RECT 430.500 344.400 435.600 345.600 ;
        RECT 410.100 342.300 411.300 344.400 ;
        RECT 407.700 341.400 411.300 342.300 ;
        RECT 404.100 337.050 405.900 338.850 ;
        RECT 407.700 337.050 408.900 341.400 ;
        RECT 410.100 337.050 411.900 338.850 ;
        RECT 425.100 337.050 426.900 338.850 ;
        RECT 431.250 337.050 433.050 338.850 ;
        RECT 434.700 337.050 435.600 344.400 ;
        RECT 449.100 341.400 450.900 351.000 ;
        RECT 455.700 342.000 457.500 350.400 ;
        RECT 473.100 345.300 474.900 350.400 ;
        RECT 476.100 346.200 477.900 351.000 ;
        RECT 479.100 345.300 480.900 350.400 ;
        RECT 473.100 343.950 480.900 345.300 ;
        RECT 482.100 344.400 483.900 350.400 ;
        RECT 500.100 345.300 501.900 350.400 ;
        RECT 503.100 346.200 504.900 351.000 ;
        RECT 506.100 345.300 507.900 350.400 ;
        RECT 482.100 342.300 483.300 344.400 ;
        RECT 500.100 343.950 507.900 345.300 ;
        RECT 509.100 344.400 510.900 350.400 ;
        RECT 509.100 342.300 510.300 344.400 ;
        RECT 455.700 340.800 459.000 342.000 ;
        RECT 449.100 337.050 450.900 338.850 ;
        RECT 455.100 337.050 456.900 338.850 ;
        RECT 458.100 337.050 459.000 340.800 ;
        RECT 479.700 341.400 483.300 342.300 ;
        RECT 506.700 341.400 510.300 342.300 ;
        RECT 526.500 342.000 528.300 350.400 ;
        RECT 476.100 337.050 477.900 338.850 ;
        RECT 479.700 337.050 480.900 341.400 ;
        RECT 482.100 337.050 483.900 338.850 ;
        RECT 503.100 337.050 504.900 338.850 ;
        RECT 506.700 337.050 507.900 341.400 ;
        RECT 525.000 340.800 528.300 342.000 ;
        RECT 533.100 341.400 534.900 351.000 ;
        RECT 548.100 341.400 549.900 351.000 ;
        RECT 554.700 342.000 556.500 350.400 ;
        RECT 575.100 344.400 576.900 350.400 ;
        RECT 575.700 342.300 576.900 344.400 ;
        RECT 578.100 345.300 579.900 350.400 ;
        RECT 581.100 346.200 582.900 351.000 ;
        RECT 584.100 345.300 585.900 350.400 ;
        RECT 578.100 343.950 585.900 345.300 ;
        RECT 599.700 343.200 601.500 350.400 ;
        RECT 604.800 344.400 606.600 351.000 ;
        RECT 624.600 346.200 626.400 350.400 ;
        RECT 623.700 344.400 626.400 346.200 ;
        RECT 627.600 344.400 629.400 351.000 ;
        RECT 599.700 342.300 603.900 343.200 ;
        RECT 554.700 340.800 558.000 342.000 ;
        RECT 575.700 341.400 579.300 342.300 ;
        RECT 509.100 337.050 510.900 338.850 ;
        RECT 525.000 337.050 525.900 340.800 ;
        RECT 527.100 337.050 528.900 338.850 ;
        RECT 533.100 337.050 534.900 338.850 ;
        RECT 548.100 337.050 549.900 338.850 ;
        RECT 554.100 337.050 555.900 338.850 ;
        RECT 557.100 337.050 558.000 340.800 ;
        RECT 570.000 339.450 574.050 340.050 ;
        RECT 569.550 337.950 574.050 339.450 ;
        RECT 160.800 334.950 162.900 337.050 ;
        RECT 175.950 334.950 178.050 337.050 ;
        RECT 178.950 334.950 181.050 337.050 ;
        RECT 181.950 334.950 184.050 337.050 ;
        RECT 184.950 334.950 187.050 337.050 ;
        RECT 158.100 330.300 159.900 330.900 ;
        RECT 123.750 329.100 135.450 329.700 ;
        RECT 95.100 315.600 96.900 321.600 ;
        RECT 98.100 315.000 99.900 321.600 ;
        RECT 101.550 315.600 103.350 327.600 ;
        RECT 104.550 315.000 106.350 327.600 ;
        RECT 110.250 327.300 115.050 328.200 ;
        RECT 117.150 328.500 135.450 329.100 ;
        RECT 117.150 328.200 125.550 328.500 ;
        RECT 110.250 326.400 111.450 327.300 ;
        RECT 108.450 324.600 111.450 326.400 ;
        RECT 112.350 326.100 114.150 326.400 ;
        RECT 117.150 326.100 118.050 328.200 ;
        RECT 134.550 327.600 135.450 328.500 ;
        RECT 112.350 325.200 118.050 326.100 ;
        RECT 118.950 326.700 120.750 327.300 ;
        RECT 118.950 325.500 126.750 326.700 ;
        RECT 112.350 324.600 114.150 325.200 ;
        RECT 124.650 324.600 126.750 325.500 ;
        RECT 109.350 321.600 111.450 323.700 ;
        RECT 115.950 323.550 117.750 324.300 ;
        RECT 120.750 323.550 122.550 324.300 ;
        RECT 115.950 322.500 122.550 323.550 ;
        RECT 109.350 315.600 111.150 321.600 ;
        RECT 113.850 315.000 115.650 321.600 ;
        RECT 116.850 315.600 118.650 322.500 ;
        RECT 119.850 315.000 121.650 321.600 ;
        RECT 124.650 315.600 126.450 324.600 ;
        RECT 130.050 315.000 131.850 327.600 ;
        RECT 133.050 325.800 135.450 327.600 ;
        RECT 152.100 329.100 159.900 330.300 ;
        RECT 152.100 327.600 153.300 329.100 ;
        RECT 160.800 327.600 162.000 334.950 ;
        RECT 176.100 333.150 177.900 334.950 ;
        RECT 169.950 330.450 172.050 331.050 ;
        RECT 178.950 330.450 181.050 331.050 ;
        RECT 169.950 329.550 181.050 330.450 ;
        RECT 169.950 328.950 172.050 329.550 ;
        RECT 178.950 328.950 181.050 329.550 ;
        RECT 182.700 327.600 183.900 334.950 ;
        RECT 190.950 334.050 193.050 337.050 ;
        RECT 202.950 334.950 205.050 337.050 ;
        RECT 205.950 334.950 208.050 337.050 ;
        RECT 208.950 334.950 211.050 337.050 ;
        RECT 211.950 334.950 214.050 337.050 ;
        RECT 229.950 334.950 232.050 337.050 ;
        RECT 232.950 334.950 235.050 337.050 ;
        RECT 235.950 334.950 238.050 337.050 ;
        RECT 253.950 334.950 256.050 337.050 ;
        RECT 256.950 334.950 259.050 337.050 ;
        RECT 259.950 334.950 262.050 337.050 ;
        RECT 274.950 334.950 277.050 337.050 ;
        RECT 277.950 334.950 280.050 337.050 ;
        RECT 280.950 334.950 283.050 337.050 ;
        RECT 295.950 334.950 298.050 337.050 ;
        RECT 298.950 334.950 301.050 337.050 ;
        RECT 301.950 334.950 304.050 337.050 ;
        RECT 316.950 334.950 319.050 337.050 ;
        RECT 319.950 334.950 322.050 337.050 ;
        RECT 322.950 334.950 325.050 337.050 ;
        RECT 325.950 334.950 328.050 337.050 ;
        RECT 328.950 334.950 331.050 337.050 ;
        RECT 346.950 334.950 349.050 337.050 ;
        RECT 349.950 334.950 352.050 337.050 ;
        RECT 367.800 334.950 369.900 337.050 ;
        RECT 373.950 334.950 376.050 337.050 ;
        RECT 376.950 334.950 379.050 337.050 ;
        RECT 382.500 334.950 384.600 337.050 ;
        RECT 400.950 334.950 403.050 337.050 ;
        RECT 403.950 334.950 406.050 337.050 ;
        RECT 406.950 334.950 409.050 337.050 ;
        RECT 409.950 334.950 412.050 337.050 ;
        RECT 424.950 334.950 427.050 337.050 ;
        RECT 427.950 334.950 430.050 337.050 ;
        RECT 430.950 334.950 433.050 337.050 ;
        RECT 433.950 334.950 436.050 337.050 ;
        RECT 448.950 334.950 451.050 337.050 ;
        RECT 451.950 334.950 454.050 337.050 ;
        RECT 454.950 334.950 457.050 337.050 ;
        RECT 457.950 334.950 460.050 337.050 ;
        RECT 472.950 334.950 475.050 337.050 ;
        RECT 475.950 334.950 478.050 337.050 ;
        RECT 478.950 334.950 481.050 337.050 ;
        RECT 481.950 334.950 484.050 337.050 ;
        RECT 499.950 334.950 502.050 337.050 ;
        RECT 502.950 334.950 505.050 337.050 ;
        RECT 505.950 334.950 508.050 337.050 ;
        RECT 508.950 334.950 511.050 337.050 ;
        RECT 523.950 334.950 526.050 337.050 ;
        RECT 526.950 334.950 529.050 337.050 ;
        RECT 529.950 334.950 532.050 337.050 ;
        RECT 532.950 334.950 535.050 337.050 ;
        RECT 547.950 334.950 550.050 337.050 ;
        RECT 550.950 334.950 553.050 337.050 ;
        RECT 553.950 334.950 556.050 337.050 ;
        RECT 556.950 334.950 559.050 337.050 ;
        RECT 187.950 333.000 193.050 334.050 ;
        RECT 187.950 332.550 192.450 333.000 ;
        RECT 187.950 331.950 192.000 332.550 ;
        RECT 133.050 315.600 134.850 325.800 ;
        RECT 152.100 315.600 153.900 327.600 ;
        RECT 156.600 315.000 158.400 327.600 ;
        RECT 159.600 326.100 162.000 327.600 ;
        RECT 159.600 315.600 161.400 326.100 ;
        RECT 176.400 315.000 178.200 327.600 ;
        RECT 181.500 326.100 183.900 327.600 ;
        RECT 206.100 327.600 207.300 334.950 ;
        RECT 212.100 333.150 213.900 334.950 ;
        RECT 206.100 326.100 208.500 327.600 ;
        RECT 181.500 315.600 183.300 326.100 ;
        RECT 184.200 323.100 186.000 324.900 ;
        RECT 204.000 323.100 205.800 324.900 ;
        RECT 184.500 315.000 186.300 321.600 ;
        RECT 203.700 315.000 205.500 321.600 ;
        RECT 206.700 315.600 208.500 326.100 ;
        RECT 211.800 315.000 213.600 327.600 ;
        RECT 233.700 321.600 234.900 334.950 ;
        RECT 257.100 321.600 258.300 334.950 ;
        RECT 275.100 333.150 276.900 334.950 ;
        RECT 278.700 327.600 279.600 334.950 ;
        RECT 280.950 333.150 282.750 334.950 ;
        RECT 276.000 326.400 279.600 327.600 ;
        RECT 230.100 315.000 231.900 321.600 ;
        RECT 233.100 315.600 234.900 321.600 ;
        RECT 236.100 315.000 237.900 321.600 ;
        RECT 254.100 315.000 255.900 321.600 ;
        RECT 257.100 315.600 258.900 321.600 ;
        RECT 260.100 315.000 261.900 321.600 ;
        RECT 276.000 315.600 277.800 326.400 ;
        RECT 281.100 315.000 282.900 327.600 ;
        RECT 299.700 321.600 300.900 334.950 ;
        RECT 320.250 333.150 322.050 334.950 ;
        RECT 323.100 329.400 324.000 334.950 ;
        RECT 326.100 333.150 327.900 334.950 ;
        RECT 347.100 333.150 348.900 334.950 ;
        RECT 323.100 328.500 327.900 329.400 ;
        RECT 317.100 326.400 324.900 327.300 ;
        RECT 296.100 315.000 297.900 321.600 ;
        RECT 299.100 315.600 300.900 321.600 ;
        RECT 302.100 315.000 303.900 321.600 ;
        RECT 317.100 315.600 318.900 326.400 ;
        RECT 320.100 315.000 321.900 325.500 ;
        RECT 323.100 316.500 324.900 326.400 ;
        RECT 326.100 317.400 327.900 328.500 ;
        RECT 329.100 316.500 330.900 327.600 ;
        RECT 350.100 321.600 351.300 334.950 ;
        RECT 368.100 333.150 369.900 334.950 ;
        RECT 377.250 333.150 379.050 334.950 ;
        RECT 365.100 325.500 372.900 326.400 ;
        RECT 323.100 315.600 330.900 316.500 ;
        RECT 347.100 315.000 348.900 321.600 ;
        RECT 350.100 315.600 351.900 321.600 ;
        RECT 365.100 315.600 366.900 325.500 ;
        RECT 368.100 315.000 369.900 324.600 ;
        RECT 371.100 316.500 372.900 325.500 ;
        RECT 374.100 325.200 381.900 326.100 ;
        RECT 374.100 317.400 375.900 325.200 ;
        RECT 377.100 316.500 378.900 324.300 ;
        RECT 371.100 315.600 378.900 316.500 ;
        RECT 380.100 316.500 381.900 325.200 ;
        RECT 383.100 325.200 384.300 334.950 ;
        RECT 401.100 333.150 402.900 334.950 ;
        RECT 407.700 327.600 408.900 334.950 ;
        RECT 428.250 333.150 430.050 334.950 ;
        RECT 434.700 327.600 435.600 334.950 ;
        RECT 452.100 333.150 453.900 334.950 ;
        RECT 383.100 317.400 384.900 325.200 ;
        RECT 386.100 316.500 387.900 325.800 ;
        RECT 380.100 315.600 387.900 316.500 ;
        RECT 401.400 315.000 403.200 327.600 ;
        RECT 406.500 326.100 408.900 327.600 ;
        RECT 425.100 326.700 432.900 327.600 ;
        RECT 406.500 315.600 408.300 326.100 ;
        RECT 409.200 323.100 411.000 324.900 ;
        RECT 409.500 315.000 411.300 321.600 ;
        RECT 425.100 315.600 426.900 326.700 ;
        RECT 428.100 315.000 429.900 325.800 ;
        RECT 431.100 315.600 432.900 326.700 ;
        RECT 434.100 315.600 435.900 327.600 ;
        RECT 458.100 322.800 459.000 334.950 ;
        RECT 473.100 333.150 474.900 334.950 ;
        RECT 479.700 327.600 480.900 334.950 ;
        RECT 484.950 333.450 487.050 334.050 ;
        RECT 493.950 333.450 496.050 334.050 ;
        RECT 484.950 332.550 496.050 333.450 ;
        RECT 500.100 333.150 501.900 334.950 ;
        RECT 484.950 331.950 487.050 332.550 ;
        RECT 493.950 331.950 496.050 332.550 ;
        RECT 506.700 327.600 507.900 334.950 ;
        RECT 452.400 321.900 459.000 322.800 ;
        RECT 452.400 321.600 453.900 321.900 ;
        RECT 449.100 315.000 450.900 321.600 ;
        RECT 452.100 315.600 453.900 321.600 ;
        RECT 458.100 321.600 459.000 321.900 ;
        RECT 455.100 315.000 456.900 321.000 ;
        RECT 458.100 315.600 459.900 321.600 ;
        RECT 473.400 315.000 475.200 327.600 ;
        RECT 478.500 326.100 480.900 327.600 ;
        RECT 478.500 315.600 480.300 326.100 ;
        RECT 481.200 323.100 483.000 324.900 ;
        RECT 481.500 315.000 483.300 321.600 ;
        RECT 500.400 315.000 502.200 327.600 ;
        RECT 505.500 326.100 507.900 327.600 ;
        RECT 505.500 315.600 507.300 326.100 ;
        RECT 508.200 323.100 510.000 324.900 ;
        RECT 525.000 322.800 525.900 334.950 ;
        RECT 530.100 333.150 531.900 334.950 ;
        RECT 551.100 333.150 552.900 334.950 ;
        RECT 557.100 322.800 558.000 334.950 ;
        RECT 569.550 334.050 570.450 337.950 ;
        RECT 575.100 337.050 576.900 338.850 ;
        RECT 578.100 337.050 579.300 341.400 ;
        RECT 581.100 337.050 582.900 338.850 ;
        RECT 599.100 337.050 600.900 338.850 ;
        RECT 602.700 337.050 603.900 342.300 ;
        RECT 604.950 337.050 606.750 338.850 ;
        RECT 623.700 337.050 624.600 344.400 ;
        RECT 625.500 342.600 627.300 343.500 ;
        RECT 632.100 342.600 633.900 350.400 ;
        RECT 647.100 347.400 648.900 350.400 ;
        RECT 647.100 343.500 648.300 347.400 ;
        RECT 650.100 344.400 651.900 351.000 ;
        RECT 653.100 344.400 654.900 350.400 ;
        RECT 647.100 342.600 652.800 343.500 ;
        RECT 625.500 341.700 633.900 342.600 ;
        RECT 651.000 341.700 652.800 342.600 ;
        RECT 574.950 334.950 577.050 337.050 ;
        RECT 577.950 334.950 580.050 337.050 ;
        RECT 580.950 334.950 583.050 337.050 ;
        RECT 583.950 334.950 586.050 337.050 ;
        RECT 598.950 334.950 601.050 337.050 ;
        RECT 601.950 334.950 604.050 337.050 ;
        RECT 604.950 334.950 607.050 337.050 ;
        RECT 623.100 334.950 625.200 337.050 ;
        RECT 626.400 334.950 628.500 337.050 ;
        RECT 569.550 332.550 574.050 334.050 ;
        RECT 570.000 331.950 574.050 332.550 ;
        RECT 578.100 327.600 579.300 334.950 ;
        RECT 584.100 333.150 585.900 334.950 ;
        RECT 578.100 326.100 580.500 327.600 ;
        RECT 576.000 323.100 577.800 324.900 ;
        RECT 525.000 321.900 531.600 322.800 ;
        RECT 525.000 321.600 525.900 321.900 ;
        RECT 508.500 315.000 510.300 321.600 ;
        RECT 524.100 315.600 525.900 321.600 ;
        RECT 530.100 321.600 531.600 321.900 ;
        RECT 551.400 321.900 558.000 322.800 ;
        RECT 551.400 321.600 552.900 321.900 ;
        RECT 527.100 315.000 528.900 321.000 ;
        RECT 530.100 315.600 531.900 321.600 ;
        RECT 533.100 315.000 534.900 321.600 ;
        RECT 548.100 315.000 549.900 321.600 ;
        RECT 551.100 315.600 552.900 321.600 ;
        RECT 557.100 321.600 558.000 321.900 ;
        RECT 554.100 315.000 555.900 321.000 ;
        RECT 557.100 315.600 558.900 321.600 ;
        RECT 575.700 315.000 577.500 321.600 ;
        RECT 578.700 315.600 580.500 326.100 ;
        RECT 583.800 315.000 585.600 327.600 ;
        RECT 602.700 321.600 603.900 334.950 ;
        RECT 623.700 327.600 624.600 334.950 ;
        RECT 627.000 333.150 628.800 334.950 ;
        RECT 599.100 315.000 600.900 321.600 ;
        RECT 602.100 315.600 603.900 321.600 ;
        RECT 605.100 315.000 606.900 321.600 ;
        RECT 623.100 315.600 624.900 327.600 ;
        RECT 626.100 315.000 627.900 327.000 ;
        RECT 630.000 321.600 630.900 341.700 ;
        RECT 631.950 337.050 633.750 338.850 ;
        RECT 631.800 334.950 633.900 337.050 ;
        RECT 647.400 334.950 649.500 337.050 ;
        RECT 647.400 333.150 649.200 334.950 ;
        RECT 651.000 330.300 651.900 341.700 ;
        RECT 653.700 337.050 654.900 344.400 ;
        RECT 671.700 343.200 673.500 350.400 ;
        RECT 676.800 344.400 678.600 351.000 ;
        RECT 696.000 344.400 697.800 351.000 ;
        RECT 700.500 345.600 702.300 350.400 ;
        RECT 703.500 347.400 705.300 351.000 ;
        RECT 719.100 347.400 720.900 350.400 ;
        RECT 722.100 347.400 723.900 351.000 ;
        RECT 700.500 344.400 705.600 345.600 ;
        RECT 671.700 342.300 675.900 343.200 ;
        RECT 671.100 337.050 672.900 338.850 ;
        RECT 674.700 337.050 675.900 342.300 ;
        RECT 676.950 337.050 678.750 338.850 ;
        RECT 695.100 337.050 696.900 338.850 ;
        RECT 701.250 337.050 703.050 338.850 ;
        RECT 704.700 337.050 705.600 344.400 ;
        RECT 719.700 337.050 720.900 347.400 ;
        RECT 737.100 344.400 738.900 350.400 ;
        RECT 737.700 342.300 738.900 344.400 ;
        RECT 740.100 345.300 741.900 350.400 ;
        RECT 743.100 346.200 744.900 351.000 ;
        RECT 746.100 345.300 747.900 350.400 ;
        RECT 740.100 343.950 747.900 345.300 ;
        RECT 761.100 345.300 762.900 350.400 ;
        RECT 764.100 346.200 765.900 351.000 ;
        RECT 767.100 345.300 768.900 350.400 ;
        RECT 761.100 343.950 768.900 345.300 ;
        RECT 770.100 344.400 771.900 350.400 ;
        RECT 770.100 342.300 771.300 344.400 ;
        RECT 737.700 341.400 741.300 342.300 ;
        RECT 737.100 337.050 738.900 338.850 ;
        RECT 740.100 337.050 741.300 341.400 ;
        RECT 767.700 341.400 771.300 342.300 ;
        RECT 785.100 341.400 786.900 351.000 ;
        RECT 791.700 342.000 793.500 350.400 ;
        RECT 809.700 343.200 811.500 350.400 ;
        RECT 814.800 344.400 816.600 351.000 ;
        RECT 830.100 344.400 831.900 350.400 ;
        RECT 809.700 342.300 813.900 343.200 ;
        RECT 743.100 337.050 744.900 338.850 ;
        RECT 764.100 337.050 765.900 338.850 ;
        RECT 767.700 337.050 768.900 341.400 ;
        RECT 791.700 340.800 795.000 342.000 ;
        RECT 772.950 339.450 777.000 340.050 ;
        RECT 770.100 337.050 771.900 338.850 ;
        RECT 772.950 337.950 777.450 339.450 ;
        RECT 652.800 334.950 654.900 337.050 ;
        RECT 670.950 334.950 673.050 337.050 ;
        RECT 673.950 334.950 676.050 337.050 ;
        RECT 676.950 334.950 679.050 337.050 ;
        RECT 694.950 334.950 697.050 337.050 ;
        RECT 697.950 334.950 700.050 337.050 ;
        RECT 700.950 334.950 703.050 337.050 ;
        RECT 703.950 334.950 706.050 337.050 ;
        RECT 718.950 334.950 721.050 337.050 ;
        RECT 721.950 334.950 724.050 337.050 ;
        RECT 736.950 334.950 739.050 337.050 ;
        RECT 739.950 334.950 742.050 337.050 ;
        RECT 742.950 334.950 745.050 337.050 ;
        RECT 745.950 334.950 748.050 337.050 ;
        RECT 760.950 334.950 763.050 337.050 ;
        RECT 763.950 334.950 766.050 337.050 ;
        RECT 766.950 334.950 769.050 337.050 ;
        RECT 769.950 334.950 772.050 337.050 ;
        RECT 651.000 329.400 652.800 330.300 ;
        RECT 647.100 328.500 652.800 329.400 ;
        RECT 647.100 321.600 648.300 328.500 ;
        RECT 653.700 327.600 654.900 334.950 ;
        RECT 629.100 315.600 630.900 321.600 ;
        RECT 632.100 315.000 633.900 321.600 ;
        RECT 647.100 315.600 648.900 321.600 ;
        RECT 650.100 315.000 651.900 325.800 ;
        RECT 653.100 315.600 654.900 327.600 ;
        RECT 674.700 321.600 675.900 334.950 ;
        RECT 698.250 333.150 700.050 334.950 ;
        RECT 704.700 327.600 705.600 334.950 ;
        RECT 695.100 326.700 702.900 327.600 ;
        RECT 671.100 315.000 672.900 321.600 ;
        RECT 674.100 315.600 675.900 321.600 ;
        RECT 677.100 315.000 678.900 321.600 ;
        RECT 695.100 315.600 696.900 326.700 ;
        RECT 698.100 315.000 699.900 325.800 ;
        RECT 701.100 315.600 702.900 326.700 ;
        RECT 704.100 315.600 705.900 327.600 ;
        RECT 719.700 321.600 720.900 334.950 ;
        RECT 722.100 333.150 723.900 334.950 ;
        RECT 740.100 327.600 741.300 334.950 ;
        RECT 746.100 333.150 747.900 334.950 ;
        RECT 761.100 333.150 762.900 334.950 ;
        RECT 745.950 330.450 748.050 331.050 ;
        RECT 754.950 330.450 757.050 331.050 ;
        RECT 745.950 329.550 757.050 330.450 ;
        RECT 745.950 328.950 748.050 329.550 ;
        RECT 754.950 328.950 757.050 329.550 ;
        RECT 767.700 327.600 768.900 334.950 ;
        RECT 776.550 333.450 777.450 337.950 ;
        RECT 785.100 337.050 786.900 338.850 ;
        RECT 791.100 337.050 792.900 338.850 ;
        RECT 794.100 337.050 795.000 340.800 ;
        RECT 809.100 337.050 810.900 338.850 ;
        RECT 812.700 337.050 813.900 342.300 ;
        RECT 830.700 342.300 831.900 344.400 ;
        RECT 833.100 345.300 834.900 350.400 ;
        RECT 836.100 346.200 837.900 351.000 ;
        RECT 839.100 345.300 840.900 350.400 ;
        RECT 854.700 347.400 856.500 351.000 ;
        RECT 857.700 345.600 859.500 350.400 ;
        RECT 833.100 343.950 840.900 345.300 ;
        RECT 854.400 344.400 859.500 345.600 ;
        RECT 862.200 344.400 864.000 351.000 ;
        RECT 830.700 341.400 834.300 342.300 ;
        RECT 814.950 337.050 816.750 338.850 ;
        RECT 830.100 337.050 831.900 338.850 ;
        RECT 833.100 337.050 834.300 341.400 ;
        RECT 836.100 337.050 837.900 338.850 ;
        RECT 854.400 337.050 855.300 344.400 ;
        RECT 856.950 342.450 859.050 343.050 ;
        RECT 856.950 341.550 870.450 342.450 ;
        RECT 880.500 342.000 882.300 350.400 ;
        RECT 856.950 340.950 859.050 341.550 ;
        RECT 856.950 337.050 858.750 338.850 ;
        RECT 863.100 337.050 864.900 338.850 ;
        RECT 784.950 334.950 787.050 337.050 ;
        RECT 787.950 334.950 790.050 337.050 ;
        RECT 790.950 334.950 793.050 337.050 ;
        RECT 793.950 334.950 796.050 337.050 ;
        RECT 808.950 334.950 811.050 337.050 ;
        RECT 811.950 334.950 814.050 337.050 ;
        RECT 814.950 334.950 817.050 337.050 ;
        RECT 829.950 334.950 832.050 337.050 ;
        RECT 832.950 334.950 835.050 337.050 ;
        RECT 835.950 334.950 838.050 337.050 ;
        RECT 838.950 334.950 841.050 337.050 ;
        RECT 853.950 334.950 856.050 337.050 ;
        RECT 856.950 334.950 859.050 337.050 ;
        RECT 859.950 334.950 862.050 337.050 ;
        RECT 862.950 334.950 865.050 337.050 ;
        RECT 781.950 333.450 784.050 334.050 ;
        RECT 776.550 332.550 784.050 333.450 ;
        RECT 788.100 333.150 789.900 334.950 ;
        RECT 781.950 331.950 784.050 332.550 ;
        RECT 740.100 326.100 742.500 327.600 ;
        RECT 738.000 323.100 739.800 324.900 ;
        RECT 719.100 315.600 720.900 321.600 ;
        RECT 722.100 315.000 723.900 321.600 ;
        RECT 737.700 315.000 739.500 321.600 ;
        RECT 740.700 315.600 742.500 326.100 ;
        RECT 745.800 315.000 747.600 327.600 ;
        RECT 761.400 315.000 763.200 327.600 ;
        RECT 766.500 326.100 768.900 327.600 ;
        RECT 766.500 315.600 768.300 326.100 ;
        RECT 769.200 323.100 771.000 324.900 ;
        RECT 794.100 322.800 795.000 334.950 ;
        RECT 788.400 321.900 795.000 322.800 ;
        RECT 788.400 321.600 789.900 321.900 ;
        RECT 769.500 315.000 771.300 321.600 ;
        RECT 785.100 315.000 786.900 321.600 ;
        RECT 788.100 315.600 789.900 321.600 ;
        RECT 794.100 321.600 795.000 321.900 ;
        RECT 812.700 321.600 813.900 334.950 ;
        RECT 833.100 327.600 834.300 334.950 ;
        RECT 839.100 333.150 840.900 334.950 ;
        RECT 854.400 327.600 855.300 334.950 ;
        RECT 859.950 333.150 861.750 334.950 ;
        RECT 869.550 333.450 870.450 341.550 ;
        RECT 879.000 340.800 882.300 342.000 ;
        RECT 887.100 341.400 888.900 351.000 ;
        RECT 873.000 339.450 877.050 340.050 ;
        RECT 866.550 332.550 870.450 333.450 ;
        RECT 872.550 337.950 877.050 339.450 ;
        RECT 856.950 330.450 859.050 330.750 ;
        RECT 866.550 330.450 867.450 332.550 ;
        RECT 872.550 331.050 873.450 337.950 ;
        RECT 879.000 337.050 879.900 340.800 ;
        RECT 881.100 337.050 882.900 338.850 ;
        RECT 887.100 337.050 888.900 338.850 ;
        RECT 877.950 334.950 880.050 337.050 ;
        RECT 880.950 334.950 883.050 337.050 ;
        RECT 883.950 334.950 886.050 337.050 ;
        RECT 886.950 334.950 889.050 337.050 ;
        RECT 856.950 329.550 867.450 330.450 ;
        RECT 868.950 329.550 873.450 331.050 ;
        RECT 856.950 328.650 859.050 329.550 ;
        RECT 868.950 328.950 873.000 329.550 ;
        RECT 833.100 326.100 835.500 327.600 ;
        RECT 831.000 323.100 832.800 324.900 ;
        RECT 791.100 315.000 792.900 321.000 ;
        RECT 794.100 315.600 795.900 321.600 ;
        RECT 809.100 315.000 810.900 321.600 ;
        RECT 812.100 315.600 813.900 321.600 ;
        RECT 815.100 315.000 816.900 321.600 ;
        RECT 830.700 315.000 832.500 321.600 ;
        RECT 833.700 315.600 835.500 326.100 ;
        RECT 838.800 315.000 840.600 327.600 ;
        RECT 854.100 315.600 855.900 327.600 ;
        RECT 857.100 326.700 864.900 327.600 ;
        RECT 857.100 315.600 858.900 326.700 ;
        RECT 860.100 315.000 861.900 325.800 ;
        RECT 863.100 315.600 864.900 326.700 ;
        RECT 879.000 322.800 879.900 334.950 ;
        RECT 884.100 333.150 885.900 334.950 ;
        RECT 879.000 321.900 885.600 322.800 ;
        RECT 879.000 321.600 879.900 321.900 ;
        RECT 878.100 315.600 879.900 321.600 ;
        RECT 884.100 321.600 885.600 321.900 ;
        RECT 881.100 315.000 882.900 321.000 ;
        RECT 884.100 315.600 885.900 321.600 ;
        RECT 887.100 315.000 888.900 321.600 ;
        RECT 14.100 300.600 15.900 311.400 ;
        RECT 17.100 301.500 18.900 312.000 ;
        RECT 14.100 299.400 18.900 300.600 ;
        RECT 16.800 298.500 18.900 299.400 ;
        RECT 21.600 299.400 23.400 311.400 ;
        RECT 26.100 301.500 27.900 312.000 ;
        RECT 29.100 300.300 30.900 311.400 ;
        RECT 47.100 305.400 48.900 312.000 ;
        RECT 50.100 305.400 51.900 311.400 ;
        RECT 53.100 305.400 54.900 312.000 ;
        RECT 26.400 299.400 30.900 300.300 ;
        RECT 21.600 298.050 22.800 299.400 ;
        RECT 21.300 297.000 22.800 298.050 ;
        RECT 26.400 297.300 28.500 299.400 ;
        RECT 21.300 295.050 22.200 297.000 ;
        RECT 14.400 292.050 16.200 293.850 ;
        RECT 20.100 292.950 22.200 295.050 ;
        RECT 23.100 295.500 25.200 295.800 ;
        RECT 23.100 293.700 27.000 295.500 ;
        RECT 14.100 289.950 16.200 292.050 ;
        RECT 20.700 292.800 22.200 292.950 ;
        RECT 20.700 291.900 23.100 292.800 ;
        RECT 18.900 289.200 20.700 291.000 ;
        RECT 18.900 287.100 21.000 289.200 ;
        RECT 21.900 286.200 23.100 291.900 ;
        RECT 24.000 292.050 25.800 292.500 ;
        RECT 50.100 292.050 51.300 305.400 ;
        RECT 56.550 299.400 58.350 311.400 ;
        RECT 59.550 299.400 61.350 312.000 ;
        RECT 64.350 305.400 66.150 311.400 ;
        RECT 68.850 305.400 70.650 312.000 ;
        RECT 64.350 303.300 66.450 305.400 ;
        RECT 71.850 304.500 73.650 311.400 ;
        RECT 74.850 305.400 76.650 312.000 ;
        RECT 70.950 303.450 77.550 304.500 ;
        RECT 70.950 302.700 72.750 303.450 ;
        RECT 75.750 302.700 77.550 303.450 ;
        RECT 79.650 302.400 81.450 311.400 ;
        RECT 63.450 300.600 66.450 302.400 ;
        RECT 67.350 301.800 69.150 302.400 ;
        RECT 67.350 300.900 73.050 301.800 ;
        RECT 79.650 301.500 81.750 302.400 ;
        RECT 67.350 300.600 69.150 300.900 ;
        RECT 65.250 299.700 66.450 300.600 ;
        RECT 56.550 292.050 57.750 299.400 ;
        RECT 65.250 298.800 70.050 299.700 ;
        RECT 58.650 296.100 60.450 296.550 ;
        RECT 64.350 296.100 66.450 296.700 ;
        RECT 58.650 294.900 66.450 296.100 ;
        RECT 58.650 294.750 60.450 294.900 ;
        RECT 64.350 294.600 66.450 294.900 ;
        RECT 24.000 290.700 30.900 292.050 ;
        RECT 28.800 289.950 30.900 290.700 ;
        RECT 46.950 289.950 49.050 292.050 ;
        RECT 49.950 289.950 52.050 292.050 ;
        RECT 52.950 289.950 55.050 292.050 ;
        RECT 56.550 291.750 61.050 292.050 ;
        RECT 56.550 289.950 62.850 291.750 ;
        RECT 16.800 283.500 18.900 284.700 ;
        RECT 20.100 284.100 23.100 286.200 ;
        RECT 24.000 287.400 25.800 289.200 ;
        RECT 28.800 288.150 30.600 289.950 ;
        RECT 47.250 288.150 49.050 289.950 ;
        RECT 24.000 285.300 26.100 287.400 ;
        RECT 24.000 284.400 30.300 285.300 ;
        RECT 14.100 282.600 18.900 283.500 ;
        RECT 21.900 282.600 23.100 284.100 ;
        RECT 29.100 282.600 30.300 284.400 ;
        RECT 50.100 284.700 51.300 289.950 ;
        RECT 53.100 288.150 54.900 289.950 ;
        RECT 50.100 283.800 54.300 284.700 ;
        RECT 14.100 276.600 15.900 282.600 ;
        RECT 17.100 276.000 18.900 281.700 ;
        RECT 21.600 276.600 23.400 282.600 ;
        RECT 26.100 276.000 27.900 281.700 ;
        RECT 29.100 276.600 30.900 282.600 ;
        RECT 47.400 276.000 49.200 282.600 ;
        RECT 52.500 276.600 54.300 283.800 ;
        RECT 56.550 282.600 57.750 289.950 ;
        RECT 69.150 286.200 70.050 298.800 ;
        RECT 72.150 298.800 73.050 300.900 ;
        RECT 73.950 300.300 81.750 301.500 ;
        RECT 73.950 299.700 75.750 300.300 ;
        RECT 85.050 299.400 86.850 312.000 ;
        RECT 88.050 301.200 89.850 311.400 ;
        RECT 104.100 305.400 105.900 312.000 ;
        RECT 107.100 305.400 108.900 311.400 ;
        RECT 110.100 305.400 111.900 312.000 ;
        RECT 125.100 305.400 126.900 312.000 ;
        RECT 128.100 305.400 129.900 311.400 ;
        RECT 88.050 299.400 90.450 301.200 ;
        RECT 72.150 298.500 80.550 298.800 ;
        RECT 89.550 298.500 90.450 299.400 ;
        RECT 72.150 297.900 90.450 298.500 ;
        RECT 78.750 297.300 90.450 297.900 ;
        RECT 78.750 297.000 80.550 297.300 ;
        RECT 76.800 290.400 78.900 292.050 ;
        RECT 76.800 289.200 84.900 290.400 ;
        RECT 85.950 289.950 88.050 292.050 ;
        RECT 83.100 288.600 84.900 289.200 ;
        RECT 80.100 287.400 81.900 288.000 ;
        RECT 86.250 287.400 88.050 289.950 ;
        RECT 80.100 286.200 88.050 287.400 ;
        RECT 69.150 285.000 81.150 286.200 ;
        RECT 69.150 284.400 70.950 285.000 ;
        RECT 80.100 283.200 81.150 285.000 ;
        RECT 56.550 276.600 58.350 282.600 ;
        RECT 59.850 276.000 61.650 282.600 ;
        RECT 64.350 279.600 66.750 281.700 ;
        RECT 76.350 281.550 78.150 282.300 ;
        RECT 73.200 280.500 78.150 281.550 ;
        RECT 79.350 281.400 81.150 283.200 ;
        RECT 89.550 282.600 90.450 297.300 ;
        RECT 107.100 292.050 108.300 305.400 ;
        RECT 103.950 289.950 106.050 292.050 ;
        RECT 106.950 289.950 109.050 292.050 ;
        RECT 109.950 289.950 112.050 292.050 ;
        RECT 125.100 289.950 127.200 292.050 ;
        RECT 104.250 288.150 106.050 289.950 ;
        RECT 107.100 284.700 108.300 289.950 ;
        RECT 110.100 288.150 111.900 289.950 ;
        RECT 125.250 288.150 127.050 289.950 ;
        RECT 128.100 285.300 129.000 305.400 ;
        RECT 131.100 300.000 132.900 312.000 ;
        RECT 134.100 299.400 135.900 311.400 ;
        RECT 149.100 299.400 150.900 312.000 ;
        RECT 154.200 300.600 156.000 311.400 ;
        RECT 152.400 299.400 156.000 300.600 ;
        RECT 170.400 299.400 172.200 312.000 ;
        RECT 175.500 300.900 177.300 311.400 ;
        RECT 178.500 305.400 180.300 312.000 ;
        RECT 197.700 305.400 199.500 312.000 ;
        RECT 178.200 302.100 180.000 303.900 ;
        RECT 198.000 302.100 199.800 303.900 ;
        RECT 200.700 300.900 202.500 311.400 ;
        RECT 175.500 299.400 177.900 300.900 ;
        RECT 130.200 292.050 132.000 293.850 ;
        RECT 134.400 292.050 135.300 299.400 ;
        RECT 149.250 292.050 151.050 293.850 ;
        RECT 152.400 292.050 153.300 299.400 ;
        RECT 155.100 292.050 156.900 293.850 ;
        RECT 170.100 292.050 171.900 293.850 ;
        RECT 176.700 292.050 177.900 299.400 ;
        RECT 200.100 299.400 202.500 300.900 ;
        RECT 205.800 299.400 207.600 312.000 ;
        RECT 221.100 305.400 222.900 312.000 ;
        RECT 224.100 305.400 225.900 311.400 ;
        RECT 227.100 305.400 228.900 312.000 ;
        RECT 242.100 305.400 243.900 311.400 ;
        RECT 245.100 305.400 246.900 312.000 ;
        RECT 200.100 292.050 201.300 299.400 ;
        RECT 206.100 292.050 207.900 293.850 ;
        RECT 224.100 292.050 225.300 305.400 ;
        RECT 242.700 292.050 243.900 305.400 ;
        RECT 261.000 300.600 262.800 311.400 ;
        RECT 261.000 299.400 264.600 300.600 ;
        RECT 266.100 299.400 267.900 312.000 ;
        RECT 284.700 305.400 286.500 312.000 ;
        RECT 285.000 302.100 286.800 303.900 ;
        RECT 287.700 300.900 289.500 311.400 ;
        RECT 287.100 299.400 289.500 300.900 ;
        RECT 292.800 299.400 294.600 312.000 ;
        RECT 311.100 305.400 312.900 312.000 ;
        RECT 314.100 305.400 315.900 311.400 ;
        RECT 329.100 305.400 330.900 312.000 ;
        RECT 332.100 305.400 333.900 311.400 ;
        RECT 245.100 292.050 246.900 293.850 ;
        RECT 260.100 292.050 261.900 293.850 ;
        RECT 263.700 292.050 264.600 299.400 ;
        RECT 265.950 292.050 267.750 293.850 ;
        RECT 287.100 292.050 288.300 299.400 ;
        RECT 293.100 292.050 294.900 293.850 ;
        RECT 311.100 292.050 312.900 293.850 ;
        RECT 314.100 292.050 315.300 305.400 ;
        RECT 329.100 292.050 330.900 293.850 ;
        RECT 332.100 292.050 333.300 305.400 ;
        RECT 350.100 300.300 351.900 311.400 ;
        RECT 353.100 301.200 354.900 312.000 ;
        RECT 356.100 300.300 357.900 311.400 ;
        RECT 350.100 299.400 357.900 300.300 ;
        RECT 359.100 299.400 360.900 311.400 ;
        RECT 374.100 305.400 375.900 312.000 ;
        RECT 377.100 305.400 378.900 311.400 ;
        RECT 380.100 306.000 381.900 312.000 ;
        RECT 377.400 305.100 378.900 305.400 ;
        RECT 383.100 305.400 384.900 311.400 ;
        RECT 383.100 305.100 384.000 305.400 ;
        RECT 377.400 304.200 384.000 305.100 ;
        RECT 353.250 292.050 355.050 293.850 ;
        RECT 359.700 292.050 360.600 299.400 ;
        RECT 377.100 292.050 378.900 293.850 ;
        RECT 383.100 292.050 384.000 304.200 ;
        RECT 401.400 299.400 403.200 312.000 ;
        RECT 406.500 300.900 408.300 311.400 ;
        RECT 409.500 305.400 411.300 312.000 ;
        RECT 425.100 305.400 426.900 312.000 ;
        RECT 428.100 305.400 429.900 311.400 ;
        RECT 446.100 305.400 447.900 312.000 ;
        RECT 449.100 305.400 450.900 311.400 ;
        RECT 409.200 302.100 411.000 303.900 ;
        RECT 406.500 299.400 408.900 300.900 ;
        RECT 401.100 292.050 402.900 293.850 ;
        RECT 407.700 292.050 408.900 299.400 ;
        RECT 425.100 292.050 426.900 293.850 ;
        RECT 428.100 292.050 429.300 305.400 ;
        RECT 130.500 289.950 132.600 292.050 ;
        RECT 133.800 289.950 135.900 292.050 ;
        RECT 148.950 289.950 151.050 292.050 ;
        RECT 151.950 289.950 154.050 292.050 ;
        RECT 154.950 289.950 157.050 292.050 ;
        RECT 169.950 289.950 172.050 292.050 ;
        RECT 172.950 289.950 175.050 292.050 ;
        RECT 175.950 289.950 178.050 292.050 ;
        RECT 178.950 289.950 181.050 292.050 ;
        RECT 196.950 289.950 199.050 292.050 ;
        RECT 199.950 289.950 202.050 292.050 ;
        RECT 202.950 289.950 205.050 292.050 ;
        RECT 205.950 289.950 208.050 292.050 ;
        RECT 220.950 289.950 223.050 292.050 ;
        RECT 223.950 289.950 226.050 292.050 ;
        RECT 226.950 289.950 229.050 292.050 ;
        RECT 241.950 289.950 244.050 292.050 ;
        RECT 244.950 289.950 247.050 292.050 ;
        RECT 259.950 289.950 262.050 292.050 ;
        RECT 262.950 289.950 265.050 292.050 ;
        RECT 265.950 289.950 268.050 292.050 ;
        RECT 283.950 289.950 286.050 292.050 ;
        RECT 286.950 289.950 289.050 292.050 ;
        RECT 289.950 289.950 292.050 292.050 ;
        RECT 292.950 289.950 295.050 292.050 ;
        RECT 310.950 289.950 313.050 292.050 ;
        RECT 313.950 289.950 316.050 292.050 ;
        RECT 328.950 289.950 331.050 292.050 ;
        RECT 331.950 289.950 334.050 292.050 ;
        RECT 349.950 289.950 352.050 292.050 ;
        RECT 352.950 289.950 355.050 292.050 ;
        RECT 355.950 289.950 358.050 292.050 ;
        RECT 358.950 289.950 361.050 292.050 ;
        RECT 373.950 289.950 376.050 292.050 ;
        RECT 376.950 289.950 379.050 292.050 ;
        RECT 379.950 289.950 382.050 292.050 ;
        RECT 382.950 289.950 385.050 292.050 ;
        RECT 400.950 289.950 403.050 292.050 ;
        RECT 403.950 289.950 406.050 292.050 ;
        RECT 406.950 289.950 409.050 292.050 ;
        RECT 409.950 289.950 412.050 292.050 ;
        RECT 424.950 289.950 427.050 292.050 ;
        RECT 427.950 289.950 430.050 292.050 ;
        RECT 446.100 289.950 448.200 292.050 ;
        RECT 107.100 283.800 111.300 284.700 ;
        RECT 73.200 279.600 74.250 280.500 ;
        RECT 82.050 280.200 84.150 281.700 ;
        RECT 80.250 279.600 84.150 280.200 ;
        RECT 64.950 276.600 66.750 279.600 ;
        RECT 69.450 276.000 71.250 279.600 ;
        RECT 72.450 276.600 74.250 279.600 ;
        RECT 75.750 276.000 77.550 279.600 ;
        RECT 80.250 278.700 83.850 279.600 ;
        RECT 80.250 276.600 82.050 278.700 ;
        RECT 85.050 276.000 86.850 282.600 ;
        RECT 88.050 280.800 90.450 282.600 ;
        RECT 88.050 276.600 89.850 280.800 ;
        RECT 104.400 276.000 106.200 282.600 ;
        RECT 109.500 276.600 111.300 283.800 ;
        RECT 125.100 284.400 133.500 285.300 ;
        RECT 125.100 276.600 126.900 284.400 ;
        RECT 131.700 283.500 133.500 284.400 ;
        RECT 134.400 282.600 135.300 289.950 ;
        RECT 129.600 276.000 131.400 282.600 ;
        RECT 132.600 280.800 135.300 282.600 ;
        RECT 132.600 276.600 134.400 280.800 ;
        RECT 152.400 279.600 153.300 289.950 ;
        RECT 160.950 288.450 163.050 289.050 ;
        RECT 166.950 288.450 169.050 289.050 ;
        RECT 160.950 287.550 169.050 288.450 ;
        RECT 173.100 288.150 174.900 289.950 ;
        RECT 160.950 286.950 163.050 287.550 ;
        RECT 166.950 286.950 169.050 287.550 ;
        RECT 154.950 285.450 157.050 286.050 ;
        RECT 163.950 285.450 166.050 286.050 ;
        RECT 154.950 284.550 166.050 285.450 ;
        RECT 176.700 285.600 177.900 289.950 ;
        RECT 179.100 288.150 180.900 289.950 ;
        RECT 197.100 288.150 198.900 289.950 ;
        RECT 200.100 285.600 201.300 289.950 ;
        RECT 203.100 288.150 204.900 289.950 ;
        RECT 221.250 288.150 223.050 289.950 ;
        RECT 176.700 284.700 180.300 285.600 ;
        RECT 154.950 283.950 157.050 284.550 ;
        RECT 163.950 283.950 166.050 284.550 ;
        RECT 170.100 281.700 177.900 283.050 ;
        RECT 149.100 276.000 150.900 279.600 ;
        RECT 152.100 276.600 153.900 279.600 ;
        RECT 155.100 276.000 156.900 279.600 ;
        RECT 170.100 276.600 171.900 281.700 ;
        RECT 173.100 276.000 174.900 280.800 ;
        RECT 176.100 276.600 177.900 281.700 ;
        RECT 179.100 282.600 180.300 284.700 ;
        RECT 197.700 284.700 201.300 285.600 ;
        RECT 224.100 284.700 225.300 289.950 ;
        RECT 227.100 288.150 228.900 289.950 ;
        RECT 197.700 282.600 198.900 284.700 ;
        RECT 224.100 283.800 228.300 284.700 ;
        RECT 179.100 276.600 180.900 282.600 ;
        RECT 197.100 276.600 198.900 282.600 ;
        RECT 200.100 281.700 207.900 283.050 ;
        RECT 200.100 276.600 201.900 281.700 ;
        RECT 203.100 276.000 204.900 280.800 ;
        RECT 206.100 276.600 207.900 281.700 ;
        RECT 221.400 276.000 223.200 282.600 ;
        RECT 226.500 276.600 228.300 283.800 ;
        RECT 242.700 279.600 243.900 289.950 ;
        RECT 263.700 279.600 264.600 289.950 ;
        RECT 284.100 288.150 285.900 289.950 ;
        RECT 287.100 285.600 288.300 289.950 ;
        RECT 290.100 288.150 291.900 289.950 ;
        RECT 284.700 284.700 288.300 285.600 ;
        RECT 268.950 282.450 271.050 283.050 ;
        RECT 277.950 282.450 280.050 283.050 ;
        RECT 284.700 282.600 285.900 284.700 ;
        RECT 268.950 281.550 280.050 282.450 ;
        RECT 268.950 280.950 271.050 281.550 ;
        RECT 277.950 280.950 280.050 281.550 ;
        RECT 242.100 276.600 243.900 279.600 ;
        RECT 245.100 276.000 246.900 279.600 ;
        RECT 260.100 276.000 261.900 279.600 ;
        RECT 263.100 276.600 264.900 279.600 ;
        RECT 266.100 276.000 267.900 279.600 ;
        RECT 284.100 276.600 285.900 282.600 ;
        RECT 287.100 281.700 294.900 283.050 ;
        RECT 287.100 276.600 288.900 281.700 ;
        RECT 290.100 276.000 291.900 280.800 ;
        RECT 293.100 276.600 294.900 281.700 ;
        RECT 314.100 279.600 315.300 289.950 ;
        RECT 332.100 279.600 333.300 289.950 ;
        RECT 350.100 288.150 351.900 289.950 ;
        RECT 356.250 288.150 358.050 289.950 ;
        RECT 359.700 282.600 360.600 289.950 ;
        RECT 374.100 288.150 375.900 289.950 ;
        RECT 380.100 288.150 381.900 289.950 ;
        RECT 383.100 286.200 384.000 289.950 ;
        RECT 404.100 288.150 405.900 289.950 ;
        RECT 311.100 276.000 312.900 279.600 ;
        RECT 314.100 276.600 315.900 279.600 ;
        RECT 329.100 276.000 330.900 279.600 ;
        RECT 332.100 276.600 333.900 279.600 ;
        RECT 351.000 276.000 352.800 282.600 ;
        RECT 355.500 281.400 360.600 282.600 ;
        RECT 355.500 276.600 357.300 281.400 ;
        RECT 358.500 276.000 360.300 279.600 ;
        RECT 374.100 276.000 375.900 285.600 ;
        RECT 380.700 285.000 384.000 286.200 ;
        RECT 407.700 285.600 408.900 289.950 ;
        RECT 410.100 288.150 411.900 289.950 ;
        RECT 380.700 276.600 382.500 285.000 ;
        RECT 407.700 284.700 411.300 285.600 ;
        RECT 401.100 281.700 408.900 283.050 ;
        RECT 401.100 276.600 402.900 281.700 ;
        RECT 404.100 276.000 405.900 280.800 ;
        RECT 407.100 276.600 408.900 281.700 ;
        RECT 410.100 282.600 411.300 284.700 ;
        RECT 410.100 276.600 411.900 282.600 ;
        RECT 428.100 279.600 429.300 289.950 ;
        RECT 446.250 288.150 448.050 289.950 ;
        RECT 449.100 285.300 450.000 305.400 ;
        RECT 452.100 300.000 453.900 312.000 ;
        RECT 455.100 299.400 456.900 311.400 ;
        RECT 470.100 305.400 471.900 312.000 ;
        RECT 473.100 305.400 474.900 311.400 ;
        RECT 476.100 306.000 477.900 312.000 ;
        RECT 473.400 305.100 474.900 305.400 ;
        RECT 479.100 305.400 480.900 311.400 ;
        RECT 479.100 305.100 480.000 305.400 ;
        RECT 473.400 304.200 480.000 305.100 ;
        RECT 469.950 300.450 472.050 301.050 ;
        RECT 475.950 300.450 478.050 301.050 ;
        RECT 469.950 299.550 478.050 300.450 ;
        RECT 451.200 292.050 453.000 293.850 ;
        RECT 455.400 292.050 456.300 299.400 ;
        RECT 469.950 298.950 472.050 299.550 ;
        RECT 475.950 298.950 478.050 299.550 ;
        RECT 473.100 292.050 474.900 293.850 ;
        RECT 479.100 292.050 480.000 304.200 ;
        RECT 494.400 299.400 496.200 312.000 ;
        RECT 499.500 300.900 501.300 311.400 ;
        RECT 502.500 305.400 504.300 312.000 ;
        RECT 521.100 310.500 528.900 311.400 ;
        RECT 502.200 302.100 504.000 303.900 ;
        RECT 499.500 299.400 501.900 300.900 ;
        RECT 521.100 299.400 522.900 310.500 ;
        RECT 494.100 292.050 495.900 293.850 ;
        RECT 500.700 292.050 501.900 299.400 ;
        RECT 524.100 298.500 525.900 309.600 ;
        RECT 527.100 300.600 528.900 310.500 ;
        RECT 530.100 301.500 531.900 312.000 ;
        RECT 533.100 300.600 534.900 311.400 ;
        RECT 548.100 305.400 549.900 312.000 ;
        RECT 551.100 305.400 552.900 311.400 ;
        RECT 554.100 305.400 555.900 312.000 ;
        RECT 569.100 305.400 570.900 312.000 ;
        RECT 572.100 305.400 573.900 311.400 ;
        RECT 575.100 306.000 576.900 312.000 ;
        RECT 527.100 299.700 534.900 300.600 ;
        RECT 524.100 297.600 528.900 298.500 ;
        RECT 524.100 292.050 525.900 293.850 ;
        RECT 528.000 292.050 528.900 297.600 ;
        RECT 529.950 292.050 531.750 293.850 ;
        RECT 551.700 292.050 552.900 305.400 ;
        RECT 572.400 305.100 573.900 305.400 ;
        RECT 578.100 305.400 579.900 311.400 ;
        RECT 593.100 305.400 594.900 311.400 ;
        RECT 596.100 305.400 597.900 312.000 ;
        RECT 611.100 305.400 612.900 312.000 ;
        RECT 614.100 305.400 615.900 311.400 ;
        RECT 578.100 305.100 579.000 305.400 ;
        RECT 572.400 304.200 579.000 305.100 ;
        RECT 553.950 300.450 556.050 301.050 ;
        RECT 568.950 300.450 571.050 301.050 ;
        RECT 553.950 299.550 571.050 300.450 ;
        RECT 553.950 298.950 556.050 299.550 ;
        RECT 568.950 298.950 571.050 299.550 ;
        RECT 574.950 297.450 577.050 298.050 ;
        RECT 566.550 296.550 577.050 297.450 ;
        RECT 566.550 294.450 567.450 296.550 ;
        RECT 574.950 295.950 577.050 296.550 ;
        RECT 563.550 293.550 567.450 294.450 ;
        RECT 451.500 289.950 453.600 292.050 ;
        RECT 454.800 289.950 456.900 292.050 ;
        RECT 469.950 289.950 472.050 292.050 ;
        RECT 472.950 289.950 475.050 292.050 ;
        RECT 475.950 289.950 478.050 292.050 ;
        RECT 478.950 289.950 481.050 292.050 ;
        RECT 493.950 289.950 496.050 292.050 ;
        RECT 496.950 289.950 499.050 292.050 ;
        RECT 499.950 289.950 502.050 292.050 ;
        RECT 502.950 289.950 505.050 292.050 ;
        RECT 520.950 289.950 523.050 292.050 ;
        RECT 523.950 289.950 526.050 292.050 ;
        RECT 526.950 289.950 529.050 292.050 ;
        RECT 529.950 289.950 532.050 292.050 ;
        RECT 532.950 289.950 535.050 292.050 ;
        RECT 547.950 289.950 550.050 292.050 ;
        RECT 550.950 289.950 553.050 292.050 ;
        RECT 553.950 289.950 556.050 292.050 ;
        RECT 446.100 284.400 454.500 285.300 ;
        RECT 425.100 276.000 426.900 279.600 ;
        RECT 428.100 276.600 429.900 279.600 ;
        RECT 446.100 276.600 447.900 284.400 ;
        RECT 452.700 283.500 454.500 284.400 ;
        RECT 455.400 282.600 456.300 289.950 ;
        RECT 470.100 288.150 471.900 289.950 ;
        RECT 476.100 288.150 477.900 289.950 ;
        RECT 479.100 286.200 480.000 289.950 ;
        RECT 497.100 288.150 498.900 289.950 ;
        RECT 450.600 276.000 452.400 282.600 ;
        RECT 453.600 280.800 456.300 282.600 ;
        RECT 453.600 276.600 455.400 280.800 ;
        RECT 470.100 276.000 471.900 285.600 ;
        RECT 476.700 285.000 480.000 286.200 ;
        RECT 500.700 285.600 501.900 289.950 ;
        RECT 503.100 288.150 504.900 289.950 ;
        RECT 521.100 288.150 522.900 289.950 ;
        RECT 476.700 276.600 478.500 285.000 ;
        RECT 500.700 284.700 504.300 285.600 ;
        RECT 494.100 281.700 501.900 283.050 ;
        RECT 494.100 276.600 495.900 281.700 ;
        RECT 497.100 276.000 498.900 280.800 ;
        RECT 500.100 276.600 501.900 281.700 ;
        RECT 503.100 282.600 504.300 284.700 ;
        RECT 527.700 282.600 528.900 289.950 ;
        RECT 532.950 288.150 534.750 289.950 ;
        RECT 548.100 288.150 549.900 289.950 ;
        RECT 551.700 284.700 552.900 289.950 ;
        RECT 553.950 288.150 555.750 289.950 ;
        RECT 563.550 288.450 564.450 293.550 ;
        RECT 572.100 292.050 573.900 293.850 ;
        RECT 578.100 292.050 579.000 304.200 ;
        RECT 593.700 292.050 594.900 305.400 ;
        RECT 596.100 292.050 597.900 293.850 ;
        RECT 568.950 289.950 571.050 292.050 ;
        RECT 571.950 289.950 574.050 292.050 ;
        RECT 574.950 289.950 577.050 292.050 ;
        RECT 577.950 289.950 580.050 292.050 ;
        RECT 592.950 289.950 595.050 292.050 ;
        RECT 595.950 289.950 598.050 292.050 ;
        RECT 611.100 289.950 613.200 292.050 ;
        RECT 557.550 288.000 564.450 288.450 ;
        RECT 569.100 288.150 570.900 289.950 ;
        RECT 575.100 288.150 576.900 289.950 ;
        RECT 548.700 283.800 552.900 284.700 ;
        RECT 556.950 287.550 564.450 288.000 ;
        RECT 556.950 283.950 559.050 287.550 ;
        RECT 578.100 286.200 579.000 289.950 ;
        RECT 503.100 276.600 504.900 282.600 ;
        RECT 523.500 276.000 525.300 282.600 ;
        RECT 528.000 276.600 529.800 282.600 ;
        RECT 532.500 276.000 534.300 282.600 ;
        RECT 538.950 282.450 541.050 282.900 ;
        RECT 544.950 282.450 547.050 283.050 ;
        RECT 538.950 281.550 547.050 282.450 ;
        RECT 538.950 280.800 541.050 281.550 ;
        RECT 544.950 280.950 547.050 281.550 ;
        RECT 548.700 276.600 550.500 283.800 ;
        RECT 553.800 276.000 555.600 282.600 ;
        RECT 556.950 279.450 559.050 280.050 ;
        RECT 562.950 279.450 565.050 280.050 ;
        RECT 556.950 278.550 565.050 279.450 ;
        RECT 556.950 277.950 559.050 278.550 ;
        RECT 562.950 277.950 565.050 278.550 ;
        RECT 569.100 276.000 570.900 285.600 ;
        RECT 575.700 285.000 579.000 286.200 ;
        RECT 575.700 276.600 577.500 285.000 ;
        RECT 593.700 279.600 594.900 289.950 ;
        RECT 611.250 288.150 613.050 289.950 ;
        RECT 614.100 285.300 615.000 305.400 ;
        RECT 617.100 300.000 618.900 312.000 ;
        RECT 620.100 299.400 621.900 311.400 ;
        RECT 638.100 305.400 639.900 312.000 ;
        RECT 641.100 305.400 642.900 311.400 ;
        RECT 644.100 305.400 645.900 312.000 ;
        RECT 659.100 305.400 660.900 312.000 ;
        RECT 662.100 305.400 663.900 311.400 ;
        RECT 665.100 306.000 666.900 312.000 ;
        RECT 616.200 292.050 618.000 293.850 ;
        RECT 620.400 292.050 621.300 299.400 ;
        RECT 641.100 292.050 642.300 305.400 ;
        RECT 662.400 305.100 663.900 305.400 ;
        RECT 668.100 305.400 669.900 311.400 ;
        RECT 683.100 305.400 684.900 312.000 ;
        RECT 686.100 305.400 687.900 311.400 ;
        RECT 689.100 306.000 690.900 312.000 ;
        RECT 668.100 305.100 669.000 305.400 ;
        RECT 662.400 304.200 669.000 305.100 ;
        RECT 686.400 305.100 687.900 305.400 ;
        RECT 692.100 305.400 693.900 311.400 ;
        RECT 707.100 305.400 708.900 312.000 ;
        RECT 710.100 305.400 711.900 311.400 ;
        RECT 713.100 306.000 714.900 312.000 ;
        RECT 692.100 305.100 693.000 305.400 ;
        RECT 686.400 304.200 693.000 305.100 ;
        RECT 710.400 305.100 711.900 305.400 ;
        RECT 716.100 305.400 717.900 311.400 ;
        RECT 734.100 305.400 735.900 312.000 ;
        RECT 737.100 305.400 738.900 311.400 ;
        RECT 740.100 305.400 741.900 312.000 ;
        RECT 716.100 305.100 717.000 305.400 ;
        RECT 710.400 304.200 717.000 305.100 ;
        RECT 662.100 292.050 663.900 293.850 ;
        RECT 668.100 292.050 669.000 304.200 ;
        RECT 686.100 292.050 687.900 293.850 ;
        RECT 692.100 292.050 693.000 304.200 ;
        RECT 710.100 292.050 711.900 293.850 ;
        RECT 716.100 292.050 717.000 304.200 ;
        RECT 737.100 292.050 738.300 305.400 ;
        RECT 755.100 299.400 756.900 311.400 ;
        RECT 758.100 300.300 759.900 311.400 ;
        RECT 761.100 301.200 762.900 312.000 ;
        RECT 764.100 300.300 765.900 311.400 ;
        RECT 779.100 305.400 780.900 312.000 ;
        RECT 782.100 305.400 783.900 311.400 ;
        RECT 785.100 306.000 786.900 312.000 ;
        RECT 782.400 305.100 783.900 305.400 ;
        RECT 788.100 305.400 789.900 311.400 ;
        RECT 803.100 305.400 804.900 311.400 ;
        RECT 806.100 306.000 807.900 312.000 ;
        RECT 788.100 305.100 789.000 305.400 ;
        RECT 782.400 304.200 789.000 305.100 ;
        RECT 758.100 299.400 765.900 300.300 ;
        RECT 750.000 294.450 754.050 295.050 ;
        RECT 749.550 292.950 754.050 294.450 ;
        RECT 616.500 289.950 618.600 292.050 ;
        RECT 619.800 289.950 621.900 292.050 ;
        RECT 637.950 289.950 640.050 292.050 ;
        RECT 640.950 289.950 643.050 292.050 ;
        RECT 643.950 289.950 646.050 292.050 ;
        RECT 658.950 289.950 661.050 292.050 ;
        RECT 661.950 289.950 664.050 292.050 ;
        RECT 664.950 289.950 667.050 292.050 ;
        RECT 667.950 289.950 670.050 292.050 ;
        RECT 682.950 289.950 685.050 292.050 ;
        RECT 685.950 289.950 688.050 292.050 ;
        RECT 688.950 289.950 691.050 292.050 ;
        RECT 691.950 289.950 694.050 292.050 ;
        RECT 706.950 289.950 709.050 292.050 ;
        RECT 709.950 289.950 712.050 292.050 ;
        RECT 712.950 289.950 715.050 292.050 ;
        RECT 715.950 289.950 718.050 292.050 ;
        RECT 733.950 289.950 736.050 292.050 ;
        RECT 736.950 289.950 739.050 292.050 ;
        RECT 739.950 289.950 742.050 292.050 ;
        RECT 611.100 284.400 619.500 285.300 ;
        RECT 593.100 276.600 594.900 279.600 ;
        RECT 596.100 276.000 597.900 279.600 ;
        RECT 611.100 276.600 612.900 284.400 ;
        RECT 617.700 283.500 619.500 284.400 ;
        RECT 620.400 282.600 621.300 289.950 ;
        RECT 625.950 288.450 628.050 289.050 ;
        RECT 625.950 288.000 636.450 288.450 ;
        RECT 638.250 288.150 640.050 289.950 ;
        RECT 625.950 287.550 637.050 288.000 ;
        RECT 625.950 286.950 628.050 287.550 ;
        RECT 634.950 283.950 637.050 287.550 ;
        RECT 641.100 284.700 642.300 289.950 ;
        RECT 644.100 288.150 645.900 289.950 ;
        RECT 659.100 288.150 660.900 289.950 ;
        RECT 665.100 288.150 666.900 289.950 ;
        RECT 668.100 286.200 669.000 289.950 ;
        RECT 683.100 288.150 684.900 289.950 ;
        RECT 689.100 288.150 690.900 289.950 ;
        RECT 692.100 286.200 693.000 289.950 ;
        RECT 707.100 288.150 708.900 289.950 ;
        RECT 713.100 288.150 714.900 289.950 ;
        RECT 716.100 286.200 717.000 289.950 ;
        RECT 734.250 288.150 736.050 289.950 ;
        RECT 641.100 283.800 645.300 284.700 ;
        RECT 615.600 276.000 617.400 282.600 ;
        RECT 618.600 280.800 621.300 282.600 ;
        RECT 618.600 276.600 620.400 280.800 ;
        RECT 638.400 276.000 640.200 282.600 ;
        RECT 643.500 276.600 645.300 283.800 ;
        RECT 659.100 276.000 660.900 285.600 ;
        RECT 665.700 285.000 669.000 286.200 ;
        RECT 665.700 276.600 667.500 285.000 ;
        RECT 683.100 276.000 684.900 285.600 ;
        RECT 689.700 285.000 693.000 286.200 ;
        RECT 689.700 276.600 691.500 285.000 ;
        RECT 707.100 276.000 708.900 285.600 ;
        RECT 713.700 285.000 717.000 286.200 ;
        RECT 713.700 276.600 715.500 285.000 ;
        RECT 737.100 284.700 738.300 289.950 ;
        RECT 740.100 288.150 741.900 289.950 ;
        RECT 749.550 289.050 750.450 292.950 ;
        RECT 755.400 292.050 756.300 299.400 ;
        RECT 760.950 292.050 762.750 293.850 ;
        RECT 782.100 292.050 783.900 293.850 ;
        RECT 788.100 292.050 789.000 304.200 ;
        RECT 804.000 305.100 804.900 305.400 ;
        RECT 809.100 305.400 810.900 311.400 ;
        RECT 812.100 305.400 813.900 312.000 ;
        RECT 827.700 305.400 829.500 312.000 ;
        RECT 809.100 305.100 810.600 305.400 ;
        RECT 804.000 304.200 810.600 305.100 ;
        RECT 804.000 292.050 804.900 304.200 ;
        RECT 828.000 302.100 829.800 303.900 ;
        RECT 830.700 300.900 832.500 311.400 ;
        RECT 830.100 299.400 832.500 300.900 ;
        RECT 835.800 299.400 837.600 312.000 ;
        RECT 854.100 300.300 855.900 311.400 ;
        RECT 857.100 301.200 858.900 312.000 ;
        RECT 860.100 300.300 861.900 311.400 ;
        RECT 854.100 299.400 861.900 300.300 ;
        RECT 863.100 299.400 864.900 311.400 ;
        RECT 878.100 305.400 879.900 311.400 ;
        RECT 881.100 306.000 882.900 312.000 ;
        RECT 879.000 305.100 879.900 305.400 ;
        RECT 884.100 305.400 885.900 311.400 ;
        RECT 887.100 305.400 888.900 312.000 ;
        RECT 884.100 305.100 885.600 305.400 ;
        RECT 879.000 304.200 885.600 305.100 ;
        RECT 809.100 292.050 810.900 293.850 ;
        RECT 830.100 292.050 831.300 299.400 ;
        RECT 832.950 297.450 835.050 298.050 ;
        RECT 856.950 297.450 859.050 298.050 ;
        RECT 832.950 296.550 859.050 297.450 ;
        RECT 832.950 295.950 835.050 296.550 ;
        RECT 856.950 295.950 859.050 296.550 ;
        RECT 850.950 294.450 853.050 295.050 ;
        RECT 836.100 292.050 837.900 293.850 ;
        RECT 842.550 293.550 853.050 294.450 ;
        RECT 754.950 289.950 757.050 292.050 ;
        RECT 757.950 289.950 760.050 292.050 ;
        RECT 760.950 289.950 763.050 292.050 ;
        RECT 763.950 289.950 766.050 292.050 ;
        RECT 778.950 289.950 781.050 292.050 ;
        RECT 781.950 289.950 784.050 292.050 ;
        RECT 784.950 289.950 787.050 292.050 ;
        RECT 787.950 289.950 790.050 292.050 ;
        RECT 802.950 289.950 805.050 292.050 ;
        RECT 805.950 289.950 808.050 292.050 ;
        RECT 808.950 289.950 811.050 292.050 ;
        RECT 811.950 289.950 814.050 292.050 ;
        RECT 826.950 289.950 829.050 292.050 ;
        RECT 829.950 289.950 832.050 292.050 ;
        RECT 832.950 289.950 835.050 292.050 ;
        RECT 835.950 289.950 838.050 292.050 ;
        RECT 749.550 287.550 754.050 289.050 ;
        RECT 750.000 286.950 754.050 287.550 ;
        RECT 737.100 283.800 741.300 284.700 ;
        RECT 718.950 279.450 721.050 280.050 ;
        RECT 727.950 279.450 730.050 280.050 ;
        RECT 718.950 278.550 730.050 279.450 ;
        RECT 718.950 277.950 721.050 278.550 ;
        RECT 727.950 277.950 730.050 278.550 ;
        RECT 734.400 276.000 736.200 282.600 ;
        RECT 739.500 276.600 741.300 283.800 ;
        RECT 755.400 282.600 756.300 289.950 ;
        RECT 757.950 288.150 759.750 289.950 ;
        RECT 764.100 288.150 765.900 289.950 ;
        RECT 779.100 288.150 780.900 289.950 ;
        RECT 785.100 288.150 786.900 289.950 ;
        RECT 788.100 286.200 789.000 289.950 ;
        RECT 755.400 281.400 760.500 282.600 ;
        RECT 755.700 276.000 757.500 279.600 ;
        RECT 758.700 276.600 760.500 281.400 ;
        RECT 763.200 276.000 765.000 282.600 ;
        RECT 779.100 276.000 780.900 285.600 ;
        RECT 785.700 285.000 789.000 286.200 ;
        RECT 804.000 286.200 804.900 289.950 ;
        RECT 806.100 288.150 807.900 289.950 ;
        RECT 812.100 288.150 813.900 289.950 ;
        RECT 827.100 288.150 828.900 289.950 ;
        RECT 804.000 285.000 807.300 286.200 ;
        RECT 830.100 285.600 831.300 289.950 ;
        RECT 833.100 288.150 834.900 289.950 ;
        RECT 842.550 289.050 843.450 293.550 ;
        RECT 850.950 292.950 853.050 293.550 ;
        RECT 857.250 292.050 859.050 293.850 ;
        RECT 863.700 292.050 864.600 299.400 ;
        RECT 879.000 292.050 879.900 304.200 ;
        RECT 886.950 297.450 889.050 298.200 ;
        RECT 892.950 297.450 895.050 297.900 ;
        RECT 886.950 296.550 895.050 297.450 ;
        RECT 886.950 296.100 889.050 296.550 ;
        RECT 892.950 295.800 895.050 296.550 ;
        RECT 884.100 292.050 885.900 293.850 ;
        RECT 853.950 289.950 856.050 292.050 ;
        RECT 856.950 289.950 859.050 292.050 ;
        RECT 859.950 289.950 862.050 292.050 ;
        RECT 862.950 289.950 865.050 292.050 ;
        RECT 877.950 289.950 880.050 292.050 ;
        RECT 880.950 289.950 883.050 292.050 ;
        RECT 883.950 289.950 886.050 292.050 ;
        RECT 886.950 289.950 889.050 292.050 ;
        RECT 838.950 287.550 843.450 289.050 ;
        RECT 854.100 288.150 855.900 289.950 ;
        RECT 860.250 288.150 862.050 289.950 ;
        RECT 838.950 286.950 843.000 287.550 ;
        RECT 785.700 276.600 787.500 285.000 ;
        RECT 805.500 276.600 807.300 285.000 ;
        RECT 812.100 276.000 813.900 285.600 ;
        RECT 827.700 284.700 831.300 285.600 ;
        RECT 839.550 285.450 840.450 286.950 ;
        RECT 853.950 285.450 856.050 286.050 ;
        RECT 827.700 282.600 828.900 284.700 ;
        RECT 839.550 284.550 856.050 285.450 ;
        RECT 853.950 283.950 856.050 284.550 ;
        RECT 827.100 276.600 828.900 282.600 ;
        RECT 830.100 281.700 837.900 283.050 ;
        RECT 863.700 282.600 864.600 289.950 ;
        RECT 879.000 286.200 879.900 289.950 ;
        RECT 881.100 288.150 882.900 289.950 ;
        RECT 887.100 288.150 888.900 289.950 ;
        RECT 879.000 285.000 882.300 286.200 ;
        RECT 830.100 276.600 831.900 281.700 ;
        RECT 833.100 276.000 834.900 280.800 ;
        RECT 836.100 276.600 837.900 281.700 ;
        RECT 855.000 276.000 856.800 282.600 ;
        RECT 859.500 281.400 864.600 282.600 ;
        RECT 859.500 276.600 861.300 281.400 ;
        RECT 862.500 276.000 864.300 279.600 ;
        RECT 880.500 276.600 882.300 285.000 ;
        RECT 887.100 276.000 888.900 285.600 ;
        RECT 17.100 267.300 18.900 272.400 ;
        RECT 20.100 268.200 21.900 273.000 ;
        RECT 23.100 267.300 24.900 272.400 ;
        RECT 17.100 265.950 24.900 267.300 ;
        RECT 26.100 266.400 27.900 272.400 ;
        RECT 41.100 269.400 42.900 273.000 ;
        RECT 44.100 269.400 45.900 272.400 ;
        RECT 26.100 264.300 27.300 266.400 ;
        RECT 23.700 263.400 27.300 264.300 ;
        RECT 20.100 259.050 21.900 260.850 ;
        RECT 23.700 259.050 24.900 263.400 ;
        RECT 28.950 261.450 33.000 262.050 ;
        RECT 26.100 259.050 27.900 260.850 ;
        RECT 28.950 259.950 33.450 261.450 ;
        RECT 16.950 256.950 19.050 259.050 ;
        RECT 19.950 256.950 22.050 259.050 ;
        RECT 22.950 256.950 25.050 259.050 ;
        RECT 25.950 256.950 28.050 259.050 ;
        RECT 17.100 255.150 18.900 256.950 ;
        RECT 23.700 249.600 24.900 256.950 ;
        RECT 32.550 252.900 33.450 259.950 ;
        RECT 44.100 259.050 45.300 269.400 ;
        RECT 59.100 267.300 60.900 272.400 ;
        RECT 62.100 268.200 63.900 273.000 ;
        RECT 65.100 267.300 66.900 272.400 ;
        RECT 59.100 265.950 66.900 267.300 ;
        RECT 68.100 266.400 69.900 272.400 ;
        RECT 86.100 269.400 87.900 272.400 ;
        RECT 89.100 269.400 90.900 273.000 ;
        RECT 68.100 264.300 69.300 266.400 ;
        RECT 65.700 263.400 69.300 264.300 ;
        RECT 62.100 259.050 63.900 260.850 ;
        RECT 65.700 259.050 66.900 263.400 ;
        RECT 68.100 259.050 69.900 260.850 ;
        RECT 86.700 259.050 87.900 269.400 ;
        RECT 104.100 263.400 105.900 273.000 ;
        RECT 110.700 264.000 112.500 272.400 ;
        RECT 116.550 266.400 118.350 272.400 ;
        RECT 119.850 266.400 121.650 273.000 ;
        RECT 124.950 269.400 126.750 272.400 ;
        RECT 129.450 269.400 131.250 273.000 ;
        RECT 132.450 269.400 134.250 272.400 ;
        RECT 135.750 269.400 137.550 273.000 ;
        RECT 140.250 270.300 142.050 272.400 ;
        RECT 140.250 269.400 143.850 270.300 ;
        RECT 124.350 267.300 126.750 269.400 ;
        RECT 133.200 268.500 134.250 269.400 ;
        RECT 140.250 268.800 144.150 269.400 ;
        RECT 133.200 267.450 138.150 268.500 ;
        RECT 136.350 266.700 138.150 267.450 ;
        RECT 110.700 262.800 114.000 264.000 ;
        RECT 104.100 259.050 105.900 260.850 ;
        RECT 110.100 259.050 111.900 260.850 ;
        RECT 113.100 259.050 114.000 262.800 ;
        RECT 116.550 259.050 117.750 266.400 ;
        RECT 139.350 265.800 141.150 267.600 ;
        RECT 142.050 267.300 144.150 268.800 ;
        RECT 145.050 266.400 146.850 273.000 ;
        RECT 148.050 268.200 149.850 272.400 ;
        RECT 167.100 269.400 168.900 272.400 ;
        RECT 170.100 269.400 171.900 273.000 ;
        RECT 148.050 266.400 150.450 268.200 ;
        RECT 129.150 264.000 130.950 264.600 ;
        RECT 140.100 264.000 141.150 265.800 ;
        RECT 129.150 262.800 141.150 264.000 ;
        RECT 40.950 256.950 43.050 259.050 ;
        RECT 43.950 256.950 46.050 259.050 ;
        RECT 58.950 256.950 61.050 259.050 ;
        RECT 61.950 256.950 64.050 259.050 ;
        RECT 64.950 256.950 67.050 259.050 ;
        RECT 67.950 256.950 70.050 259.050 ;
        RECT 85.950 256.950 88.050 259.050 ;
        RECT 88.950 256.950 91.050 259.050 ;
        RECT 103.950 256.950 106.050 259.050 ;
        RECT 106.950 256.950 109.050 259.050 ;
        RECT 109.950 256.950 112.050 259.050 ;
        RECT 112.950 256.950 115.050 259.050 ;
        RECT 116.550 257.250 122.850 259.050 ;
        RECT 116.550 256.950 121.050 257.250 ;
        RECT 41.100 255.150 42.900 256.950 ;
        RECT 31.950 250.800 34.050 252.900 ;
        RECT 17.400 237.000 19.200 249.600 ;
        RECT 22.500 248.100 24.900 249.600 ;
        RECT 22.500 237.600 24.300 248.100 ;
        RECT 25.200 245.100 27.000 246.900 ;
        RECT 44.100 243.600 45.300 256.950 ;
        RECT 59.100 255.150 60.900 256.950 ;
        RECT 65.700 249.600 66.900 256.950 ;
        RECT 73.950 255.450 76.050 256.050 ;
        RECT 82.950 255.450 85.050 256.050 ;
        RECT 73.950 254.550 85.050 255.450 ;
        RECT 73.950 253.950 76.050 254.550 ;
        RECT 82.950 253.950 85.050 254.550 ;
        RECT 25.500 237.000 27.300 243.600 ;
        RECT 41.100 237.000 42.900 243.600 ;
        RECT 44.100 237.600 45.900 243.600 ;
        RECT 59.400 237.000 61.200 249.600 ;
        RECT 64.500 248.100 66.900 249.600 ;
        RECT 64.500 237.600 66.300 248.100 ;
        RECT 67.200 245.100 69.000 246.900 ;
        RECT 86.700 243.600 87.900 256.950 ;
        RECT 89.100 255.150 90.900 256.950 ;
        RECT 107.100 255.150 108.900 256.950 ;
        RECT 113.100 244.800 114.000 256.950 ;
        RECT 107.400 243.900 114.000 244.800 ;
        RECT 107.400 243.600 108.900 243.900 ;
        RECT 67.500 237.000 69.300 243.600 ;
        RECT 86.100 237.600 87.900 243.600 ;
        RECT 89.100 237.000 90.900 243.600 ;
        RECT 104.100 237.000 105.900 243.600 ;
        RECT 107.100 237.600 108.900 243.600 ;
        RECT 113.100 243.600 114.000 243.900 ;
        RECT 116.550 249.600 117.750 256.950 ;
        RECT 118.650 254.100 120.450 254.250 ;
        RECT 124.350 254.100 126.450 254.400 ;
        RECT 118.650 252.900 126.450 254.100 ;
        RECT 118.650 252.450 120.450 252.900 ;
        RECT 124.350 252.300 126.450 252.900 ;
        RECT 129.150 250.200 130.050 262.800 ;
        RECT 140.100 261.600 148.050 262.800 ;
        RECT 140.100 261.000 141.900 261.600 ;
        RECT 143.100 259.800 144.900 260.400 ;
        RECT 136.800 258.600 144.900 259.800 ;
        RECT 146.250 259.050 148.050 261.600 ;
        RECT 136.800 256.950 138.900 258.600 ;
        RECT 145.950 256.950 148.050 259.050 ;
        RECT 138.750 251.700 140.550 252.000 ;
        RECT 149.550 251.700 150.450 266.400 ;
        RECT 167.700 259.050 168.900 269.400 ;
        RECT 185.100 266.400 186.900 272.400 ;
        RECT 185.700 264.300 186.900 266.400 ;
        RECT 188.100 267.300 189.900 272.400 ;
        RECT 191.100 268.200 192.900 273.000 ;
        RECT 194.100 267.300 195.900 272.400 ;
        RECT 209.100 269.400 210.900 273.000 ;
        RECT 212.100 269.400 213.900 272.400 ;
        RECT 215.100 269.400 216.900 273.000 ;
        RECT 233.100 269.400 234.900 273.000 ;
        RECT 236.100 269.400 237.900 272.400 ;
        RECT 251.100 269.400 252.900 272.400 ;
        RECT 254.100 269.400 255.900 273.000 ;
        RECT 277.200 269.400 279.900 272.400 ;
        RECT 281.100 269.400 282.900 273.000 ;
        RECT 284.100 269.400 285.900 272.400 ;
        RECT 287.100 269.400 289.200 273.000 ;
        RECT 188.100 265.950 195.900 267.300 ;
        RECT 185.700 263.400 189.300 264.300 ;
        RECT 185.100 259.050 186.900 260.850 ;
        RECT 188.100 259.050 189.300 263.400 ;
        RECT 191.100 259.050 192.900 260.850 ;
        RECT 212.400 259.050 213.300 269.400 ;
        RECT 236.100 259.050 237.300 269.400 ;
        RECT 251.700 259.050 252.900 269.400 ;
        RECT 277.200 268.500 278.100 269.400 ;
        RECT 284.400 268.500 285.300 269.400 ;
        RECT 272.700 267.600 285.300 268.500 ;
        RECT 272.700 259.050 273.900 267.600 ;
        RECT 286.950 267.450 289.050 268.050 ;
        RECT 295.950 267.450 298.050 268.050 ;
        RECT 286.950 266.550 298.050 267.450 ;
        RECT 286.950 265.950 289.050 266.550 ;
        RECT 295.950 265.950 298.050 266.550 ;
        RECT 308.100 267.300 309.900 272.400 ;
        RECT 311.100 268.200 312.900 273.000 ;
        RECT 314.100 267.300 315.900 272.400 ;
        RECT 308.100 265.950 315.900 267.300 ;
        RECT 317.100 266.400 318.900 272.400 ;
        RECT 332.100 267.300 333.900 272.400 ;
        RECT 335.100 268.200 336.900 273.000 ;
        RECT 338.100 267.300 339.900 272.400 ;
        RECT 317.100 264.300 318.300 266.400 ;
        RECT 332.100 265.950 339.900 267.300 ;
        RECT 341.100 266.400 342.900 272.400 ;
        RECT 356.700 266.400 358.500 273.000 ;
        RECT 361.200 266.400 363.000 272.400 ;
        RECT 365.700 266.400 367.500 273.000 ;
        RECT 341.100 264.300 342.300 266.400 ;
        RECT 314.700 263.400 318.300 264.300 ;
        RECT 338.700 263.400 342.300 264.300 ;
        RECT 281.250 259.050 283.050 260.850 ;
        RECT 311.100 259.050 312.900 260.850 ;
        RECT 314.700 259.050 315.900 263.400 ;
        RECT 317.100 259.050 318.900 260.850 ;
        RECT 335.100 259.050 336.900 260.850 ;
        RECT 338.700 259.050 339.900 263.400 ;
        RECT 343.950 261.450 348.000 262.050 ;
        RECT 341.100 259.050 342.900 260.850 ;
        RECT 343.950 259.950 348.450 261.450 ;
        RECT 166.950 256.950 169.050 259.050 ;
        RECT 169.950 256.950 172.050 259.050 ;
        RECT 184.950 256.950 187.050 259.050 ;
        RECT 187.950 256.950 190.050 259.050 ;
        RECT 190.950 256.950 193.050 259.050 ;
        RECT 193.950 256.950 196.050 259.050 ;
        RECT 208.950 256.950 211.050 259.050 ;
        RECT 211.950 256.950 214.050 259.050 ;
        RECT 214.950 256.950 217.050 259.050 ;
        RECT 232.950 256.950 235.050 259.050 ;
        RECT 235.950 256.950 238.050 259.050 ;
        RECT 250.950 256.950 253.050 259.050 ;
        RECT 253.950 256.950 256.050 259.050 ;
        RECT 272.400 256.950 274.500 259.050 ;
        RECT 277.950 256.950 280.050 259.050 ;
        RECT 280.950 256.950 283.050 259.050 ;
        RECT 287.100 256.950 289.200 259.050 ;
        RECT 307.950 256.950 310.050 259.050 ;
        RECT 310.950 256.950 313.050 259.050 ;
        RECT 313.950 256.950 316.050 259.050 ;
        RECT 316.950 256.950 319.050 259.050 ;
        RECT 331.950 256.950 334.050 259.050 ;
        RECT 334.950 256.950 337.050 259.050 ;
        RECT 337.950 256.950 340.050 259.050 ;
        RECT 340.950 256.950 343.050 259.050 ;
        RECT 138.750 251.100 150.450 251.700 ;
        RECT 110.100 237.000 111.900 243.000 ;
        RECT 113.100 237.600 114.900 243.600 ;
        RECT 116.550 237.600 118.350 249.600 ;
        RECT 119.550 237.000 121.350 249.600 ;
        RECT 125.250 249.300 130.050 250.200 ;
        RECT 132.150 250.500 150.450 251.100 ;
        RECT 132.150 250.200 140.550 250.500 ;
        RECT 125.250 248.400 126.450 249.300 ;
        RECT 123.450 246.600 126.450 248.400 ;
        RECT 127.350 248.100 129.150 248.400 ;
        RECT 132.150 248.100 133.050 250.200 ;
        RECT 149.550 249.600 150.450 250.500 ;
        RECT 127.350 247.200 133.050 248.100 ;
        RECT 133.950 248.700 135.750 249.300 ;
        RECT 133.950 247.500 141.750 248.700 ;
        RECT 127.350 246.600 129.150 247.200 ;
        RECT 139.650 246.600 141.750 247.500 ;
        RECT 124.350 243.600 126.450 245.700 ;
        RECT 130.950 245.550 132.750 246.300 ;
        RECT 135.750 245.550 137.550 246.300 ;
        RECT 130.950 244.500 137.550 245.550 ;
        RECT 124.350 237.600 126.150 243.600 ;
        RECT 128.850 237.000 130.650 243.600 ;
        RECT 131.850 237.600 133.650 244.500 ;
        RECT 134.850 237.000 136.650 243.600 ;
        RECT 139.650 237.600 141.450 246.600 ;
        RECT 145.050 237.000 146.850 249.600 ;
        RECT 148.050 247.800 150.450 249.600 ;
        RECT 148.050 237.600 149.850 247.800 ;
        RECT 167.700 243.600 168.900 256.950 ;
        RECT 170.100 255.150 171.900 256.950 ;
        RECT 188.100 249.600 189.300 256.950 ;
        RECT 194.100 255.150 195.900 256.950 ;
        RECT 209.250 255.150 211.050 256.950 ;
        RECT 212.400 249.600 213.300 256.950 ;
        RECT 215.100 255.150 216.900 256.950 ;
        RECT 233.100 255.150 234.900 256.950 ;
        RECT 188.100 248.100 190.500 249.600 ;
        RECT 186.000 245.100 187.800 246.900 ;
        RECT 167.100 237.600 168.900 243.600 ;
        RECT 170.100 237.000 171.900 243.600 ;
        RECT 185.700 237.000 187.500 243.600 ;
        RECT 188.700 237.600 190.500 248.100 ;
        RECT 193.800 237.000 195.600 249.600 ;
        RECT 209.100 237.000 210.900 249.600 ;
        RECT 212.400 248.400 216.000 249.600 ;
        RECT 214.200 237.600 216.000 248.400 ;
        RECT 236.100 243.600 237.300 256.950 ;
        RECT 251.700 243.600 252.900 256.950 ;
        RECT 254.100 255.150 255.900 256.950 ;
        RECT 233.100 237.000 234.900 243.600 ;
        RECT 236.100 237.600 237.900 243.600 ;
        RECT 251.100 237.600 252.900 243.600 ;
        RECT 254.100 237.000 255.900 243.600 ;
        RECT 269.100 238.500 270.900 247.800 ;
        RECT 272.700 247.200 273.900 256.950 ;
        RECT 277.950 255.150 279.750 256.950 ;
        RECT 287.100 255.150 288.900 256.950 ;
        RECT 308.100 255.150 309.900 256.950 ;
        RECT 314.700 249.600 315.900 256.950 ;
        RECT 332.100 255.150 333.900 256.950 ;
        RECT 338.700 249.600 339.900 256.950 ;
        RECT 347.550 256.050 348.450 259.950 ;
        RECT 356.250 259.050 358.050 260.850 ;
        RECT 362.100 259.050 363.300 266.400 ;
        RECT 383.100 263.400 384.900 273.000 ;
        RECT 389.700 264.000 391.500 272.400 ;
        RECT 407.100 269.400 408.900 273.000 ;
        RECT 410.100 269.400 411.900 272.400 ;
        RECT 389.700 262.800 393.000 264.000 ;
        RECT 368.100 259.050 369.900 260.850 ;
        RECT 383.100 259.050 384.900 260.850 ;
        RECT 389.100 259.050 390.900 260.850 ;
        RECT 392.100 259.050 393.000 262.800 ;
        RECT 410.100 259.050 411.300 269.400 ;
        RECT 426.600 268.200 428.400 272.400 ;
        RECT 425.700 266.400 428.400 268.200 ;
        RECT 429.600 266.400 431.400 273.000 ;
        RECT 425.700 259.050 426.600 266.400 ;
        RECT 427.500 264.600 429.300 265.500 ;
        RECT 434.100 264.600 435.900 272.400 ;
        RECT 449.100 267.000 450.900 272.400 ;
        RECT 452.100 267.900 453.900 273.000 ;
        RECT 455.100 271.500 462.900 272.400 ;
        RECT 455.100 267.000 456.900 271.500 ;
        RECT 449.100 266.100 456.900 267.000 ;
        RECT 458.100 266.400 459.900 270.600 ;
        RECT 461.100 266.400 462.900 271.500 ;
        RECT 476.100 267.300 477.900 272.400 ;
        RECT 479.100 268.200 480.900 273.000 ;
        RECT 482.100 267.300 483.900 272.400 ;
        RECT 458.400 264.900 459.300 266.400 ;
        RECT 476.100 265.950 483.900 267.300 ;
        RECT 485.100 266.400 486.900 272.400 ;
        RECT 500.100 267.300 501.900 272.400 ;
        RECT 503.100 268.200 504.900 273.000 ;
        RECT 506.100 267.300 507.900 272.400 ;
        RECT 427.500 263.700 435.900 264.600 ;
        RECT 454.950 263.700 459.300 264.900 ;
        RECT 485.100 264.300 486.300 266.400 ;
        RECT 500.100 265.950 507.900 267.300 ;
        RECT 509.100 266.400 510.900 272.400 ;
        RECT 524.100 266.400 525.900 272.400 ;
        RECT 527.100 266.400 528.900 273.000 ;
        RECT 509.100 264.300 510.300 266.400 ;
        RECT 355.950 256.950 358.050 259.050 ;
        RECT 358.950 256.950 361.050 259.050 ;
        RECT 361.950 256.950 364.050 259.050 ;
        RECT 364.950 256.950 367.050 259.050 ;
        RECT 367.950 256.950 370.050 259.050 ;
        RECT 382.950 256.950 385.050 259.050 ;
        RECT 385.950 256.950 388.050 259.050 ;
        RECT 388.950 256.950 391.050 259.050 ;
        RECT 391.950 256.950 394.050 259.050 ;
        RECT 406.950 256.950 409.050 259.050 ;
        RECT 409.950 256.950 412.050 259.050 ;
        RECT 425.100 256.950 427.200 259.050 ;
        RECT 428.400 256.950 430.500 259.050 ;
        RECT 343.950 254.550 348.450 256.050 ;
        RECT 359.250 255.150 361.050 256.950 ;
        RECT 343.950 253.950 348.000 254.550 ;
        RECT 362.100 251.400 363.000 256.950 ;
        RECT 365.100 255.150 366.900 256.950 ;
        RECT 386.100 255.150 387.900 256.950 ;
        RECT 362.100 250.500 366.900 251.400 ;
        RECT 272.100 239.400 273.900 247.200 ;
        RECT 275.100 247.200 282.900 248.100 ;
        RECT 275.100 238.500 276.900 247.200 ;
        RECT 269.100 237.600 276.900 238.500 ;
        RECT 278.100 238.500 279.900 246.300 ;
        RECT 281.100 239.400 282.900 247.200 ;
        RECT 284.100 247.500 291.900 248.400 ;
        RECT 284.100 238.500 285.900 247.500 ;
        RECT 278.100 237.600 285.900 238.500 ;
        RECT 287.100 237.000 288.900 246.600 ;
        RECT 290.100 237.600 291.900 247.500 ;
        RECT 308.400 237.000 310.200 249.600 ;
        RECT 313.500 248.100 315.900 249.600 ;
        RECT 313.500 237.600 315.300 248.100 ;
        RECT 316.200 245.100 318.000 246.900 ;
        RECT 316.500 237.000 318.300 243.600 ;
        RECT 332.400 237.000 334.200 249.600 ;
        RECT 337.500 248.100 339.900 249.600 ;
        RECT 356.100 248.400 363.900 249.300 ;
        RECT 337.500 237.600 339.300 248.100 ;
        RECT 340.200 245.100 342.000 246.900 ;
        RECT 340.500 237.000 342.300 243.600 ;
        RECT 356.100 237.600 357.900 248.400 ;
        RECT 359.100 237.000 360.900 247.500 ;
        RECT 362.100 238.500 363.900 248.400 ;
        RECT 365.100 239.400 366.900 250.500 ;
        RECT 368.100 238.500 369.900 249.600 ;
        RECT 392.100 244.800 393.000 256.950 ;
        RECT 407.100 255.150 408.900 256.950 ;
        RECT 386.400 243.900 393.000 244.800 ;
        RECT 386.400 243.600 387.900 243.900 ;
        RECT 362.100 237.600 369.900 238.500 ;
        RECT 383.100 237.000 384.900 243.600 ;
        RECT 386.100 237.600 387.900 243.600 ;
        RECT 392.100 243.600 393.000 243.900 ;
        RECT 410.100 243.600 411.300 256.950 ;
        RECT 425.700 249.600 426.600 256.950 ;
        RECT 429.000 255.150 430.800 256.950 ;
        RECT 389.100 237.000 390.900 243.000 ;
        RECT 392.100 237.600 393.900 243.600 ;
        RECT 407.100 237.000 408.900 243.600 ;
        RECT 410.100 237.600 411.900 243.600 ;
        RECT 425.100 237.600 426.900 249.600 ;
        RECT 428.100 237.000 429.900 249.000 ;
        RECT 432.000 243.600 432.900 263.700 ;
        RECT 433.950 259.050 435.750 260.850 ;
        RECT 452.250 259.050 454.050 260.850 ;
        RECT 433.800 256.950 435.900 259.050 ;
        RECT 448.950 256.950 451.050 259.050 ;
        RECT 451.950 256.950 454.050 259.050 ;
        RECT 454.950 259.050 456.000 263.700 ;
        RECT 482.700 263.400 486.300 264.300 ;
        RECT 506.700 263.400 510.300 264.300 ;
        RECT 472.950 261.450 475.050 262.050 ;
        RECT 457.950 259.050 459.750 260.850 ;
        RECT 467.550 260.550 475.050 261.450 ;
        RECT 454.950 256.950 457.050 259.050 ;
        RECT 457.950 256.950 460.050 259.050 ;
        RECT 460.950 256.950 463.050 259.050 ;
        RECT 449.100 255.150 450.900 256.950 ;
        RECT 454.950 249.600 456.000 256.950 ;
        RECT 460.950 255.150 462.750 256.950 ;
        RECT 467.550 255.450 468.450 260.550 ;
        RECT 472.950 259.950 475.050 260.550 ;
        RECT 479.100 259.050 480.900 260.850 ;
        RECT 482.700 259.050 483.900 263.400 ;
        RECT 487.950 261.450 492.000 262.050 ;
        RECT 485.100 259.050 486.900 260.850 ;
        RECT 487.950 259.950 492.450 261.450 ;
        RECT 475.950 256.950 478.050 259.050 ;
        RECT 478.950 256.950 481.050 259.050 ;
        RECT 481.950 256.950 484.050 259.050 ;
        RECT 484.950 256.950 487.050 259.050 ;
        RECT 464.550 254.550 468.450 255.450 ;
        RECT 476.100 255.150 477.900 256.950 ;
        RECT 457.950 252.450 460.050 253.050 ;
        RECT 464.550 252.450 465.450 254.550 ;
        RECT 457.950 251.550 465.450 252.450 ;
        RECT 457.950 250.950 460.050 251.550 ;
        RECT 482.700 249.600 483.900 256.950 ;
        RECT 491.550 256.050 492.450 259.950 ;
        RECT 503.100 259.050 504.900 260.850 ;
        RECT 506.700 259.050 507.900 263.400 ;
        RECT 509.100 259.050 510.900 260.850 ;
        RECT 524.700 259.050 525.900 266.400 ;
        RECT 545.700 265.200 547.500 272.400 ;
        RECT 550.800 266.400 552.600 273.000 ;
        RECT 566.100 269.400 567.900 273.000 ;
        RECT 569.100 269.400 570.900 272.400 ;
        RECT 572.100 269.400 573.900 273.000 ;
        RECT 545.700 264.300 549.900 265.200 ;
        RECT 529.950 261.450 532.050 262.050 ;
        RECT 535.950 261.450 538.050 262.050 ;
        RECT 527.100 259.050 528.900 260.850 ;
        RECT 529.950 260.550 538.050 261.450 ;
        RECT 529.950 259.950 532.050 260.550 ;
        RECT 535.950 259.950 538.050 260.550 ;
        RECT 545.100 259.050 546.900 260.850 ;
        RECT 548.700 259.050 549.900 264.300 ;
        RECT 550.950 259.050 552.750 260.850 ;
        RECT 569.700 259.050 570.600 269.400 ;
        RECT 587.400 266.400 589.200 273.000 ;
        RECT 592.500 265.200 594.300 272.400 ;
        RECT 608.100 267.300 609.900 272.400 ;
        RECT 611.100 268.200 612.900 273.000 ;
        RECT 614.100 267.300 615.900 272.400 ;
        RECT 608.100 265.950 615.900 267.300 ;
        RECT 617.100 266.400 618.900 272.400 ;
        RECT 632.400 266.400 634.200 273.000 ;
        RECT 590.100 264.300 594.300 265.200 ;
        RECT 617.100 264.300 618.300 266.400 ;
        RECT 637.500 265.200 639.300 272.400 ;
        RECT 656.100 269.400 657.900 272.400 ;
        RECT 659.100 269.400 660.900 273.000 ;
        RECT 587.250 259.050 589.050 260.850 ;
        RECT 590.100 259.050 591.300 264.300 ;
        RECT 614.700 263.400 618.300 264.300 ;
        RECT 635.100 264.300 639.300 265.200 ;
        RECT 593.100 259.050 594.900 260.850 ;
        RECT 611.100 259.050 612.900 260.850 ;
        RECT 614.700 259.050 615.900 263.400 ;
        RECT 617.100 259.050 618.900 260.850 ;
        RECT 632.250 259.050 634.050 260.850 ;
        RECT 635.100 259.050 636.300 264.300 ;
        RECT 638.100 259.050 639.900 260.850 ;
        RECT 656.700 259.050 657.900 269.400 ;
        RECT 676.500 264.000 678.300 272.400 ;
        RECT 675.000 262.800 678.300 264.000 ;
        RECT 683.100 263.400 684.900 273.000 ;
        RECT 700.500 264.000 702.300 272.400 ;
        RECT 699.000 262.800 702.300 264.000 ;
        RECT 707.100 263.400 708.900 273.000 ;
        RECT 722.100 264.600 723.900 272.400 ;
        RECT 726.600 266.400 728.400 273.000 ;
        RECT 729.600 268.200 731.400 272.400 ;
        RECT 729.600 266.400 732.300 268.200 ;
        RECT 749.700 266.400 751.500 273.000 ;
        RECT 754.200 266.400 756.000 272.400 ;
        RECT 758.700 266.400 760.500 273.000 ;
        RECT 728.700 264.600 730.500 265.500 ;
        RECT 722.100 263.700 730.500 264.600 ;
        RECT 675.000 259.050 675.900 262.800 ;
        RECT 677.100 259.050 678.900 260.850 ;
        RECT 683.100 259.050 684.900 260.850 ;
        RECT 699.000 259.050 699.900 262.800 ;
        RECT 701.100 259.050 702.900 260.850 ;
        RECT 707.100 259.050 708.900 260.850 ;
        RECT 722.250 259.050 724.050 260.850 ;
        RECT 499.950 256.950 502.050 259.050 ;
        RECT 502.950 256.950 505.050 259.050 ;
        RECT 505.950 256.950 508.050 259.050 ;
        RECT 508.950 256.950 511.050 259.050 ;
        RECT 523.950 256.950 526.050 259.050 ;
        RECT 526.950 256.950 529.050 259.050 ;
        RECT 544.950 256.950 547.050 259.050 ;
        RECT 547.950 256.950 550.050 259.050 ;
        RECT 550.950 256.950 553.050 259.050 ;
        RECT 565.950 256.950 568.050 259.050 ;
        RECT 568.950 256.950 571.050 259.050 ;
        RECT 571.950 256.950 574.050 259.050 ;
        RECT 586.950 256.950 589.050 259.050 ;
        RECT 589.950 256.950 592.050 259.050 ;
        RECT 592.950 256.950 595.050 259.050 ;
        RECT 607.950 256.950 610.050 259.050 ;
        RECT 610.950 256.950 613.050 259.050 ;
        RECT 613.950 256.950 616.050 259.050 ;
        RECT 616.950 256.950 619.050 259.050 ;
        RECT 631.950 256.950 634.050 259.050 ;
        RECT 634.950 256.950 637.050 259.050 ;
        RECT 637.950 256.950 640.050 259.050 ;
        RECT 655.950 256.950 658.050 259.050 ;
        RECT 658.950 256.950 661.050 259.050 ;
        RECT 673.950 256.950 676.050 259.050 ;
        RECT 676.950 256.950 679.050 259.050 ;
        RECT 679.950 256.950 682.050 259.050 ;
        RECT 682.950 256.950 685.050 259.050 ;
        RECT 697.950 256.950 700.050 259.050 ;
        RECT 700.950 256.950 703.050 259.050 ;
        RECT 703.950 256.950 706.050 259.050 ;
        RECT 706.950 256.950 709.050 259.050 ;
        RECT 722.100 256.950 724.200 259.050 ;
        RECT 487.950 254.550 492.450 256.050 ;
        RECT 500.100 255.150 501.900 256.950 ;
        RECT 487.950 253.950 492.000 254.550 ;
        RECT 493.950 252.450 496.050 253.050 ;
        RECT 502.950 252.450 505.050 253.050 ;
        RECT 493.950 251.550 505.050 252.450 ;
        RECT 493.950 250.950 496.050 251.550 ;
        RECT 502.950 250.950 505.050 251.550 ;
        RECT 506.700 249.600 507.900 256.950 ;
        RECT 524.700 249.600 525.900 256.950 ;
        RECT 431.100 237.600 432.900 243.600 ;
        RECT 434.100 237.000 435.900 243.600 ;
        RECT 449.100 237.000 450.900 249.600 ;
        RECT 453.600 237.600 456.900 249.600 ;
        RECT 459.600 237.000 461.400 249.600 ;
        RECT 476.400 237.000 478.200 249.600 ;
        RECT 481.500 248.100 483.900 249.600 ;
        RECT 481.500 237.600 483.300 248.100 ;
        RECT 484.200 245.100 486.000 246.900 ;
        RECT 484.500 237.000 486.300 243.600 ;
        RECT 500.400 237.000 502.200 249.600 ;
        RECT 505.500 248.100 507.900 249.600 ;
        RECT 505.500 237.600 507.300 248.100 ;
        RECT 508.200 245.100 510.000 246.900 ;
        RECT 508.500 237.000 510.300 243.600 ;
        RECT 524.100 237.600 525.900 249.600 ;
        RECT 527.100 237.000 528.900 249.600 ;
        RECT 548.700 243.600 549.900 256.950 ;
        RECT 566.100 255.150 567.900 256.950 ;
        RECT 569.700 249.600 570.600 256.950 ;
        RECT 571.950 255.150 573.750 256.950 ;
        RECT 567.000 248.400 570.600 249.600 ;
        RECT 545.100 237.000 546.900 243.600 ;
        RECT 548.100 237.600 549.900 243.600 ;
        RECT 551.100 237.000 552.900 243.600 ;
        RECT 567.000 237.600 568.800 248.400 ;
        RECT 572.100 237.000 573.900 249.600 ;
        RECT 590.100 243.600 591.300 256.950 ;
        RECT 608.100 255.150 609.900 256.950 ;
        RECT 614.700 249.600 615.900 256.950 ;
        RECT 616.950 252.450 619.050 253.050 ;
        RECT 631.950 252.450 634.050 253.050 ;
        RECT 616.950 251.550 634.050 252.450 ;
        RECT 616.950 250.950 619.050 251.550 ;
        RECT 631.950 250.950 634.050 251.550 ;
        RECT 587.100 237.000 588.900 243.600 ;
        RECT 590.100 237.600 591.900 243.600 ;
        RECT 593.100 237.000 594.900 243.600 ;
        RECT 608.400 237.000 610.200 249.600 ;
        RECT 613.500 248.100 615.900 249.600 ;
        RECT 613.500 237.600 615.300 248.100 ;
        RECT 616.200 245.100 618.000 246.900 ;
        RECT 635.100 243.600 636.300 256.950 ;
        RECT 640.950 249.450 643.050 250.050 ;
        RECT 652.950 249.450 655.050 250.050 ;
        RECT 640.950 248.550 655.050 249.450 ;
        RECT 640.950 247.950 643.050 248.550 ;
        RECT 652.950 247.950 655.050 248.550 ;
        RECT 656.700 243.600 657.900 256.950 ;
        RECT 659.100 255.150 660.900 256.950 ;
        RECT 675.000 244.800 675.900 256.950 ;
        RECT 680.100 255.150 681.900 256.950 ;
        RECT 699.000 244.800 699.900 256.950 ;
        RECT 704.100 255.150 705.900 256.950 ;
        RECT 675.000 243.900 681.600 244.800 ;
        RECT 675.000 243.600 675.900 243.900 ;
        RECT 616.500 237.000 618.300 243.600 ;
        RECT 632.100 237.000 633.900 243.600 ;
        RECT 635.100 237.600 636.900 243.600 ;
        RECT 638.100 237.000 639.900 243.600 ;
        RECT 656.100 237.600 657.900 243.600 ;
        RECT 659.100 237.000 660.900 243.600 ;
        RECT 674.100 237.600 675.900 243.600 ;
        RECT 680.100 243.600 681.600 243.900 ;
        RECT 699.000 243.900 705.600 244.800 ;
        RECT 699.000 243.600 699.900 243.900 ;
        RECT 677.100 237.000 678.900 243.000 ;
        RECT 680.100 237.600 681.900 243.600 ;
        RECT 683.100 237.000 684.900 243.600 ;
        RECT 698.100 237.600 699.900 243.600 ;
        RECT 704.100 243.600 705.600 243.900 ;
        RECT 725.100 243.600 726.000 263.700 ;
        RECT 731.400 259.050 732.300 266.400 ;
        RECT 749.250 259.050 751.050 260.850 ;
        RECT 755.100 259.050 756.300 266.400 ;
        RECT 779.100 263.400 780.900 273.000 ;
        RECT 785.700 264.000 787.500 272.400 ;
        RECT 804.000 266.400 805.800 273.000 ;
        RECT 808.500 267.600 810.300 272.400 ;
        RECT 811.500 269.400 813.300 273.000 ;
        RECT 808.500 266.400 813.600 267.600 ;
        RECT 785.700 262.800 789.000 264.000 ;
        RECT 761.100 259.050 762.900 260.850 ;
        RECT 779.100 259.050 780.900 260.850 ;
        RECT 785.100 259.050 786.900 260.850 ;
        RECT 788.100 259.050 789.000 262.800 ;
        RECT 803.100 259.050 804.900 260.850 ;
        RECT 809.250 259.050 811.050 260.850 ;
        RECT 812.700 259.050 813.600 266.400 ;
        RECT 829.500 264.000 831.300 272.400 ;
        RECT 828.000 262.800 831.300 264.000 ;
        RECT 836.100 263.400 837.900 273.000 ;
        RECT 851.700 269.400 853.500 273.000 ;
        RECT 854.700 267.600 856.500 272.400 ;
        RECT 851.400 266.400 856.500 267.600 ;
        RECT 859.200 266.400 861.000 273.000 ;
        RECT 828.000 259.050 828.900 262.800 ;
        RECT 830.100 259.050 831.900 260.850 ;
        RECT 836.100 259.050 837.900 260.850 ;
        RECT 851.400 259.050 852.300 266.400 ;
        RECT 875.700 265.200 877.500 272.400 ;
        RECT 880.800 266.400 882.600 273.000 ;
        RECT 875.700 264.300 879.900 265.200 ;
        RECT 865.950 261.450 868.050 262.050 ;
        RECT 871.950 261.450 874.050 262.050 ;
        RECT 853.950 259.050 855.750 260.850 ;
        RECT 860.100 259.050 861.900 260.850 ;
        RECT 865.950 260.550 874.050 261.450 ;
        RECT 865.950 259.950 868.050 260.550 ;
        RECT 871.950 259.950 874.050 260.550 ;
        RECT 875.100 259.050 876.900 260.850 ;
        RECT 878.700 259.050 879.900 264.300 ;
        RECT 880.950 259.050 882.750 260.850 ;
        RECT 727.500 256.950 729.600 259.050 ;
        RECT 730.800 256.950 732.900 259.050 ;
        RECT 748.950 256.950 751.050 259.050 ;
        RECT 751.950 256.950 754.050 259.050 ;
        RECT 754.950 256.950 757.050 259.050 ;
        RECT 757.950 256.950 760.050 259.050 ;
        RECT 760.950 256.950 763.050 259.050 ;
        RECT 778.950 256.950 781.050 259.050 ;
        RECT 781.950 256.950 784.050 259.050 ;
        RECT 784.950 256.950 787.050 259.050 ;
        RECT 787.950 256.950 790.050 259.050 ;
        RECT 802.950 256.950 805.050 259.050 ;
        RECT 805.950 256.950 808.050 259.050 ;
        RECT 808.950 256.950 811.050 259.050 ;
        RECT 811.950 256.950 814.050 259.050 ;
        RECT 826.950 256.950 829.050 259.050 ;
        RECT 829.950 256.950 832.050 259.050 ;
        RECT 832.950 256.950 835.050 259.050 ;
        RECT 835.950 256.950 838.050 259.050 ;
        RECT 850.950 256.950 853.050 259.050 ;
        RECT 853.950 256.950 856.050 259.050 ;
        RECT 856.950 256.950 859.050 259.050 ;
        RECT 859.950 256.950 862.050 259.050 ;
        RECT 874.950 256.950 877.050 259.050 ;
        RECT 877.950 256.950 880.050 259.050 ;
        RECT 880.950 256.950 883.050 259.050 ;
        RECT 727.200 255.150 729.000 256.950 ;
        RECT 731.400 249.600 732.300 256.950 ;
        RECT 752.250 255.150 754.050 256.950 ;
        RECT 733.950 252.450 736.050 253.050 ;
        RECT 751.950 252.450 754.050 253.050 ;
        RECT 733.950 251.550 754.050 252.450 ;
        RECT 733.950 250.950 736.050 251.550 ;
        RECT 751.950 250.950 754.050 251.550 ;
        RECT 755.100 251.400 756.000 256.950 ;
        RECT 758.100 255.150 759.900 256.950 ;
        RECT 782.100 255.150 783.900 256.950 ;
        RECT 755.100 250.500 759.900 251.400 ;
        RECT 701.100 237.000 702.900 243.000 ;
        RECT 704.100 237.600 705.900 243.600 ;
        RECT 707.100 237.000 708.900 243.600 ;
        RECT 722.100 237.000 723.900 243.600 ;
        RECT 725.100 237.600 726.900 243.600 ;
        RECT 728.100 237.000 729.900 249.000 ;
        RECT 731.100 237.600 732.900 249.600 ;
        RECT 749.100 248.400 756.900 249.300 ;
        RECT 749.100 237.600 750.900 248.400 ;
        RECT 752.100 237.000 753.900 247.500 ;
        RECT 755.100 238.500 756.900 248.400 ;
        RECT 758.100 239.400 759.900 250.500 ;
        RECT 761.100 238.500 762.900 249.600 ;
        RECT 788.100 244.800 789.000 256.950 ;
        RECT 806.250 255.150 808.050 256.950 ;
        RECT 812.700 249.600 813.600 256.950 ;
        RECT 782.400 243.900 789.000 244.800 ;
        RECT 782.400 243.600 783.900 243.900 ;
        RECT 755.100 237.600 762.900 238.500 ;
        RECT 779.100 237.000 780.900 243.600 ;
        RECT 782.100 237.600 783.900 243.600 ;
        RECT 788.100 243.600 789.000 243.900 ;
        RECT 803.100 248.700 810.900 249.600 ;
        RECT 785.100 237.000 786.900 243.000 ;
        RECT 788.100 237.600 789.900 243.600 ;
        RECT 803.100 237.600 804.900 248.700 ;
        RECT 806.100 237.000 807.900 247.800 ;
        RECT 809.100 237.600 810.900 248.700 ;
        RECT 812.100 237.600 813.900 249.600 ;
        RECT 828.000 244.800 828.900 256.950 ;
        RECT 833.100 255.150 834.900 256.950 ;
        RECT 838.950 255.450 841.050 256.050 ;
        RECT 844.950 255.450 847.050 256.050 ;
        RECT 838.950 254.550 847.050 255.450 ;
        RECT 838.950 253.950 841.050 254.550 ;
        RECT 844.950 253.950 847.050 254.550 ;
        RECT 851.400 249.600 852.300 256.950 ;
        RECT 856.950 255.150 858.750 256.950 ;
        RECT 828.000 243.900 834.600 244.800 ;
        RECT 828.000 243.600 828.900 243.900 ;
        RECT 827.100 237.600 828.900 243.600 ;
        RECT 833.100 243.600 834.600 243.900 ;
        RECT 830.100 237.000 831.900 243.000 ;
        RECT 833.100 237.600 834.900 243.600 ;
        RECT 836.100 237.000 837.900 243.600 ;
        RECT 851.100 237.600 852.900 249.600 ;
        RECT 854.100 248.700 861.900 249.600 ;
        RECT 854.100 237.600 855.900 248.700 ;
        RECT 857.100 237.000 858.900 247.800 ;
        RECT 860.100 237.600 861.900 248.700 ;
        RECT 878.700 243.600 879.900 256.950 ;
        RECT 880.950 252.450 883.050 253.050 ;
        RECT 889.950 252.450 892.050 253.050 ;
        RECT 880.950 251.550 892.050 252.450 ;
        RECT 880.950 250.950 883.050 251.550 ;
        RECT 889.950 250.950 892.050 251.550 ;
        RECT 875.100 237.000 876.900 243.600 ;
        RECT 878.100 237.600 879.900 243.600 ;
        RECT 881.100 237.000 882.900 243.600 ;
        RECT 14.100 222.600 15.900 233.400 ;
        RECT 17.100 223.500 19.200 234.000 ;
        RECT 14.100 221.400 19.200 222.600 ;
        RECT 21.600 222.300 23.400 233.400 ;
        RECT 26.100 223.500 27.900 234.000 ;
        RECT 29.100 222.300 30.900 233.400 ;
        RECT 44.100 227.400 45.900 234.000 ;
        RECT 47.100 227.400 48.900 233.400 ;
        RECT 50.100 227.400 51.900 234.000 ;
        RECT 17.100 220.500 19.200 221.400 ;
        RECT 20.100 221.400 23.400 222.300 ;
        RECT 20.100 217.050 21.300 221.400 ;
        RECT 26.100 221.100 30.900 222.300 ;
        RECT 26.100 220.200 28.200 221.100 ;
        RECT 22.800 219.300 28.200 220.200 ;
        RECT 22.800 217.500 24.600 219.300 ;
        RECT 19.800 216.300 21.900 217.050 ;
        RECT 14.400 214.050 16.200 215.850 ;
        RECT 19.800 214.950 22.800 216.300 ;
        RECT 14.100 211.950 16.200 214.050 ;
        RECT 19.200 212.100 21.000 213.900 ;
        RECT 18.900 210.000 21.000 212.100 ;
        RECT 21.900 208.200 22.800 214.950 ;
        RECT 24.300 214.200 26.100 216.000 ;
        RECT 24.000 212.100 26.100 214.200 ;
        RECT 47.700 214.050 48.900 227.400 ;
        RECT 65.100 222.600 66.900 233.400 ;
        RECT 68.100 223.500 69.900 234.000 ;
        RECT 65.100 221.400 69.900 222.600 ;
        RECT 67.800 220.500 69.900 221.400 ;
        RECT 72.600 221.400 74.400 233.400 ;
        RECT 77.100 223.500 78.900 234.000 ;
        RECT 80.100 222.300 81.900 233.400 ;
        RECT 95.100 227.400 96.900 233.400 ;
        RECT 98.100 228.000 99.900 234.000 ;
        RECT 77.400 221.400 81.900 222.300 ;
        RECT 96.000 227.100 96.900 227.400 ;
        RECT 101.100 227.400 102.900 233.400 ;
        RECT 104.100 227.400 105.900 234.000 ;
        RECT 119.100 227.400 120.900 234.000 ;
        RECT 122.100 227.400 123.900 233.400 ;
        RECT 125.100 227.400 126.900 234.000 ;
        RECT 101.100 227.100 102.600 227.400 ;
        RECT 96.000 226.200 102.600 227.100 ;
        RECT 72.600 220.050 73.800 221.400 ;
        RECT 72.300 219.000 73.800 220.050 ;
        RECT 77.400 219.300 79.500 221.400 ;
        RECT 72.300 217.050 73.200 219.000 ;
        RECT 82.950 217.950 85.050 220.050 ;
        RECT 65.400 214.050 67.200 215.850 ;
        RECT 71.100 214.950 73.200 217.050 ;
        RECT 74.100 217.500 76.200 217.800 ;
        RECT 74.100 215.700 78.000 217.500 ;
        RECT 28.800 211.800 30.900 214.050 ;
        RECT 43.950 211.950 46.050 214.050 ;
        RECT 46.950 211.950 49.050 214.050 ;
        RECT 49.950 211.950 52.050 214.050 ;
        RECT 65.100 211.950 67.200 214.050 ;
        RECT 71.700 214.800 73.200 214.950 ;
        RECT 71.700 213.900 74.100 214.800 ;
        RECT 28.800 211.200 30.600 211.800 ;
        RECT 24.000 210.000 30.600 211.200 ;
        RECT 44.100 210.150 45.900 211.950 ;
        RECT 24.000 209.100 26.100 210.000 ;
        RECT 16.500 205.500 18.600 207.900 ;
        RECT 19.800 206.100 22.800 208.200 ;
        RECT 23.700 207.300 25.500 209.100 ;
        RECT 14.100 204.600 18.600 205.500 ;
        RECT 14.100 198.600 15.900 204.600 ;
        RECT 21.900 204.000 22.800 206.100 ;
        RECT 26.400 207.000 28.500 207.600 ;
        RECT 26.400 205.500 30.900 207.000 ;
        RECT 47.700 206.700 48.900 211.950 ;
        RECT 49.950 210.150 51.750 211.950 ;
        RECT 69.900 211.200 71.700 213.000 ;
        RECT 69.900 209.100 72.000 211.200 ;
        RECT 72.900 208.200 74.100 213.900 ;
        RECT 75.000 214.050 76.800 214.500 ;
        RECT 75.000 212.700 81.900 214.050 ;
        RECT 79.800 211.950 81.900 212.700 ;
        RECT 29.400 204.600 30.900 205.500 ;
        RECT 17.400 198.000 19.200 203.700 ;
        RECT 21.900 198.600 23.700 204.000 ;
        RECT 26.100 198.000 27.900 203.700 ;
        RECT 29.100 198.600 30.900 204.600 ;
        RECT 44.700 205.800 48.900 206.700 ;
        RECT 44.700 198.600 46.500 205.800 ;
        RECT 67.800 205.500 69.900 206.700 ;
        RECT 71.100 206.100 74.100 208.200 ;
        RECT 75.000 209.400 76.800 211.200 ;
        RECT 79.800 210.150 81.600 211.950 ;
        RECT 75.000 207.300 77.100 209.400 ;
        RECT 83.550 207.900 84.450 217.950 ;
        RECT 96.000 214.050 96.900 226.200 ;
        RECT 101.100 214.050 102.900 215.850 ;
        RECT 122.100 214.050 123.300 227.400 ;
        RECT 140.100 222.300 141.900 233.400 ;
        RECT 143.100 223.500 144.900 234.000 ;
        RECT 147.600 222.300 149.400 233.400 ;
        RECT 151.800 223.500 153.900 234.000 ;
        RECT 155.100 222.600 156.900 233.400 ;
        RECT 170.100 227.400 171.900 233.400 ;
        RECT 173.100 228.000 174.900 234.000 ;
        RECT 140.100 221.100 144.900 222.300 ;
        RECT 147.600 221.400 150.900 222.300 ;
        RECT 142.800 220.200 144.900 221.100 ;
        RECT 142.800 219.300 148.200 220.200 ;
        RECT 146.400 217.500 148.200 219.300 ;
        RECT 149.700 217.050 150.900 221.400 ;
        RECT 151.800 221.400 156.900 222.600 ;
        RECT 171.000 227.100 171.900 227.400 ;
        RECT 176.100 227.400 177.900 233.400 ;
        RECT 179.100 227.400 180.900 234.000 ;
        RECT 176.100 227.100 177.600 227.400 ;
        RECT 171.000 226.200 177.600 227.100 ;
        RECT 151.800 220.500 153.900 221.400 ;
        RECT 149.100 216.300 151.200 217.050 ;
        RECT 144.900 214.200 146.700 216.000 ;
        RECT 148.200 214.950 151.200 216.300 ;
        RECT 94.950 211.950 97.050 214.050 ;
        RECT 97.950 211.950 100.050 214.050 ;
        RECT 100.950 211.950 103.050 214.050 ;
        RECT 103.950 211.950 106.050 214.050 ;
        RECT 118.950 211.950 121.050 214.050 ;
        RECT 121.950 211.950 124.050 214.050 ;
        RECT 124.950 211.950 127.050 214.050 ;
        RECT 96.000 208.200 96.900 211.950 ;
        RECT 98.100 210.150 99.900 211.950 ;
        RECT 104.100 210.150 105.900 211.950 ;
        RECT 119.250 210.150 121.050 211.950 ;
        RECT 75.000 206.400 81.300 207.300 ;
        RECT 65.100 204.600 69.900 205.500 ;
        RECT 72.900 204.600 74.100 206.100 ;
        RECT 80.100 204.600 81.300 206.400 ;
        RECT 82.950 205.800 85.050 207.900 ;
        RECT 96.000 207.000 99.300 208.200 ;
        RECT 49.800 198.000 51.600 204.600 ;
        RECT 65.100 198.600 66.900 204.600 ;
        RECT 68.100 198.000 69.900 203.700 ;
        RECT 72.600 198.600 74.400 204.600 ;
        RECT 77.100 198.000 78.900 203.700 ;
        RECT 80.100 198.600 81.900 204.600 ;
        RECT 97.500 198.600 99.300 207.000 ;
        RECT 104.100 198.000 105.900 207.600 ;
        RECT 122.100 206.700 123.300 211.950 ;
        RECT 125.100 210.150 126.900 211.950 ;
        RECT 140.100 211.800 142.200 214.050 ;
        RECT 144.900 212.100 147.000 214.200 ;
        RECT 140.400 211.200 142.200 211.800 ;
        RECT 140.400 210.000 147.000 211.200 ;
        RECT 144.900 209.100 147.000 210.000 ;
        RECT 142.500 207.000 144.600 207.600 ;
        RECT 145.500 207.300 147.300 209.100 ;
        RECT 148.200 208.200 149.100 214.950 ;
        RECT 154.800 214.050 156.600 215.850 ;
        RECT 171.000 214.050 171.900 226.200 ;
        RECT 194.100 222.300 195.900 233.400 ;
        RECT 197.100 223.200 198.900 234.000 ;
        RECT 200.100 222.300 201.900 233.400 ;
        RECT 194.100 221.400 201.900 222.300 ;
        RECT 203.100 221.400 204.900 233.400 ;
        RECT 218.400 221.400 220.200 234.000 ;
        RECT 223.500 222.900 225.300 233.400 ;
        RECT 226.500 227.400 228.300 234.000 ;
        RECT 226.200 224.100 228.000 225.900 ;
        RECT 223.500 221.400 225.900 222.900 ;
        RECT 242.100 221.400 243.900 233.400 ;
        RECT 245.100 222.300 246.900 233.400 ;
        RECT 248.100 223.200 249.900 234.000 ;
        RECT 251.100 222.300 252.900 233.400 ;
        RECT 266.100 227.400 267.900 234.000 ;
        RECT 269.100 227.400 270.900 233.400 ;
        RECT 272.100 228.000 273.900 234.000 ;
        RECT 269.400 227.100 270.900 227.400 ;
        RECT 275.100 227.400 276.900 233.400 ;
        RECT 293.100 227.400 294.900 234.000 ;
        RECT 296.100 227.400 297.900 233.400 ;
        RECT 299.100 228.000 300.900 234.000 ;
        RECT 275.100 227.100 276.000 227.400 ;
        RECT 269.400 226.200 276.000 227.100 ;
        RECT 296.400 227.100 297.900 227.400 ;
        RECT 302.100 227.400 303.900 233.400 ;
        RECT 317.100 227.400 318.900 233.400 ;
        RECT 320.100 228.000 321.900 234.000 ;
        RECT 302.100 227.100 303.000 227.400 ;
        RECT 296.400 226.200 303.000 227.100 ;
        RECT 245.100 221.400 252.900 222.300 ;
        RECT 178.950 219.450 181.050 219.900 ;
        RECT 199.950 219.450 202.050 220.050 ;
        RECT 178.950 218.550 202.050 219.450 ;
        RECT 178.950 217.800 181.050 218.550 ;
        RECT 199.950 217.950 202.050 218.550 ;
        RECT 176.100 214.050 177.900 215.850 ;
        RECT 197.250 214.050 199.050 215.850 ;
        RECT 203.700 214.050 204.600 221.400 ;
        RECT 218.100 214.050 219.900 215.850 ;
        RECT 224.700 214.050 225.900 221.400 ;
        RECT 226.950 219.450 229.050 220.050 ;
        RECT 235.950 219.450 238.050 220.050 ;
        RECT 226.950 218.550 238.050 219.450 ;
        RECT 226.950 217.950 229.050 218.550 ;
        RECT 235.950 217.950 238.050 218.550 ;
        RECT 242.400 214.050 243.300 221.400 ;
        RECT 244.950 219.450 247.050 220.050 ;
        RECT 259.950 219.450 262.050 220.050 ;
        RECT 244.950 218.550 262.050 219.450 ;
        RECT 244.950 217.950 247.050 218.550 ;
        RECT 259.950 217.950 262.050 218.550 ;
        RECT 247.950 214.050 249.750 215.850 ;
        RECT 269.100 214.050 270.900 215.850 ;
        RECT 275.100 214.050 276.000 226.200 ;
        RECT 296.100 214.050 297.900 215.850 ;
        RECT 302.100 214.050 303.000 226.200 ;
        RECT 318.000 227.100 318.900 227.400 ;
        RECT 323.100 227.400 324.900 233.400 ;
        RECT 326.100 227.400 327.900 234.000 ;
        RECT 341.100 227.400 342.900 233.400 ;
        RECT 344.100 227.400 345.900 234.000 ;
        RECT 323.100 227.100 324.600 227.400 ;
        RECT 318.000 226.200 324.600 227.100 ;
        RECT 318.000 214.050 318.900 226.200 ;
        RECT 323.100 214.050 324.900 215.850 ;
        RECT 341.700 214.050 342.900 227.400 ;
        RECT 346.950 225.450 349.050 226.050 ;
        RECT 352.950 225.450 355.050 226.050 ;
        RECT 346.950 224.550 355.050 225.450 ;
        RECT 346.950 223.950 349.050 224.550 ;
        RECT 352.950 223.950 355.050 224.550 ;
        RECT 362.400 221.400 364.200 234.000 ;
        RECT 367.500 222.900 369.300 233.400 ;
        RECT 370.500 227.400 372.300 234.000 ;
        RECT 370.200 224.100 372.000 225.900 ;
        RECT 367.500 221.400 369.900 222.900 ;
        RECT 386.400 221.400 388.200 234.000 ;
        RECT 391.500 222.900 393.300 233.400 ;
        RECT 394.500 227.400 396.300 234.000 ;
        RECT 410.100 227.400 411.900 234.000 ;
        RECT 413.100 227.400 414.900 233.400 ;
        RECT 416.100 228.000 417.900 234.000 ;
        RECT 413.400 227.100 414.900 227.400 ;
        RECT 419.100 227.400 420.900 233.400 ;
        RECT 434.100 227.400 435.900 234.000 ;
        RECT 437.100 227.400 438.900 233.400 ;
        RECT 440.100 228.000 441.900 234.000 ;
        RECT 419.100 227.100 420.000 227.400 ;
        RECT 413.400 226.200 420.000 227.100 ;
        RECT 437.400 227.100 438.900 227.400 ;
        RECT 443.100 227.400 444.900 233.400 ;
        RECT 461.100 227.400 462.900 234.000 ;
        RECT 464.100 227.400 465.900 233.400 ;
        RECT 467.100 228.000 468.900 234.000 ;
        RECT 443.100 227.100 444.000 227.400 ;
        RECT 437.400 226.200 444.000 227.100 ;
        RECT 464.400 227.100 465.900 227.400 ;
        RECT 470.100 227.400 471.900 233.400 ;
        RECT 470.100 227.100 471.000 227.400 ;
        RECT 464.400 226.200 471.000 227.100 ;
        RECT 394.200 224.100 396.000 225.900 ;
        RECT 391.500 221.400 393.900 222.900 ;
        RECT 344.100 214.050 345.900 215.850 ;
        RECT 362.100 214.050 363.900 215.850 ;
        RECT 368.700 214.050 369.900 221.400 ;
        RECT 370.950 219.450 373.050 220.200 ;
        RECT 370.950 218.550 378.450 219.450 ;
        RECT 370.950 218.100 373.050 218.550 ;
        RECT 150.000 212.100 151.800 213.900 ;
        RECT 150.000 210.000 152.100 212.100 ;
        RECT 154.800 211.950 156.900 214.050 ;
        RECT 169.950 211.950 172.050 214.050 ;
        RECT 172.950 211.950 175.050 214.050 ;
        RECT 175.950 211.950 178.050 214.050 ;
        RECT 178.950 211.950 181.050 214.050 ;
        RECT 193.950 211.950 196.050 214.050 ;
        RECT 196.950 211.950 199.050 214.050 ;
        RECT 199.950 211.950 202.050 214.050 ;
        RECT 202.950 211.950 205.050 214.050 ;
        RECT 217.950 211.950 220.050 214.050 ;
        RECT 220.950 211.950 223.050 214.050 ;
        RECT 223.950 211.950 226.050 214.050 ;
        RECT 226.950 211.950 229.050 214.050 ;
        RECT 241.950 211.950 244.050 214.050 ;
        RECT 244.950 211.950 247.050 214.050 ;
        RECT 247.950 211.950 250.050 214.050 ;
        RECT 250.950 211.950 253.050 214.050 ;
        RECT 265.950 211.950 268.050 214.050 ;
        RECT 268.950 211.950 271.050 214.050 ;
        RECT 271.950 211.950 274.050 214.050 ;
        RECT 274.950 211.950 277.050 214.050 ;
        RECT 292.950 211.950 295.050 214.050 ;
        RECT 295.950 211.950 298.050 214.050 ;
        RECT 298.950 211.950 301.050 214.050 ;
        RECT 301.950 211.950 304.050 214.050 ;
        RECT 316.950 211.950 319.050 214.050 ;
        RECT 319.950 211.950 322.050 214.050 ;
        RECT 322.950 211.950 325.050 214.050 ;
        RECT 325.950 211.950 328.050 214.050 ;
        RECT 340.950 211.950 343.050 214.050 ;
        RECT 343.950 211.950 346.050 214.050 ;
        RECT 361.950 211.950 364.050 214.050 ;
        RECT 364.950 211.950 367.050 214.050 ;
        RECT 367.950 211.950 370.050 214.050 ;
        RECT 370.950 211.950 373.050 214.050 ;
        RECT 171.000 208.200 171.900 211.950 ;
        RECT 173.100 210.150 174.900 211.950 ;
        RECT 179.100 210.150 180.900 211.950 ;
        RECT 194.100 210.150 195.900 211.950 ;
        RECT 200.250 210.150 202.050 211.950 ;
        RECT 122.100 205.800 126.300 206.700 ;
        RECT 119.400 198.000 121.200 204.600 ;
        RECT 124.500 198.600 126.300 205.800 ;
        RECT 140.100 205.500 144.600 207.000 ;
        RECT 148.200 206.100 151.200 208.200 ;
        RECT 140.100 204.600 141.600 205.500 ;
        RECT 140.100 198.600 141.900 204.600 ;
        RECT 148.200 204.000 149.100 206.100 ;
        RECT 152.400 205.500 154.500 207.900 ;
        RECT 171.000 207.000 174.300 208.200 ;
        RECT 152.400 204.600 156.900 205.500 ;
        RECT 143.100 198.000 144.900 203.700 ;
        RECT 147.300 198.600 149.100 204.000 ;
        RECT 151.800 198.000 153.600 203.700 ;
        RECT 155.100 198.600 156.900 204.600 ;
        RECT 172.500 198.600 174.300 207.000 ;
        RECT 179.100 198.000 180.900 207.600 ;
        RECT 203.700 204.600 204.600 211.950 ;
        RECT 221.100 210.150 222.900 211.950 ;
        RECT 224.700 207.600 225.900 211.950 ;
        RECT 227.100 210.150 228.900 211.950 ;
        RECT 224.700 206.700 228.300 207.600 ;
        RECT 195.000 198.000 196.800 204.600 ;
        RECT 199.500 203.400 204.600 204.600 ;
        RECT 218.100 203.700 225.900 205.050 ;
        RECT 199.500 198.600 201.300 203.400 ;
        RECT 202.500 198.000 204.300 201.600 ;
        RECT 218.100 198.600 219.900 203.700 ;
        RECT 221.100 198.000 222.900 202.800 ;
        RECT 224.100 198.600 225.900 203.700 ;
        RECT 227.100 204.600 228.300 206.700 ;
        RECT 242.400 204.600 243.300 211.950 ;
        RECT 244.950 210.150 246.750 211.950 ;
        RECT 251.100 210.150 252.900 211.950 ;
        RECT 266.100 210.150 267.900 211.950 ;
        RECT 272.100 210.150 273.900 211.950 ;
        RECT 275.100 208.200 276.000 211.950 ;
        RECT 277.950 210.450 280.050 211.050 ;
        RECT 286.950 210.450 289.050 211.050 ;
        RECT 277.950 209.550 289.050 210.450 ;
        RECT 293.100 210.150 294.900 211.950 ;
        RECT 299.100 210.150 300.900 211.950 ;
        RECT 277.950 208.950 280.050 209.550 ;
        RECT 286.950 208.950 289.050 209.550 ;
        RECT 302.100 208.200 303.000 211.950 ;
        RECT 227.100 198.600 228.900 204.600 ;
        RECT 242.400 203.400 247.500 204.600 ;
        RECT 242.700 198.000 244.500 201.600 ;
        RECT 245.700 198.600 247.500 203.400 ;
        RECT 250.200 198.000 252.000 204.600 ;
        RECT 266.100 198.000 267.900 207.600 ;
        RECT 272.700 207.000 276.000 208.200 ;
        RECT 272.700 198.600 274.500 207.000 ;
        RECT 293.100 198.000 294.900 207.600 ;
        RECT 299.700 207.000 303.000 208.200 ;
        RECT 318.000 208.200 318.900 211.950 ;
        RECT 320.100 210.150 321.900 211.950 ;
        RECT 326.100 210.150 327.900 211.950 ;
        RECT 328.950 210.450 331.050 211.050 ;
        RECT 334.950 210.450 337.050 211.050 ;
        RECT 328.950 209.550 337.050 210.450 ;
        RECT 328.950 208.950 331.050 209.550 ;
        RECT 334.950 208.950 337.050 209.550 ;
        RECT 318.000 207.000 321.300 208.200 ;
        RECT 299.700 198.600 301.500 207.000 ;
        RECT 319.500 198.600 321.300 207.000 ;
        RECT 326.100 198.000 327.900 207.600 ;
        RECT 341.700 201.600 342.900 211.950 ;
        RECT 365.100 210.150 366.900 211.950 ;
        RECT 368.700 207.600 369.900 211.950 ;
        RECT 371.100 210.150 372.900 211.950 ;
        RECT 377.550 211.050 378.450 218.550 ;
        RECT 386.100 214.050 387.900 215.850 ;
        RECT 392.700 214.050 393.900 221.400 ;
        RECT 413.100 214.050 414.900 215.850 ;
        RECT 419.100 214.050 420.000 226.200 ;
        RECT 437.100 214.050 438.900 215.850 ;
        RECT 443.100 214.050 444.000 226.200 ;
        RECT 457.950 219.450 460.050 220.050 ;
        RECT 466.950 219.450 469.050 219.900 ;
        RECT 457.950 218.550 469.050 219.450 ;
        RECT 457.950 217.950 460.050 218.550 ;
        RECT 466.950 217.800 469.050 218.550 ;
        RECT 464.100 214.050 465.900 215.850 ;
        RECT 470.100 214.050 471.000 226.200 ;
        RECT 485.100 221.400 486.900 233.400 ;
        RECT 488.100 222.300 489.900 233.400 ;
        RECT 491.100 223.200 492.900 234.000 ;
        RECT 494.100 222.300 495.900 233.400 ;
        RECT 488.100 221.400 495.900 222.300 ;
        RECT 509.100 221.400 510.900 233.400 ;
        RECT 512.100 222.000 513.900 234.000 ;
        RECT 515.100 227.400 516.900 233.400 ;
        RECT 518.100 227.400 519.900 234.000 ;
        RECT 536.100 227.400 537.900 234.000 ;
        RECT 539.100 227.400 540.900 233.400 ;
        RECT 542.100 228.000 543.900 234.000 ;
        RECT 485.400 214.050 486.300 221.400 ;
        RECT 490.950 214.050 492.750 215.850 ;
        RECT 509.700 214.050 510.600 221.400 ;
        RECT 513.000 214.050 514.800 215.850 ;
        RECT 385.950 211.950 388.050 214.050 ;
        RECT 388.950 211.950 391.050 214.050 ;
        RECT 391.950 211.950 394.050 214.050 ;
        RECT 394.950 211.950 397.050 214.050 ;
        RECT 409.950 211.950 412.050 214.050 ;
        RECT 412.950 211.950 415.050 214.050 ;
        RECT 415.950 211.950 418.050 214.050 ;
        RECT 418.950 211.950 421.050 214.050 ;
        RECT 433.950 211.950 436.050 214.050 ;
        RECT 436.950 211.950 439.050 214.050 ;
        RECT 439.950 211.950 442.050 214.050 ;
        RECT 442.950 211.950 445.050 214.050 ;
        RECT 460.950 211.950 463.050 214.050 ;
        RECT 463.950 211.950 466.050 214.050 ;
        RECT 466.950 211.950 469.050 214.050 ;
        RECT 469.950 211.950 472.050 214.050 ;
        RECT 484.950 211.950 487.050 214.050 ;
        RECT 487.950 211.950 490.050 214.050 ;
        RECT 490.950 211.950 493.050 214.050 ;
        RECT 493.950 211.950 496.050 214.050 ;
        RECT 509.100 211.950 511.200 214.050 ;
        RECT 512.400 211.950 514.500 214.050 ;
        RECT 373.950 209.550 378.450 211.050 ;
        RECT 389.100 210.150 390.900 211.950 ;
        RECT 373.950 208.950 378.000 209.550 ;
        RECT 392.700 207.600 393.900 211.950 ;
        RECT 395.100 210.150 396.900 211.950 ;
        RECT 410.100 210.150 411.900 211.950 ;
        RECT 416.100 210.150 417.900 211.950 ;
        RECT 419.100 208.200 420.000 211.950 ;
        RECT 434.100 210.150 435.900 211.950 ;
        RECT 440.100 210.150 441.900 211.950 ;
        RECT 443.100 208.200 444.000 211.950 ;
        RECT 461.100 210.150 462.900 211.950 ;
        RECT 467.100 210.150 468.900 211.950 ;
        RECT 470.100 208.200 471.000 211.950 ;
        RECT 368.700 206.700 372.300 207.600 ;
        RECT 392.700 206.700 396.300 207.600 ;
        RECT 362.100 203.700 369.900 205.050 ;
        RECT 341.100 198.600 342.900 201.600 ;
        RECT 344.100 198.000 345.900 201.600 ;
        RECT 362.100 198.600 363.900 203.700 ;
        RECT 365.100 198.000 366.900 202.800 ;
        RECT 368.100 198.600 369.900 203.700 ;
        RECT 371.100 204.600 372.300 206.700 ;
        RECT 371.100 198.600 372.900 204.600 ;
        RECT 386.100 203.700 393.900 205.050 ;
        RECT 386.100 198.600 387.900 203.700 ;
        RECT 389.100 198.000 390.900 202.800 ;
        RECT 392.100 198.600 393.900 203.700 ;
        RECT 395.100 204.600 396.300 206.700 ;
        RECT 395.100 198.600 396.900 204.600 ;
        RECT 410.100 198.000 411.900 207.600 ;
        RECT 416.700 207.000 420.000 208.200 ;
        RECT 416.700 198.600 418.500 207.000 ;
        RECT 434.100 198.000 435.900 207.600 ;
        RECT 440.700 207.000 444.000 208.200 ;
        RECT 440.700 198.600 442.500 207.000 ;
        RECT 461.100 198.000 462.900 207.600 ;
        RECT 467.700 207.000 471.000 208.200 ;
        RECT 467.700 198.600 469.500 207.000 ;
        RECT 485.400 204.600 486.300 211.950 ;
        RECT 487.950 210.150 489.750 211.950 ;
        RECT 494.100 210.150 495.900 211.950 ;
        RECT 509.700 204.600 510.600 211.950 ;
        RECT 516.000 207.300 516.900 227.400 ;
        RECT 539.400 227.100 540.900 227.400 ;
        RECT 545.100 227.400 546.900 233.400 ;
        RECT 545.100 227.100 546.000 227.400 ;
        RECT 539.400 226.200 546.000 227.100 ;
        RECT 539.100 214.050 540.900 215.850 ;
        RECT 545.100 214.050 546.000 226.200 ;
        RECT 563.100 221.400 564.900 233.400 ;
        RECT 566.100 223.200 567.900 234.000 ;
        RECT 569.100 227.400 570.900 233.400 ;
        RECT 563.100 214.050 564.300 221.400 ;
        RECT 569.700 220.500 570.900 227.400 ;
        RECT 565.200 219.600 570.900 220.500 ;
        RECT 572.550 221.400 574.350 233.400 ;
        RECT 575.550 221.400 577.350 234.000 ;
        RECT 580.350 227.400 582.150 233.400 ;
        RECT 584.850 227.400 586.650 234.000 ;
        RECT 580.350 225.300 582.450 227.400 ;
        RECT 587.850 226.500 589.650 233.400 ;
        RECT 590.850 227.400 592.650 234.000 ;
        RECT 586.950 225.450 593.550 226.500 ;
        RECT 586.950 224.700 588.750 225.450 ;
        RECT 591.750 224.700 593.550 225.450 ;
        RECT 595.650 224.400 597.450 233.400 ;
        RECT 579.450 222.600 582.450 224.400 ;
        RECT 583.350 223.800 585.150 224.400 ;
        RECT 583.350 222.900 589.050 223.800 ;
        RECT 595.650 223.500 597.750 224.400 ;
        RECT 583.350 222.600 585.150 222.900 ;
        RECT 581.250 221.700 582.450 222.600 ;
        RECT 565.200 218.700 567.000 219.600 ;
        RECT 517.800 211.950 519.900 214.050 ;
        RECT 535.950 211.950 538.050 214.050 ;
        RECT 538.950 211.950 541.050 214.050 ;
        RECT 541.950 211.950 544.050 214.050 ;
        RECT 544.950 211.950 547.050 214.050 ;
        RECT 563.100 211.950 565.200 214.050 ;
        RECT 517.950 210.150 519.750 211.950 ;
        RECT 536.100 210.150 537.900 211.950 ;
        RECT 542.100 210.150 543.900 211.950 ;
        RECT 545.100 208.200 546.000 211.950 ;
        RECT 511.500 206.400 519.900 207.300 ;
        RECT 511.500 205.500 513.300 206.400 ;
        RECT 485.400 203.400 490.500 204.600 ;
        RECT 485.700 198.000 487.500 201.600 ;
        RECT 488.700 198.600 490.500 203.400 ;
        RECT 493.200 198.000 495.000 204.600 ;
        RECT 509.700 202.800 512.400 204.600 ;
        RECT 510.600 198.600 512.400 202.800 ;
        RECT 513.600 198.000 515.400 204.600 ;
        RECT 518.100 198.600 519.900 206.400 ;
        RECT 536.100 198.000 537.900 207.600 ;
        RECT 542.700 207.000 546.000 208.200 ;
        RECT 542.700 198.600 544.500 207.000 ;
        RECT 563.100 204.600 564.300 211.950 ;
        RECT 566.100 207.300 567.000 218.700 ;
        RECT 568.800 214.050 570.600 215.850 ;
        RECT 568.500 211.950 570.600 214.050 ;
        RECT 572.550 214.050 573.750 221.400 ;
        RECT 581.250 220.800 586.050 221.700 ;
        RECT 574.650 218.100 576.450 218.550 ;
        RECT 580.350 218.100 582.450 218.700 ;
        RECT 574.650 216.900 582.450 218.100 ;
        RECT 574.650 216.750 576.450 216.900 ;
        RECT 580.350 216.600 582.450 216.900 ;
        RECT 572.550 213.750 577.050 214.050 ;
        RECT 572.550 211.950 578.850 213.750 ;
        RECT 565.200 206.400 567.000 207.300 ;
        RECT 565.200 205.500 570.900 206.400 ;
        RECT 563.100 198.600 564.900 204.600 ;
        RECT 566.100 198.000 567.900 204.600 ;
        RECT 569.700 201.600 570.900 205.500 ;
        RECT 569.100 198.600 570.900 201.600 ;
        RECT 572.550 204.600 573.750 211.950 ;
        RECT 585.150 208.200 586.050 220.800 ;
        RECT 588.150 220.800 589.050 222.900 ;
        RECT 589.950 222.300 597.750 223.500 ;
        RECT 589.950 221.700 591.750 222.300 ;
        RECT 601.050 221.400 602.850 234.000 ;
        RECT 604.050 223.200 605.850 233.400 ;
        RECT 604.050 221.400 606.450 223.200 ;
        RECT 588.150 220.500 596.550 220.800 ;
        RECT 605.550 220.500 606.450 221.400 ;
        RECT 588.150 219.900 606.450 220.500 ;
        RECT 594.750 219.300 606.450 219.900 ;
        RECT 594.750 219.000 596.550 219.300 ;
        RECT 592.800 212.400 594.900 214.050 ;
        RECT 592.800 211.200 600.900 212.400 ;
        RECT 601.950 211.950 604.050 214.050 ;
        RECT 599.100 210.600 600.900 211.200 ;
        RECT 596.100 209.400 597.900 210.000 ;
        RECT 602.250 209.400 604.050 211.950 ;
        RECT 596.100 208.200 604.050 209.400 ;
        RECT 585.150 207.000 597.150 208.200 ;
        RECT 585.150 206.400 586.950 207.000 ;
        RECT 596.100 205.200 597.150 207.000 ;
        RECT 572.550 198.600 574.350 204.600 ;
        RECT 575.850 198.000 577.650 204.600 ;
        RECT 580.350 201.600 582.750 203.700 ;
        RECT 592.350 203.550 594.150 204.300 ;
        RECT 589.200 202.500 594.150 203.550 ;
        RECT 595.350 203.400 597.150 205.200 ;
        RECT 605.550 204.600 606.450 219.300 ;
        RECT 589.200 201.600 590.250 202.500 ;
        RECT 598.050 202.200 600.150 203.700 ;
        RECT 596.250 201.600 600.150 202.200 ;
        RECT 580.950 198.600 582.750 201.600 ;
        RECT 585.450 198.000 587.250 201.600 ;
        RECT 588.450 198.600 590.250 201.600 ;
        RECT 591.750 198.000 593.550 201.600 ;
        RECT 596.250 200.700 599.850 201.600 ;
        RECT 596.250 198.600 598.050 200.700 ;
        RECT 601.050 198.000 602.850 204.600 ;
        RECT 604.050 202.800 606.450 204.600 ;
        RECT 608.550 221.400 610.350 233.400 ;
        RECT 611.550 221.400 613.350 234.000 ;
        RECT 616.350 227.400 618.150 233.400 ;
        RECT 620.850 227.400 622.650 234.000 ;
        RECT 616.350 225.300 618.450 227.400 ;
        RECT 623.850 226.500 625.650 233.400 ;
        RECT 626.850 227.400 628.650 234.000 ;
        RECT 622.950 225.450 629.550 226.500 ;
        RECT 622.950 224.700 624.750 225.450 ;
        RECT 627.750 224.700 629.550 225.450 ;
        RECT 631.650 224.400 633.450 233.400 ;
        RECT 615.450 222.600 618.450 224.400 ;
        RECT 619.350 223.800 621.150 224.400 ;
        RECT 619.350 222.900 625.050 223.800 ;
        RECT 631.650 223.500 633.750 224.400 ;
        RECT 619.350 222.600 621.150 222.900 ;
        RECT 617.250 221.700 618.450 222.600 ;
        RECT 608.550 214.050 609.750 221.400 ;
        RECT 617.250 220.800 622.050 221.700 ;
        RECT 610.650 218.100 612.450 218.550 ;
        RECT 616.350 218.100 618.450 218.700 ;
        RECT 610.650 216.900 618.450 218.100 ;
        RECT 610.650 216.750 612.450 216.900 ;
        RECT 616.350 216.600 618.450 216.900 ;
        RECT 608.550 213.750 613.050 214.050 ;
        RECT 608.550 211.950 614.850 213.750 ;
        RECT 608.550 204.600 609.750 211.950 ;
        RECT 621.150 208.200 622.050 220.800 ;
        RECT 624.150 220.800 625.050 222.900 ;
        RECT 625.950 222.300 633.750 223.500 ;
        RECT 625.950 221.700 627.750 222.300 ;
        RECT 637.050 221.400 638.850 234.000 ;
        RECT 640.050 223.200 641.850 233.400 ;
        RECT 656.700 227.400 658.500 234.000 ;
        RECT 657.000 224.100 658.800 225.900 ;
        RECT 640.050 221.400 642.450 223.200 ;
        RECT 659.700 222.900 661.500 233.400 ;
        RECT 624.150 220.500 632.550 220.800 ;
        RECT 641.550 220.500 642.450 221.400 ;
        RECT 624.150 219.900 642.450 220.500 ;
        RECT 630.750 219.300 642.450 219.900 ;
        RECT 630.750 219.000 632.550 219.300 ;
        RECT 628.800 212.400 630.900 214.050 ;
        RECT 628.800 211.200 636.900 212.400 ;
        RECT 637.950 211.950 640.050 214.050 ;
        RECT 635.100 210.600 636.900 211.200 ;
        RECT 632.100 209.400 633.900 210.000 ;
        RECT 638.250 209.400 640.050 211.950 ;
        RECT 632.100 208.200 640.050 209.400 ;
        RECT 621.150 207.000 633.150 208.200 ;
        RECT 621.150 206.400 622.950 207.000 ;
        RECT 632.100 205.200 633.150 207.000 ;
        RECT 604.050 198.600 605.850 202.800 ;
        RECT 608.550 198.600 610.350 204.600 ;
        RECT 611.850 198.000 613.650 204.600 ;
        RECT 616.350 201.600 618.750 203.700 ;
        RECT 628.350 203.550 630.150 204.300 ;
        RECT 625.200 202.500 630.150 203.550 ;
        RECT 631.350 203.400 633.150 205.200 ;
        RECT 641.550 204.600 642.450 219.300 ;
        RECT 659.100 221.400 661.500 222.900 ;
        RECT 664.800 221.400 666.600 234.000 ;
        RECT 680.100 221.400 681.900 233.400 ;
        RECT 683.100 222.300 684.900 233.400 ;
        RECT 686.100 223.200 687.900 234.000 ;
        RECT 689.100 222.300 690.900 233.400 ;
        RECT 704.100 227.400 705.900 234.000 ;
        RECT 707.100 227.400 708.900 233.400 ;
        RECT 725.700 227.400 727.500 234.000 ;
        RECT 683.100 221.400 690.900 222.300 ;
        RECT 659.100 214.050 660.300 221.400 ;
        RECT 661.950 219.450 664.050 220.050 ;
        RECT 661.950 218.550 669.450 219.450 ;
        RECT 661.950 217.950 664.050 218.550 ;
        RECT 668.550 216.450 669.450 218.550 ;
        RECT 665.100 214.050 666.900 215.850 ;
        RECT 668.550 215.550 672.450 216.450 ;
        RECT 655.950 211.950 658.050 214.050 ;
        RECT 658.950 211.950 661.050 214.050 ;
        RECT 661.950 211.950 664.050 214.050 ;
        RECT 664.950 211.950 667.050 214.050 ;
        RECT 656.100 210.150 657.900 211.950 ;
        RECT 659.100 207.600 660.300 211.950 ;
        RECT 662.100 210.150 663.900 211.950 ;
        RECT 671.550 210.450 672.450 215.550 ;
        RECT 680.400 214.050 681.300 221.400 ;
        RECT 685.950 214.050 687.750 215.850 ;
        RECT 704.100 214.050 705.900 215.850 ;
        RECT 707.100 214.050 708.300 227.400 ;
        RECT 726.000 224.100 727.800 225.900 ;
        RECT 728.700 222.900 730.500 233.400 ;
        RECT 728.100 221.400 730.500 222.900 ;
        RECT 733.800 221.400 735.600 234.000 ;
        RECT 749.100 227.400 750.900 233.400 ;
        RECT 752.100 228.000 753.900 234.000 ;
        RECT 750.000 227.100 750.900 227.400 ;
        RECT 755.100 227.400 756.900 233.400 ;
        RECT 758.100 227.400 759.900 234.000 ;
        RECT 755.100 227.100 756.600 227.400 ;
        RECT 750.000 226.200 756.600 227.100 ;
        RECT 728.100 214.050 729.300 221.400 ;
        RECT 734.100 214.050 735.900 215.850 ;
        RECT 750.000 214.050 750.900 226.200 ;
        RECT 776.100 221.400 777.900 233.400 ;
        RECT 779.100 222.300 780.900 233.400 ;
        RECT 782.100 223.200 783.900 234.000 ;
        RECT 785.100 222.300 786.900 233.400 ;
        RECT 779.100 221.400 786.900 222.300 ;
        RECT 800.400 221.400 802.200 234.000 ;
        RECT 805.500 222.900 807.300 233.400 ;
        RECT 808.500 227.400 810.300 234.000 ;
        RECT 808.200 224.100 810.000 225.900 ;
        RECT 805.500 221.400 807.900 222.900 ;
        RECT 763.950 216.450 766.050 217.050 ;
        RECT 769.950 216.450 772.050 217.050 ;
        RECT 755.100 214.050 756.900 215.850 ;
        RECT 763.950 215.550 772.050 216.450 ;
        RECT 763.950 214.950 766.050 215.550 ;
        RECT 769.950 214.950 772.050 215.550 ;
        RECT 776.400 214.050 777.300 221.400 ;
        RECT 793.950 219.450 796.050 220.050 ;
        RECT 799.950 219.450 802.050 220.050 ;
        RECT 793.950 218.550 802.050 219.450 ;
        RECT 793.950 217.950 796.050 218.550 ;
        RECT 799.950 217.950 802.050 218.550 ;
        RECT 781.950 214.050 783.750 215.850 ;
        RECT 800.100 214.050 801.900 215.850 ;
        RECT 806.700 214.050 807.900 221.400 ;
        RECT 808.950 222.450 811.050 223.050 ;
        RECT 814.950 222.450 817.050 223.050 ;
        RECT 808.950 221.550 817.050 222.450 ;
        RECT 808.950 220.950 811.050 221.550 ;
        RECT 814.950 220.950 817.050 221.550 ;
        RECT 824.400 221.400 826.200 234.000 ;
        RECT 829.500 222.900 831.300 233.400 ;
        RECT 832.500 227.400 834.300 234.000 ;
        RECT 832.200 224.100 834.000 225.900 ;
        RECT 829.500 221.400 831.900 222.900 ;
        RECT 849.000 222.600 850.800 233.400 ;
        RECT 849.000 221.400 852.600 222.600 ;
        RECT 854.100 221.400 855.900 234.000 ;
        RECT 872.100 227.400 873.900 234.000 ;
        RECT 875.100 227.400 876.900 233.400 ;
        RECT 878.100 227.400 879.900 234.000 ;
        RECT 817.950 219.450 820.050 219.900 ;
        RECT 823.950 219.450 826.050 220.050 ;
        RECT 817.950 218.550 826.050 219.450 ;
        RECT 817.950 217.800 820.050 218.550 ;
        RECT 823.950 217.950 826.050 218.550 ;
        RECT 824.100 214.050 825.900 215.850 ;
        RECT 830.700 214.050 831.900 221.400 ;
        RECT 835.950 219.450 838.050 220.050 ;
        RECT 847.950 219.450 850.050 220.050 ;
        RECT 835.950 218.550 850.050 219.450 ;
        RECT 835.950 217.950 838.050 218.550 ;
        RECT 847.950 217.950 850.050 218.550 ;
        RECT 835.950 216.450 838.050 216.900 ;
        RECT 841.950 216.450 844.050 217.050 ;
        RECT 835.950 215.550 844.050 216.450 ;
        RECT 835.950 214.800 838.050 215.550 ;
        RECT 841.950 214.950 844.050 215.550 ;
        RECT 848.100 214.050 849.900 215.850 ;
        RECT 851.700 214.050 852.600 221.400 ;
        RECT 865.950 219.450 868.050 220.050 ;
        RECT 871.950 219.450 874.050 220.050 ;
        RECT 865.950 218.550 874.050 219.450 ;
        RECT 865.950 217.950 868.050 218.550 ;
        RECT 871.950 217.950 874.050 218.550 ;
        RECT 853.950 214.050 855.750 215.850 ;
        RECT 875.100 214.050 876.300 227.400 ;
        RECT 679.950 211.950 682.050 214.050 ;
        RECT 682.950 211.950 685.050 214.050 ;
        RECT 685.950 211.950 688.050 214.050 ;
        RECT 688.950 211.950 691.050 214.050 ;
        RECT 703.950 211.950 706.050 214.050 ;
        RECT 706.950 211.950 709.050 214.050 ;
        RECT 724.950 211.950 727.050 214.050 ;
        RECT 727.950 211.950 730.050 214.050 ;
        RECT 730.950 211.950 733.050 214.050 ;
        RECT 733.950 211.950 736.050 214.050 ;
        RECT 748.950 211.950 751.050 214.050 ;
        RECT 751.950 211.950 754.050 214.050 ;
        RECT 754.950 211.950 757.050 214.050 ;
        RECT 757.950 211.950 760.050 214.050 ;
        RECT 775.950 211.950 778.050 214.050 ;
        RECT 778.950 211.950 781.050 214.050 ;
        RECT 781.950 211.950 784.050 214.050 ;
        RECT 784.950 211.950 787.050 214.050 ;
        RECT 799.950 211.950 802.050 214.050 ;
        RECT 802.950 211.950 805.050 214.050 ;
        RECT 805.950 211.950 808.050 214.050 ;
        RECT 808.950 211.950 811.050 214.050 ;
        RECT 823.950 211.950 826.050 214.050 ;
        RECT 826.950 211.950 829.050 214.050 ;
        RECT 829.950 211.950 832.050 214.050 ;
        RECT 832.950 211.950 835.050 214.050 ;
        RECT 847.950 211.950 850.050 214.050 ;
        RECT 850.950 211.950 853.050 214.050 ;
        RECT 853.950 211.950 856.050 214.050 ;
        RECT 871.950 211.950 874.050 214.050 ;
        RECT 874.950 211.950 877.050 214.050 ;
        RECT 877.950 211.950 880.050 214.050 ;
        RECT 676.950 210.450 679.050 211.050 ;
        RECT 671.550 209.550 679.050 210.450 ;
        RECT 676.950 208.950 679.050 209.550 ;
        RECT 656.700 206.700 660.300 207.600 ;
        RECT 656.700 204.600 657.900 206.700 ;
        RECT 625.200 201.600 626.250 202.500 ;
        RECT 634.050 202.200 636.150 203.700 ;
        RECT 632.250 201.600 636.150 202.200 ;
        RECT 616.950 198.600 618.750 201.600 ;
        RECT 621.450 198.000 623.250 201.600 ;
        RECT 624.450 198.600 626.250 201.600 ;
        RECT 627.750 198.000 629.550 201.600 ;
        RECT 632.250 200.700 635.850 201.600 ;
        RECT 632.250 198.600 634.050 200.700 ;
        RECT 637.050 198.000 638.850 204.600 ;
        RECT 640.050 202.800 642.450 204.600 ;
        RECT 640.050 198.600 641.850 202.800 ;
        RECT 656.100 198.600 657.900 204.600 ;
        RECT 659.100 203.700 666.900 205.050 ;
        RECT 659.100 198.600 660.900 203.700 ;
        RECT 662.100 198.000 663.900 202.800 ;
        RECT 665.100 198.600 666.900 203.700 ;
        RECT 680.400 204.600 681.300 211.950 ;
        RECT 682.950 210.150 684.750 211.950 ;
        RECT 689.100 210.150 690.900 211.950 ;
        RECT 680.400 203.400 685.500 204.600 ;
        RECT 680.700 198.000 682.500 201.600 ;
        RECT 683.700 198.600 685.500 203.400 ;
        RECT 688.200 198.000 690.000 204.600 ;
        RECT 707.100 201.600 708.300 211.950 ;
        RECT 725.100 210.150 726.900 211.950 ;
        RECT 728.100 207.600 729.300 211.950 ;
        RECT 731.100 210.150 732.900 211.950 ;
        RECT 725.700 206.700 729.300 207.600 ;
        RECT 750.000 208.200 750.900 211.950 ;
        RECT 752.100 210.150 753.900 211.950 ;
        RECT 758.100 210.150 759.900 211.950 ;
        RECT 769.950 210.450 772.050 211.050 ;
        RECT 761.550 210.000 772.050 210.450 ;
        RECT 760.950 209.550 772.050 210.000 ;
        RECT 750.000 207.000 753.300 208.200 ;
        RECT 709.950 204.450 712.050 205.050 ;
        RECT 718.950 204.450 721.050 205.050 ;
        RECT 725.700 204.600 726.900 206.700 ;
        RECT 709.950 203.550 721.050 204.450 ;
        RECT 709.950 202.950 712.050 203.550 ;
        RECT 718.950 202.950 721.050 203.550 ;
        RECT 704.100 198.000 705.900 201.600 ;
        RECT 707.100 198.600 708.900 201.600 ;
        RECT 725.100 198.600 726.900 204.600 ;
        RECT 728.100 203.700 735.900 205.050 ;
        RECT 728.100 198.600 729.900 203.700 ;
        RECT 731.100 198.000 732.900 202.800 ;
        RECT 734.100 198.600 735.900 203.700 ;
        RECT 751.500 198.600 753.300 207.000 ;
        RECT 758.100 198.000 759.900 207.600 ;
        RECT 760.950 205.950 763.050 209.550 ;
        RECT 769.950 208.950 772.050 209.550 ;
        RECT 776.400 204.600 777.300 211.950 ;
        RECT 778.950 210.150 780.750 211.950 ;
        RECT 785.100 210.150 786.900 211.950 ;
        RECT 803.100 210.150 804.900 211.950 ;
        RECT 806.700 207.600 807.900 211.950 ;
        RECT 809.100 210.150 810.900 211.950 ;
        RECT 827.100 210.150 828.900 211.950 ;
        RECT 830.700 207.600 831.900 211.950 ;
        RECT 833.100 210.150 834.900 211.950 ;
        RECT 806.700 206.700 810.300 207.600 ;
        RECT 830.700 206.700 834.300 207.600 ;
        RECT 776.400 203.400 781.500 204.600 ;
        RECT 776.700 198.000 778.500 201.600 ;
        RECT 779.700 198.600 781.500 203.400 ;
        RECT 784.200 198.000 786.000 204.600 ;
        RECT 800.100 203.700 807.900 205.050 ;
        RECT 800.100 198.600 801.900 203.700 ;
        RECT 803.100 198.000 804.900 202.800 ;
        RECT 806.100 198.600 807.900 203.700 ;
        RECT 809.100 204.600 810.300 206.700 ;
        RECT 809.100 198.600 810.900 204.600 ;
        RECT 824.100 203.700 831.900 205.050 ;
        RECT 824.100 198.600 825.900 203.700 ;
        RECT 827.100 198.000 828.900 202.800 ;
        RECT 830.100 198.600 831.900 203.700 ;
        RECT 833.100 204.600 834.300 206.700 ;
        RECT 833.100 198.600 834.900 204.600 ;
        RECT 851.700 201.600 852.600 211.950 ;
        RECT 872.250 210.150 874.050 211.950 ;
        RECT 853.950 207.450 856.050 208.050 ;
        RECT 865.950 207.450 868.050 208.050 ;
        RECT 853.950 206.550 868.050 207.450 ;
        RECT 853.950 205.950 856.050 206.550 ;
        RECT 865.950 205.950 868.050 206.550 ;
        RECT 875.100 206.700 876.300 211.950 ;
        RECT 878.100 210.150 879.900 211.950 ;
        RECT 875.100 205.800 879.300 206.700 ;
        RECT 848.100 198.000 849.900 201.600 ;
        RECT 851.100 198.600 852.900 201.600 ;
        RECT 854.100 198.000 855.900 201.600 ;
        RECT 872.400 198.000 874.200 204.600 ;
        RECT 877.500 198.600 879.300 205.800 ;
        RECT 14.400 188.400 16.200 195.000 ;
        RECT 19.500 187.200 21.300 194.400 ;
        RECT 35.100 191.400 36.900 194.400 ;
        RECT 38.100 191.400 39.900 195.000 ;
        RECT 17.100 186.300 21.300 187.200 ;
        RECT 14.250 181.050 16.050 182.850 ;
        RECT 17.100 181.050 18.300 186.300 ;
        RECT 20.100 181.050 21.900 182.850 ;
        RECT 35.700 181.050 36.900 191.400 ;
        RECT 53.400 188.400 55.200 195.000 ;
        RECT 58.500 187.200 60.300 194.400 ;
        RECT 56.100 186.300 60.300 187.200 ;
        RECT 74.700 187.200 76.500 194.400 ;
        RECT 79.800 188.400 81.600 195.000 ;
        RECT 74.700 186.300 78.900 187.200 ;
        RECT 53.250 181.050 55.050 182.850 ;
        RECT 56.100 181.050 57.300 186.300 ;
        RECT 59.100 181.050 60.900 182.850 ;
        RECT 74.100 181.050 75.900 182.850 ;
        RECT 77.700 181.050 78.900 186.300 ;
        RECT 100.500 186.000 102.300 194.400 ;
        RECT 99.000 184.800 102.300 186.000 ;
        RECT 107.100 185.400 108.900 195.000 ;
        RECT 122.100 188.400 123.900 194.400 ;
        RECT 122.700 186.300 123.900 188.400 ;
        RECT 125.100 189.300 126.900 194.400 ;
        RECT 128.100 190.200 129.900 195.000 ;
        RECT 131.100 189.300 132.900 194.400 ;
        RECT 125.100 187.950 132.900 189.300 ;
        RECT 146.100 188.400 147.900 194.400 ;
        RECT 149.100 189.300 150.900 195.000 ;
        RECT 153.600 188.400 155.400 194.400 ;
        RECT 158.100 189.300 159.900 195.000 ;
        RECT 161.100 188.400 162.900 194.400 ;
        RECT 179.100 191.400 180.900 195.000 ;
        RECT 182.100 191.400 183.900 194.400 ;
        RECT 185.100 191.400 186.900 195.000 ;
        RECT 200.100 191.400 201.900 195.000 ;
        RECT 203.100 191.400 204.900 194.400 ;
        RECT 146.100 187.500 150.900 188.400 ;
        RECT 148.800 186.300 150.900 187.500 ;
        RECT 153.900 186.900 155.100 188.400 ;
        RECT 122.700 185.400 126.300 186.300 ;
        RECT 79.950 181.050 81.750 182.850 ;
        RECT 99.000 181.050 99.900 184.800 ;
        RECT 101.100 181.050 102.900 182.850 ;
        RECT 107.100 181.050 108.900 182.850 ;
        RECT 122.100 181.050 123.900 182.850 ;
        RECT 125.100 181.050 126.300 185.400 ;
        RECT 152.100 184.800 155.100 186.900 ;
        RECT 161.100 186.600 162.300 188.400 ;
        RECT 128.100 181.050 129.900 182.850 ;
        RECT 150.900 181.800 153.000 183.900 ;
        RECT 13.950 178.950 16.050 181.050 ;
        RECT 16.950 178.950 19.050 181.050 ;
        RECT 19.950 178.950 22.050 181.050 ;
        RECT 34.950 178.950 37.050 181.050 ;
        RECT 37.950 178.950 40.050 181.050 ;
        RECT 52.950 178.950 55.050 181.050 ;
        RECT 55.950 178.950 58.050 181.050 ;
        RECT 58.950 178.950 61.050 181.050 ;
        RECT 73.950 178.950 76.050 181.050 ;
        RECT 76.950 178.950 79.050 181.050 ;
        RECT 79.950 178.950 82.050 181.050 ;
        RECT 97.950 178.950 100.050 181.050 ;
        RECT 100.950 178.950 103.050 181.050 ;
        RECT 103.950 178.950 106.050 181.050 ;
        RECT 106.950 178.950 109.050 181.050 ;
        RECT 121.950 178.950 124.050 181.050 ;
        RECT 124.950 178.950 127.050 181.050 ;
        RECT 127.950 178.950 130.050 181.050 ;
        RECT 130.950 178.950 133.050 181.050 ;
        RECT 146.100 178.950 148.200 181.050 ;
        RECT 150.900 180.000 152.700 181.800 ;
        RECT 153.900 179.100 155.100 184.800 ;
        RECT 156.000 185.700 162.300 186.600 ;
        RECT 156.000 183.600 158.100 185.700 ;
        RECT 156.000 181.800 157.800 183.600 ;
        RECT 160.800 181.050 162.600 182.850 ;
        RECT 182.700 181.050 183.600 191.400 ;
        RECT 203.100 181.050 204.300 191.400 ;
        RECT 218.100 189.300 219.900 194.400 ;
        RECT 221.100 190.200 222.900 195.000 ;
        RECT 224.100 189.300 225.900 194.400 ;
        RECT 218.100 187.950 225.900 189.300 ;
        RECT 227.100 188.400 228.900 194.400 ;
        RECT 242.100 189.300 243.900 194.400 ;
        RECT 245.100 190.200 246.900 195.000 ;
        RECT 248.100 189.300 249.900 194.400 ;
        RECT 227.100 186.300 228.300 188.400 ;
        RECT 242.100 187.950 249.900 189.300 ;
        RECT 251.100 188.400 252.900 194.400 ;
        RECT 266.100 191.400 267.900 194.400 ;
        RECT 269.100 191.400 270.900 195.000 ;
        RECT 251.100 186.300 252.300 188.400 ;
        RECT 224.700 185.400 228.300 186.300 ;
        RECT 248.700 185.400 252.300 186.300 ;
        RECT 221.100 181.050 222.900 182.850 ;
        RECT 224.700 181.050 225.900 185.400 ;
        RECT 227.100 181.050 228.900 182.850 ;
        RECT 245.100 181.050 246.900 182.850 ;
        RECT 248.700 181.050 249.900 185.400 ;
        RECT 251.100 181.050 252.900 182.850 ;
        RECT 266.700 181.050 267.900 191.400 ;
        RECT 286.500 186.000 288.300 194.400 ;
        RECT 285.000 184.800 288.300 186.000 ;
        RECT 293.100 185.400 294.900 195.000 ;
        RECT 309.000 188.400 310.800 195.000 ;
        RECT 313.500 189.600 315.300 194.400 ;
        RECT 316.500 191.400 318.300 195.000 ;
        RECT 313.500 188.400 318.600 189.600 ;
        RECT 285.000 181.050 285.900 184.800 ;
        RECT 287.100 181.050 288.900 182.850 ;
        RECT 293.100 181.050 294.900 182.850 ;
        RECT 308.100 181.050 309.900 182.850 ;
        RECT 314.250 181.050 316.050 182.850 ;
        RECT 317.700 181.050 318.600 188.400 ;
        RECT 335.100 186.600 336.900 194.400 ;
        RECT 339.600 188.400 341.400 195.000 ;
        RECT 342.600 190.200 344.400 194.400 ;
        RECT 363.600 190.200 365.400 194.400 ;
        RECT 342.600 188.400 345.300 190.200 ;
        RECT 341.700 186.600 343.500 187.500 ;
        RECT 335.100 185.700 343.500 186.600 ;
        RECT 335.250 181.050 337.050 182.850 ;
        RECT 160.800 180.300 162.900 181.050 ;
        RECT 17.100 165.600 18.300 178.950 ;
        RECT 35.700 165.600 36.900 178.950 ;
        RECT 38.100 177.150 39.900 178.950 ;
        RECT 43.950 174.450 46.050 175.050 ;
        RECT 52.950 174.450 55.050 175.050 ;
        RECT 43.950 173.550 55.050 174.450 ;
        RECT 43.950 172.950 46.050 173.550 ;
        RECT 52.950 172.950 55.050 173.550 ;
        RECT 56.100 165.600 57.300 178.950 ;
        RECT 77.700 165.600 78.900 178.950 ;
        RECT 82.950 177.450 85.050 178.050 ;
        RECT 88.950 177.450 91.050 178.050 ;
        RECT 82.950 176.550 91.050 177.450 ;
        RECT 82.950 175.950 85.050 176.550 ;
        RECT 88.950 175.950 91.050 176.550 ;
        RECT 99.000 166.800 99.900 178.950 ;
        RECT 104.100 177.150 105.900 178.950 ;
        RECT 125.100 171.600 126.300 178.950 ;
        RECT 131.100 177.150 132.900 178.950 ;
        RECT 146.400 177.150 148.200 178.950 ;
        RECT 152.700 178.200 155.100 179.100 ;
        RECT 156.000 178.950 162.900 180.300 ;
        RECT 178.950 178.950 181.050 181.050 ;
        RECT 181.950 178.950 184.050 181.050 ;
        RECT 184.950 178.950 187.050 181.050 ;
        RECT 199.950 178.950 202.050 181.050 ;
        RECT 202.950 178.950 205.050 181.050 ;
        RECT 217.950 178.950 220.050 181.050 ;
        RECT 220.950 178.950 223.050 181.050 ;
        RECT 223.950 178.950 226.050 181.050 ;
        RECT 226.950 178.950 229.050 181.050 ;
        RECT 241.950 178.950 244.050 181.050 ;
        RECT 244.950 178.950 247.050 181.050 ;
        RECT 247.950 178.950 250.050 181.050 ;
        RECT 250.950 178.950 253.050 181.050 ;
        RECT 265.950 178.950 268.050 181.050 ;
        RECT 268.950 178.950 271.050 181.050 ;
        RECT 283.950 178.950 286.050 181.050 ;
        RECT 286.950 178.950 289.050 181.050 ;
        RECT 289.950 178.950 292.050 181.050 ;
        RECT 292.950 178.950 295.050 181.050 ;
        RECT 307.950 178.950 310.050 181.050 ;
        RECT 310.950 178.950 313.050 181.050 ;
        RECT 313.950 178.950 316.050 181.050 ;
        RECT 316.950 178.950 319.050 181.050 ;
        RECT 335.100 178.950 337.200 181.050 ;
        RECT 156.000 178.500 157.800 178.950 ;
        RECT 152.700 178.050 154.200 178.200 ;
        RECT 152.100 175.950 154.200 178.050 ;
        RECT 153.300 174.000 154.200 175.950 ;
        RECT 155.100 175.500 159.000 177.300 ;
        RECT 179.100 177.150 180.900 178.950 ;
        RECT 155.100 175.200 157.200 175.500 ;
        RECT 153.300 172.950 154.800 174.000 ;
        RECT 148.800 171.600 150.900 172.500 ;
        RECT 125.100 170.100 127.500 171.600 ;
        RECT 123.000 167.100 124.800 168.900 ;
        RECT 99.000 165.900 105.600 166.800 ;
        RECT 99.000 165.600 99.900 165.900 ;
        RECT 14.100 159.000 15.900 165.600 ;
        RECT 17.100 159.600 18.900 165.600 ;
        RECT 20.100 159.000 21.900 165.600 ;
        RECT 35.100 159.600 36.900 165.600 ;
        RECT 38.100 159.000 39.900 165.600 ;
        RECT 53.100 159.000 54.900 165.600 ;
        RECT 56.100 159.600 57.900 165.600 ;
        RECT 59.100 159.000 60.900 165.600 ;
        RECT 74.100 159.000 75.900 165.600 ;
        RECT 77.100 159.600 78.900 165.600 ;
        RECT 80.100 159.000 81.900 165.600 ;
        RECT 98.100 159.600 99.900 165.600 ;
        RECT 104.100 165.600 105.600 165.900 ;
        RECT 101.100 159.000 102.900 165.000 ;
        RECT 104.100 159.600 105.900 165.600 ;
        RECT 107.100 159.000 108.900 165.600 ;
        RECT 122.700 159.000 124.500 165.600 ;
        RECT 125.700 159.600 127.500 170.100 ;
        RECT 130.800 159.000 132.600 171.600 ;
        RECT 146.100 170.400 150.900 171.600 ;
        RECT 153.600 171.600 154.800 172.950 ;
        RECT 158.400 171.600 160.500 173.700 ;
        RECT 182.700 171.600 183.600 178.950 ;
        RECT 184.950 177.150 186.750 178.950 ;
        RECT 200.100 177.150 201.900 178.950 ;
        RECT 146.100 159.600 147.900 170.400 ;
        RECT 149.100 159.000 150.900 169.500 ;
        RECT 153.600 159.600 155.400 171.600 ;
        RECT 158.400 170.700 162.900 171.600 ;
        RECT 158.100 159.000 159.900 169.500 ;
        RECT 161.100 159.600 162.900 170.700 ;
        RECT 180.000 170.400 183.600 171.600 ;
        RECT 180.000 159.600 181.800 170.400 ;
        RECT 185.100 159.000 186.900 171.600 ;
        RECT 203.100 165.600 204.300 178.950 ;
        RECT 218.100 177.150 219.900 178.950 ;
        RECT 224.700 171.600 225.900 178.950 ;
        RECT 242.100 177.150 243.900 178.950 ;
        RECT 248.700 171.600 249.900 178.950 ;
        RECT 250.950 174.450 253.050 175.050 ;
        RECT 262.950 174.450 265.050 175.050 ;
        RECT 250.950 173.550 265.050 174.450 ;
        RECT 250.950 172.950 253.050 173.550 ;
        RECT 262.950 172.950 265.050 173.550 ;
        RECT 200.100 159.000 201.900 165.600 ;
        RECT 203.100 159.600 204.900 165.600 ;
        RECT 218.400 159.000 220.200 171.600 ;
        RECT 223.500 170.100 225.900 171.600 ;
        RECT 223.500 159.600 225.300 170.100 ;
        RECT 226.200 167.100 228.000 168.900 ;
        RECT 226.500 159.000 228.300 165.600 ;
        RECT 242.400 159.000 244.200 171.600 ;
        RECT 247.500 170.100 249.900 171.600 ;
        RECT 247.500 159.600 249.300 170.100 ;
        RECT 250.200 167.100 252.000 168.900 ;
        RECT 266.700 165.600 267.900 178.950 ;
        RECT 269.100 177.150 270.900 178.950 ;
        RECT 285.000 166.800 285.900 178.950 ;
        RECT 290.100 177.150 291.900 178.950 ;
        RECT 311.250 177.150 313.050 178.950 ;
        RECT 317.700 171.600 318.600 178.950 ;
        RECT 308.100 170.700 315.900 171.600 ;
        RECT 285.000 165.900 291.600 166.800 ;
        RECT 285.000 165.600 285.900 165.900 ;
        RECT 250.500 159.000 252.300 165.600 ;
        RECT 266.100 159.600 267.900 165.600 ;
        RECT 269.100 159.000 270.900 165.600 ;
        RECT 284.100 159.600 285.900 165.600 ;
        RECT 290.100 165.600 291.600 165.900 ;
        RECT 287.100 159.000 288.900 165.000 ;
        RECT 290.100 159.600 291.900 165.600 ;
        RECT 293.100 159.000 294.900 165.600 ;
        RECT 308.100 159.600 309.900 170.700 ;
        RECT 311.100 159.000 312.900 169.800 ;
        RECT 314.100 159.600 315.900 170.700 ;
        RECT 317.100 159.600 318.900 171.600 ;
        RECT 338.100 165.600 339.000 185.700 ;
        RECT 344.400 181.050 345.300 188.400 ;
        RECT 362.700 188.400 365.400 190.200 ;
        RECT 366.600 188.400 368.400 195.000 ;
        RECT 362.700 181.050 363.600 188.400 ;
        RECT 364.500 186.600 366.300 187.500 ;
        RECT 371.100 186.600 372.900 194.400 ;
        RECT 387.000 188.400 388.800 195.000 ;
        RECT 391.500 189.600 393.300 194.400 ;
        RECT 394.500 191.400 396.300 195.000 ;
        RECT 410.100 191.400 411.900 195.000 ;
        RECT 413.100 191.400 414.900 194.400 ;
        RECT 416.100 191.400 417.900 195.000 ;
        RECT 391.500 188.400 396.600 189.600 ;
        RECT 364.500 185.700 372.900 186.600 ;
        RECT 340.500 178.950 342.600 181.050 ;
        RECT 343.800 178.950 345.900 181.050 ;
        RECT 362.100 178.950 364.200 181.050 ;
        RECT 365.400 178.950 367.500 181.050 ;
        RECT 340.200 177.150 342.000 178.950 ;
        RECT 344.400 171.600 345.300 178.950 ;
        RECT 362.700 171.600 363.600 178.950 ;
        RECT 366.000 177.150 367.800 178.950 ;
        RECT 335.100 159.000 336.900 165.600 ;
        RECT 338.100 159.600 339.900 165.600 ;
        RECT 341.100 159.000 342.900 171.000 ;
        RECT 344.100 159.600 345.900 171.600 ;
        RECT 362.100 159.600 363.900 171.600 ;
        RECT 365.100 159.000 366.900 171.000 ;
        RECT 369.000 165.600 369.900 185.700 ;
        RECT 370.950 181.050 372.750 182.850 ;
        RECT 386.100 181.050 387.900 182.850 ;
        RECT 392.250 181.050 394.050 182.850 ;
        RECT 395.700 181.050 396.600 188.400 ;
        RECT 413.400 181.050 414.300 191.400 ;
        RECT 431.100 189.300 432.900 194.400 ;
        RECT 434.100 190.200 435.900 195.000 ;
        RECT 437.100 189.300 438.900 194.400 ;
        RECT 431.100 187.950 438.900 189.300 ;
        RECT 440.100 188.400 441.900 194.400 ;
        RECT 440.100 186.300 441.300 188.400 ;
        RECT 455.700 187.200 457.500 194.400 ;
        RECT 460.800 188.400 462.600 195.000 ;
        RECT 476.100 191.400 477.900 195.000 ;
        RECT 479.100 191.400 480.900 194.400 ;
        RECT 455.700 186.300 459.900 187.200 ;
        RECT 437.700 185.400 441.300 186.300 ;
        RECT 434.100 181.050 435.900 182.850 ;
        RECT 437.700 181.050 438.900 185.400 ;
        RECT 442.950 183.450 447.000 184.050 ;
        RECT 440.100 181.050 441.900 182.850 ;
        RECT 442.950 181.950 447.450 183.450 ;
        RECT 370.800 178.950 372.900 181.050 ;
        RECT 385.950 178.950 388.050 181.050 ;
        RECT 388.950 178.950 391.050 181.050 ;
        RECT 391.950 178.950 394.050 181.050 ;
        RECT 394.950 178.950 397.050 181.050 ;
        RECT 409.950 178.950 412.050 181.050 ;
        RECT 412.950 178.950 415.050 181.050 ;
        RECT 415.950 178.950 418.050 181.050 ;
        RECT 430.950 178.950 433.050 181.050 ;
        RECT 433.950 178.950 436.050 181.050 ;
        RECT 436.950 178.950 439.050 181.050 ;
        RECT 439.950 178.950 442.050 181.050 ;
        RECT 389.250 177.150 391.050 178.950 ;
        RECT 373.950 174.450 376.050 175.050 ;
        RECT 391.950 174.450 394.050 175.050 ;
        RECT 373.950 173.550 394.050 174.450 ;
        RECT 373.950 172.950 376.050 173.550 ;
        RECT 391.950 172.950 394.050 173.550 ;
        RECT 395.700 171.600 396.600 178.950 ;
        RECT 410.250 177.150 412.050 178.950 ;
        RECT 413.400 171.600 414.300 178.950 ;
        RECT 416.100 177.150 417.900 178.950 ;
        RECT 431.100 177.150 432.900 178.950 ;
        RECT 437.700 171.600 438.900 178.950 ;
        RECT 446.550 178.050 447.450 181.950 ;
        RECT 455.100 181.050 456.900 182.850 ;
        RECT 458.700 181.050 459.900 186.300 ;
        RECT 460.950 181.050 462.750 182.850 ;
        RECT 479.100 181.050 480.300 191.400 ;
        RECT 494.100 185.400 495.900 195.000 ;
        RECT 500.700 186.000 502.500 194.400 ;
        RECT 520.500 186.000 522.300 194.400 ;
        RECT 500.700 184.800 504.000 186.000 ;
        RECT 494.100 181.050 495.900 182.850 ;
        RECT 500.100 181.050 501.900 182.850 ;
        RECT 503.100 181.050 504.000 184.800 ;
        RECT 519.000 184.800 522.300 186.000 ;
        RECT 527.100 185.400 528.900 195.000 ;
        RECT 545.100 191.400 546.900 195.000 ;
        RECT 548.100 191.400 549.900 194.400 ;
        RECT 563.100 191.400 564.900 195.000 ;
        RECT 566.100 191.400 567.900 194.400 ;
        RECT 569.100 191.400 570.900 195.000 ;
        RECT 519.000 181.050 519.900 184.800 ;
        RECT 521.100 181.050 522.900 182.850 ;
        RECT 527.100 181.050 528.900 182.850 ;
        RECT 548.100 181.050 549.300 191.400 ;
        RECT 566.400 181.050 567.300 191.400 ;
        RECT 585.000 188.400 586.800 195.000 ;
        RECT 589.500 189.600 591.300 194.400 ;
        RECT 592.500 191.400 594.300 195.000 ;
        RECT 589.500 188.400 594.600 189.600 ;
        RECT 608.100 188.400 609.900 194.400 ;
        RECT 611.100 189.300 612.900 195.000 ;
        RECT 615.600 188.400 617.400 194.400 ;
        RECT 620.100 189.300 621.900 195.000 ;
        RECT 623.100 188.400 624.900 194.400 ;
        RECT 639.000 188.400 640.800 195.000 ;
        RECT 643.500 189.600 645.300 194.400 ;
        RECT 646.500 191.400 648.300 195.000 ;
        RECT 673.200 191.400 675.900 194.400 ;
        RECT 677.100 191.400 678.900 195.000 ;
        RECT 680.100 191.400 681.900 194.400 ;
        RECT 683.100 191.400 685.200 195.000 ;
        RECT 673.200 190.500 674.100 191.400 ;
        RECT 680.400 190.500 681.300 191.400 ;
        RECT 668.700 189.600 681.300 190.500 ;
        RECT 643.500 188.400 648.600 189.600 ;
        RECT 571.950 183.450 574.050 184.050 ;
        RECT 577.950 183.450 580.050 184.050 ;
        RECT 571.950 182.550 580.050 183.450 ;
        RECT 571.950 181.950 574.050 182.550 ;
        RECT 577.950 181.950 580.050 182.550 ;
        RECT 584.100 181.050 585.900 182.850 ;
        RECT 590.250 181.050 592.050 182.850 ;
        RECT 593.700 181.050 594.600 188.400 ;
        RECT 608.700 186.600 609.900 188.400 ;
        RECT 615.900 186.900 617.100 188.400 ;
        RECT 620.100 187.500 624.900 188.400 ;
        RECT 608.700 185.700 615.000 186.600 ;
        RECT 612.900 183.600 615.000 185.700 ;
        RECT 608.400 181.050 610.200 182.850 ;
        RECT 613.200 181.800 615.000 183.600 ;
        RECT 615.900 184.800 618.900 186.900 ;
        RECT 620.100 186.300 622.200 187.500 ;
        RECT 454.950 178.950 457.050 181.050 ;
        RECT 457.950 178.950 460.050 181.050 ;
        RECT 460.950 178.950 463.050 181.050 ;
        RECT 475.950 178.950 478.050 181.050 ;
        RECT 478.950 178.950 481.050 181.050 ;
        RECT 493.950 178.950 496.050 181.050 ;
        RECT 496.950 178.950 499.050 181.050 ;
        RECT 499.950 178.950 502.050 181.050 ;
        RECT 502.950 178.950 505.050 181.050 ;
        RECT 517.950 178.950 520.050 181.050 ;
        RECT 520.950 178.950 523.050 181.050 ;
        RECT 523.950 178.950 526.050 181.050 ;
        RECT 526.950 178.950 529.050 181.050 ;
        RECT 544.950 178.950 547.050 181.050 ;
        RECT 547.950 178.950 550.050 181.050 ;
        RECT 562.950 178.950 565.050 181.050 ;
        RECT 565.950 178.950 568.050 181.050 ;
        RECT 568.950 178.950 571.050 181.050 ;
        RECT 583.950 178.950 586.050 181.050 ;
        RECT 586.950 178.950 589.050 181.050 ;
        RECT 589.950 178.950 592.050 181.050 ;
        RECT 592.950 178.950 595.050 181.050 ;
        RECT 608.100 180.300 610.200 181.050 ;
        RECT 608.100 178.950 615.000 180.300 ;
        RECT 442.950 176.550 447.450 178.050 ;
        RECT 442.950 175.950 447.000 176.550 ;
        RECT 448.950 174.450 451.050 175.050 ;
        RECT 454.950 174.450 457.050 175.050 ;
        RECT 448.950 173.550 457.050 174.450 ;
        RECT 448.950 172.950 451.050 173.550 ;
        RECT 454.950 172.950 457.050 173.550 ;
        RECT 386.100 170.700 393.900 171.600 ;
        RECT 368.100 159.600 369.900 165.600 ;
        RECT 371.100 159.000 372.900 165.600 ;
        RECT 386.100 159.600 387.900 170.700 ;
        RECT 389.100 159.000 390.900 169.800 ;
        RECT 392.100 159.600 393.900 170.700 ;
        RECT 395.100 159.600 396.900 171.600 ;
        RECT 410.100 159.000 411.900 171.600 ;
        RECT 413.400 170.400 417.000 171.600 ;
        RECT 415.200 159.600 417.000 170.400 ;
        RECT 431.400 159.000 433.200 171.600 ;
        RECT 436.500 170.100 438.900 171.600 ;
        RECT 436.500 159.600 438.300 170.100 ;
        RECT 439.200 167.100 441.000 168.900 ;
        RECT 458.700 165.600 459.900 178.950 ;
        RECT 476.100 177.150 477.900 178.950 ;
        RECT 460.950 174.450 463.050 175.050 ;
        RECT 466.950 174.450 469.050 175.050 ;
        RECT 460.950 173.550 469.050 174.450 ;
        RECT 460.950 172.950 463.050 173.550 ;
        RECT 466.950 172.950 469.050 173.550 ;
        RECT 479.100 165.600 480.300 178.950 ;
        RECT 497.100 177.150 498.900 178.950 ;
        RECT 484.950 174.450 487.050 175.050 ;
        RECT 499.950 174.450 502.050 175.050 ;
        RECT 484.950 173.550 502.050 174.450 ;
        RECT 484.950 172.950 487.050 173.550 ;
        RECT 499.950 172.950 502.050 173.550 ;
        RECT 503.100 166.800 504.000 178.950 ;
        RECT 497.400 165.900 504.000 166.800 ;
        RECT 497.400 165.600 498.900 165.900 ;
        RECT 439.500 159.000 441.300 165.600 ;
        RECT 455.100 159.000 456.900 165.600 ;
        RECT 458.100 159.600 459.900 165.600 ;
        RECT 461.100 159.000 462.900 165.600 ;
        RECT 476.100 159.000 477.900 165.600 ;
        RECT 479.100 159.600 480.900 165.600 ;
        RECT 494.100 159.000 495.900 165.600 ;
        RECT 497.100 159.600 498.900 165.600 ;
        RECT 503.100 165.600 504.000 165.900 ;
        RECT 519.000 166.800 519.900 178.950 ;
        RECT 524.100 177.150 525.900 178.950 ;
        RECT 545.100 177.150 546.900 178.950 ;
        RECT 519.000 165.900 525.600 166.800 ;
        RECT 519.000 165.600 519.900 165.900 ;
        RECT 500.100 159.000 501.900 165.000 ;
        RECT 503.100 159.600 504.900 165.600 ;
        RECT 518.100 159.600 519.900 165.600 ;
        RECT 524.100 165.600 525.600 165.900 ;
        RECT 548.100 165.600 549.300 178.950 ;
        RECT 563.250 177.150 565.050 178.950 ;
        RECT 566.400 171.600 567.300 178.950 ;
        RECT 569.100 177.150 570.900 178.950 ;
        RECT 587.250 177.150 589.050 178.950 ;
        RECT 593.700 171.600 594.600 178.950 ;
        RECT 613.200 178.500 615.000 178.950 ;
        RECT 615.900 179.100 617.100 184.800 ;
        RECT 618.000 181.800 620.100 183.900 ;
        RECT 618.300 180.000 620.100 181.800 ;
        RECT 638.100 181.050 639.900 182.850 ;
        RECT 644.250 181.050 646.050 182.850 ;
        RECT 647.700 181.050 648.600 188.400 ;
        RECT 668.700 181.050 669.900 189.600 ;
        RECT 682.950 189.450 685.050 190.050 ;
        RECT 691.950 189.450 694.050 190.050 ;
        RECT 682.950 188.550 694.050 189.450 ;
        RECT 682.950 187.950 685.050 188.550 ;
        RECT 691.950 187.950 694.050 188.550 ;
        RECT 701.100 188.400 702.900 194.400 ;
        RECT 673.950 186.450 676.050 187.050 ;
        RECT 694.950 186.450 697.050 187.050 ;
        RECT 673.950 185.550 697.050 186.450 ;
        RECT 673.950 184.950 676.050 185.550 ;
        RECT 694.950 184.950 697.050 185.550 ;
        RECT 701.700 186.300 702.900 188.400 ;
        RECT 704.100 189.300 705.900 194.400 ;
        RECT 707.100 190.200 708.900 195.000 ;
        RECT 710.100 189.300 711.900 194.400 ;
        RECT 704.100 187.950 711.900 189.300 ;
        RECT 701.700 185.400 705.300 186.300 ;
        RECT 730.500 186.000 732.300 194.400 ;
        RECT 677.250 181.050 679.050 182.850 ;
        RECT 701.100 181.050 702.900 182.850 ;
        RECT 704.100 181.050 705.300 185.400 ;
        RECT 729.000 184.800 732.300 186.000 ;
        RECT 737.100 185.400 738.900 195.000 ;
        RECT 754.500 186.000 756.300 194.400 ;
        RECT 753.000 184.800 756.300 186.000 ;
        RECT 761.100 185.400 762.900 195.000 ;
        RECT 776.700 191.400 778.500 195.000 ;
        RECT 779.700 189.600 781.500 194.400 ;
        RECT 776.400 188.400 781.500 189.600 ;
        RECT 784.200 188.400 786.000 195.000 ;
        RECT 715.950 183.450 718.050 184.050 ;
        RECT 724.950 183.450 727.050 184.050 ;
        RECT 707.100 181.050 708.900 182.850 ;
        RECT 715.950 182.550 727.050 183.450 ;
        RECT 715.950 181.950 718.050 182.550 ;
        RECT 724.950 181.950 727.050 182.550 ;
        RECT 729.000 181.050 729.900 184.800 ;
        RECT 747.000 183.450 751.050 184.050 ;
        RECT 731.100 181.050 732.900 182.850 ;
        RECT 737.100 181.050 738.900 182.850 ;
        RECT 746.550 181.950 751.050 183.450 ;
        RECT 615.900 178.200 618.300 179.100 ;
        RECT 616.800 178.050 618.300 178.200 ;
        RECT 622.800 178.950 624.900 181.050 ;
        RECT 637.950 178.950 640.050 181.050 ;
        RECT 640.950 178.950 643.050 181.050 ;
        RECT 643.950 178.950 646.050 181.050 ;
        RECT 646.950 178.950 649.050 181.050 ;
        RECT 668.400 178.950 670.500 181.050 ;
        RECT 673.950 178.950 676.050 181.050 ;
        RECT 676.950 178.950 679.050 181.050 ;
        RECT 683.100 178.950 685.200 181.050 ;
        RECT 700.950 178.950 703.050 181.050 ;
        RECT 703.950 178.950 706.050 181.050 ;
        RECT 706.950 178.950 709.050 181.050 ;
        RECT 709.950 178.950 712.050 181.050 ;
        RECT 727.950 178.950 730.050 181.050 ;
        RECT 730.950 178.950 733.050 181.050 ;
        RECT 733.950 178.950 736.050 181.050 ;
        RECT 736.950 178.950 739.050 181.050 ;
        RECT 612.000 175.500 615.900 177.300 ;
        RECT 613.800 175.200 615.900 175.500 ;
        RECT 616.800 175.950 618.900 178.050 ;
        RECT 622.800 177.150 624.600 178.950 ;
        RECT 641.250 177.150 643.050 178.950 ;
        RECT 616.800 174.000 617.700 175.950 ;
        RECT 610.500 171.600 612.600 173.700 ;
        RECT 616.200 172.950 617.700 174.000 ;
        RECT 616.200 171.600 617.400 172.950 ;
        RECT 521.100 159.000 522.900 165.000 ;
        RECT 524.100 159.600 525.900 165.600 ;
        RECT 527.100 159.000 528.900 165.600 ;
        RECT 545.100 159.000 546.900 165.600 ;
        RECT 548.100 159.600 549.900 165.600 ;
        RECT 563.100 159.000 564.900 171.600 ;
        RECT 566.400 170.400 570.000 171.600 ;
        RECT 568.200 159.600 570.000 170.400 ;
        RECT 584.100 170.700 591.900 171.600 ;
        RECT 584.100 159.600 585.900 170.700 ;
        RECT 587.100 159.000 588.900 169.800 ;
        RECT 590.100 159.600 591.900 170.700 ;
        RECT 593.100 159.600 594.900 171.600 ;
        RECT 608.100 170.700 612.600 171.600 ;
        RECT 608.100 159.600 609.900 170.700 ;
        RECT 611.100 159.000 612.900 169.500 ;
        RECT 615.600 159.600 617.400 171.600 ;
        RECT 620.100 171.600 622.200 172.500 ;
        RECT 647.700 171.600 648.600 178.950 ;
        RECT 620.100 170.400 624.900 171.600 ;
        RECT 620.100 159.000 621.900 169.500 ;
        RECT 623.100 159.600 624.900 170.400 ;
        RECT 638.100 170.700 645.900 171.600 ;
        RECT 638.100 159.600 639.900 170.700 ;
        RECT 641.100 159.000 642.900 169.800 ;
        RECT 644.100 159.600 645.900 170.700 ;
        RECT 647.100 159.600 648.900 171.600 ;
        RECT 665.100 160.500 666.900 169.800 ;
        RECT 668.700 169.200 669.900 178.950 ;
        RECT 673.950 177.150 675.750 178.950 ;
        RECT 683.100 177.150 684.900 178.950 ;
        RECT 688.950 174.450 691.050 175.050 ;
        RECT 700.950 174.450 703.050 175.050 ;
        RECT 688.950 173.550 703.050 174.450 ;
        RECT 688.950 172.950 691.050 173.550 ;
        RECT 700.950 172.950 703.050 173.550 ;
        RECT 704.100 171.600 705.300 178.950 ;
        RECT 710.100 177.150 711.900 178.950 ;
        RECT 668.100 161.400 669.900 169.200 ;
        RECT 671.100 169.200 678.900 170.100 ;
        RECT 671.100 160.500 672.900 169.200 ;
        RECT 665.100 159.600 672.900 160.500 ;
        RECT 674.100 160.500 675.900 168.300 ;
        RECT 677.100 161.400 678.900 169.200 ;
        RECT 680.100 169.500 687.900 170.400 ;
        RECT 704.100 170.100 706.500 171.600 ;
        RECT 680.100 160.500 681.900 169.500 ;
        RECT 674.100 159.600 681.900 160.500 ;
        RECT 683.100 159.000 684.900 168.600 ;
        RECT 686.100 159.600 687.900 169.500 ;
        RECT 702.000 167.100 703.800 168.900 ;
        RECT 701.700 159.000 703.500 165.600 ;
        RECT 704.700 159.600 706.500 170.100 ;
        RECT 709.800 159.000 711.600 171.600 ;
        RECT 729.000 166.800 729.900 178.950 ;
        RECT 734.100 177.150 735.900 178.950 ;
        RECT 746.550 178.050 747.450 181.950 ;
        RECT 753.000 181.050 753.900 184.800 ;
        RECT 755.100 181.050 756.900 182.850 ;
        RECT 761.100 181.050 762.900 182.850 ;
        RECT 776.400 181.050 777.300 188.400 ;
        RECT 802.500 186.000 804.300 194.400 ;
        RECT 801.000 184.800 804.300 186.000 ;
        RECT 809.100 185.400 810.900 195.000 ;
        RECT 824.700 187.200 826.500 194.400 ;
        RECT 829.800 188.400 831.600 195.000 ;
        RECT 845.700 187.200 847.500 194.400 ;
        RECT 850.800 188.400 852.600 195.000 ;
        RECT 866.100 188.400 867.900 194.400 ;
        RECT 869.400 189.300 871.200 195.000 ;
        RECT 873.900 189.000 875.700 194.400 ;
        RECT 878.100 189.300 879.900 195.000 ;
        RECT 866.100 187.500 870.600 188.400 ;
        RECT 824.700 186.300 828.900 187.200 ;
        RECT 778.950 181.050 780.750 182.850 ;
        RECT 785.100 181.050 786.900 182.850 ;
        RECT 801.000 181.050 801.900 184.800 ;
        RECT 819.000 183.450 823.050 184.050 ;
        RECT 803.100 181.050 804.900 182.850 ;
        RECT 809.100 181.050 810.900 182.850 ;
        RECT 818.550 181.950 823.050 183.450 ;
        RECT 751.950 178.950 754.050 181.050 ;
        RECT 754.950 178.950 757.050 181.050 ;
        RECT 757.950 178.950 760.050 181.050 ;
        RECT 760.950 178.950 763.050 181.050 ;
        RECT 775.950 178.950 778.050 181.050 ;
        RECT 778.950 178.950 781.050 181.050 ;
        RECT 781.950 178.950 784.050 181.050 ;
        RECT 784.950 178.950 787.050 181.050 ;
        RECT 799.950 178.950 802.050 181.050 ;
        RECT 802.950 178.950 805.050 181.050 ;
        RECT 805.950 178.950 808.050 181.050 ;
        RECT 808.950 178.950 811.050 181.050 ;
        RECT 746.550 176.550 751.050 178.050 ;
        RECT 747.000 175.950 751.050 176.550 ;
        RECT 753.000 166.800 753.900 178.950 ;
        RECT 758.100 177.150 759.900 178.950 ;
        RECT 757.950 174.450 760.050 175.050 ;
        RECT 766.950 174.450 769.050 175.050 ;
        RECT 757.950 173.550 769.050 174.450 ;
        RECT 757.950 172.950 760.050 173.550 ;
        RECT 766.950 172.950 769.050 173.550 ;
        RECT 776.400 171.600 777.300 178.950 ;
        RECT 781.950 177.150 783.750 178.950 ;
        RECT 729.000 165.900 735.600 166.800 ;
        RECT 729.000 165.600 729.900 165.900 ;
        RECT 728.100 159.600 729.900 165.600 ;
        RECT 734.100 165.600 735.600 165.900 ;
        RECT 753.000 165.900 759.600 166.800 ;
        RECT 753.000 165.600 753.900 165.900 ;
        RECT 731.100 159.000 732.900 165.000 ;
        RECT 734.100 159.600 735.900 165.600 ;
        RECT 737.100 159.000 738.900 165.600 ;
        RECT 752.100 159.600 753.900 165.600 ;
        RECT 758.100 165.600 759.600 165.900 ;
        RECT 755.100 159.000 756.900 165.000 ;
        RECT 758.100 159.600 759.900 165.600 ;
        RECT 761.100 159.000 762.900 165.600 ;
        RECT 776.100 159.600 777.900 171.600 ;
        RECT 779.100 170.700 786.900 171.600 ;
        RECT 779.100 159.600 780.900 170.700 ;
        RECT 782.100 159.000 783.900 169.800 ;
        RECT 785.100 159.600 786.900 170.700 ;
        RECT 801.000 166.800 801.900 178.950 ;
        RECT 806.100 177.150 807.900 178.950 ;
        RECT 818.550 178.050 819.450 181.950 ;
        RECT 824.100 181.050 825.900 182.850 ;
        RECT 827.700 181.050 828.900 186.300 ;
        RECT 829.950 186.450 832.050 187.050 ;
        RECT 838.950 186.450 841.050 187.050 ;
        RECT 829.950 185.550 841.050 186.450 ;
        RECT 845.700 186.300 849.900 187.200 ;
        RECT 829.950 184.950 832.050 185.550 ;
        RECT 838.950 184.950 841.050 185.550 ;
        RECT 832.950 183.450 837.000 184.050 ;
        RECT 829.950 181.050 831.750 182.850 ;
        RECT 832.950 181.950 837.450 183.450 ;
        RECT 823.950 178.950 826.050 181.050 ;
        RECT 826.950 178.950 829.050 181.050 ;
        RECT 829.950 178.950 832.050 181.050 ;
        RECT 818.550 176.550 823.050 178.050 ;
        RECT 819.000 175.950 823.050 176.550 ;
        RECT 802.950 174.450 805.050 175.050 ;
        RECT 814.950 174.450 817.050 175.050 ;
        RECT 823.950 174.450 826.050 175.050 ;
        RECT 802.950 173.550 826.050 174.450 ;
        RECT 802.950 172.950 805.050 173.550 ;
        RECT 814.950 172.950 817.050 173.550 ;
        RECT 823.950 172.950 826.050 173.550 ;
        RECT 801.000 165.900 807.600 166.800 ;
        RECT 801.000 165.600 801.900 165.900 ;
        RECT 800.100 159.600 801.900 165.600 ;
        RECT 806.100 165.600 807.600 165.900 ;
        RECT 827.700 165.600 828.900 178.950 ;
        RECT 836.550 177.450 837.450 181.950 ;
        RECT 845.100 181.050 846.900 182.850 ;
        RECT 848.700 181.050 849.900 186.300 ;
        RECT 868.500 185.100 870.600 187.500 ;
        RECT 873.900 186.900 874.800 189.000 ;
        RECT 881.100 188.400 882.900 194.400 ;
        RECT 881.400 187.500 882.900 188.400 ;
        RECT 871.800 184.800 874.800 186.900 ;
        RECT 878.400 186.000 882.900 187.500 ;
        RECT 850.950 181.050 852.750 182.850 ;
        RECT 856.950 181.950 859.050 184.050 ;
        RECT 844.950 178.950 847.050 181.050 ;
        RECT 847.950 178.950 850.050 181.050 ;
        RECT 850.950 178.950 853.050 181.050 ;
        RECT 841.950 177.450 844.050 178.050 ;
        RECT 836.550 176.550 844.050 177.450 ;
        RECT 841.950 175.950 844.050 176.550 ;
        RECT 848.700 165.600 849.900 178.950 ;
        RECT 857.550 178.050 858.450 181.950 ;
        RECT 866.100 178.950 868.200 181.050 ;
        RECT 870.900 180.900 873.000 183.000 ;
        RECT 871.200 179.100 873.000 180.900 ;
        RECT 853.950 176.550 858.450 178.050 ;
        RECT 866.400 177.150 868.200 178.950 ;
        RECT 873.900 178.050 874.800 184.800 ;
        RECT 875.700 183.900 877.500 185.700 ;
        RECT 878.400 185.400 880.500 186.000 ;
        RECT 876.000 183.000 878.100 183.900 ;
        RECT 876.000 181.800 882.600 183.000 ;
        RECT 880.800 181.200 882.600 181.800 ;
        RECT 876.000 178.800 878.100 180.900 ;
        RECT 880.800 178.950 882.900 181.200 ;
        RECT 871.800 176.700 874.800 178.050 ;
        RECT 876.300 177.000 878.100 178.800 ;
        RECT 853.950 175.950 858.000 176.550 ;
        RECT 871.800 175.950 873.900 176.700 ;
        RECT 869.100 171.600 871.200 172.500 ;
        RECT 866.100 170.400 871.200 171.600 ;
        RECT 872.100 171.600 873.300 175.950 ;
        RECT 874.800 173.700 876.600 175.500 ;
        RECT 874.800 172.800 880.200 173.700 ;
        RECT 878.100 171.900 880.200 172.800 ;
        RECT 872.100 170.700 875.400 171.600 ;
        RECT 878.100 170.700 882.900 171.900 ;
        RECT 803.100 159.000 804.900 165.000 ;
        RECT 806.100 159.600 807.900 165.600 ;
        RECT 809.100 159.000 810.900 165.600 ;
        RECT 824.100 159.000 825.900 165.600 ;
        RECT 827.100 159.600 828.900 165.600 ;
        RECT 830.100 159.000 831.900 165.600 ;
        RECT 845.100 159.000 846.900 165.600 ;
        RECT 848.100 159.600 849.900 165.600 ;
        RECT 851.100 159.000 852.900 165.600 ;
        RECT 866.100 159.600 867.900 170.400 ;
        RECT 869.100 159.000 871.200 169.500 ;
        RECT 873.600 159.600 875.400 170.700 ;
        RECT 878.100 159.000 879.900 169.500 ;
        RECT 881.100 159.600 882.900 170.700 ;
        RECT 14.100 144.600 15.900 155.400 ;
        RECT 17.100 145.500 19.200 156.000 ;
        RECT 14.100 143.400 19.200 144.600 ;
        RECT 21.600 144.300 23.400 155.400 ;
        RECT 26.100 145.500 27.900 156.000 ;
        RECT 29.100 144.300 30.900 155.400 ;
        RECT 47.100 149.400 48.900 156.000 ;
        RECT 50.100 149.400 51.900 155.400 ;
        RECT 65.100 149.400 66.900 156.000 ;
        RECT 68.100 149.400 69.900 155.400 ;
        RECT 71.100 149.400 72.900 156.000 ;
        RECT 86.100 149.400 87.900 156.000 ;
        RECT 89.100 149.400 90.900 155.400 ;
        RECT 17.100 142.500 19.200 143.400 ;
        RECT 20.100 143.400 23.400 144.300 ;
        RECT 20.100 139.050 21.300 143.400 ;
        RECT 26.100 143.100 30.900 144.300 ;
        RECT 26.100 142.200 28.200 143.100 ;
        RECT 22.800 141.300 28.200 142.200 ;
        RECT 22.800 139.500 24.600 141.300 ;
        RECT 19.800 138.300 21.900 139.050 ;
        RECT 14.400 136.050 16.200 137.850 ;
        RECT 19.800 136.950 22.800 138.300 ;
        RECT 14.100 133.950 16.200 136.050 ;
        RECT 19.200 134.100 21.000 135.900 ;
        RECT 18.900 132.000 21.000 134.100 ;
        RECT 21.900 130.200 22.800 136.950 ;
        RECT 24.300 136.200 26.100 138.000 ;
        RECT 24.000 134.100 26.100 136.200 ;
        RECT 47.100 136.050 48.900 137.850 ;
        RECT 50.100 136.050 51.300 149.400 ;
        RECT 52.950 141.450 55.050 142.050 ;
        RECT 64.950 141.450 67.050 142.050 ;
        RECT 52.950 140.550 67.050 141.450 ;
        RECT 52.950 139.950 55.050 140.550 ;
        RECT 64.950 139.950 67.050 140.550 ;
        RECT 68.700 136.050 69.900 149.400 ;
        RECT 86.100 136.050 87.900 137.850 ;
        RECT 89.100 136.050 90.300 149.400 ;
        RECT 104.400 143.400 106.200 156.000 ;
        RECT 109.500 144.900 111.300 155.400 ;
        RECT 112.500 149.400 114.300 156.000 ;
        RECT 112.200 146.100 114.000 147.900 ;
        RECT 109.500 143.400 111.900 144.900 ;
        RECT 129.000 144.600 130.800 155.400 ;
        RECT 129.000 143.400 132.600 144.600 ;
        RECT 134.100 143.400 135.900 156.000 ;
        RECT 152.100 149.400 153.900 155.400 ;
        RECT 155.100 149.400 156.900 156.000 ;
        RECT 170.700 149.400 172.500 156.000 ;
        RECT 104.100 136.050 105.900 137.850 ;
        RECT 110.700 136.050 111.900 143.400 ;
        RECT 128.100 136.050 129.900 137.850 ;
        RECT 131.700 136.050 132.600 143.400 ;
        RECT 133.950 136.050 135.750 137.850 ;
        RECT 152.700 136.050 153.900 149.400 ;
        RECT 171.000 146.100 172.800 147.900 ;
        RECT 173.700 144.900 175.500 155.400 ;
        RECT 173.100 143.400 175.500 144.900 ;
        RECT 178.800 143.400 180.600 156.000 ;
        RECT 194.100 144.600 195.900 155.400 ;
        RECT 197.100 145.500 198.900 156.000 ;
        RECT 200.100 154.500 207.900 155.400 ;
        RECT 200.100 144.600 201.900 154.500 ;
        RECT 194.100 143.700 201.900 144.600 ;
        RECT 155.100 136.050 156.900 137.850 ;
        RECT 173.100 136.050 174.300 143.400 ;
        RECT 203.100 142.500 204.900 153.600 ;
        RECT 206.100 143.400 207.900 154.500 ;
        RECT 221.100 149.400 222.900 155.400 ;
        RECT 224.100 149.400 225.900 156.000 ;
        RECT 187.950 141.450 190.050 142.050 ;
        RECT 193.950 141.450 196.050 142.200 ;
        RECT 187.950 140.550 196.050 141.450 ;
        RECT 187.950 139.950 190.050 140.550 ;
        RECT 193.950 140.100 196.050 140.550 ;
        RECT 200.100 141.600 204.900 142.500 ;
        RECT 179.100 136.050 180.900 137.850 ;
        RECT 197.250 136.050 199.050 137.850 ;
        RECT 200.100 136.050 201.000 141.600 ;
        RECT 208.950 138.450 211.050 139.050 ;
        RECT 214.950 138.450 217.050 139.050 ;
        RECT 203.100 136.050 204.900 137.850 ;
        RECT 208.950 137.550 217.050 138.450 ;
        RECT 208.950 136.950 211.050 137.550 ;
        RECT 214.950 136.950 217.050 137.550 ;
        RECT 221.700 136.050 222.900 149.400 ;
        RECT 239.100 143.400 240.900 155.400 ;
        RECT 242.100 144.300 243.900 155.400 ;
        RECT 245.100 145.200 246.900 156.000 ;
        RECT 248.100 144.300 249.900 155.400 ;
        RECT 266.100 149.400 267.900 156.000 ;
        RECT 269.100 149.400 270.900 155.400 ;
        RECT 272.100 149.400 273.900 156.000 ;
        RECT 287.100 149.400 288.900 155.400 ;
        RECT 290.100 150.000 291.900 156.000 ;
        RECT 242.100 143.400 249.900 144.300 ;
        RECT 224.100 136.050 225.900 137.850 ;
        RECT 239.400 136.050 240.300 143.400 ;
        RECT 244.950 136.050 246.750 137.850 ;
        RECT 269.100 136.050 270.300 149.400 ;
        RECT 288.000 149.100 288.900 149.400 ;
        RECT 293.100 149.400 294.900 155.400 ;
        RECT 296.100 149.400 297.900 156.000 ;
        RECT 293.100 149.100 294.600 149.400 ;
        RECT 288.000 148.200 294.600 149.100 ;
        RECT 274.950 144.450 277.050 145.050 ;
        RECT 283.950 144.450 286.050 145.050 ;
        RECT 274.950 143.550 286.050 144.450 ;
        RECT 274.950 142.950 277.050 143.550 ;
        RECT 283.950 142.950 286.050 143.550 ;
        RECT 288.000 136.050 288.900 148.200 ;
        RECT 314.100 144.300 315.900 155.400 ;
        RECT 317.100 145.200 318.900 156.000 ;
        RECT 320.100 144.300 321.900 155.400 ;
        RECT 314.100 143.400 321.900 144.300 ;
        RECT 323.100 143.400 324.900 155.400 ;
        RECT 338.100 149.400 339.900 156.000 ;
        RECT 341.100 149.400 342.900 155.400 ;
        RECT 344.100 150.000 345.900 156.000 ;
        RECT 341.400 149.100 342.900 149.400 ;
        RECT 347.100 149.400 348.900 155.400 ;
        RECT 347.100 149.100 348.000 149.400 ;
        RECT 341.400 148.200 348.000 149.100 ;
        RECT 331.950 144.450 334.050 145.050 ;
        RECT 340.950 144.450 343.050 145.050 ;
        RECT 331.950 143.550 343.050 144.450 ;
        RECT 293.100 136.050 294.900 137.850 ;
        RECT 317.250 136.050 319.050 137.850 ;
        RECT 323.700 136.050 324.600 143.400 ;
        RECT 331.950 142.950 334.050 143.550 ;
        RECT 340.950 142.950 343.050 143.550 ;
        RECT 341.100 136.050 342.900 137.850 ;
        RECT 347.100 136.050 348.000 148.200 ;
        RECT 362.400 143.400 364.200 156.000 ;
        RECT 367.500 144.900 369.300 155.400 ;
        RECT 370.500 149.400 372.300 156.000 ;
        RECT 386.100 149.400 387.900 155.400 ;
        RECT 389.100 149.400 390.900 156.000 ;
        RECT 404.100 149.400 405.900 155.400 ;
        RECT 407.100 150.000 408.900 156.000 ;
        RECT 370.200 146.100 372.000 147.900 ;
        RECT 367.500 143.400 369.900 144.900 ;
        RECT 352.950 138.450 355.050 139.050 ;
        RECT 358.950 138.450 361.050 139.050 ;
        RECT 352.950 137.550 361.050 138.450 ;
        RECT 352.950 136.950 355.050 137.550 ;
        RECT 358.950 136.950 361.050 137.550 ;
        RECT 362.100 136.050 363.900 137.850 ;
        RECT 368.700 136.050 369.900 143.400 ;
        RECT 386.700 136.050 387.900 149.400 ;
        RECT 405.000 149.100 405.900 149.400 ;
        RECT 410.100 149.400 411.900 155.400 ;
        RECT 413.100 149.400 414.900 156.000 ;
        RECT 428.100 149.400 429.900 156.000 ;
        RECT 431.100 149.400 432.900 155.400 ;
        RECT 434.100 149.400 435.900 156.000 ;
        RECT 449.100 149.400 450.900 156.000 ;
        RECT 452.100 149.400 453.900 155.400 ;
        RECT 455.100 149.400 456.900 156.000 ;
        RECT 410.100 149.100 411.600 149.400 ;
        RECT 405.000 148.200 411.600 149.100 ;
        RECT 389.100 136.050 390.900 137.850 ;
        RECT 405.000 136.050 405.900 148.200 ;
        RECT 410.100 136.050 411.900 137.850 ;
        RECT 431.100 136.050 432.300 149.400 ;
        RECT 452.100 136.050 453.300 149.400 ;
        RECT 473.100 144.600 474.900 155.400 ;
        RECT 476.100 145.500 477.900 156.000 ;
        RECT 479.100 154.500 486.900 155.400 ;
        RECT 479.100 144.600 480.900 154.500 ;
        RECT 473.100 143.700 480.900 144.600 ;
        RECT 482.100 142.500 483.900 153.600 ;
        RECT 485.100 143.400 486.900 154.500 ;
        RECT 503.100 149.400 504.900 156.000 ;
        RECT 506.100 149.400 507.900 155.400 ;
        RECT 524.100 149.400 525.900 155.400 ;
        RECT 527.100 150.000 528.900 156.000 ;
        RECT 479.100 141.600 483.900 142.500 ;
        RECT 476.250 136.050 478.050 137.850 ;
        RECT 479.100 136.050 480.000 141.600 ;
        RECT 482.100 136.050 483.900 137.850 ;
        RECT 503.100 136.050 504.900 137.850 ;
        RECT 506.100 136.050 507.300 149.400 ;
        RECT 525.000 149.100 525.900 149.400 ;
        RECT 530.100 149.400 531.900 155.400 ;
        RECT 533.100 149.400 534.900 156.000 ;
        RECT 548.100 149.400 549.900 156.000 ;
        RECT 551.100 149.400 552.900 155.400 ;
        RECT 554.100 149.400 555.900 156.000 ;
        RECT 569.100 149.400 570.900 156.000 ;
        RECT 572.100 149.400 573.900 155.400 ;
        RECT 575.100 149.400 576.900 156.000 ;
        RECT 593.700 149.400 595.500 156.000 ;
        RECT 530.100 149.100 531.600 149.400 ;
        RECT 525.000 148.200 531.600 149.100 ;
        RECT 525.000 136.050 525.900 148.200 ;
        RECT 532.950 141.450 535.050 142.050 ;
        RECT 547.950 141.450 550.050 142.200 ;
        RECT 532.950 140.550 550.050 141.450 ;
        RECT 532.950 139.950 535.050 140.550 ;
        RECT 547.950 140.100 550.050 140.550 ;
        RECT 530.100 136.050 531.900 137.850 ;
        RECT 551.100 136.050 552.300 149.400 ;
        RECT 572.100 136.050 573.300 149.400 ;
        RECT 594.000 146.100 595.800 147.900 ;
        RECT 596.700 144.900 598.500 155.400 ;
        RECT 596.100 143.400 598.500 144.900 ;
        RECT 601.800 143.400 603.600 156.000 ;
        RECT 617.100 144.300 618.900 155.400 ;
        RECT 620.100 145.500 621.900 156.000 ;
        RECT 617.100 143.400 621.600 144.300 ;
        RECT 624.600 143.400 626.400 155.400 ;
        RECT 629.100 145.500 630.900 156.000 ;
        RECT 632.100 144.600 633.900 155.400 ;
        RECT 647.100 149.400 648.900 156.000 ;
        RECT 650.100 149.400 651.900 155.400 ;
        RECT 653.100 149.400 654.900 156.000 ;
        RECT 668.700 149.400 670.500 156.000 ;
        RECT 596.100 136.050 597.300 143.400 ;
        RECT 619.500 141.300 621.600 143.400 ;
        RECT 625.200 142.050 626.400 143.400 ;
        RECT 629.100 143.400 633.900 144.600 ;
        RECT 629.100 142.500 631.200 143.400 ;
        RECT 625.200 141.000 626.700 142.050 ;
        RECT 622.800 139.500 624.900 139.800 ;
        RECT 602.100 136.050 603.900 137.850 ;
        RECT 621.000 137.700 624.900 139.500 ;
        RECT 625.800 139.050 626.700 141.000 ;
        RECT 625.800 136.950 627.900 139.050 ;
        RECT 625.800 136.800 627.300 136.950 ;
        RECT 622.200 136.050 624.000 136.500 ;
        RECT 28.800 133.800 30.900 136.050 ;
        RECT 46.950 133.950 49.050 136.050 ;
        RECT 49.950 133.950 52.050 136.050 ;
        RECT 64.950 133.950 67.050 136.050 ;
        RECT 67.950 133.950 70.050 136.050 ;
        RECT 70.950 133.950 73.050 136.050 ;
        RECT 85.950 133.950 88.050 136.050 ;
        RECT 88.950 133.950 91.050 136.050 ;
        RECT 103.950 133.950 106.050 136.050 ;
        RECT 106.950 133.950 109.050 136.050 ;
        RECT 109.950 133.950 112.050 136.050 ;
        RECT 112.950 133.950 115.050 136.050 ;
        RECT 127.950 133.950 130.050 136.050 ;
        RECT 130.950 133.950 133.050 136.050 ;
        RECT 133.950 133.950 136.050 136.050 ;
        RECT 151.950 133.950 154.050 136.050 ;
        RECT 154.950 133.950 157.050 136.050 ;
        RECT 169.950 133.950 172.050 136.050 ;
        RECT 172.950 133.950 175.050 136.050 ;
        RECT 175.950 133.950 178.050 136.050 ;
        RECT 178.950 133.950 181.050 136.050 ;
        RECT 193.950 133.950 196.050 136.050 ;
        RECT 196.950 133.950 199.050 136.050 ;
        RECT 199.950 133.950 202.050 136.050 ;
        RECT 202.950 133.950 205.050 136.050 ;
        RECT 205.950 133.950 208.050 136.050 ;
        RECT 220.950 133.950 223.050 136.050 ;
        RECT 223.950 133.950 226.050 136.050 ;
        RECT 238.950 133.950 241.050 136.050 ;
        RECT 241.950 133.950 244.050 136.050 ;
        RECT 244.950 133.950 247.050 136.050 ;
        RECT 247.950 133.950 250.050 136.050 ;
        RECT 265.950 133.950 268.050 136.050 ;
        RECT 268.950 133.950 271.050 136.050 ;
        RECT 271.950 133.950 274.050 136.050 ;
        RECT 286.950 133.950 289.050 136.050 ;
        RECT 289.950 133.950 292.050 136.050 ;
        RECT 292.950 133.950 295.050 136.050 ;
        RECT 295.950 133.950 298.050 136.050 ;
        RECT 313.950 133.950 316.050 136.050 ;
        RECT 316.950 133.950 319.050 136.050 ;
        RECT 319.950 133.950 322.050 136.050 ;
        RECT 322.950 133.950 325.050 136.050 ;
        RECT 337.950 133.950 340.050 136.050 ;
        RECT 340.950 133.950 343.050 136.050 ;
        RECT 343.950 133.950 346.050 136.050 ;
        RECT 346.950 133.950 349.050 136.050 ;
        RECT 361.950 133.950 364.050 136.050 ;
        RECT 364.950 133.950 367.050 136.050 ;
        RECT 367.950 133.950 370.050 136.050 ;
        RECT 370.950 133.950 373.050 136.050 ;
        RECT 385.950 133.950 388.050 136.050 ;
        RECT 388.950 133.950 391.050 136.050 ;
        RECT 403.950 133.950 406.050 136.050 ;
        RECT 406.950 133.950 409.050 136.050 ;
        RECT 409.950 133.950 412.050 136.050 ;
        RECT 412.950 133.950 415.050 136.050 ;
        RECT 427.950 133.950 430.050 136.050 ;
        RECT 430.950 133.950 433.050 136.050 ;
        RECT 433.950 133.950 436.050 136.050 ;
        RECT 448.950 133.950 451.050 136.050 ;
        RECT 451.950 133.950 454.050 136.050 ;
        RECT 454.950 133.950 457.050 136.050 ;
        RECT 472.950 133.950 475.050 136.050 ;
        RECT 475.950 133.950 478.050 136.050 ;
        RECT 478.950 133.950 481.050 136.050 ;
        RECT 481.950 133.950 484.050 136.050 ;
        RECT 484.950 133.950 487.050 136.050 ;
        RECT 502.950 133.950 505.050 136.050 ;
        RECT 505.950 133.950 508.050 136.050 ;
        RECT 523.950 133.950 526.050 136.050 ;
        RECT 526.950 133.950 529.050 136.050 ;
        RECT 529.950 133.950 532.050 136.050 ;
        RECT 532.950 133.950 535.050 136.050 ;
        RECT 547.950 133.950 550.050 136.050 ;
        RECT 550.950 133.950 553.050 136.050 ;
        RECT 553.950 133.950 556.050 136.050 ;
        RECT 568.950 133.950 571.050 136.050 ;
        RECT 571.950 133.950 574.050 136.050 ;
        RECT 574.950 133.950 577.050 136.050 ;
        RECT 592.950 133.950 595.050 136.050 ;
        RECT 595.950 133.950 598.050 136.050 ;
        RECT 598.950 133.950 601.050 136.050 ;
        RECT 601.950 133.950 604.050 136.050 ;
        RECT 617.100 134.700 624.000 136.050 ;
        RECT 624.900 135.900 627.300 136.800 ;
        RECT 631.800 136.050 633.600 137.850 ;
        RECT 650.100 136.050 651.300 149.400 ;
        RECT 669.000 146.100 670.800 147.900 ;
        RECT 671.700 144.900 673.500 155.400 ;
        RECT 671.100 143.400 673.500 144.900 ;
        RECT 676.800 143.400 678.600 156.000 ;
        RECT 695.100 143.400 696.900 155.400 ;
        RECT 698.100 144.300 699.900 155.400 ;
        RECT 701.100 145.200 702.900 156.000 ;
        RECT 704.100 144.300 705.900 155.400 ;
        RECT 719.100 149.400 720.900 155.400 ;
        RECT 722.100 150.000 723.900 156.000 ;
        RECT 698.100 143.400 705.900 144.300 ;
        RECT 720.000 149.100 720.900 149.400 ;
        RECT 725.100 149.400 726.900 155.400 ;
        RECT 728.100 149.400 729.900 156.000 ;
        RECT 743.100 149.400 744.900 156.000 ;
        RECT 746.100 149.400 747.900 155.400 ;
        RECT 725.100 149.100 726.600 149.400 ;
        RECT 720.000 148.200 726.600 149.100 ;
        RECT 671.100 136.050 672.300 143.400 ;
        RECT 677.100 136.050 678.900 137.850 ;
        RECT 695.400 136.050 696.300 143.400 ;
        RECT 697.950 141.450 700.050 142.050 ;
        RECT 712.950 141.450 715.050 142.050 ;
        RECT 697.950 140.550 715.050 141.450 ;
        RECT 697.950 139.950 700.050 140.550 ;
        RECT 712.950 139.950 715.050 140.550 ;
        RECT 700.950 136.050 702.750 137.850 ;
        RECT 720.000 136.050 720.900 148.200 ;
        RECT 725.100 136.050 726.900 137.850 ;
        RECT 617.100 133.950 619.200 134.700 ;
        RECT 28.800 133.200 30.600 133.800 ;
        RECT 24.000 132.000 30.600 133.200 ;
        RECT 24.000 131.100 26.100 132.000 ;
        RECT 16.500 127.500 18.600 129.900 ;
        RECT 19.800 128.100 22.800 130.200 ;
        RECT 23.700 129.300 25.500 131.100 ;
        RECT 14.100 126.600 18.600 127.500 ;
        RECT 14.100 120.600 15.900 126.600 ;
        RECT 21.900 126.000 22.800 128.100 ;
        RECT 26.400 129.000 28.500 129.600 ;
        RECT 26.400 127.500 30.900 129.000 ;
        RECT 29.400 126.600 30.900 127.500 ;
        RECT 17.400 120.000 19.200 125.700 ;
        RECT 21.900 120.600 23.700 126.000 ;
        RECT 26.100 120.000 27.900 125.700 ;
        RECT 29.100 120.600 30.900 126.600 ;
        RECT 50.100 123.600 51.300 133.950 ;
        RECT 65.100 132.150 66.900 133.950 ;
        RECT 68.700 128.700 69.900 133.950 ;
        RECT 70.950 132.150 72.750 133.950 ;
        RECT 65.700 127.800 69.900 128.700 ;
        RECT 47.100 120.000 48.900 123.600 ;
        RECT 50.100 120.600 51.900 123.600 ;
        RECT 65.700 120.600 67.500 127.800 ;
        RECT 70.800 120.000 72.600 126.600 ;
        RECT 89.100 123.600 90.300 133.950 ;
        RECT 107.100 132.150 108.900 133.950 ;
        RECT 110.700 129.600 111.900 133.950 ;
        RECT 113.100 132.150 114.900 133.950 ;
        RECT 110.700 128.700 114.300 129.600 ;
        RECT 104.100 125.700 111.900 127.050 ;
        RECT 86.100 120.000 87.900 123.600 ;
        RECT 89.100 120.600 90.900 123.600 ;
        RECT 104.100 120.600 105.900 125.700 ;
        RECT 107.100 120.000 108.900 124.800 ;
        RECT 110.100 120.600 111.900 125.700 ;
        RECT 113.100 126.600 114.300 128.700 ;
        RECT 121.950 129.450 124.050 130.050 ;
        RECT 127.950 129.450 130.050 130.050 ;
        RECT 121.950 128.550 130.050 129.450 ;
        RECT 121.950 127.950 124.050 128.550 ;
        RECT 127.950 127.950 130.050 128.550 ;
        RECT 113.100 120.600 114.900 126.600 ;
        RECT 131.700 123.600 132.600 133.950 ;
        RECT 152.700 123.600 153.900 133.950 ;
        RECT 170.100 132.150 171.900 133.950 ;
        RECT 173.100 129.600 174.300 133.950 ;
        RECT 176.100 132.150 177.900 133.950 ;
        RECT 194.250 132.150 196.050 133.950 ;
        RECT 170.700 128.700 174.300 129.600 ;
        RECT 170.700 126.600 171.900 128.700 ;
        RECT 128.100 120.000 129.900 123.600 ;
        RECT 131.100 120.600 132.900 123.600 ;
        RECT 134.100 120.000 135.900 123.600 ;
        RECT 152.100 120.600 153.900 123.600 ;
        RECT 155.100 120.000 156.900 123.600 ;
        RECT 170.100 120.600 171.900 126.600 ;
        RECT 173.100 125.700 180.900 127.050 ;
        RECT 200.100 126.600 201.300 133.950 ;
        RECT 206.100 132.150 207.900 133.950 ;
        RECT 202.950 129.450 205.050 130.050 ;
        RECT 211.950 129.450 214.050 130.050 ;
        RECT 202.950 128.550 214.050 129.450 ;
        RECT 202.950 127.950 205.050 128.550 ;
        RECT 211.950 127.950 214.050 128.550 ;
        RECT 173.100 120.600 174.900 125.700 ;
        RECT 176.100 120.000 177.900 124.800 ;
        RECT 179.100 120.600 180.900 125.700 ;
        RECT 194.700 120.000 196.500 126.600 ;
        RECT 199.200 120.600 201.000 126.600 ;
        RECT 203.700 120.000 205.500 126.600 ;
        RECT 221.700 123.600 222.900 133.950 ;
        RECT 239.400 126.600 240.300 133.950 ;
        RECT 241.950 132.150 243.750 133.950 ;
        RECT 248.100 132.150 249.900 133.950 ;
        RECT 266.250 132.150 268.050 133.950 ;
        RECT 269.100 128.700 270.300 133.950 ;
        RECT 272.100 132.150 273.900 133.950 ;
        RECT 277.950 132.450 280.050 133.050 ;
        RECT 283.950 132.450 286.050 133.050 ;
        RECT 277.950 131.550 286.050 132.450 ;
        RECT 277.950 130.950 280.050 131.550 ;
        RECT 283.950 130.950 286.050 131.550 ;
        RECT 288.000 130.200 288.900 133.950 ;
        RECT 290.100 132.150 291.900 133.950 ;
        RECT 296.100 132.150 297.900 133.950 ;
        RECT 314.100 132.150 315.900 133.950 ;
        RECT 320.250 132.150 322.050 133.950 ;
        RECT 288.000 129.000 291.300 130.200 ;
        RECT 269.100 127.800 273.300 128.700 ;
        RECT 239.400 125.400 244.500 126.600 ;
        RECT 221.100 120.600 222.900 123.600 ;
        RECT 224.100 120.000 225.900 123.600 ;
        RECT 239.700 120.000 241.500 123.600 ;
        RECT 242.700 120.600 244.500 125.400 ;
        RECT 247.200 120.000 249.000 126.600 ;
        RECT 266.400 120.000 268.200 126.600 ;
        RECT 271.500 120.600 273.300 127.800 ;
        RECT 289.500 120.600 291.300 129.000 ;
        RECT 296.100 120.000 297.900 129.600 ;
        RECT 323.700 126.600 324.600 133.950 ;
        RECT 338.100 132.150 339.900 133.950 ;
        RECT 344.100 132.150 345.900 133.950 ;
        RECT 347.100 130.200 348.000 133.950 ;
        RECT 365.100 132.150 366.900 133.950 ;
        RECT 315.000 120.000 316.800 126.600 ;
        RECT 319.500 125.400 324.600 126.600 ;
        RECT 319.500 120.600 321.300 125.400 ;
        RECT 322.500 120.000 324.300 123.600 ;
        RECT 338.100 120.000 339.900 129.600 ;
        RECT 344.700 129.000 348.000 130.200 ;
        RECT 368.700 129.600 369.900 133.950 ;
        RECT 371.100 132.150 372.900 133.950 ;
        RECT 344.700 120.600 346.500 129.000 ;
        RECT 368.700 128.700 372.300 129.600 ;
        RECT 362.100 125.700 369.900 127.050 ;
        RECT 362.100 120.600 363.900 125.700 ;
        RECT 365.100 120.000 366.900 124.800 ;
        RECT 368.100 120.600 369.900 125.700 ;
        RECT 371.100 126.600 372.300 128.700 ;
        RECT 371.100 120.600 372.900 126.600 ;
        RECT 386.700 123.600 387.900 133.950 ;
        RECT 405.000 130.200 405.900 133.950 ;
        RECT 407.100 132.150 408.900 133.950 ;
        RECT 413.100 132.150 414.900 133.950 ;
        RECT 428.250 132.150 430.050 133.950 ;
        RECT 405.000 129.000 408.300 130.200 ;
        RECT 386.100 120.600 387.900 123.600 ;
        RECT 389.100 120.000 390.900 123.600 ;
        RECT 406.500 120.600 408.300 129.000 ;
        RECT 413.100 120.000 414.900 129.600 ;
        RECT 431.100 128.700 432.300 133.950 ;
        RECT 434.100 132.150 435.900 133.950 ;
        RECT 449.250 132.150 451.050 133.950 ;
        RECT 452.100 128.700 453.300 133.950 ;
        RECT 455.100 132.150 456.900 133.950 ;
        RECT 473.250 132.150 475.050 133.950 ;
        RECT 460.950 129.450 463.050 130.050 ;
        RECT 475.950 129.450 478.050 130.050 ;
        RECT 431.100 127.800 435.300 128.700 ;
        RECT 452.100 127.800 456.300 128.700 ;
        RECT 460.950 128.550 478.050 129.450 ;
        RECT 460.950 127.950 463.050 128.550 ;
        RECT 475.950 127.950 478.050 128.550 ;
        RECT 428.400 120.000 430.200 126.600 ;
        RECT 433.500 120.600 435.300 127.800 ;
        RECT 449.400 120.000 451.200 126.600 ;
        RECT 454.500 120.600 456.300 127.800 ;
        RECT 479.100 126.600 480.300 133.950 ;
        RECT 485.100 132.150 486.900 133.950 ;
        RECT 473.700 120.000 475.500 126.600 ;
        RECT 478.200 120.600 480.000 126.600 ;
        RECT 482.700 120.000 484.500 126.600 ;
        RECT 506.100 123.600 507.300 133.950 ;
        RECT 525.000 130.200 525.900 133.950 ;
        RECT 527.100 132.150 528.900 133.950 ;
        RECT 533.100 132.150 534.900 133.950 ;
        RECT 548.250 132.150 550.050 133.950 ;
        RECT 525.000 129.000 528.300 130.200 ;
        RECT 503.100 120.000 504.900 123.600 ;
        RECT 506.100 120.600 507.900 123.600 ;
        RECT 526.500 120.600 528.300 129.000 ;
        RECT 533.100 120.000 534.900 129.600 ;
        RECT 551.100 128.700 552.300 133.950 ;
        RECT 554.100 132.150 555.900 133.950 ;
        RECT 569.250 132.150 571.050 133.950 ;
        RECT 572.100 128.700 573.300 133.950 ;
        RECT 575.100 132.150 576.900 133.950 ;
        RECT 593.100 132.150 594.900 133.950 ;
        RECT 596.100 129.600 597.300 133.950 ;
        RECT 599.100 132.150 600.900 133.950 ;
        RECT 617.400 132.150 619.200 133.950 ;
        RECT 622.200 131.400 624.000 133.200 ;
        RECT 593.700 128.700 597.300 129.600 ;
        RECT 621.900 129.300 624.000 131.400 ;
        RECT 551.100 127.800 555.300 128.700 ;
        RECT 572.100 127.800 576.300 128.700 ;
        RECT 548.400 120.000 550.200 126.600 ;
        RECT 553.500 120.600 555.300 127.800 ;
        RECT 569.400 120.000 571.200 126.600 ;
        RECT 574.500 120.600 576.300 127.800 ;
        RECT 593.700 126.600 594.900 128.700 ;
        RECT 617.700 128.400 624.000 129.300 ;
        RECT 624.900 130.200 626.100 135.900 ;
        RECT 627.300 133.200 629.100 135.000 ;
        RECT 631.800 133.950 633.900 136.050 ;
        RECT 646.950 133.950 649.050 136.050 ;
        RECT 649.950 133.950 652.050 136.050 ;
        RECT 652.950 133.950 655.050 136.050 ;
        RECT 667.950 133.950 670.050 136.050 ;
        RECT 670.950 133.950 673.050 136.050 ;
        RECT 673.950 133.950 676.050 136.050 ;
        RECT 676.950 133.950 679.050 136.050 ;
        RECT 694.950 133.950 697.050 136.050 ;
        RECT 697.950 133.950 700.050 136.050 ;
        RECT 700.950 133.950 703.050 136.050 ;
        RECT 703.950 133.950 706.050 136.050 ;
        RECT 718.950 133.950 721.050 136.050 ;
        RECT 721.950 133.950 724.050 136.050 ;
        RECT 724.950 133.950 727.050 136.050 ;
        RECT 727.950 133.950 730.050 136.050 ;
        RECT 743.100 133.950 745.200 136.050 ;
        RECT 627.000 131.100 629.100 133.200 ;
        RECT 647.250 132.150 649.050 133.950 ;
        RECT 593.100 120.600 594.900 126.600 ;
        RECT 596.100 125.700 603.900 127.050 ;
        RECT 617.700 126.600 618.900 128.400 ;
        RECT 624.900 128.100 627.900 130.200 ;
        RECT 650.100 128.700 651.300 133.950 ;
        RECT 653.100 132.150 654.900 133.950 ;
        RECT 668.100 132.150 669.900 133.950 ;
        RECT 671.100 129.600 672.300 133.950 ;
        RECT 674.100 132.150 675.900 133.950 ;
        RECT 668.700 128.700 672.300 129.600 ;
        RECT 624.900 126.600 626.100 128.100 ;
        RECT 629.100 127.500 631.200 128.700 ;
        RECT 650.100 127.800 654.300 128.700 ;
        RECT 629.100 126.600 633.900 127.500 ;
        RECT 596.100 120.600 597.900 125.700 ;
        RECT 599.100 120.000 600.900 124.800 ;
        RECT 602.100 120.600 603.900 125.700 ;
        RECT 617.100 120.600 618.900 126.600 ;
        RECT 620.100 120.000 621.900 125.700 ;
        RECT 624.600 120.600 626.400 126.600 ;
        RECT 629.100 120.000 630.900 125.700 ;
        RECT 632.100 120.600 633.900 126.600 ;
        RECT 647.400 120.000 649.200 126.600 ;
        RECT 652.500 120.600 654.300 127.800 ;
        RECT 668.700 126.600 669.900 128.700 ;
        RECT 668.100 120.600 669.900 126.600 ;
        RECT 671.100 125.700 678.900 127.050 ;
        RECT 671.100 120.600 672.900 125.700 ;
        RECT 674.100 120.000 675.900 124.800 ;
        RECT 677.100 120.600 678.900 125.700 ;
        RECT 695.400 126.600 696.300 133.950 ;
        RECT 697.950 132.150 699.750 133.950 ;
        RECT 704.100 132.150 705.900 133.950 ;
        RECT 720.000 130.200 720.900 133.950 ;
        RECT 722.100 132.150 723.900 133.950 ;
        RECT 728.100 132.150 729.900 133.950 ;
        RECT 743.250 132.150 745.050 133.950 ;
        RECT 720.000 129.000 723.300 130.200 ;
        RECT 695.400 125.400 700.500 126.600 ;
        RECT 695.700 120.000 697.500 123.600 ;
        RECT 698.700 120.600 700.500 125.400 ;
        RECT 703.200 120.000 705.000 126.600 ;
        RECT 721.500 120.600 723.300 129.000 ;
        RECT 728.100 120.000 729.900 129.600 ;
        RECT 746.100 129.300 747.000 149.400 ;
        RECT 749.100 144.000 750.900 156.000 ;
        RECT 752.100 143.400 753.900 155.400 ;
        RECT 767.100 149.400 768.900 156.000 ;
        RECT 770.100 149.400 771.900 155.400 ;
        RECT 773.100 149.400 774.900 156.000 ;
        RECT 748.200 136.050 750.000 137.850 ;
        RECT 752.400 136.050 753.300 143.400 ;
        RECT 770.100 136.050 771.300 149.400 ;
        RECT 788.100 144.600 789.900 155.400 ;
        RECT 791.100 145.500 792.900 156.000 ;
        RECT 794.100 154.500 801.900 155.400 ;
        RECT 794.100 144.600 795.900 154.500 ;
        RECT 788.100 143.700 795.900 144.600 ;
        RECT 797.100 142.500 798.900 153.600 ;
        RECT 800.100 143.400 801.900 154.500 ;
        RECT 815.100 143.400 816.900 155.400 ;
        RECT 818.100 144.300 819.900 155.400 ;
        RECT 821.100 145.200 822.900 156.000 ;
        RECT 824.100 144.300 825.900 155.400 ;
        RECT 839.100 149.400 840.900 155.400 ;
        RECT 842.100 150.000 843.900 156.000 ;
        RECT 818.100 143.400 825.900 144.300 ;
        RECT 840.000 149.100 840.900 149.400 ;
        RECT 845.100 149.400 846.900 155.400 ;
        RECT 848.100 149.400 849.900 156.000 ;
        RECT 863.100 149.400 864.900 156.000 ;
        RECT 866.100 149.400 867.900 155.400 ;
        RECT 869.100 149.400 870.900 156.000 ;
        RECT 887.100 149.400 888.900 156.000 ;
        RECT 890.100 149.400 891.900 155.400 ;
        RECT 845.100 149.100 846.600 149.400 ;
        RECT 840.000 148.200 846.600 149.100 ;
        RECT 781.950 141.450 784.050 142.050 ;
        RECT 790.950 141.450 793.050 142.050 ;
        RECT 781.950 140.550 793.050 141.450 ;
        RECT 781.950 139.950 784.050 140.550 ;
        RECT 790.950 139.950 793.050 140.550 ;
        RECT 794.100 141.600 798.900 142.500 ;
        RECT 791.250 136.050 793.050 137.850 ;
        RECT 794.100 136.050 795.000 141.600 ;
        RECT 797.100 136.050 798.900 137.850 ;
        RECT 815.400 136.050 816.300 143.400 ;
        RECT 820.950 141.450 823.050 142.050 ;
        RECT 820.950 140.550 831.450 141.450 ;
        RECT 820.950 139.950 823.050 140.550 ;
        RECT 820.950 136.050 822.750 137.850 ;
        RECT 748.500 133.950 750.600 136.050 ;
        RECT 751.800 133.950 753.900 136.050 ;
        RECT 766.950 133.950 769.050 136.050 ;
        RECT 769.950 133.950 772.050 136.050 ;
        RECT 772.950 133.950 775.050 136.050 ;
        RECT 787.950 133.950 790.050 136.050 ;
        RECT 790.950 133.950 793.050 136.050 ;
        RECT 793.950 133.950 796.050 136.050 ;
        RECT 796.950 133.950 799.050 136.050 ;
        RECT 799.950 133.950 802.050 136.050 ;
        RECT 814.950 133.950 817.050 136.050 ;
        RECT 817.950 133.950 820.050 136.050 ;
        RECT 820.950 133.950 823.050 136.050 ;
        RECT 823.950 133.950 826.050 136.050 ;
        RECT 743.100 128.400 751.500 129.300 ;
        RECT 743.100 120.600 744.900 128.400 ;
        RECT 749.700 127.500 751.500 128.400 ;
        RECT 752.400 126.600 753.300 133.950 ;
        RECT 767.250 132.150 769.050 133.950 ;
        RECT 770.100 128.700 771.300 133.950 ;
        RECT 773.100 132.150 774.900 133.950 ;
        RECT 788.250 132.150 790.050 133.950 ;
        RECT 770.100 127.800 774.300 128.700 ;
        RECT 747.600 120.000 749.400 126.600 ;
        RECT 750.600 124.800 753.300 126.600 ;
        RECT 750.600 120.600 752.400 124.800 ;
        RECT 767.400 120.000 769.200 126.600 ;
        RECT 772.500 120.600 774.300 127.800 ;
        RECT 794.100 126.600 795.300 133.950 ;
        RECT 800.100 132.150 801.900 133.950 ;
        RECT 815.400 126.600 816.300 133.950 ;
        RECT 817.950 132.150 819.750 133.950 ;
        RECT 824.100 132.150 825.900 133.950 ;
        RECT 830.550 132.450 831.450 140.550 ;
        RECT 840.000 136.050 840.900 148.200 ;
        RECT 841.950 141.450 844.050 142.050 ;
        RECT 853.950 141.450 856.050 142.050 ;
        RECT 841.950 140.550 856.050 141.450 ;
        RECT 841.950 139.950 844.050 140.550 ;
        RECT 853.950 139.950 856.050 140.550 ;
        RECT 845.100 136.050 846.900 137.850 ;
        RECT 866.700 136.050 867.900 149.400 ;
        RECT 887.100 136.050 888.900 137.850 ;
        RECT 890.100 136.050 891.300 149.400 ;
        RECT 838.950 133.950 841.050 136.050 ;
        RECT 841.950 133.950 844.050 136.050 ;
        RECT 844.950 133.950 847.050 136.050 ;
        RECT 847.950 133.950 850.050 136.050 ;
        RECT 862.950 133.950 865.050 136.050 ;
        RECT 865.950 133.950 868.050 136.050 ;
        RECT 868.950 133.950 871.050 136.050 ;
        RECT 886.950 133.950 889.050 136.050 ;
        RECT 889.950 133.950 892.050 136.050 ;
        RECT 827.550 131.550 831.450 132.450 ;
        RECT 820.950 129.450 823.050 129.750 ;
        RECT 827.550 129.450 828.450 131.550 ;
        RECT 820.950 128.550 828.450 129.450 ;
        RECT 840.000 130.200 840.900 133.950 ;
        RECT 842.100 132.150 843.900 133.950 ;
        RECT 848.100 132.150 849.900 133.950 ;
        RECT 863.100 132.150 864.900 133.950 ;
        RECT 840.000 129.000 843.300 130.200 ;
        RECT 820.950 127.650 823.050 128.550 ;
        RECT 788.700 120.000 790.500 126.600 ;
        RECT 793.200 120.600 795.000 126.600 ;
        RECT 797.700 120.000 799.500 126.600 ;
        RECT 815.400 125.400 820.500 126.600 ;
        RECT 815.700 120.000 817.500 123.600 ;
        RECT 818.700 120.600 820.500 125.400 ;
        RECT 823.200 120.000 825.000 126.600 ;
        RECT 841.500 120.600 843.300 129.000 ;
        RECT 848.100 120.000 849.900 129.600 ;
        RECT 866.700 128.700 867.900 133.950 ;
        RECT 868.950 132.150 870.750 133.950 ;
        RECT 863.700 127.800 867.900 128.700 ;
        RECT 863.700 120.600 865.500 127.800 ;
        RECT 868.800 120.000 870.600 126.600 ;
        RECT 890.100 123.600 891.300 133.950 ;
        RECT 887.100 120.000 888.900 123.600 ;
        RECT 890.100 120.600 891.900 123.600 ;
        RECT 19.500 108.000 21.300 116.400 ;
        RECT 18.000 106.800 21.300 108.000 ;
        RECT 26.100 107.400 27.900 117.000 ;
        RECT 42.000 110.400 43.800 117.000 ;
        RECT 46.500 111.600 48.300 116.400 ;
        RECT 49.500 113.400 51.300 117.000 ;
        RECT 46.500 110.400 51.600 111.600 ;
        RECT 18.000 103.050 18.900 106.800 ;
        RECT 20.100 103.050 21.900 104.850 ;
        RECT 26.100 103.050 27.900 104.850 ;
        RECT 41.100 103.050 42.900 104.850 ;
        RECT 47.250 103.050 49.050 104.850 ;
        RECT 50.700 103.050 51.600 110.400 ;
        RECT 58.950 106.950 61.050 109.050 ;
        RECT 65.100 107.400 66.900 117.000 ;
        RECT 71.700 108.000 73.500 116.400 ;
        RECT 89.100 113.400 90.900 117.000 ;
        RECT 92.100 113.400 93.900 116.400 ;
        RECT 16.950 100.950 19.050 103.050 ;
        RECT 19.950 100.950 22.050 103.050 ;
        RECT 22.950 100.950 25.050 103.050 ;
        RECT 25.950 100.950 28.050 103.050 ;
        RECT 40.950 100.950 43.050 103.050 ;
        RECT 43.950 100.950 46.050 103.050 ;
        RECT 46.950 100.950 49.050 103.050 ;
        RECT 49.950 100.950 52.050 103.050 ;
        RECT 18.000 88.800 18.900 100.950 ;
        RECT 23.100 99.150 24.900 100.950 ;
        RECT 44.250 99.150 46.050 100.950 ;
        RECT 19.950 96.450 22.050 97.050 ;
        RECT 34.950 96.450 37.050 97.050 ;
        RECT 46.950 96.450 49.050 97.050 ;
        RECT 19.950 95.550 49.050 96.450 ;
        RECT 19.950 94.950 22.050 95.550 ;
        RECT 34.950 94.950 37.050 95.550 ;
        RECT 46.950 94.950 49.050 95.550 ;
        RECT 50.700 93.600 51.600 100.950 ;
        RECT 59.550 100.050 60.450 106.950 ;
        RECT 71.700 106.800 75.000 108.000 ;
        RECT 65.100 103.050 66.900 104.850 ;
        RECT 71.100 103.050 72.900 104.850 ;
        RECT 74.100 103.050 75.000 106.800 ;
        RECT 92.100 103.050 93.300 113.400 ;
        RECT 107.100 111.300 108.900 116.400 ;
        RECT 110.100 112.200 111.900 117.000 ;
        RECT 113.100 111.300 114.900 116.400 ;
        RECT 107.100 109.950 114.900 111.300 ;
        RECT 116.100 110.400 117.900 116.400 ;
        RECT 116.100 108.300 117.300 110.400 ;
        RECT 131.700 109.200 133.500 116.400 ;
        RECT 136.800 110.400 138.600 117.000 ;
        RECT 152.100 110.400 153.900 116.400 ;
        RECT 155.400 111.300 157.200 117.000 ;
        RECT 159.900 111.000 161.700 116.400 ;
        RECT 164.100 111.300 165.900 117.000 ;
        RECT 152.100 109.500 156.600 110.400 ;
        RECT 131.700 108.300 135.900 109.200 ;
        RECT 113.700 107.400 117.300 108.300 ;
        RECT 110.100 103.050 111.900 104.850 ;
        RECT 113.700 103.050 114.900 107.400 ;
        RECT 116.100 103.050 117.900 104.850 ;
        RECT 131.100 103.050 132.900 104.850 ;
        RECT 134.700 103.050 135.900 108.300 ;
        RECT 154.500 107.100 156.600 109.500 ;
        RECT 159.900 108.900 160.800 111.000 ;
        RECT 167.100 110.400 168.900 116.400 ;
        RECT 183.600 112.200 185.400 116.400 ;
        RECT 167.400 109.500 168.900 110.400 ;
        RECT 157.800 106.800 160.800 108.900 ;
        RECT 164.400 108.000 168.900 109.500 ;
        RECT 182.700 110.400 185.400 112.200 ;
        RECT 186.600 110.400 188.400 117.000 ;
        RECT 136.950 103.050 138.750 104.850 ;
        RECT 64.950 100.950 67.050 103.050 ;
        RECT 67.950 100.950 70.050 103.050 ;
        RECT 70.950 100.950 73.050 103.050 ;
        RECT 73.950 100.950 76.050 103.050 ;
        RECT 88.950 100.950 91.050 103.050 ;
        RECT 91.950 100.950 94.050 103.050 ;
        RECT 106.950 100.950 109.050 103.050 ;
        RECT 109.950 100.950 112.050 103.050 ;
        RECT 112.950 100.950 115.050 103.050 ;
        RECT 115.950 100.950 118.050 103.050 ;
        RECT 130.950 100.950 133.050 103.050 ;
        RECT 133.950 100.950 136.050 103.050 ;
        RECT 136.950 100.950 139.050 103.050 ;
        RECT 152.100 100.950 154.200 103.050 ;
        RECT 156.900 102.900 159.000 105.000 ;
        RECT 157.200 101.100 159.000 102.900 ;
        RECT 59.550 98.550 64.050 100.050 ;
        RECT 68.100 99.150 69.900 100.950 ;
        RECT 60.000 97.950 64.050 98.550 ;
        RECT 41.100 92.700 48.900 93.600 ;
        RECT 18.000 87.900 24.600 88.800 ;
        RECT 18.000 87.600 18.900 87.900 ;
        RECT 17.100 81.600 18.900 87.600 ;
        RECT 23.100 87.600 24.600 87.900 ;
        RECT 20.100 81.000 21.900 87.000 ;
        RECT 23.100 81.600 24.900 87.600 ;
        RECT 26.100 81.000 27.900 87.600 ;
        RECT 41.100 81.600 42.900 92.700 ;
        RECT 44.100 81.000 45.900 91.800 ;
        RECT 47.100 81.600 48.900 92.700 ;
        RECT 50.100 81.600 51.900 93.600 ;
        RECT 61.950 93.450 64.050 94.050 ;
        RECT 70.950 93.450 73.050 93.900 ;
        RECT 61.950 92.550 73.050 93.450 ;
        RECT 61.950 91.950 64.050 92.550 ;
        RECT 70.950 91.800 73.050 92.550 ;
        RECT 74.100 88.800 75.000 100.950 ;
        RECT 89.100 99.150 90.900 100.950 ;
        RECT 68.400 87.900 75.000 88.800 ;
        RECT 68.400 87.600 69.900 87.900 ;
        RECT 65.100 81.000 66.900 87.600 ;
        RECT 68.100 81.600 69.900 87.600 ;
        RECT 74.100 87.600 75.000 87.900 ;
        RECT 92.100 87.600 93.300 100.950 ;
        RECT 107.100 99.150 108.900 100.950 ;
        RECT 113.700 93.600 114.900 100.950 ;
        RECT 71.100 81.000 72.900 87.000 ;
        RECT 74.100 81.600 75.900 87.600 ;
        RECT 89.100 81.000 90.900 87.600 ;
        RECT 92.100 81.600 93.900 87.600 ;
        RECT 107.400 81.000 109.200 93.600 ;
        RECT 112.500 92.100 114.900 93.600 ;
        RECT 112.500 81.600 114.300 92.100 ;
        RECT 115.200 89.100 117.000 90.900 ;
        RECT 134.700 87.600 135.900 100.950 ;
        RECT 152.400 99.150 154.200 100.950 ;
        RECT 159.900 100.050 160.800 106.800 ;
        RECT 161.700 105.900 163.500 107.700 ;
        RECT 164.400 107.400 166.500 108.000 ;
        RECT 162.000 105.000 164.100 105.900 ;
        RECT 162.000 103.800 168.600 105.000 ;
        RECT 166.800 103.200 168.600 103.800 ;
        RECT 162.000 100.800 164.100 102.900 ;
        RECT 166.800 100.950 168.900 103.200 ;
        RECT 182.700 103.050 183.600 110.400 ;
        RECT 184.500 108.600 186.300 109.500 ;
        RECT 191.100 108.600 192.900 116.400 ;
        RECT 184.500 107.700 192.900 108.600 ;
        RECT 206.700 109.200 208.500 116.400 ;
        RECT 211.800 110.400 213.600 117.000 ;
        RECT 230.100 111.300 231.900 116.400 ;
        RECT 233.100 112.200 234.900 117.000 ;
        RECT 236.100 111.300 237.900 116.400 ;
        RECT 230.100 109.950 237.900 111.300 ;
        RECT 239.100 110.400 240.900 116.400 ;
        RECT 206.700 108.300 210.900 109.200 ;
        RECT 239.100 108.300 240.300 110.400 ;
        RECT 182.100 100.950 184.200 103.050 ;
        RECT 185.400 100.950 187.500 103.050 ;
        RECT 157.800 98.700 160.800 100.050 ;
        RECT 162.300 99.000 164.100 100.800 ;
        RECT 157.800 97.950 159.900 98.700 ;
        RECT 136.950 96.450 139.050 97.050 ;
        RECT 142.950 96.450 145.050 97.050 ;
        RECT 136.950 95.550 145.050 96.450 ;
        RECT 136.950 94.950 139.050 95.550 ;
        RECT 142.950 94.950 145.050 95.550 ;
        RECT 155.100 93.600 157.200 94.500 ;
        RECT 152.100 92.400 157.200 93.600 ;
        RECT 158.100 93.600 159.300 97.950 ;
        RECT 160.800 95.700 162.600 97.500 ;
        RECT 160.800 94.800 166.200 95.700 ;
        RECT 164.100 93.900 166.200 94.800 ;
        RECT 158.100 92.700 161.400 93.600 ;
        RECT 164.100 92.700 168.900 93.900 ;
        RECT 182.700 93.600 183.600 100.950 ;
        RECT 186.000 99.150 187.800 100.950 ;
        RECT 115.500 81.000 117.300 87.600 ;
        RECT 131.100 81.000 132.900 87.600 ;
        RECT 134.100 81.600 135.900 87.600 ;
        RECT 137.100 81.000 138.900 87.600 ;
        RECT 152.100 81.600 153.900 92.400 ;
        RECT 155.100 81.000 157.200 91.500 ;
        RECT 159.600 81.600 161.400 92.700 ;
        RECT 164.100 81.000 165.900 91.500 ;
        RECT 167.100 81.600 168.900 92.700 ;
        RECT 182.100 81.600 183.900 93.600 ;
        RECT 185.100 81.000 186.900 93.000 ;
        RECT 189.000 87.600 189.900 107.700 ;
        RECT 190.950 103.050 192.750 104.850 ;
        RECT 206.100 103.050 207.900 104.850 ;
        RECT 209.700 103.050 210.900 108.300 ;
        RECT 236.700 107.400 240.300 108.300 ;
        RECT 256.500 108.000 258.300 116.400 ;
        RECT 211.950 103.050 213.750 104.850 ;
        RECT 233.100 103.050 234.900 104.850 ;
        RECT 236.700 103.050 237.900 107.400 ;
        RECT 255.000 106.800 258.300 108.000 ;
        RECT 263.100 107.400 264.900 117.000 ;
        RECT 278.400 110.400 280.200 117.000 ;
        RECT 283.500 109.200 285.300 116.400 ;
        RECT 299.100 110.400 300.900 116.400 ;
        RECT 302.400 111.300 304.200 117.000 ;
        RECT 306.900 111.000 308.700 116.400 ;
        RECT 311.100 111.300 312.900 117.000 ;
        RECT 299.100 109.500 303.600 110.400 ;
        RECT 281.100 108.300 285.300 109.200 ;
        RECT 239.100 103.050 240.900 104.850 ;
        RECT 255.000 103.050 255.900 106.800 ;
        RECT 257.100 103.050 258.900 104.850 ;
        RECT 263.100 103.050 264.900 104.850 ;
        RECT 278.250 103.050 280.050 104.850 ;
        RECT 281.100 103.050 282.300 108.300 ;
        RECT 301.500 107.100 303.600 109.500 ;
        RECT 306.900 108.900 307.800 111.000 ;
        RECT 314.100 110.400 315.900 116.400 ;
        RECT 318.150 112.200 319.950 116.400 ;
        RECT 314.400 109.500 315.900 110.400 ;
        RECT 304.800 106.800 307.800 108.900 ;
        RECT 311.400 108.000 315.900 109.500 ;
        RECT 317.550 110.400 319.950 112.200 ;
        RECT 321.150 110.400 322.950 117.000 ;
        RECT 325.950 114.300 327.750 116.400 ;
        RECT 324.150 113.400 327.750 114.300 ;
        RECT 330.450 113.400 332.250 117.000 ;
        RECT 333.750 113.400 335.550 116.400 ;
        RECT 336.750 113.400 338.550 117.000 ;
        RECT 341.250 113.400 343.050 116.400 ;
        RECT 323.850 112.800 327.750 113.400 ;
        RECT 323.850 111.300 325.950 112.800 ;
        RECT 333.750 112.500 334.800 113.400 ;
        RECT 284.100 103.050 285.900 104.850 ;
        RECT 190.800 100.950 192.900 103.050 ;
        RECT 205.950 100.950 208.050 103.050 ;
        RECT 208.950 100.950 211.050 103.050 ;
        RECT 211.950 100.950 214.050 103.050 ;
        RECT 229.950 100.950 232.050 103.050 ;
        RECT 232.950 100.950 235.050 103.050 ;
        RECT 235.950 100.950 238.050 103.050 ;
        RECT 238.950 100.950 241.050 103.050 ;
        RECT 253.950 100.950 256.050 103.050 ;
        RECT 256.950 100.950 259.050 103.050 ;
        RECT 259.950 100.950 262.050 103.050 ;
        RECT 262.950 100.950 265.050 103.050 ;
        RECT 277.950 100.950 280.050 103.050 ;
        RECT 280.950 100.950 283.050 103.050 ;
        RECT 283.950 100.950 286.050 103.050 ;
        RECT 299.100 100.950 301.200 103.050 ;
        RECT 303.900 102.900 306.000 105.000 ;
        RECT 304.200 101.100 306.000 102.900 ;
        RECT 209.700 87.600 210.900 100.950 ;
        RECT 230.100 99.150 231.900 100.950 ;
        RECT 236.700 93.600 237.900 100.950 ;
        RECT 188.100 81.600 189.900 87.600 ;
        RECT 191.100 81.000 192.900 87.600 ;
        RECT 206.100 81.000 207.900 87.600 ;
        RECT 209.100 81.600 210.900 87.600 ;
        RECT 212.100 81.000 213.900 87.600 ;
        RECT 230.400 81.000 232.200 93.600 ;
        RECT 235.500 92.100 237.900 93.600 ;
        RECT 235.500 81.600 237.300 92.100 ;
        RECT 238.200 89.100 240.000 90.900 ;
        RECT 255.000 88.800 255.900 100.950 ;
        RECT 260.100 99.150 261.900 100.950 ;
        RECT 255.000 87.900 261.600 88.800 ;
        RECT 255.000 87.600 255.900 87.900 ;
        RECT 238.500 81.000 240.300 87.600 ;
        RECT 254.100 81.600 255.900 87.600 ;
        RECT 260.100 87.600 261.600 87.900 ;
        RECT 281.100 87.600 282.300 100.950 ;
        RECT 299.400 99.150 301.200 100.950 ;
        RECT 306.900 100.050 307.800 106.800 ;
        RECT 308.700 105.900 310.500 107.700 ;
        RECT 311.400 107.400 313.500 108.000 ;
        RECT 309.000 105.000 311.100 105.900 ;
        RECT 309.000 103.800 315.600 105.000 ;
        RECT 313.800 103.200 315.600 103.800 ;
        RECT 309.000 100.800 311.100 102.900 ;
        RECT 313.800 100.950 315.900 103.200 ;
        RECT 304.800 98.700 307.800 100.050 ;
        RECT 309.300 99.000 311.100 100.800 ;
        RECT 304.800 97.950 306.900 98.700 ;
        RECT 302.100 93.600 304.200 94.500 ;
        RECT 299.100 92.400 304.200 93.600 ;
        RECT 305.100 93.600 306.300 97.950 ;
        RECT 307.800 95.700 309.600 97.500 ;
        RECT 317.550 95.700 318.450 110.400 ;
        RECT 326.850 109.800 328.650 111.600 ;
        RECT 329.850 111.450 334.800 112.500 ;
        RECT 329.850 110.700 331.650 111.450 ;
        RECT 341.250 111.300 343.650 113.400 ;
        RECT 346.350 110.400 348.150 117.000 ;
        RECT 349.650 110.400 351.450 116.400 ;
        RECT 365.100 113.400 366.900 116.400 ;
        RECT 368.100 113.400 369.900 117.000 ;
        RECT 326.850 108.000 327.900 109.800 ;
        RECT 337.050 108.000 338.850 108.600 ;
        RECT 326.850 106.800 338.850 108.000 ;
        RECT 319.950 105.600 327.900 106.800 ;
        RECT 319.950 103.050 321.750 105.600 ;
        RECT 326.100 105.000 327.900 105.600 ;
        RECT 323.100 103.800 324.900 104.400 ;
        RECT 319.950 100.950 322.050 103.050 ;
        RECT 323.100 102.600 331.200 103.800 ;
        RECT 329.100 100.950 331.200 102.600 ;
        RECT 327.450 95.700 329.250 96.000 ;
        RECT 307.800 94.800 313.200 95.700 ;
        RECT 311.100 93.900 313.200 94.800 ;
        RECT 317.550 95.100 329.250 95.700 ;
        RECT 317.550 94.500 335.850 95.100 ;
        RECT 305.100 92.700 308.400 93.600 ;
        RECT 311.100 92.700 315.900 93.900 ;
        RECT 257.100 81.000 258.900 87.000 ;
        RECT 260.100 81.600 261.900 87.600 ;
        RECT 263.100 81.000 264.900 87.600 ;
        RECT 278.100 81.000 279.900 87.600 ;
        RECT 281.100 81.600 282.900 87.600 ;
        RECT 284.100 81.000 285.900 87.600 ;
        RECT 299.100 81.600 300.900 92.400 ;
        RECT 302.100 81.000 304.200 91.500 ;
        RECT 306.600 81.600 308.400 92.700 ;
        RECT 311.100 81.000 312.900 91.500 ;
        RECT 314.100 81.600 315.900 92.700 ;
        RECT 317.550 93.600 318.450 94.500 ;
        RECT 327.450 94.200 335.850 94.500 ;
        RECT 317.550 91.800 319.950 93.600 ;
        RECT 318.150 81.600 319.950 91.800 ;
        RECT 321.150 81.000 322.950 93.600 ;
        RECT 332.250 92.700 334.050 93.300 ;
        RECT 326.250 91.500 334.050 92.700 ;
        RECT 334.950 92.100 335.850 94.200 ;
        RECT 337.950 94.200 338.850 106.800 ;
        RECT 350.250 103.050 351.450 110.400 ;
        RECT 365.700 103.050 366.900 113.400 ;
        RECT 383.100 111.300 384.900 116.400 ;
        RECT 386.100 112.200 387.900 117.000 ;
        RECT 389.100 111.300 390.900 116.400 ;
        RECT 383.100 109.950 390.900 111.300 ;
        RECT 392.100 110.400 393.900 116.400 ;
        RECT 392.100 108.300 393.300 110.400 ;
        RECT 389.700 107.400 393.300 108.300 ;
        RECT 409.500 108.000 411.300 116.400 ;
        RECT 386.100 103.050 387.900 104.850 ;
        RECT 389.700 103.050 390.900 107.400 ;
        RECT 408.000 106.800 411.300 108.000 ;
        RECT 416.100 107.400 417.900 117.000 ;
        RECT 431.100 107.400 432.900 117.000 ;
        RECT 437.700 108.000 439.500 116.400 ;
        RECT 437.700 106.800 441.000 108.000 ;
        RECT 455.100 107.400 456.900 117.000 ;
        RECT 461.700 108.000 463.500 116.400 ;
        RECT 481.500 108.000 483.300 116.400 ;
        RECT 461.700 106.800 465.000 108.000 ;
        RECT 392.100 103.050 393.900 104.850 ;
        RECT 408.000 103.050 408.900 106.800 ;
        RECT 410.100 103.050 411.900 104.850 ;
        RECT 416.100 103.050 417.900 104.850 ;
        RECT 431.100 103.050 432.900 104.850 ;
        RECT 437.100 103.050 438.900 104.850 ;
        RECT 440.100 103.050 441.000 106.800 ;
        RECT 455.100 103.050 456.900 104.850 ;
        RECT 461.100 103.050 462.900 104.850 ;
        RECT 464.100 103.050 465.000 106.800 ;
        RECT 480.000 106.800 483.300 108.000 ;
        RECT 488.100 107.400 489.900 117.000 ;
        RECT 504.000 110.400 505.800 117.000 ;
        RECT 508.500 111.600 510.300 116.400 ;
        RECT 511.500 113.400 513.300 117.000 ;
        RECT 508.500 110.400 513.600 111.600 ;
        RECT 480.000 103.050 480.900 106.800 ;
        RECT 482.100 103.050 483.900 104.850 ;
        RECT 488.100 103.050 489.900 104.850 ;
        RECT 503.100 103.050 504.900 104.850 ;
        RECT 509.250 103.050 511.050 104.850 ;
        RECT 512.700 103.050 513.600 110.400 ;
        RECT 517.950 108.450 520.050 109.050 ;
        RECT 523.950 108.450 526.050 109.050 ;
        RECT 517.950 107.550 526.050 108.450 ;
        RECT 517.950 106.950 520.050 107.550 ;
        RECT 523.950 106.950 526.050 107.550 ;
        RECT 527.100 107.400 528.900 117.000 ;
        RECT 533.700 108.000 535.500 116.400 ;
        RECT 552.000 110.400 553.800 117.000 ;
        RECT 556.500 111.600 558.300 116.400 ;
        RECT 559.500 113.400 561.300 117.000 ;
        RECT 556.500 110.400 561.600 111.600 ;
        RECT 533.700 106.800 537.000 108.000 ;
        RECT 527.100 103.050 528.900 104.850 ;
        RECT 533.100 103.050 534.900 104.850 ;
        RECT 536.100 103.050 537.000 106.800 ;
        RECT 551.100 103.050 552.900 104.850 ;
        RECT 557.250 103.050 559.050 104.850 ;
        RECT 560.700 103.050 561.600 110.400 ;
        RECT 575.100 111.300 576.900 116.400 ;
        RECT 578.100 112.200 579.900 117.000 ;
        RECT 581.100 111.300 582.900 116.400 ;
        RECT 575.100 109.950 582.900 111.300 ;
        RECT 584.100 110.400 585.900 116.400 ;
        RECT 584.100 108.300 585.300 110.400 ;
        RECT 581.700 107.400 585.300 108.300 ;
        RECT 601.500 108.000 603.300 116.400 ;
        RECT 578.100 103.050 579.900 104.850 ;
        RECT 581.700 103.050 582.900 107.400 ;
        RECT 600.000 106.800 603.300 108.000 ;
        RECT 608.100 107.400 609.900 117.000 ;
        RECT 623.100 113.400 624.900 116.400 ;
        RECT 626.100 113.400 627.900 117.000 ;
        RECT 641.700 113.400 643.500 117.000 ;
        RECT 584.100 103.050 585.900 104.850 ;
        RECT 600.000 103.050 600.900 106.800 ;
        RECT 602.100 103.050 603.900 104.850 ;
        RECT 608.100 103.050 609.900 104.850 ;
        RECT 623.700 103.050 624.900 113.400 ;
        RECT 644.700 111.600 646.500 116.400 ;
        RECT 641.400 110.400 646.500 111.600 ;
        RECT 649.200 110.400 651.000 117.000 ;
        RECT 665.100 113.400 666.900 116.400 ;
        RECT 668.100 113.400 669.900 117.000 ;
        RECT 625.950 108.450 628.050 109.200 ;
        RECT 631.950 108.450 634.050 109.050 ;
        RECT 625.950 107.550 634.050 108.450 ;
        RECT 625.950 107.100 628.050 107.550 ;
        RECT 631.950 106.950 634.050 107.550 ;
        RECT 641.400 103.050 642.300 110.400 ;
        RECT 643.950 103.050 645.750 104.850 ;
        RECT 650.100 103.050 651.900 104.850 ;
        RECT 665.700 103.050 666.900 113.400 ;
        RECT 686.100 110.400 687.900 116.400 ;
        RECT 686.700 108.300 687.900 110.400 ;
        RECT 689.100 111.300 690.900 116.400 ;
        RECT 692.100 112.200 693.900 117.000 ;
        RECT 695.100 111.300 696.900 116.400 ;
        RECT 689.100 109.950 696.900 111.300 ;
        RECT 686.700 107.400 690.300 108.300 ;
        RECT 713.100 107.400 714.900 117.000 ;
        RECT 719.700 108.000 721.500 116.400 ;
        RECT 737.100 113.400 738.900 117.000 ;
        RECT 740.100 113.400 741.900 116.400 ;
        RECT 686.100 103.050 687.900 104.850 ;
        RECT 689.100 103.050 690.300 107.400 ;
        RECT 719.700 106.800 723.000 108.000 ;
        RECT 692.100 103.050 693.900 104.850 ;
        RECT 713.100 103.050 714.900 104.850 ;
        RECT 719.100 103.050 720.900 104.850 ;
        RECT 722.100 103.050 723.000 106.800 ;
        RECT 740.100 103.050 741.300 113.400 ;
        RECT 757.500 108.000 759.300 116.400 ;
        RECT 756.000 106.800 759.300 108.000 ;
        RECT 764.100 107.400 765.900 117.000 ;
        RECT 779.700 113.400 781.500 117.000 ;
        RECT 782.700 111.600 784.500 116.400 ;
        RECT 779.400 110.400 784.500 111.600 ;
        RECT 787.200 110.400 789.000 117.000 ;
        RECT 803.700 113.400 805.500 117.000 ;
        RECT 806.700 111.600 808.500 116.400 ;
        RECT 803.400 110.400 808.500 111.600 ;
        RECT 811.200 110.400 813.000 117.000 ;
        RECT 756.000 103.050 756.900 106.800 ;
        RECT 758.100 103.050 759.900 104.850 ;
        RECT 764.100 103.050 765.900 104.850 ;
        RECT 779.400 103.050 780.300 110.400 ;
        RECT 781.950 108.450 784.050 109.050 ;
        RECT 793.950 108.450 796.050 109.050 ;
        RECT 781.950 107.550 796.050 108.450 ;
        RECT 781.950 106.950 784.050 107.550 ;
        RECT 793.950 106.950 796.050 107.550 ;
        RECT 781.950 103.050 783.750 104.850 ;
        RECT 788.100 103.050 789.900 104.850 ;
        RECT 803.400 103.050 804.300 110.400 ;
        RECT 829.500 108.000 831.300 116.400 ;
        RECT 828.000 106.800 831.300 108.000 ;
        RECT 836.100 107.400 837.900 117.000 ;
        RECT 851.400 110.400 853.200 117.000 ;
        RECT 856.500 109.200 858.300 116.400 ;
        RECT 872.400 110.400 874.200 117.000 ;
        RECT 877.500 109.200 879.300 116.400 ;
        RECT 854.100 108.300 858.300 109.200 ;
        RECT 875.100 108.300 879.300 109.200 ;
        RECT 805.950 103.050 807.750 104.850 ;
        RECT 812.100 103.050 813.900 104.850 ;
        RECT 828.000 103.050 828.900 106.800 ;
        RECT 830.100 103.050 831.900 104.850 ;
        RECT 836.100 103.050 837.900 104.850 ;
        RECT 851.250 103.050 853.050 104.850 ;
        RECT 854.100 103.050 855.300 108.300 ;
        RECT 857.100 103.050 858.900 104.850 ;
        RECT 872.250 103.050 874.050 104.850 ;
        RECT 875.100 103.050 876.300 108.300 ;
        RECT 878.100 103.050 879.900 104.850 ;
        RECT 345.150 101.250 351.450 103.050 ;
        RECT 346.950 100.950 351.450 101.250 ;
        RECT 364.950 100.950 367.050 103.050 ;
        RECT 367.950 100.950 370.050 103.050 ;
        RECT 382.950 100.950 385.050 103.050 ;
        RECT 385.950 100.950 388.050 103.050 ;
        RECT 388.950 100.950 391.050 103.050 ;
        RECT 391.950 100.950 394.050 103.050 ;
        RECT 406.950 100.950 409.050 103.050 ;
        RECT 409.950 100.950 412.050 103.050 ;
        RECT 412.950 100.950 415.050 103.050 ;
        RECT 415.950 100.950 418.050 103.050 ;
        RECT 430.950 100.950 433.050 103.050 ;
        RECT 433.950 100.950 436.050 103.050 ;
        RECT 436.950 100.950 439.050 103.050 ;
        RECT 439.950 100.950 442.050 103.050 ;
        RECT 454.950 100.950 457.050 103.050 ;
        RECT 457.950 100.950 460.050 103.050 ;
        RECT 460.950 100.950 463.050 103.050 ;
        RECT 463.950 100.950 466.050 103.050 ;
        RECT 478.950 100.950 481.050 103.050 ;
        RECT 481.950 100.950 484.050 103.050 ;
        RECT 484.950 100.950 487.050 103.050 ;
        RECT 487.950 100.950 490.050 103.050 ;
        RECT 502.950 100.950 505.050 103.050 ;
        RECT 505.950 100.950 508.050 103.050 ;
        RECT 508.950 100.950 511.050 103.050 ;
        RECT 511.950 100.950 514.050 103.050 ;
        RECT 526.950 100.950 529.050 103.050 ;
        RECT 529.950 100.950 532.050 103.050 ;
        RECT 532.950 100.950 535.050 103.050 ;
        RECT 535.950 100.950 538.050 103.050 ;
        RECT 550.950 100.950 553.050 103.050 ;
        RECT 553.950 100.950 556.050 103.050 ;
        RECT 556.950 100.950 559.050 103.050 ;
        RECT 559.950 100.950 562.050 103.050 ;
        RECT 574.950 100.950 577.050 103.050 ;
        RECT 577.950 100.950 580.050 103.050 ;
        RECT 580.950 100.950 583.050 103.050 ;
        RECT 583.950 100.950 586.050 103.050 ;
        RECT 598.950 100.950 601.050 103.050 ;
        RECT 601.950 100.950 604.050 103.050 ;
        RECT 604.950 100.950 607.050 103.050 ;
        RECT 607.950 100.950 610.050 103.050 ;
        RECT 622.950 100.950 625.050 103.050 ;
        RECT 625.950 100.950 628.050 103.050 ;
        RECT 640.950 100.950 643.050 103.050 ;
        RECT 643.950 100.950 646.050 103.050 ;
        RECT 646.950 100.950 649.050 103.050 ;
        RECT 649.950 100.950 652.050 103.050 ;
        RECT 664.950 100.950 667.050 103.050 ;
        RECT 667.950 100.950 670.050 103.050 ;
        RECT 685.950 100.950 688.050 103.050 ;
        RECT 688.950 100.950 691.050 103.050 ;
        RECT 691.950 100.950 694.050 103.050 ;
        RECT 694.950 100.950 697.050 103.050 ;
        RECT 712.950 100.950 715.050 103.050 ;
        RECT 715.950 100.950 718.050 103.050 ;
        RECT 718.950 100.950 721.050 103.050 ;
        RECT 721.950 100.950 724.050 103.050 ;
        RECT 736.950 100.950 739.050 103.050 ;
        RECT 739.950 100.950 742.050 103.050 ;
        RECT 754.950 100.950 757.050 103.050 ;
        RECT 757.950 100.950 760.050 103.050 ;
        RECT 760.950 100.950 763.050 103.050 ;
        RECT 763.950 100.950 766.050 103.050 ;
        RECT 778.950 100.950 781.050 103.050 ;
        RECT 781.950 100.950 784.050 103.050 ;
        RECT 784.950 100.950 787.050 103.050 ;
        RECT 787.950 100.950 790.050 103.050 ;
        RECT 802.950 100.950 805.050 103.050 ;
        RECT 805.950 100.950 808.050 103.050 ;
        RECT 808.950 100.950 811.050 103.050 ;
        RECT 811.950 100.950 814.050 103.050 ;
        RECT 826.950 100.950 829.050 103.050 ;
        RECT 829.950 100.950 832.050 103.050 ;
        RECT 832.950 100.950 835.050 103.050 ;
        RECT 835.950 100.950 838.050 103.050 ;
        RECT 850.950 100.950 853.050 103.050 ;
        RECT 853.950 100.950 856.050 103.050 ;
        RECT 856.950 100.950 859.050 103.050 ;
        RECT 341.550 98.100 343.650 98.400 ;
        RECT 347.550 98.100 349.350 98.250 ;
        RECT 341.550 96.900 349.350 98.100 ;
        RECT 341.550 96.300 343.650 96.900 ;
        RECT 347.550 96.450 349.350 96.900 ;
        RECT 337.950 93.300 342.750 94.200 ;
        RECT 350.250 93.600 351.450 100.950 ;
        RECT 341.550 92.400 342.750 93.300 ;
        RECT 338.850 92.100 340.650 92.400 ;
        RECT 326.250 90.600 328.350 91.500 ;
        RECT 334.950 91.200 340.650 92.100 ;
        RECT 338.850 90.600 340.650 91.200 ;
        RECT 341.550 90.600 344.550 92.400 ;
        RECT 326.550 81.600 328.350 90.600 ;
        RECT 330.450 89.550 332.250 90.300 ;
        RECT 335.250 89.550 337.050 90.300 ;
        RECT 330.450 88.500 337.050 89.550 ;
        RECT 331.350 81.000 333.150 87.600 ;
        RECT 334.350 81.600 336.150 88.500 ;
        RECT 341.550 87.600 343.650 89.700 ;
        RECT 337.350 81.000 339.150 87.600 ;
        RECT 341.850 81.600 343.650 87.600 ;
        RECT 346.650 81.000 348.450 93.600 ;
        RECT 349.650 81.600 351.450 93.600 ;
        RECT 365.700 87.600 366.900 100.950 ;
        RECT 368.100 99.150 369.900 100.950 ;
        RECT 383.100 99.150 384.900 100.950 ;
        RECT 389.700 93.600 390.900 100.950 ;
        RECT 365.100 81.600 366.900 87.600 ;
        RECT 368.100 81.000 369.900 87.600 ;
        RECT 383.400 81.000 385.200 93.600 ;
        RECT 388.500 92.100 390.900 93.600 ;
        RECT 388.500 81.600 390.300 92.100 ;
        RECT 391.200 89.100 393.000 90.900 ;
        RECT 408.000 88.800 408.900 100.950 ;
        RECT 413.100 99.150 414.900 100.950 ;
        RECT 434.100 99.150 435.900 100.950 ;
        RECT 440.100 88.800 441.000 100.950 ;
        RECT 458.100 99.150 459.900 100.950 ;
        RECT 464.100 88.800 465.000 100.950 ;
        RECT 408.000 87.900 414.600 88.800 ;
        RECT 408.000 87.600 408.900 87.900 ;
        RECT 391.500 81.000 393.300 87.600 ;
        RECT 407.100 81.600 408.900 87.600 ;
        RECT 413.100 87.600 414.600 87.900 ;
        RECT 434.400 87.900 441.000 88.800 ;
        RECT 434.400 87.600 435.900 87.900 ;
        RECT 410.100 81.000 411.900 87.000 ;
        RECT 413.100 81.600 414.900 87.600 ;
        RECT 416.100 81.000 417.900 87.600 ;
        RECT 431.100 81.000 432.900 87.600 ;
        RECT 434.100 81.600 435.900 87.600 ;
        RECT 440.100 87.600 441.000 87.900 ;
        RECT 458.400 87.900 465.000 88.800 ;
        RECT 458.400 87.600 459.900 87.900 ;
        RECT 437.100 81.000 438.900 87.000 ;
        RECT 440.100 81.600 441.900 87.600 ;
        RECT 455.100 81.000 456.900 87.600 ;
        RECT 458.100 81.600 459.900 87.600 ;
        RECT 464.100 87.600 465.000 87.900 ;
        RECT 480.000 88.800 480.900 100.950 ;
        RECT 485.100 99.150 486.900 100.950 ;
        RECT 506.250 99.150 508.050 100.950 ;
        RECT 487.950 93.450 490.050 94.050 ;
        RECT 496.950 93.450 499.050 94.050 ;
        RECT 512.700 93.600 513.600 100.950 ;
        RECT 530.100 99.150 531.900 100.950 ;
        RECT 517.950 96.450 520.050 97.050 ;
        RECT 526.950 96.450 529.050 96.750 ;
        RECT 517.950 95.550 529.050 96.450 ;
        RECT 517.950 94.950 520.050 95.550 ;
        RECT 526.950 94.650 529.050 95.550 ;
        RECT 487.950 92.550 499.050 93.450 ;
        RECT 487.950 91.950 490.050 92.550 ;
        RECT 496.950 91.950 499.050 92.550 ;
        RECT 503.100 92.700 510.900 93.600 ;
        RECT 480.000 87.900 486.600 88.800 ;
        RECT 480.000 87.600 480.900 87.900 ;
        RECT 461.100 81.000 462.900 87.000 ;
        RECT 464.100 81.600 465.900 87.600 ;
        RECT 479.100 81.600 480.900 87.600 ;
        RECT 485.100 87.600 486.600 87.900 ;
        RECT 482.100 81.000 483.900 87.000 ;
        RECT 485.100 81.600 486.900 87.600 ;
        RECT 488.100 81.000 489.900 87.600 ;
        RECT 503.100 81.600 504.900 92.700 ;
        RECT 506.100 81.000 507.900 91.800 ;
        RECT 509.100 81.600 510.900 92.700 ;
        RECT 512.100 81.600 513.900 93.600 ;
        RECT 536.100 88.800 537.000 100.950 ;
        RECT 554.250 99.150 556.050 100.950 ;
        RECT 560.700 93.600 561.600 100.950 ;
        RECT 575.100 99.150 576.900 100.950 ;
        RECT 581.700 93.600 582.900 100.950 ;
        RECT 530.400 87.900 537.000 88.800 ;
        RECT 530.400 87.600 531.900 87.900 ;
        RECT 527.100 81.000 528.900 87.600 ;
        RECT 530.100 81.600 531.900 87.600 ;
        RECT 536.100 87.600 537.000 87.900 ;
        RECT 551.100 92.700 558.900 93.600 ;
        RECT 533.100 81.000 534.900 87.000 ;
        RECT 536.100 81.600 537.900 87.600 ;
        RECT 551.100 81.600 552.900 92.700 ;
        RECT 554.100 81.000 555.900 91.800 ;
        RECT 557.100 81.600 558.900 92.700 ;
        RECT 560.100 81.600 561.900 93.600 ;
        RECT 575.400 81.000 577.200 93.600 ;
        RECT 580.500 92.100 582.900 93.600 ;
        RECT 580.500 81.600 582.300 92.100 ;
        RECT 583.200 89.100 585.000 90.900 ;
        RECT 600.000 88.800 600.900 100.950 ;
        RECT 605.100 99.150 606.900 100.950 ;
        RECT 600.000 87.900 606.600 88.800 ;
        RECT 600.000 87.600 600.900 87.900 ;
        RECT 583.500 81.000 585.300 87.600 ;
        RECT 599.100 81.600 600.900 87.600 ;
        RECT 605.100 87.600 606.600 87.900 ;
        RECT 623.700 87.600 624.900 100.950 ;
        RECT 626.100 99.150 627.900 100.950 ;
        RECT 641.400 93.600 642.300 100.950 ;
        RECT 646.950 99.150 648.750 100.950 ;
        RECT 643.950 96.450 646.050 97.050 ;
        RECT 661.950 96.450 664.050 97.050 ;
        RECT 643.950 95.550 664.050 96.450 ;
        RECT 643.950 94.950 646.050 95.550 ;
        RECT 661.950 94.950 664.050 95.550 ;
        RECT 602.100 81.000 603.900 87.000 ;
        RECT 605.100 81.600 606.900 87.600 ;
        RECT 608.100 81.000 609.900 87.600 ;
        RECT 623.100 81.600 624.900 87.600 ;
        RECT 626.100 81.000 627.900 87.600 ;
        RECT 641.100 81.600 642.900 93.600 ;
        RECT 644.100 92.700 651.900 93.600 ;
        RECT 644.100 81.600 645.900 92.700 ;
        RECT 647.100 81.000 648.900 91.800 ;
        RECT 650.100 81.600 651.900 92.700 ;
        RECT 665.700 87.600 666.900 100.950 ;
        RECT 668.100 99.150 669.900 100.950 ;
        RECT 689.100 93.600 690.300 100.950 ;
        RECT 695.100 99.150 696.900 100.950 ;
        RECT 716.100 99.150 717.900 100.950 ;
        RECT 689.100 92.100 691.500 93.600 ;
        RECT 687.000 89.100 688.800 90.900 ;
        RECT 665.100 81.600 666.900 87.600 ;
        RECT 668.100 81.000 669.900 87.600 ;
        RECT 686.700 81.000 688.500 87.600 ;
        RECT 689.700 81.600 691.500 92.100 ;
        RECT 694.800 81.000 696.600 93.600 ;
        RECT 722.100 88.800 723.000 100.950 ;
        RECT 737.100 99.150 738.900 100.950 ;
        RECT 716.400 87.900 723.000 88.800 ;
        RECT 716.400 87.600 717.900 87.900 ;
        RECT 713.100 81.000 714.900 87.600 ;
        RECT 716.100 81.600 717.900 87.600 ;
        RECT 722.100 87.600 723.000 87.900 ;
        RECT 740.100 87.600 741.300 100.950 ;
        RECT 756.000 88.800 756.900 100.950 ;
        RECT 761.100 99.150 762.900 100.950 ;
        RECT 779.400 93.600 780.300 100.950 ;
        RECT 784.950 99.150 786.750 100.950 ;
        RECT 803.400 93.600 804.300 100.950 ;
        RECT 808.950 99.150 810.750 100.950 ;
        RECT 756.000 87.900 762.600 88.800 ;
        RECT 756.000 87.600 756.900 87.900 ;
        RECT 719.100 81.000 720.900 87.000 ;
        RECT 722.100 81.600 723.900 87.600 ;
        RECT 737.100 81.000 738.900 87.600 ;
        RECT 740.100 81.600 741.900 87.600 ;
        RECT 755.100 81.600 756.900 87.600 ;
        RECT 761.100 87.600 762.600 87.900 ;
        RECT 758.100 81.000 759.900 87.000 ;
        RECT 761.100 81.600 762.900 87.600 ;
        RECT 764.100 81.000 765.900 87.600 ;
        RECT 779.100 81.600 780.900 93.600 ;
        RECT 782.100 92.700 789.900 93.600 ;
        RECT 782.100 81.600 783.900 92.700 ;
        RECT 785.100 81.000 786.900 91.800 ;
        RECT 788.100 81.600 789.900 92.700 ;
        RECT 803.100 81.600 804.900 93.600 ;
        RECT 806.100 92.700 813.900 93.600 ;
        RECT 806.100 81.600 807.900 92.700 ;
        RECT 809.100 81.000 810.900 91.800 ;
        RECT 812.100 81.600 813.900 92.700 ;
        RECT 828.000 88.800 828.900 100.950 ;
        RECT 833.100 99.150 834.900 100.950 ;
        RECT 828.000 87.900 834.600 88.800 ;
        RECT 828.000 87.600 828.900 87.900 ;
        RECT 827.100 81.600 828.900 87.600 ;
        RECT 833.100 87.600 834.600 87.900 ;
        RECT 854.100 87.600 855.300 100.950 ;
        RECT 862.950 100.050 865.050 103.050 ;
        RECT 871.950 100.950 874.050 103.050 ;
        RECT 874.950 100.950 877.050 103.050 ;
        RECT 877.950 100.950 880.050 103.050 ;
        RECT 859.950 99.000 865.050 100.050 ;
        RECT 859.950 98.550 864.450 99.000 ;
        RECT 859.950 97.950 864.000 98.550 ;
        RECT 875.100 87.600 876.300 100.950 ;
        RECT 830.100 81.000 831.900 87.000 ;
        RECT 833.100 81.600 834.900 87.600 ;
        RECT 836.100 81.000 837.900 87.600 ;
        RECT 851.100 81.000 852.900 87.600 ;
        RECT 854.100 81.600 855.900 87.600 ;
        RECT 857.100 81.000 858.900 87.600 ;
        RECT 872.100 81.000 873.900 87.600 ;
        RECT 875.100 81.600 876.900 87.600 ;
        RECT 878.100 81.000 879.900 87.600 ;
        RECT 17.100 71.400 18.900 77.400 ;
        RECT 20.100 71.400 21.900 78.000 ;
        RECT 35.100 71.400 36.900 78.000 ;
        RECT 38.100 71.400 39.900 77.400 ;
        RECT 41.100 71.400 42.900 78.000 ;
        RECT 17.700 58.050 18.900 71.400 ;
        RECT 20.100 58.050 21.900 59.850 ;
        RECT 38.100 58.050 39.300 71.400 ;
        RECT 56.400 65.400 58.200 78.000 ;
        RECT 61.500 66.900 63.300 77.400 ;
        RECT 64.500 71.400 66.300 78.000 ;
        RECT 64.200 68.100 66.000 69.900 ;
        RECT 61.500 65.400 63.900 66.900 ;
        RECT 81.000 66.600 82.800 77.400 ;
        RECT 81.000 65.400 84.600 66.600 ;
        RECT 86.100 65.400 87.900 78.000 ;
        RECT 101.700 71.400 103.500 78.000 ;
        RECT 102.000 68.100 103.800 69.900 ;
        RECT 104.700 66.900 106.500 77.400 ;
        RECT 104.100 65.400 106.500 66.900 ;
        RECT 109.800 65.400 111.600 78.000 ;
        RECT 125.100 71.400 126.900 77.400 ;
        RECT 128.100 71.400 129.900 78.000 ;
        RECT 146.100 71.400 147.900 78.000 ;
        RECT 149.100 71.400 150.900 77.400 ;
        RECT 152.100 71.400 153.900 78.000 ;
        RECT 56.100 58.050 57.900 59.850 ;
        RECT 62.700 58.050 63.900 65.400 ;
        RECT 80.100 58.050 81.900 59.850 ;
        RECT 83.700 58.050 84.600 65.400 ;
        RECT 85.950 58.050 87.750 59.850 ;
        RECT 104.100 58.050 105.300 65.400 ;
        RECT 110.100 58.050 111.900 59.850 ;
        RECT 125.700 58.050 126.900 71.400 ;
        RECT 128.100 58.050 129.900 59.850 ;
        RECT 149.700 58.050 150.900 71.400 ;
        RECT 167.100 65.400 168.900 77.400 ;
        RECT 171.600 65.400 173.400 78.000 ;
        RECT 174.600 66.900 176.400 77.400 ;
        RECT 194.100 71.400 195.900 78.000 ;
        RECT 197.100 71.400 198.900 77.400 ;
        RECT 200.100 72.000 201.900 78.000 ;
        RECT 197.400 71.100 198.900 71.400 ;
        RECT 203.100 71.400 204.900 77.400 ;
        RECT 203.100 71.100 204.000 71.400 ;
        RECT 197.400 70.200 204.000 71.100 ;
        RECT 174.600 65.400 177.000 66.900 ;
        RECT 167.100 63.900 168.300 65.400 ;
        RECT 167.100 62.700 174.900 63.900 ;
        RECT 173.100 62.100 174.900 62.700 ;
        RECT 171.000 58.050 172.800 59.850 ;
        RECT 16.950 55.950 19.050 58.050 ;
        RECT 19.950 55.950 22.050 58.050 ;
        RECT 34.950 55.950 37.050 58.050 ;
        RECT 37.950 55.950 40.050 58.050 ;
        RECT 40.950 55.950 43.050 58.050 ;
        RECT 55.950 55.950 58.050 58.050 ;
        RECT 58.950 55.950 61.050 58.050 ;
        RECT 61.950 55.950 64.050 58.050 ;
        RECT 64.950 55.950 67.050 58.050 ;
        RECT 79.950 55.950 82.050 58.050 ;
        RECT 82.950 55.950 85.050 58.050 ;
        RECT 85.950 55.950 88.050 58.050 ;
        RECT 100.950 55.950 103.050 58.050 ;
        RECT 103.950 55.950 106.050 58.050 ;
        RECT 106.950 55.950 109.050 58.050 ;
        RECT 109.950 55.950 112.050 58.050 ;
        RECT 124.950 55.950 127.050 58.050 ;
        RECT 127.950 55.950 130.050 58.050 ;
        RECT 145.950 55.950 148.050 58.050 ;
        RECT 148.950 55.950 151.050 58.050 ;
        RECT 151.950 55.950 154.050 58.050 ;
        RECT 167.100 55.950 169.200 58.050 ;
        RECT 170.400 55.950 172.500 58.050 ;
        RECT 17.700 45.600 18.900 55.950 ;
        RECT 35.250 54.150 37.050 55.950 ;
        RECT 38.100 50.700 39.300 55.950 ;
        RECT 41.100 54.150 42.900 55.950 ;
        RECT 59.100 54.150 60.900 55.950 ;
        RECT 62.700 51.600 63.900 55.950 ;
        RECT 65.100 54.150 66.900 55.950 ;
        RECT 62.700 50.700 66.300 51.600 ;
        RECT 38.100 49.800 42.300 50.700 ;
        RECT 17.100 42.600 18.900 45.600 ;
        RECT 20.100 42.000 21.900 45.600 ;
        RECT 35.400 42.000 37.200 48.600 ;
        RECT 40.500 42.600 42.300 49.800 ;
        RECT 56.100 47.700 63.900 49.050 ;
        RECT 56.100 42.600 57.900 47.700 ;
        RECT 59.100 42.000 60.900 46.800 ;
        RECT 62.100 42.600 63.900 47.700 ;
        RECT 65.100 48.600 66.300 50.700 ;
        RECT 65.100 42.600 66.900 48.600 ;
        RECT 83.700 45.600 84.600 55.950 ;
        RECT 101.100 54.150 102.900 55.950 ;
        RECT 104.100 51.600 105.300 55.950 ;
        RECT 107.100 54.150 108.900 55.950 ;
        RECT 101.700 50.700 105.300 51.600 ;
        RECT 101.700 48.600 102.900 50.700 ;
        RECT 80.100 42.000 81.900 45.600 ;
        RECT 83.100 42.600 84.900 45.600 ;
        RECT 86.100 42.000 87.900 45.600 ;
        RECT 101.100 42.600 102.900 48.600 ;
        RECT 104.100 47.700 111.900 49.050 ;
        RECT 104.100 42.600 105.900 47.700 ;
        RECT 107.100 42.000 108.900 46.800 ;
        RECT 110.100 42.600 111.900 47.700 ;
        RECT 125.700 45.600 126.900 55.950 ;
        RECT 146.100 54.150 147.900 55.950 ;
        RECT 149.700 50.700 150.900 55.950 ;
        RECT 151.950 54.150 153.750 55.950 ;
        RECT 167.400 54.150 169.200 55.950 ;
        RECT 173.700 51.600 174.600 62.100 ;
        RECT 175.800 58.050 177.000 65.400 ;
        RECT 178.950 63.450 181.050 64.050 ;
        RECT 199.950 63.450 202.050 64.050 ;
        RECT 178.950 62.550 202.050 63.450 ;
        RECT 178.950 61.950 181.050 62.550 ;
        RECT 199.950 61.950 202.050 62.550 ;
        RECT 197.100 58.050 198.900 59.850 ;
        RECT 203.100 58.050 204.000 70.200 ;
        RECT 218.100 66.600 219.900 77.400 ;
        RECT 221.100 67.500 222.900 78.000 ;
        RECT 218.100 65.400 222.900 66.600 ;
        RECT 220.800 64.500 222.900 65.400 ;
        RECT 225.600 65.400 227.400 77.400 ;
        RECT 230.100 67.500 231.900 78.000 ;
        RECT 233.100 66.300 234.900 77.400 ;
        RECT 248.700 71.400 250.500 78.000 ;
        RECT 249.000 68.100 250.800 69.900 ;
        RECT 251.700 66.900 253.500 77.400 ;
        RECT 230.400 65.400 234.900 66.300 ;
        RECT 251.100 65.400 253.500 66.900 ;
        RECT 256.800 65.400 258.600 78.000 ;
        RECT 272.100 71.400 273.900 78.000 ;
        RECT 275.100 71.400 276.900 77.400 ;
        RECT 293.100 71.400 294.900 77.400 ;
        RECT 296.100 72.000 297.900 78.000 ;
        RECT 225.600 64.050 226.800 65.400 ;
        RECT 225.300 63.000 226.800 64.050 ;
        RECT 230.400 63.300 232.500 65.400 ;
        RECT 225.300 61.050 226.200 63.000 ;
        RECT 218.400 58.050 220.200 59.850 ;
        RECT 224.100 58.950 226.200 61.050 ;
        RECT 227.100 61.500 229.200 61.800 ;
        RECT 227.100 59.700 231.000 61.500 ;
        RECT 175.800 55.950 177.900 58.050 ;
        RECT 193.950 55.950 196.050 58.050 ;
        RECT 196.950 55.950 199.050 58.050 ;
        RECT 199.950 55.950 202.050 58.050 ;
        RECT 202.950 55.950 205.050 58.050 ;
        RECT 218.100 55.950 220.200 58.050 ;
        RECT 224.700 58.800 226.200 58.950 ;
        RECT 224.700 57.900 227.100 58.800 ;
        RECT 173.700 50.700 175.800 51.600 ;
        RECT 146.700 49.800 150.900 50.700 ;
        RECT 170.400 49.800 175.800 50.700 ;
        RECT 125.100 42.600 126.900 45.600 ;
        RECT 128.100 42.000 129.900 45.600 ;
        RECT 146.700 42.600 148.500 49.800 ;
        RECT 151.800 42.000 153.600 48.600 ;
        RECT 170.400 45.600 171.300 49.800 ;
        RECT 177.000 48.600 177.900 55.950 ;
        RECT 194.100 54.150 195.900 55.950 ;
        RECT 200.100 54.150 201.900 55.950 ;
        RECT 203.100 52.200 204.000 55.950 ;
        RECT 222.900 55.200 224.700 57.000 ;
        RECT 222.900 53.100 225.000 55.200 ;
        RECT 225.900 52.200 227.100 57.900 ;
        RECT 228.000 58.050 229.800 58.500 ;
        RECT 251.100 58.050 252.300 65.400 ;
        RECT 257.100 58.050 258.900 59.850 ;
        RECT 272.100 58.050 273.900 59.850 ;
        RECT 275.100 58.050 276.300 71.400 ;
        RECT 294.000 71.100 294.900 71.400 ;
        RECT 299.100 71.400 300.900 77.400 ;
        RECT 302.100 71.400 303.900 78.000 ;
        RECT 317.100 71.400 318.900 78.000 ;
        RECT 320.100 71.400 321.900 77.400 ;
        RECT 323.100 71.400 324.900 78.000 ;
        RECT 299.100 71.100 300.600 71.400 ;
        RECT 294.000 70.200 300.600 71.100 ;
        RECT 294.000 58.050 294.900 70.200 ;
        RECT 304.950 60.450 307.050 61.050 ;
        RECT 310.950 60.450 313.050 61.050 ;
        RECT 299.100 58.050 300.900 59.850 ;
        RECT 304.950 59.550 313.050 60.450 ;
        RECT 304.950 58.950 307.050 59.550 ;
        RECT 310.950 58.950 313.050 59.550 ;
        RECT 320.700 58.050 321.900 71.400 ;
        RECT 327.150 67.200 328.950 77.400 ;
        RECT 326.550 65.400 328.950 67.200 ;
        RECT 330.150 65.400 331.950 78.000 ;
        RECT 335.550 68.400 337.350 77.400 ;
        RECT 340.350 71.400 342.150 78.000 ;
        RECT 343.350 70.500 345.150 77.400 ;
        RECT 346.350 71.400 348.150 78.000 ;
        RECT 350.850 71.400 352.650 77.400 ;
        RECT 339.450 69.450 346.050 70.500 ;
        RECT 339.450 68.700 341.250 69.450 ;
        RECT 344.250 68.700 346.050 69.450 ;
        RECT 350.550 69.300 352.650 71.400 ;
        RECT 335.250 67.500 337.350 68.400 ;
        RECT 347.850 67.800 349.650 68.400 ;
        RECT 335.250 66.300 343.050 67.500 ;
        RECT 341.250 65.700 343.050 66.300 ;
        RECT 343.950 66.900 349.650 67.800 ;
        RECT 326.550 64.500 327.450 65.400 ;
        RECT 343.950 64.800 344.850 66.900 ;
        RECT 347.850 66.600 349.650 66.900 ;
        RECT 350.550 66.600 353.550 68.400 ;
        RECT 350.550 65.700 351.750 66.600 ;
        RECT 336.450 64.500 344.850 64.800 ;
        RECT 326.550 63.900 344.850 64.500 ;
        RECT 346.950 64.800 351.750 65.700 ;
        RECT 355.650 65.400 357.450 78.000 ;
        RECT 358.650 65.400 360.450 77.400 ;
        RECT 374.100 71.400 375.900 78.000 ;
        RECT 377.100 71.400 378.900 77.400 ;
        RECT 380.100 71.400 381.900 78.000 ;
        RECT 326.550 63.300 338.250 63.900 ;
        RECT 228.000 56.700 234.900 58.050 ;
        RECT 232.800 55.950 234.900 56.700 ;
        RECT 247.950 55.950 250.050 58.050 ;
        RECT 250.950 55.950 253.050 58.050 ;
        RECT 253.950 55.950 256.050 58.050 ;
        RECT 256.950 55.950 259.050 58.050 ;
        RECT 271.950 55.950 274.050 58.050 ;
        RECT 274.950 55.950 277.050 58.050 ;
        RECT 292.950 55.950 295.050 58.050 ;
        RECT 295.950 55.950 298.050 58.050 ;
        RECT 298.950 55.950 301.050 58.050 ;
        RECT 301.950 55.950 304.050 58.050 ;
        RECT 316.950 55.950 319.050 58.050 ;
        RECT 319.950 55.950 322.050 58.050 ;
        RECT 322.950 55.950 325.050 58.050 ;
        RECT 167.100 42.600 168.900 45.600 ;
        RECT 170.100 42.600 171.900 45.600 ;
        RECT 167.100 42.000 168.300 42.600 ;
        RECT 173.100 42.000 174.900 48.000 ;
        RECT 176.100 42.600 177.900 48.600 ;
        RECT 194.100 42.000 195.900 51.600 ;
        RECT 200.700 51.000 204.000 52.200 ;
        RECT 200.700 42.600 202.500 51.000 ;
        RECT 220.800 49.500 222.900 50.700 ;
        RECT 224.100 50.100 227.100 52.200 ;
        RECT 228.000 53.400 229.800 55.200 ;
        RECT 232.800 54.150 234.600 55.950 ;
        RECT 248.100 54.150 249.900 55.950 ;
        RECT 228.000 51.300 230.100 53.400 ;
        RECT 251.100 51.600 252.300 55.950 ;
        RECT 254.100 54.150 255.900 55.950 ;
        RECT 228.000 50.400 234.300 51.300 ;
        RECT 218.100 48.600 222.900 49.500 ;
        RECT 225.900 48.600 227.100 50.100 ;
        RECT 233.100 48.600 234.300 50.400 ;
        RECT 248.700 50.700 252.300 51.600 ;
        RECT 248.700 48.600 249.900 50.700 ;
        RECT 218.100 42.600 219.900 48.600 ;
        RECT 221.100 42.000 222.900 47.700 ;
        RECT 225.600 42.600 227.400 48.600 ;
        RECT 230.100 42.000 231.900 47.700 ;
        RECT 233.100 42.600 234.900 48.600 ;
        RECT 248.100 42.600 249.900 48.600 ;
        RECT 251.100 47.700 258.900 49.050 ;
        RECT 251.100 42.600 252.900 47.700 ;
        RECT 254.100 42.000 255.900 46.800 ;
        RECT 257.100 42.600 258.900 47.700 ;
        RECT 275.100 45.600 276.300 55.950 ;
        RECT 294.000 52.200 294.900 55.950 ;
        RECT 296.100 54.150 297.900 55.950 ;
        RECT 302.100 54.150 303.900 55.950 ;
        RECT 317.100 54.150 318.900 55.950 ;
        RECT 294.000 51.000 297.300 52.200 ;
        RECT 272.100 42.000 273.900 45.600 ;
        RECT 275.100 42.600 276.900 45.600 ;
        RECT 295.500 42.600 297.300 51.000 ;
        RECT 302.100 42.000 303.900 51.600 ;
        RECT 320.700 50.700 321.900 55.950 ;
        RECT 322.950 54.150 324.750 55.950 ;
        RECT 317.700 49.800 321.900 50.700 ;
        RECT 317.700 42.600 319.500 49.800 ;
        RECT 326.550 48.600 327.450 63.300 ;
        RECT 336.450 63.000 338.250 63.300 ;
        RECT 328.950 55.950 331.050 58.050 ;
        RECT 338.100 56.400 340.200 58.050 ;
        RECT 328.950 53.400 330.750 55.950 ;
        RECT 332.100 55.200 340.200 56.400 ;
        RECT 332.100 54.600 333.900 55.200 ;
        RECT 335.100 53.400 336.900 54.000 ;
        RECT 328.950 52.200 336.900 53.400 ;
        RECT 346.950 52.200 347.850 64.800 ;
        RECT 350.550 62.100 352.650 62.700 ;
        RECT 356.550 62.100 358.350 62.550 ;
        RECT 350.550 60.900 358.350 62.100 ;
        RECT 350.550 60.600 352.650 60.900 ;
        RECT 356.550 60.750 358.350 60.900 ;
        RECT 359.250 58.050 360.450 65.400 ;
        RECT 377.700 58.050 378.900 71.400 ;
        RECT 395.100 66.300 396.900 77.400 ;
        RECT 398.100 67.500 399.900 78.000 ;
        RECT 402.600 66.300 404.400 77.400 ;
        RECT 406.800 67.500 408.900 78.000 ;
        RECT 410.100 66.600 411.900 77.400 ;
        RECT 425.700 71.400 427.500 78.000 ;
        RECT 426.000 68.100 427.800 69.900 ;
        RECT 428.700 66.900 430.500 77.400 ;
        RECT 395.100 65.100 399.900 66.300 ;
        RECT 402.600 65.400 405.900 66.300 ;
        RECT 397.800 64.200 399.900 65.100 ;
        RECT 397.800 63.300 403.200 64.200 ;
        RECT 401.400 61.500 403.200 63.300 ;
        RECT 404.700 61.050 405.900 65.400 ;
        RECT 406.800 65.400 411.900 66.600 ;
        RECT 428.100 65.400 430.500 66.900 ;
        RECT 433.800 65.400 435.600 78.000 ;
        RECT 449.100 71.400 450.900 78.000 ;
        RECT 452.100 71.400 453.900 77.400 ;
        RECT 455.100 71.400 456.900 78.000 ;
        RECT 473.100 71.400 474.900 78.000 ;
        RECT 476.100 71.400 477.900 77.400 ;
        RECT 479.100 71.400 480.900 78.000 ;
        RECT 494.100 71.400 495.900 78.000 ;
        RECT 497.100 71.400 498.900 77.400 ;
        RECT 500.100 71.400 501.900 78.000 ;
        RECT 518.100 71.400 519.900 78.000 ;
        RECT 521.100 71.400 522.900 77.400 ;
        RECT 406.800 64.500 408.900 65.400 ;
        RECT 404.100 60.300 406.200 61.050 ;
        RECT 399.900 58.200 401.700 60.000 ;
        RECT 403.200 58.950 406.200 60.300 ;
        RECT 355.950 57.750 360.450 58.050 ;
        RECT 354.150 55.950 360.450 57.750 ;
        RECT 373.950 55.950 376.050 58.050 ;
        RECT 376.950 55.950 379.050 58.050 ;
        RECT 379.950 55.950 382.050 58.050 ;
        RECT 335.850 51.000 347.850 52.200 ;
        RECT 335.850 49.200 336.900 51.000 ;
        RECT 346.050 50.400 347.850 51.000 ;
        RECT 322.800 42.000 324.600 48.600 ;
        RECT 326.550 46.800 328.950 48.600 ;
        RECT 327.150 42.600 328.950 46.800 ;
        RECT 330.150 42.000 331.950 48.600 ;
        RECT 332.850 46.200 334.950 47.700 ;
        RECT 335.850 47.400 337.650 49.200 ;
        RECT 359.250 48.600 360.450 55.950 ;
        RECT 374.100 54.150 375.900 55.950 ;
        RECT 377.700 50.700 378.900 55.950 ;
        RECT 379.950 54.150 381.750 55.950 ;
        RECT 395.100 55.800 397.200 58.050 ;
        RECT 399.900 56.100 402.000 58.200 ;
        RECT 395.400 55.200 397.200 55.800 ;
        RECT 395.400 54.000 402.000 55.200 ;
        RECT 399.900 53.100 402.000 54.000 ;
        RECT 397.500 51.000 399.600 51.600 ;
        RECT 400.500 51.300 402.300 53.100 ;
        RECT 403.200 52.200 404.100 58.950 ;
        RECT 409.800 58.050 411.600 59.850 ;
        RECT 428.100 58.050 429.300 65.400 ;
        RECT 434.100 58.050 435.900 59.850 ;
        RECT 452.700 58.050 453.900 71.400 ;
        RECT 476.700 58.050 477.900 71.400 ;
        RECT 497.700 58.050 498.900 71.400 ;
        RECT 405.000 56.100 406.800 57.900 ;
        RECT 405.000 54.000 407.100 56.100 ;
        RECT 409.800 55.950 411.900 58.050 ;
        RECT 424.950 55.950 427.050 58.050 ;
        RECT 427.950 55.950 430.050 58.050 ;
        RECT 430.950 55.950 433.050 58.050 ;
        RECT 433.950 55.950 436.050 58.050 ;
        RECT 448.950 55.950 451.050 58.050 ;
        RECT 451.950 55.950 454.050 58.050 ;
        RECT 454.950 55.950 457.050 58.050 ;
        RECT 472.950 55.950 475.050 58.050 ;
        RECT 475.950 55.950 478.050 58.050 ;
        RECT 478.950 55.950 481.050 58.050 ;
        RECT 493.950 55.950 496.050 58.050 ;
        RECT 496.950 55.950 499.050 58.050 ;
        RECT 499.950 55.950 502.050 58.050 ;
        RECT 518.100 55.950 520.200 58.050 ;
        RECT 425.100 54.150 426.900 55.950 ;
        RECT 338.850 47.550 340.650 48.300 ;
        RECT 338.850 46.500 343.800 47.550 ;
        RECT 332.850 45.600 336.750 46.200 ;
        RECT 342.750 45.600 343.800 46.500 ;
        RECT 350.250 45.600 352.650 47.700 ;
        RECT 333.150 44.700 336.750 45.600 ;
        RECT 334.950 42.600 336.750 44.700 ;
        RECT 339.450 42.000 341.250 45.600 ;
        RECT 342.750 42.600 344.550 45.600 ;
        RECT 345.750 42.000 347.550 45.600 ;
        RECT 350.250 42.600 352.050 45.600 ;
        RECT 355.350 42.000 357.150 48.600 ;
        RECT 358.650 42.600 360.450 48.600 ;
        RECT 374.700 49.800 378.900 50.700 ;
        RECT 374.700 42.600 376.500 49.800 ;
        RECT 395.100 49.500 399.600 51.000 ;
        RECT 403.200 50.100 406.200 52.200 ;
        RECT 395.100 48.600 396.600 49.500 ;
        RECT 379.800 42.000 381.600 48.600 ;
        RECT 395.100 42.600 396.900 48.600 ;
        RECT 403.200 48.000 404.100 50.100 ;
        RECT 407.400 49.500 409.500 51.900 ;
        RECT 428.100 51.600 429.300 55.950 ;
        RECT 431.100 54.150 432.900 55.950 ;
        RECT 449.100 54.150 450.900 55.950 ;
        RECT 425.700 50.700 429.300 51.600 ;
        RECT 452.700 50.700 453.900 55.950 ;
        RECT 454.950 54.150 456.750 55.950 ;
        RECT 473.100 54.150 474.900 55.950 ;
        RECT 476.700 50.700 477.900 55.950 ;
        RECT 478.950 54.150 480.750 55.950 ;
        RECT 494.100 54.150 495.900 55.950 ;
        RECT 497.700 50.700 498.900 55.950 ;
        RECT 499.950 54.150 501.750 55.950 ;
        RECT 518.250 54.150 520.050 55.950 ;
        RECT 521.100 51.300 522.000 71.400 ;
        RECT 524.100 66.000 525.900 78.000 ;
        RECT 527.100 65.400 528.900 77.400 ;
        RECT 542.100 71.400 543.900 78.000 ;
        RECT 545.100 71.400 546.900 77.400 ;
        RECT 548.100 71.400 549.900 78.000 ;
        RECT 563.100 71.400 564.900 78.000 ;
        RECT 566.100 71.400 567.900 77.400 ;
        RECT 569.100 72.000 570.900 78.000 ;
        RECT 523.200 58.050 525.000 59.850 ;
        RECT 527.400 58.050 528.300 65.400 ;
        RECT 545.700 58.050 546.900 71.400 ;
        RECT 566.400 71.100 567.900 71.400 ;
        RECT 572.100 71.400 573.900 77.400 ;
        RECT 590.100 71.400 591.900 78.000 ;
        RECT 593.100 71.400 594.900 77.400 ;
        RECT 596.100 71.400 597.900 78.000 ;
        RECT 572.100 71.100 573.000 71.400 ;
        RECT 566.400 70.200 573.000 71.100 ;
        RECT 566.100 58.050 567.900 59.850 ;
        RECT 572.100 58.050 573.000 70.200 ;
        RECT 593.700 58.050 594.900 71.400 ;
        RECT 611.100 65.400 612.900 78.000 ;
        RECT 616.200 66.600 618.000 77.400 ;
        RECT 614.400 65.400 618.000 66.600 ;
        RECT 633.000 66.600 634.800 77.400 ;
        RECT 633.000 65.400 636.600 66.600 ;
        RECT 638.100 65.400 639.900 78.000 ;
        RECT 653.100 71.400 654.900 78.000 ;
        RECT 656.100 71.400 657.900 77.400 ;
        RECT 659.100 72.000 660.900 78.000 ;
        RECT 656.400 71.100 657.900 71.400 ;
        RECT 662.100 71.400 663.900 77.400 ;
        RECT 662.100 71.100 663.000 71.400 ;
        RECT 656.400 70.200 663.000 71.100 ;
        RECT 652.950 66.450 655.050 67.050 ;
        RECT 658.950 66.450 661.050 67.050 ;
        RECT 652.950 65.550 661.050 66.450 ;
        RECT 611.250 58.050 613.050 59.850 ;
        RECT 614.400 58.050 615.300 65.400 ;
        RECT 617.100 58.050 618.900 59.850 ;
        RECT 632.100 58.050 633.900 59.850 ;
        RECT 635.700 58.050 636.600 65.400 ;
        RECT 652.950 64.950 655.050 65.550 ;
        RECT 658.950 64.950 661.050 65.550 ;
        RECT 637.950 58.050 639.750 59.850 ;
        RECT 656.100 58.050 657.900 59.850 ;
        RECT 662.100 58.050 663.000 70.200 ;
        RECT 677.100 66.300 678.900 77.400 ;
        RECT 680.100 67.200 681.900 78.000 ;
        RECT 683.100 66.300 684.900 77.400 ;
        RECT 677.100 65.400 684.900 66.300 ;
        RECT 686.100 65.400 687.900 77.400 ;
        RECT 701.100 71.400 702.900 78.000 ;
        RECT 704.100 71.400 705.900 77.400 ;
        RECT 707.100 72.000 708.900 78.000 ;
        RECT 704.400 71.100 705.900 71.400 ;
        RECT 710.100 71.400 711.900 77.400 ;
        RECT 725.700 71.400 727.500 78.000 ;
        RECT 710.100 71.100 711.000 71.400 ;
        RECT 704.400 70.200 711.000 71.100 ;
        RECT 680.250 58.050 682.050 59.850 ;
        RECT 686.700 58.050 687.600 65.400 ;
        RECT 704.100 58.050 705.900 59.850 ;
        RECT 710.100 58.050 711.000 70.200 ;
        RECT 726.000 68.100 727.800 69.900 ;
        RECT 728.700 66.900 730.500 77.400 ;
        RECT 728.100 65.400 730.500 66.900 ;
        RECT 733.800 65.400 735.600 78.000 ;
        RECT 749.400 65.400 751.200 78.000 ;
        RECT 754.500 66.900 756.300 77.400 ;
        RECT 757.500 71.400 759.300 78.000 ;
        RECT 773.700 71.400 775.500 78.000 ;
        RECT 757.200 68.100 759.000 69.900 ;
        RECT 774.000 68.100 775.800 69.900 ;
        RECT 776.700 66.900 778.500 77.400 ;
        RECT 754.500 65.400 756.900 66.900 ;
        RECT 728.100 58.050 729.300 65.400 ;
        RECT 734.100 58.050 735.900 59.850 ;
        RECT 749.100 58.050 750.900 59.850 ;
        RECT 755.700 58.050 756.900 65.400 ;
        RECT 776.100 65.400 778.500 66.900 ;
        RECT 781.800 65.400 783.600 78.000 ;
        RECT 797.700 71.400 799.500 78.000 ;
        RECT 798.000 68.100 799.800 69.900 ;
        RECT 800.700 66.900 802.500 77.400 ;
        RECT 800.100 65.400 802.500 66.900 ;
        RECT 805.800 65.400 807.600 78.000 ;
        RECT 824.100 65.400 825.900 77.400 ;
        RECT 827.100 66.300 828.900 77.400 ;
        RECT 830.100 67.200 831.900 78.000 ;
        RECT 833.100 66.300 834.900 77.400 ;
        RECT 848.100 71.400 849.900 77.400 ;
        RECT 851.100 72.000 852.900 78.000 ;
        RECT 827.100 65.400 834.900 66.300 ;
        RECT 849.000 71.100 849.900 71.400 ;
        RECT 854.100 71.400 855.900 77.400 ;
        RECT 857.100 71.400 858.900 78.000 ;
        RECT 875.100 71.400 876.900 78.000 ;
        RECT 878.100 71.400 879.900 77.400 ;
        RECT 881.100 71.400 882.900 78.000 ;
        RECT 854.100 71.100 855.600 71.400 ;
        RECT 849.000 70.200 855.600 71.100 ;
        RECT 776.100 58.050 777.300 65.400 ;
        RECT 782.100 58.050 783.900 59.850 ;
        RECT 800.100 58.050 801.300 65.400 ;
        RECT 806.100 58.050 807.900 59.850 ;
        RECT 824.400 58.050 825.300 65.400 ;
        RECT 829.950 58.050 831.750 59.850 ;
        RECT 849.000 58.050 849.900 70.200 ;
        RECT 854.100 58.050 855.900 59.850 ;
        RECT 878.700 58.050 879.900 71.400 ;
        RECT 523.500 55.950 525.600 58.050 ;
        RECT 526.800 55.950 528.900 58.050 ;
        RECT 541.950 55.950 544.050 58.050 ;
        RECT 544.950 55.950 547.050 58.050 ;
        RECT 547.950 55.950 550.050 58.050 ;
        RECT 562.950 55.950 565.050 58.050 ;
        RECT 565.950 55.950 568.050 58.050 ;
        RECT 568.950 55.950 571.050 58.050 ;
        RECT 571.950 55.950 574.050 58.050 ;
        RECT 589.950 55.950 592.050 58.050 ;
        RECT 592.950 55.950 595.050 58.050 ;
        RECT 595.950 55.950 598.050 58.050 ;
        RECT 610.950 55.950 613.050 58.050 ;
        RECT 613.950 55.950 616.050 58.050 ;
        RECT 616.950 55.950 619.050 58.050 ;
        RECT 631.950 55.950 634.050 58.050 ;
        RECT 634.950 55.950 637.050 58.050 ;
        RECT 637.950 55.950 640.050 58.050 ;
        RECT 652.950 55.950 655.050 58.050 ;
        RECT 655.950 55.950 658.050 58.050 ;
        RECT 658.950 55.950 661.050 58.050 ;
        RECT 661.950 55.950 664.050 58.050 ;
        RECT 676.950 55.950 679.050 58.050 ;
        RECT 679.950 55.950 682.050 58.050 ;
        RECT 682.950 55.950 685.050 58.050 ;
        RECT 685.950 55.950 688.050 58.050 ;
        RECT 700.950 55.950 703.050 58.050 ;
        RECT 703.950 55.950 706.050 58.050 ;
        RECT 706.950 55.950 709.050 58.050 ;
        RECT 709.950 55.950 712.050 58.050 ;
        RECT 724.950 55.950 727.050 58.050 ;
        RECT 727.950 55.950 730.050 58.050 ;
        RECT 730.950 55.950 733.050 58.050 ;
        RECT 733.950 55.950 736.050 58.050 ;
        RECT 748.950 55.950 751.050 58.050 ;
        RECT 751.950 55.950 754.050 58.050 ;
        RECT 754.950 55.950 757.050 58.050 ;
        RECT 757.950 55.950 760.050 58.050 ;
        RECT 772.950 55.950 775.050 58.050 ;
        RECT 775.950 55.950 778.050 58.050 ;
        RECT 778.950 55.950 781.050 58.050 ;
        RECT 781.950 55.950 784.050 58.050 ;
        RECT 796.950 55.950 799.050 58.050 ;
        RECT 799.950 55.950 802.050 58.050 ;
        RECT 802.950 55.950 805.050 58.050 ;
        RECT 805.950 55.950 808.050 58.050 ;
        RECT 823.950 55.950 826.050 58.050 ;
        RECT 826.950 55.950 829.050 58.050 ;
        RECT 829.950 55.950 832.050 58.050 ;
        RECT 832.950 55.950 835.050 58.050 ;
        RECT 847.950 55.950 850.050 58.050 ;
        RECT 850.950 55.950 853.050 58.050 ;
        RECT 853.950 55.950 856.050 58.050 ;
        RECT 856.950 55.950 859.050 58.050 ;
        RECT 874.950 55.950 877.050 58.050 ;
        RECT 877.950 55.950 880.050 58.050 ;
        RECT 880.950 55.950 883.050 58.050 ;
        RECT 407.400 48.600 411.900 49.500 ;
        RECT 425.700 48.600 426.900 50.700 ;
        RECT 449.700 49.800 453.900 50.700 ;
        RECT 473.700 49.800 477.900 50.700 ;
        RECT 494.700 49.800 498.900 50.700 ;
        RECT 518.100 50.400 526.500 51.300 ;
        RECT 398.100 42.000 399.900 47.700 ;
        RECT 402.300 42.600 404.100 48.000 ;
        RECT 406.800 42.000 408.600 47.700 ;
        RECT 410.100 42.600 411.900 48.600 ;
        RECT 425.100 42.600 426.900 48.600 ;
        RECT 428.100 47.700 435.900 49.050 ;
        RECT 428.100 42.600 429.900 47.700 ;
        RECT 431.100 42.000 432.900 46.800 ;
        RECT 434.100 42.600 435.900 47.700 ;
        RECT 449.700 42.600 451.500 49.800 ;
        RECT 454.800 42.000 456.600 48.600 ;
        RECT 473.700 42.600 475.500 49.800 ;
        RECT 478.800 42.000 480.600 48.600 ;
        RECT 494.700 42.600 496.500 49.800 ;
        RECT 499.800 42.000 501.600 48.600 ;
        RECT 518.100 42.600 519.900 50.400 ;
        RECT 524.700 49.500 526.500 50.400 ;
        RECT 527.400 48.600 528.300 55.950 ;
        RECT 542.100 54.150 543.900 55.950 ;
        RECT 545.700 50.700 546.900 55.950 ;
        RECT 547.950 54.150 549.750 55.950 ;
        RECT 563.100 54.150 564.900 55.950 ;
        RECT 569.100 54.150 570.900 55.950 ;
        RECT 572.100 52.200 573.000 55.950 ;
        RECT 590.100 54.150 591.900 55.950 ;
        RECT 522.600 42.000 524.400 48.600 ;
        RECT 525.600 46.800 528.300 48.600 ;
        RECT 542.700 49.800 546.900 50.700 ;
        RECT 525.600 42.600 527.400 46.800 ;
        RECT 542.700 42.600 544.500 49.800 ;
        RECT 547.800 42.000 549.600 48.600 ;
        RECT 563.100 42.000 564.900 51.600 ;
        RECT 569.700 51.000 573.000 52.200 ;
        RECT 569.700 42.600 571.500 51.000 ;
        RECT 593.700 50.700 594.900 55.950 ;
        RECT 595.950 54.150 597.750 55.950 ;
        RECT 590.700 49.800 594.900 50.700 ;
        RECT 590.700 42.600 592.500 49.800 ;
        RECT 595.800 42.000 597.600 48.600 ;
        RECT 614.400 45.600 615.300 55.950 ;
        RECT 635.700 45.600 636.600 55.950 ;
        RECT 653.100 54.150 654.900 55.950 ;
        RECT 659.100 54.150 660.900 55.950 ;
        RECT 662.100 52.200 663.000 55.950 ;
        RECT 677.100 54.150 678.900 55.950 ;
        RECT 683.250 54.150 685.050 55.950 ;
        RECT 611.100 42.000 612.900 45.600 ;
        RECT 614.100 42.600 615.900 45.600 ;
        RECT 617.100 42.000 618.900 45.600 ;
        RECT 632.100 42.000 633.900 45.600 ;
        RECT 635.100 42.600 636.900 45.600 ;
        RECT 638.100 42.000 639.900 45.600 ;
        RECT 653.100 42.000 654.900 51.600 ;
        RECT 659.700 51.000 663.000 52.200 ;
        RECT 670.950 51.450 673.050 52.050 ;
        RECT 679.950 51.450 682.050 52.050 ;
        RECT 659.700 42.600 661.500 51.000 ;
        RECT 670.950 50.550 682.050 51.450 ;
        RECT 670.950 49.950 673.050 50.550 ;
        RECT 679.950 49.950 682.050 50.550 ;
        RECT 686.700 48.600 687.600 55.950 ;
        RECT 701.100 54.150 702.900 55.950 ;
        RECT 707.100 54.150 708.900 55.950 ;
        RECT 710.100 52.200 711.000 55.950 ;
        RECT 725.100 54.150 726.900 55.950 ;
        RECT 678.000 42.000 679.800 48.600 ;
        RECT 682.500 47.400 687.600 48.600 ;
        RECT 682.500 42.600 684.300 47.400 ;
        RECT 685.500 42.000 687.300 45.600 ;
        RECT 701.100 42.000 702.900 51.600 ;
        RECT 707.700 51.000 711.000 52.200 ;
        RECT 728.100 51.600 729.300 55.950 ;
        RECT 731.100 54.150 732.900 55.950 ;
        RECT 752.100 54.150 753.900 55.950 ;
        RECT 707.700 42.600 709.500 51.000 ;
        RECT 725.700 50.700 729.300 51.600 ;
        RECT 755.700 51.600 756.900 55.950 ;
        RECT 758.100 54.150 759.900 55.950 ;
        RECT 773.100 54.150 774.900 55.950 ;
        RECT 776.100 51.600 777.300 55.950 ;
        RECT 779.100 54.150 780.900 55.950 ;
        RECT 797.100 54.150 798.900 55.950 ;
        RECT 800.100 51.600 801.300 55.950 ;
        RECT 803.100 54.150 804.900 55.950 ;
        RECT 755.700 50.700 759.300 51.600 ;
        RECT 725.700 48.600 726.900 50.700 ;
        RECT 725.100 42.600 726.900 48.600 ;
        RECT 728.100 47.700 735.900 49.050 ;
        RECT 728.100 42.600 729.900 47.700 ;
        RECT 731.100 42.000 732.900 46.800 ;
        RECT 734.100 42.600 735.900 47.700 ;
        RECT 749.100 47.700 756.900 49.050 ;
        RECT 749.100 42.600 750.900 47.700 ;
        RECT 752.100 42.000 753.900 46.800 ;
        RECT 755.100 42.600 756.900 47.700 ;
        RECT 758.100 48.600 759.300 50.700 ;
        RECT 773.700 50.700 777.300 51.600 ;
        RECT 797.700 50.700 801.300 51.600 ;
        RECT 773.700 48.600 774.900 50.700 ;
        RECT 758.100 42.600 759.900 48.600 ;
        RECT 773.100 42.600 774.900 48.600 ;
        RECT 776.100 47.700 783.900 49.050 ;
        RECT 797.700 48.600 798.900 50.700 ;
        RECT 776.100 42.600 777.900 47.700 ;
        RECT 779.100 42.000 780.900 46.800 ;
        RECT 782.100 42.600 783.900 47.700 ;
        RECT 797.100 42.600 798.900 48.600 ;
        RECT 800.100 47.700 807.900 49.050 ;
        RECT 800.100 42.600 801.900 47.700 ;
        RECT 803.100 42.000 804.900 46.800 ;
        RECT 806.100 42.600 807.900 47.700 ;
        RECT 824.400 48.600 825.300 55.950 ;
        RECT 826.950 54.150 828.750 55.950 ;
        RECT 833.100 54.150 834.900 55.950 ;
        RECT 849.000 52.200 849.900 55.950 ;
        RECT 851.100 54.150 852.900 55.950 ;
        RECT 857.100 54.150 858.900 55.950 ;
        RECT 875.100 54.150 876.900 55.950 ;
        RECT 849.000 51.000 852.300 52.200 ;
        RECT 824.400 47.400 829.500 48.600 ;
        RECT 824.700 42.000 826.500 45.600 ;
        RECT 827.700 42.600 829.500 47.400 ;
        RECT 832.200 42.000 834.000 48.600 ;
        RECT 850.500 42.600 852.300 51.000 ;
        RECT 857.100 42.000 858.900 51.600 ;
        RECT 878.700 50.700 879.900 55.950 ;
        RECT 880.950 54.150 882.750 55.950 ;
        RECT 875.700 49.800 879.900 50.700 ;
        RECT 875.700 42.600 877.500 49.800 ;
        RECT 880.800 42.000 882.600 48.600 ;
        RECT 17.100 35.400 18.900 39.000 ;
        RECT 20.100 35.400 21.900 38.400 ;
        RECT 20.100 25.050 21.300 35.400 ;
        RECT 35.100 32.400 36.900 38.400 ;
        RECT 38.100 33.000 39.900 39.000 ;
        RECT 44.700 38.400 45.900 39.000 ;
        RECT 41.100 35.400 42.900 38.400 ;
        RECT 44.100 35.400 45.900 38.400 ;
        RECT 35.100 25.050 36.000 32.400 ;
        RECT 41.700 31.200 42.600 35.400 ;
        RECT 37.200 30.300 42.600 31.200 ;
        RECT 59.700 31.200 61.500 38.400 ;
        RECT 64.800 32.400 66.600 39.000 ;
        RECT 80.400 32.400 82.200 39.000 ;
        RECT 85.500 31.200 87.300 38.400 ;
        RECT 59.700 30.300 63.900 31.200 ;
        RECT 37.200 29.400 39.300 30.300 ;
        RECT 16.950 22.950 19.050 25.050 ;
        RECT 19.950 22.950 22.050 25.050 ;
        RECT 35.100 22.950 37.200 25.050 ;
        RECT 17.100 21.150 18.900 22.950 ;
        RECT 20.100 9.600 21.300 22.950 ;
        RECT 36.000 15.600 37.200 22.950 ;
        RECT 38.400 18.900 39.300 29.400 ;
        RECT 43.800 25.050 45.600 26.850 ;
        RECT 59.100 25.050 60.900 26.850 ;
        RECT 62.700 25.050 63.900 30.300 ;
        RECT 70.950 30.450 73.050 31.050 ;
        RECT 79.950 30.450 82.050 31.050 ;
        RECT 70.950 29.550 82.050 30.450 ;
        RECT 70.950 28.950 73.050 29.550 ;
        RECT 79.950 28.950 82.050 29.550 ;
        RECT 83.100 30.300 87.300 31.200 ;
        RECT 101.700 31.200 103.500 38.400 ;
        RECT 106.800 32.400 108.600 39.000 ;
        RECT 122.100 35.400 123.900 39.000 ;
        RECT 125.100 35.400 126.900 38.400 ;
        RECT 128.100 35.400 129.900 39.000 ;
        RECT 143.100 35.400 144.900 38.400 ;
        RECT 146.100 35.400 147.900 39.000 ;
        RECT 101.700 30.300 105.900 31.200 ;
        RECT 64.950 25.050 66.750 26.850 ;
        RECT 80.250 25.050 82.050 26.850 ;
        RECT 83.100 25.050 84.300 30.300 ;
        RECT 86.100 25.050 87.900 26.850 ;
        RECT 101.100 25.050 102.900 26.850 ;
        RECT 104.700 25.050 105.900 30.300 ;
        RECT 106.950 25.050 108.750 26.850 ;
        RECT 125.700 25.050 126.600 35.400 ;
        RECT 143.700 25.050 144.900 35.400 ;
        RECT 161.100 33.300 162.900 38.400 ;
        RECT 164.100 34.200 165.900 39.000 ;
        RECT 167.100 33.300 168.900 38.400 ;
        RECT 161.100 31.950 168.900 33.300 ;
        RECT 170.100 32.400 171.900 38.400 ;
        RECT 185.100 35.400 186.900 38.400 ;
        RECT 188.100 35.400 189.900 39.000 ;
        RECT 170.100 30.300 171.300 32.400 ;
        RECT 167.700 29.400 171.300 30.300 ;
        RECT 164.100 25.050 165.900 26.850 ;
        RECT 167.700 25.050 168.900 29.400 ;
        RECT 170.100 25.050 171.900 26.850 ;
        RECT 185.700 25.050 186.900 35.400 ;
        RECT 207.000 32.400 208.800 39.000 ;
        RECT 211.500 33.600 213.300 38.400 ;
        RECT 214.500 35.400 216.300 39.000 ;
        RECT 211.500 32.400 216.600 33.600 ;
        RECT 206.100 25.050 207.900 26.850 ;
        RECT 212.250 25.050 214.050 26.850 ;
        RECT 215.700 25.050 216.600 32.400 ;
        RECT 233.100 32.400 234.900 38.400 ;
        RECT 236.100 33.300 237.900 39.000 ;
        RECT 240.600 32.400 242.400 38.400 ;
        RECT 245.100 33.300 246.900 39.000 ;
        RECT 248.100 32.400 249.900 38.400 ;
        RECT 252.150 34.200 253.950 38.400 ;
        RECT 251.550 32.400 253.950 34.200 ;
        RECT 255.150 32.400 256.950 39.000 ;
        RECT 259.950 36.300 261.750 38.400 ;
        RECT 258.150 35.400 261.750 36.300 ;
        RECT 264.450 35.400 266.250 39.000 ;
        RECT 267.750 35.400 269.550 38.400 ;
        RECT 270.750 35.400 272.550 39.000 ;
        RECT 275.250 35.400 277.050 38.400 ;
        RECT 257.850 34.800 261.750 35.400 ;
        RECT 257.850 33.300 259.950 34.800 ;
        RECT 267.750 34.500 268.800 35.400 ;
        RECT 233.100 31.500 237.900 32.400 ;
        RECT 235.800 30.300 237.900 31.500 ;
        RECT 240.900 30.900 242.100 32.400 ;
        RECT 239.100 28.800 242.100 30.900 ;
        RECT 248.100 30.600 249.300 32.400 ;
        RECT 223.950 27.450 226.050 28.050 ;
        RECT 229.950 27.450 232.050 28.050 ;
        RECT 223.950 26.550 232.050 27.450 ;
        RECT 223.950 25.950 226.050 26.550 ;
        RECT 229.950 25.950 232.050 26.550 ;
        RECT 237.900 25.800 240.000 27.900 ;
        RECT 40.500 22.950 42.600 25.050 ;
        RECT 43.800 22.950 45.900 25.050 ;
        RECT 58.950 22.950 61.050 25.050 ;
        RECT 61.950 22.950 64.050 25.050 ;
        RECT 64.950 22.950 67.050 25.050 ;
        RECT 79.950 22.950 82.050 25.050 ;
        RECT 82.950 22.950 85.050 25.050 ;
        RECT 85.950 22.950 88.050 25.050 ;
        RECT 100.950 22.950 103.050 25.050 ;
        RECT 103.950 22.950 106.050 25.050 ;
        RECT 106.950 22.950 109.050 25.050 ;
        RECT 121.950 22.950 124.050 25.050 ;
        RECT 124.950 22.950 127.050 25.050 ;
        RECT 127.950 22.950 130.050 25.050 ;
        RECT 142.950 22.950 145.050 25.050 ;
        RECT 145.950 22.950 148.050 25.050 ;
        RECT 160.950 22.950 163.050 25.050 ;
        RECT 163.950 22.950 166.050 25.050 ;
        RECT 166.950 22.950 169.050 25.050 ;
        RECT 169.950 22.950 172.050 25.050 ;
        RECT 184.950 22.950 187.050 25.050 ;
        RECT 187.950 22.950 190.050 25.050 ;
        RECT 205.950 22.950 208.050 25.050 ;
        RECT 208.950 22.950 211.050 25.050 ;
        RECT 211.950 22.950 214.050 25.050 ;
        RECT 214.950 22.950 217.050 25.050 ;
        RECT 233.100 22.950 235.200 25.050 ;
        RECT 237.900 24.000 239.700 25.800 ;
        RECT 240.900 23.100 242.100 28.800 ;
        RECT 243.000 29.700 249.300 30.600 ;
        RECT 243.000 27.600 245.100 29.700 ;
        RECT 243.000 25.800 244.800 27.600 ;
        RECT 247.800 25.050 249.600 26.850 ;
        RECT 247.800 24.300 249.900 25.050 ;
        RECT 40.200 21.150 42.000 22.950 ;
        RECT 38.100 18.300 39.900 18.900 ;
        RECT 38.100 17.100 45.900 18.300 ;
        RECT 44.700 15.600 45.900 17.100 ;
        RECT 36.000 14.100 38.400 15.600 ;
        RECT 17.100 3.000 18.900 9.600 ;
        RECT 20.100 3.600 21.900 9.600 ;
        RECT 36.600 3.600 38.400 14.100 ;
        RECT 39.600 3.000 41.400 15.600 ;
        RECT 44.100 3.600 45.900 15.600 ;
        RECT 62.700 9.600 63.900 22.950 ;
        RECT 83.100 9.600 84.300 22.950 ;
        RECT 104.700 9.600 105.900 22.950 ;
        RECT 122.100 21.150 123.900 22.950 ;
        RECT 125.700 15.600 126.600 22.950 ;
        RECT 127.950 21.150 129.750 22.950 ;
        RECT 123.000 14.400 126.600 15.600 ;
        RECT 59.100 3.000 60.900 9.600 ;
        RECT 62.100 3.600 63.900 9.600 ;
        RECT 65.100 3.000 66.900 9.600 ;
        RECT 80.100 3.000 81.900 9.600 ;
        RECT 83.100 3.600 84.900 9.600 ;
        RECT 86.100 3.000 87.900 9.600 ;
        RECT 101.100 3.000 102.900 9.600 ;
        RECT 104.100 3.600 105.900 9.600 ;
        RECT 107.100 3.000 108.900 9.600 ;
        RECT 123.000 3.600 124.800 14.400 ;
        RECT 128.100 3.000 129.900 15.600 ;
        RECT 143.700 9.600 144.900 22.950 ;
        RECT 146.100 21.150 147.900 22.950 ;
        RECT 161.100 21.150 162.900 22.950 ;
        RECT 167.700 15.600 168.900 22.950 ;
        RECT 143.100 3.600 144.900 9.600 ;
        RECT 146.100 3.000 147.900 9.600 ;
        RECT 161.400 3.000 163.200 15.600 ;
        RECT 166.500 14.100 168.900 15.600 ;
        RECT 166.500 3.600 168.300 14.100 ;
        RECT 169.200 11.100 171.000 12.900 ;
        RECT 185.700 9.600 186.900 22.950 ;
        RECT 188.100 21.150 189.900 22.950 ;
        RECT 209.250 21.150 211.050 22.950 ;
        RECT 193.950 18.450 196.050 19.050 ;
        RECT 211.950 18.450 214.050 19.050 ;
        RECT 193.950 17.550 214.050 18.450 ;
        RECT 193.950 16.950 196.050 17.550 ;
        RECT 211.950 16.950 214.050 17.550 ;
        RECT 215.700 15.600 216.600 22.950 ;
        RECT 233.400 21.150 235.200 22.950 ;
        RECT 239.700 22.200 242.100 23.100 ;
        RECT 243.000 22.950 249.900 24.300 ;
        RECT 243.000 22.500 244.800 22.950 ;
        RECT 239.700 22.050 241.200 22.200 ;
        RECT 239.100 19.950 241.200 22.050 ;
        RECT 240.300 18.000 241.200 19.950 ;
        RECT 242.100 19.500 246.000 21.300 ;
        RECT 242.100 19.200 244.200 19.500 ;
        RECT 240.300 16.950 241.800 18.000 ;
        RECT 251.550 17.700 252.450 32.400 ;
        RECT 260.850 31.800 262.650 33.600 ;
        RECT 263.850 33.450 268.800 34.500 ;
        RECT 263.850 32.700 265.650 33.450 ;
        RECT 275.250 33.300 277.650 35.400 ;
        RECT 280.350 32.400 282.150 39.000 ;
        RECT 283.650 32.400 285.450 38.400 ;
        RECT 288.150 34.200 289.950 38.400 ;
        RECT 260.850 30.000 261.900 31.800 ;
        RECT 271.050 30.000 272.850 30.600 ;
        RECT 260.850 28.800 272.850 30.000 ;
        RECT 253.950 27.600 261.900 28.800 ;
        RECT 253.950 25.050 255.750 27.600 ;
        RECT 260.100 27.000 261.900 27.600 ;
        RECT 257.100 25.800 258.900 26.400 ;
        RECT 253.950 22.950 256.050 25.050 ;
        RECT 257.100 24.600 265.200 25.800 ;
        RECT 263.100 22.950 265.200 24.600 ;
        RECT 261.450 17.700 263.250 18.000 ;
        RECT 235.800 15.600 237.900 16.500 ;
        RECT 206.100 14.700 213.900 15.600 ;
        RECT 169.500 3.000 171.300 9.600 ;
        RECT 185.100 3.600 186.900 9.600 ;
        RECT 188.100 3.000 189.900 9.600 ;
        RECT 206.100 3.600 207.900 14.700 ;
        RECT 209.100 3.000 210.900 13.800 ;
        RECT 212.100 3.600 213.900 14.700 ;
        RECT 215.100 3.600 216.900 15.600 ;
        RECT 233.100 14.400 237.900 15.600 ;
        RECT 240.600 15.600 241.800 16.950 ;
        RECT 245.400 15.600 247.500 17.700 ;
        RECT 251.550 17.100 263.250 17.700 ;
        RECT 251.550 16.500 269.850 17.100 ;
        RECT 251.550 15.600 252.450 16.500 ;
        RECT 261.450 16.200 269.850 16.500 ;
        RECT 233.100 3.600 234.900 14.400 ;
        RECT 236.100 3.000 237.900 13.500 ;
        RECT 240.600 3.600 242.400 15.600 ;
        RECT 245.400 14.700 249.900 15.600 ;
        RECT 245.100 3.000 246.900 13.500 ;
        RECT 248.100 3.600 249.900 14.700 ;
        RECT 251.550 13.800 253.950 15.600 ;
        RECT 252.150 3.600 253.950 13.800 ;
        RECT 255.150 3.000 256.950 15.600 ;
        RECT 266.250 14.700 268.050 15.300 ;
        RECT 260.250 13.500 268.050 14.700 ;
        RECT 268.950 14.100 269.850 16.200 ;
        RECT 271.950 16.200 272.850 28.800 ;
        RECT 284.250 25.050 285.450 32.400 ;
        RECT 279.150 23.250 285.450 25.050 ;
        RECT 280.950 22.950 285.450 23.250 ;
        RECT 275.550 20.100 277.650 20.400 ;
        RECT 281.550 20.100 283.350 20.250 ;
        RECT 275.550 18.900 283.350 20.100 ;
        RECT 275.550 18.300 277.650 18.900 ;
        RECT 281.550 18.450 283.350 18.900 ;
        RECT 271.950 15.300 276.750 16.200 ;
        RECT 284.250 15.600 285.450 22.950 ;
        RECT 275.550 14.400 276.750 15.300 ;
        RECT 272.850 14.100 274.650 14.400 ;
        RECT 260.250 12.600 262.350 13.500 ;
        RECT 268.950 13.200 274.650 14.100 ;
        RECT 272.850 12.600 274.650 13.200 ;
        RECT 275.550 12.600 278.550 14.400 ;
        RECT 260.550 3.600 262.350 12.600 ;
        RECT 264.450 11.550 266.250 12.300 ;
        RECT 269.250 11.550 271.050 12.300 ;
        RECT 264.450 10.500 271.050 11.550 ;
        RECT 265.350 3.000 267.150 9.600 ;
        RECT 268.350 3.600 270.150 10.500 ;
        RECT 275.550 9.600 277.650 11.700 ;
        RECT 271.350 3.000 273.150 9.600 ;
        RECT 275.850 3.600 277.650 9.600 ;
        RECT 280.650 3.000 282.450 15.600 ;
        RECT 283.650 3.600 285.450 15.600 ;
        RECT 287.550 32.400 289.950 34.200 ;
        RECT 291.150 32.400 292.950 39.000 ;
        RECT 295.950 36.300 297.750 38.400 ;
        RECT 294.150 35.400 297.750 36.300 ;
        RECT 300.450 35.400 302.250 39.000 ;
        RECT 303.750 35.400 305.550 38.400 ;
        RECT 306.750 35.400 308.550 39.000 ;
        RECT 311.250 35.400 313.050 38.400 ;
        RECT 293.850 34.800 297.750 35.400 ;
        RECT 293.850 33.300 295.950 34.800 ;
        RECT 303.750 34.500 304.800 35.400 ;
        RECT 287.550 17.700 288.450 32.400 ;
        RECT 296.850 31.800 298.650 33.600 ;
        RECT 299.850 33.450 304.800 34.500 ;
        RECT 299.850 32.700 301.650 33.450 ;
        RECT 311.250 33.300 313.650 35.400 ;
        RECT 316.350 32.400 318.150 39.000 ;
        RECT 319.650 32.400 321.450 38.400 ;
        RECT 296.850 30.000 297.900 31.800 ;
        RECT 307.050 30.000 308.850 30.600 ;
        RECT 296.850 28.800 308.850 30.000 ;
        RECT 289.950 27.600 297.900 28.800 ;
        RECT 289.950 25.050 291.750 27.600 ;
        RECT 296.100 27.000 297.900 27.600 ;
        RECT 293.100 25.800 294.900 26.400 ;
        RECT 289.950 22.950 292.050 25.050 ;
        RECT 293.100 24.600 301.200 25.800 ;
        RECT 299.100 22.950 301.200 24.600 ;
        RECT 297.450 17.700 299.250 18.000 ;
        RECT 287.550 17.100 299.250 17.700 ;
        RECT 287.550 16.500 305.850 17.100 ;
        RECT 287.550 15.600 288.450 16.500 ;
        RECT 297.450 16.200 305.850 16.500 ;
        RECT 287.550 13.800 289.950 15.600 ;
        RECT 288.150 3.600 289.950 13.800 ;
        RECT 291.150 3.000 292.950 15.600 ;
        RECT 302.250 14.700 304.050 15.300 ;
        RECT 296.250 13.500 304.050 14.700 ;
        RECT 304.950 14.100 305.850 16.200 ;
        RECT 307.950 16.200 308.850 28.800 ;
        RECT 320.250 25.050 321.450 32.400 ;
        RECT 335.100 35.400 336.900 38.400 ;
        RECT 335.100 31.500 336.300 35.400 ;
        RECT 338.100 32.400 339.900 39.000 ;
        RECT 341.100 32.400 342.900 38.400 ;
        RECT 335.100 30.600 340.800 31.500 ;
        RECT 339.000 29.700 340.800 30.600 ;
        RECT 315.150 23.250 321.450 25.050 ;
        RECT 316.950 22.950 321.450 23.250 ;
        RECT 311.550 20.100 313.650 20.400 ;
        RECT 317.550 20.100 319.350 20.250 ;
        RECT 311.550 18.900 319.350 20.100 ;
        RECT 311.550 18.300 313.650 18.900 ;
        RECT 317.550 18.450 319.350 18.900 ;
        RECT 307.950 15.300 312.750 16.200 ;
        RECT 320.250 15.600 321.450 22.950 ;
        RECT 335.400 22.950 337.500 25.050 ;
        RECT 335.400 21.150 337.200 22.950 ;
        RECT 339.000 18.300 339.900 29.700 ;
        RECT 341.700 25.050 342.900 32.400 ;
        RECT 340.800 22.950 342.900 25.050 ;
        RECT 339.000 17.400 340.800 18.300 ;
        RECT 311.550 14.400 312.750 15.300 ;
        RECT 308.850 14.100 310.650 14.400 ;
        RECT 296.250 12.600 298.350 13.500 ;
        RECT 304.950 13.200 310.650 14.100 ;
        RECT 308.850 12.600 310.650 13.200 ;
        RECT 311.550 12.600 314.550 14.400 ;
        RECT 296.550 3.600 298.350 12.600 ;
        RECT 300.450 11.550 302.250 12.300 ;
        RECT 305.250 11.550 307.050 12.300 ;
        RECT 300.450 10.500 307.050 11.550 ;
        RECT 301.350 3.000 303.150 9.600 ;
        RECT 304.350 3.600 306.150 10.500 ;
        RECT 311.550 9.600 313.650 11.700 ;
        RECT 307.350 3.000 309.150 9.600 ;
        RECT 311.850 3.600 313.650 9.600 ;
        RECT 316.650 3.000 318.450 15.600 ;
        RECT 319.650 3.600 321.450 15.600 ;
        RECT 335.100 16.500 340.800 17.400 ;
        RECT 335.100 9.600 336.300 16.500 ;
        RECT 341.700 15.600 342.900 22.950 ;
        RECT 335.100 3.600 336.900 9.600 ;
        RECT 338.100 3.000 339.900 13.800 ;
        RECT 341.100 3.600 342.900 15.600 ;
        RECT 356.100 32.400 357.900 38.400 ;
        RECT 359.100 32.400 360.900 39.000 ;
        RECT 362.100 35.400 363.900 38.400 ;
        RECT 356.100 25.050 357.300 32.400 ;
        RECT 362.700 31.500 363.900 35.400 ;
        RECT 378.600 34.200 380.400 38.400 ;
        RECT 358.200 30.600 363.900 31.500 ;
        RECT 377.700 32.400 380.400 34.200 ;
        RECT 381.600 32.400 383.400 39.000 ;
        RECT 358.200 29.700 360.000 30.600 ;
        RECT 356.100 22.950 358.200 25.050 ;
        RECT 356.100 15.600 357.300 22.950 ;
        RECT 359.100 18.300 360.000 29.700 ;
        RECT 377.700 25.050 378.600 32.400 ;
        RECT 379.500 30.600 381.300 31.500 ;
        RECT 386.100 30.600 387.900 38.400 ;
        RECT 379.500 29.700 387.900 30.600 ;
        RECT 401.700 31.200 403.500 38.400 ;
        RECT 406.800 32.400 408.600 39.000 ;
        RECT 425.100 32.400 426.900 38.400 ;
        RECT 428.100 33.000 429.900 39.000 ;
        RECT 434.700 38.400 435.900 39.000 ;
        RECT 431.100 35.400 432.900 38.400 ;
        RECT 434.100 35.400 435.900 38.400 ;
        RECT 401.700 30.300 405.900 31.200 ;
        RECT 361.500 22.950 363.600 25.050 ;
        RECT 377.100 22.950 379.200 25.050 ;
        RECT 380.400 22.950 382.500 25.050 ;
        RECT 361.800 21.150 363.600 22.950 ;
        RECT 358.200 17.400 360.000 18.300 ;
        RECT 358.200 16.500 363.900 17.400 ;
        RECT 356.100 3.600 357.900 15.600 ;
        RECT 359.100 3.000 360.900 13.800 ;
        RECT 362.700 9.600 363.900 16.500 ;
        RECT 377.700 15.600 378.600 22.950 ;
        RECT 381.000 21.150 382.800 22.950 ;
        RECT 362.100 3.600 363.900 9.600 ;
        RECT 377.100 3.600 378.900 15.600 ;
        RECT 380.100 3.000 381.900 15.000 ;
        RECT 384.000 9.600 384.900 29.700 ;
        RECT 385.950 25.050 387.750 26.850 ;
        RECT 401.100 25.050 402.900 26.850 ;
        RECT 404.700 25.050 405.900 30.300 ;
        RECT 406.950 25.050 408.750 26.850 ;
        RECT 425.100 25.050 426.000 32.400 ;
        RECT 431.700 31.200 432.600 35.400 ;
        RECT 449.400 32.400 451.200 39.000 ;
        RECT 454.500 31.200 456.300 38.400 ;
        RECT 427.200 30.300 432.600 31.200 ;
        RECT 452.100 30.300 456.300 31.200 ;
        RECT 470.700 31.200 472.500 38.400 ;
        RECT 475.800 32.400 477.600 39.000 ;
        RECT 491.400 32.400 493.200 39.000 ;
        RECT 496.500 31.200 498.300 38.400 ;
        RECT 470.700 30.300 474.900 31.200 ;
        RECT 427.200 29.400 429.300 30.300 ;
        RECT 385.800 22.950 387.900 25.050 ;
        RECT 400.950 22.950 403.050 25.050 ;
        RECT 403.950 22.950 406.050 25.050 ;
        RECT 406.950 22.950 409.050 25.050 ;
        RECT 425.100 22.950 427.200 25.050 ;
        RECT 404.700 9.600 405.900 22.950 ;
        RECT 406.950 18.450 409.050 19.050 ;
        RECT 415.950 18.450 418.050 19.050 ;
        RECT 406.950 17.550 418.050 18.450 ;
        RECT 406.950 16.950 409.050 17.550 ;
        RECT 415.950 16.950 418.050 17.550 ;
        RECT 426.000 15.600 427.200 22.950 ;
        RECT 428.400 18.900 429.300 29.400 ;
        RECT 433.800 25.050 435.600 26.850 ;
        RECT 449.250 25.050 451.050 26.850 ;
        RECT 452.100 25.050 453.300 30.300 ;
        RECT 455.100 25.050 456.900 26.850 ;
        RECT 470.100 25.050 471.900 26.850 ;
        RECT 473.700 25.050 474.900 30.300 ;
        RECT 494.100 30.300 498.300 31.200 ;
        RECT 512.100 30.600 513.900 38.400 ;
        RECT 516.600 32.400 518.400 39.000 ;
        RECT 519.600 34.200 521.400 38.400 ;
        RECT 536.700 35.400 538.500 39.000 ;
        RECT 519.600 32.400 522.300 34.200 ;
        RECT 539.700 33.600 541.500 38.400 ;
        RECT 518.700 30.600 520.500 31.500 ;
        RECT 475.950 25.050 477.750 26.850 ;
        RECT 491.250 25.050 493.050 26.850 ;
        RECT 494.100 25.050 495.300 30.300 ;
        RECT 512.100 29.700 520.500 30.600 ;
        RECT 497.100 25.050 498.900 26.850 ;
        RECT 512.250 25.050 514.050 26.850 ;
        RECT 430.500 22.950 432.600 25.050 ;
        RECT 433.800 22.950 435.900 25.050 ;
        RECT 448.950 22.950 451.050 25.050 ;
        RECT 451.950 22.950 454.050 25.050 ;
        RECT 454.950 22.950 457.050 25.050 ;
        RECT 469.950 22.950 472.050 25.050 ;
        RECT 472.950 22.950 475.050 25.050 ;
        RECT 475.950 22.950 478.050 25.050 ;
        RECT 490.950 22.950 493.050 25.050 ;
        RECT 493.950 22.950 496.050 25.050 ;
        RECT 496.950 22.950 499.050 25.050 ;
        RECT 512.100 22.950 514.200 25.050 ;
        RECT 430.200 21.150 432.000 22.950 ;
        RECT 428.100 18.300 429.900 18.900 ;
        RECT 428.100 17.100 435.900 18.300 ;
        RECT 434.700 15.600 435.900 17.100 ;
        RECT 426.000 14.100 428.400 15.600 ;
        RECT 383.100 3.600 384.900 9.600 ;
        RECT 386.100 3.000 387.900 9.600 ;
        RECT 401.100 3.000 402.900 9.600 ;
        RECT 404.100 3.600 405.900 9.600 ;
        RECT 407.100 3.000 408.900 9.600 ;
        RECT 426.600 3.600 428.400 14.100 ;
        RECT 429.600 3.000 431.400 15.600 ;
        RECT 434.100 3.600 435.900 15.600 ;
        RECT 452.100 9.600 453.300 22.950 ;
        RECT 473.700 9.600 474.900 22.950 ;
        RECT 494.100 9.600 495.300 22.950 ;
        RECT 515.100 9.600 516.000 29.700 ;
        RECT 521.400 25.050 522.300 32.400 ;
        RECT 536.400 32.400 541.500 33.600 ;
        RECT 544.200 32.400 546.000 39.000 ;
        RECT 563.100 35.400 564.900 38.400 ;
        RECT 566.100 35.400 567.900 39.000 ;
        RECT 536.400 25.050 537.300 32.400 ;
        RECT 538.950 25.050 540.750 26.850 ;
        RECT 545.100 25.050 546.900 26.850 ;
        RECT 563.700 25.050 564.900 35.400 ;
        RECT 581.100 32.400 582.900 38.400 ;
        RECT 581.700 30.300 582.900 32.400 ;
        RECT 584.100 33.300 585.900 38.400 ;
        RECT 587.100 34.200 588.900 39.000 ;
        RECT 590.100 33.300 591.900 38.400 ;
        RECT 584.100 31.950 591.900 33.300 ;
        RECT 605.400 32.400 607.200 39.000 ;
        RECT 610.500 31.200 612.300 38.400 ;
        RECT 626.100 32.400 627.900 38.400 ;
        RECT 629.100 33.300 630.900 39.000 ;
        RECT 633.600 32.400 635.400 38.400 ;
        RECT 638.100 33.300 639.900 39.000 ;
        RECT 641.100 32.400 642.900 38.400 ;
        RECT 656.400 32.400 658.200 39.000 ;
        RECT 626.100 31.500 630.900 32.400 ;
        RECT 608.100 30.300 612.300 31.200 ;
        RECT 628.800 30.300 630.900 31.500 ;
        RECT 633.900 30.900 635.100 32.400 ;
        RECT 581.700 29.400 585.300 30.300 ;
        RECT 581.100 25.050 582.900 26.850 ;
        RECT 584.100 25.050 585.300 29.400 ;
        RECT 587.100 25.050 588.900 26.850 ;
        RECT 605.250 25.050 607.050 26.850 ;
        RECT 608.100 25.050 609.300 30.300 ;
        RECT 632.100 28.800 635.100 30.900 ;
        RECT 641.100 30.600 642.300 32.400 ;
        RECT 661.500 31.200 663.300 38.400 ;
        RECT 680.400 32.400 682.200 39.000 ;
        RECT 685.500 31.200 687.300 38.400 ;
        RECT 690.150 34.200 691.950 38.400 ;
        RECT 611.100 25.050 612.900 26.850 ;
        RECT 630.900 25.800 633.000 27.900 ;
        RECT 517.500 22.950 519.600 25.050 ;
        RECT 520.800 22.950 522.900 25.050 ;
        RECT 535.950 22.950 538.050 25.050 ;
        RECT 538.950 22.950 541.050 25.050 ;
        RECT 541.950 22.950 544.050 25.050 ;
        RECT 544.950 22.950 547.050 25.050 ;
        RECT 562.950 22.950 565.050 25.050 ;
        RECT 565.950 22.950 568.050 25.050 ;
        RECT 580.950 22.950 583.050 25.050 ;
        RECT 583.950 22.950 586.050 25.050 ;
        RECT 586.950 22.950 589.050 25.050 ;
        RECT 589.950 22.950 592.050 25.050 ;
        RECT 604.950 22.950 607.050 25.050 ;
        RECT 607.950 22.950 610.050 25.050 ;
        RECT 610.950 22.950 613.050 25.050 ;
        RECT 626.100 22.950 628.200 25.050 ;
        RECT 630.900 24.000 632.700 25.800 ;
        RECT 633.900 23.100 635.100 28.800 ;
        RECT 636.000 29.700 642.300 30.600 ;
        RECT 659.100 30.300 663.300 31.200 ;
        RECT 683.100 30.300 687.300 31.200 ;
        RECT 689.550 32.400 691.950 34.200 ;
        RECT 693.150 32.400 694.950 39.000 ;
        RECT 697.950 36.300 699.750 38.400 ;
        RECT 696.150 35.400 699.750 36.300 ;
        RECT 702.450 35.400 704.250 39.000 ;
        RECT 705.750 35.400 707.550 38.400 ;
        RECT 708.750 35.400 710.550 39.000 ;
        RECT 713.250 35.400 715.050 38.400 ;
        RECT 695.850 34.800 699.750 35.400 ;
        RECT 695.850 33.300 697.950 34.800 ;
        RECT 705.750 34.500 706.800 35.400 ;
        RECT 636.000 27.600 638.100 29.700 ;
        RECT 636.000 25.800 637.800 27.600 ;
        RECT 640.800 25.050 642.600 26.850 ;
        RECT 656.250 25.050 658.050 26.850 ;
        RECT 659.100 25.050 660.300 30.300 ;
        RECT 662.100 25.050 663.900 26.850 ;
        RECT 680.250 25.050 682.050 26.850 ;
        RECT 683.100 25.050 684.300 30.300 ;
        RECT 686.100 25.050 687.900 26.850 ;
        RECT 640.800 24.300 642.900 25.050 ;
        RECT 517.200 21.150 519.000 22.950 ;
        RECT 521.400 15.600 522.300 22.950 ;
        RECT 536.400 15.600 537.300 22.950 ;
        RECT 541.950 21.150 543.750 22.950 ;
        RECT 449.100 3.000 450.900 9.600 ;
        RECT 452.100 3.600 453.900 9.600 ;
        RECT 455.100 3.000 456.900 9.600 ;
        RECT 470.100 3.000 471.900 9.600 ;
        RECT 473.100 3.600 474.900 9.600 ;
        RECT 476.100 3.000 477.900 9.600 ;
        RECT 491.100 3.000 492.900 9.600 ;
        RECT 494.100 3.600 495.900 9.600 ;
        RECT 497.100 3.000 498.900 9.600 ;
        RECT 512.100 3.000 513.900 9.600 ;
        RECT 515.100 3.600 516.900 9.600 ;
        RECT 518.100 3.000 519.900 15.000 ;
        RECT 521.100 3.600 522.900 15.600 ;
        RECT 536.100 3.600 537.900 15.600 ;
        RECT 539.100 14.700 546.900 15.600 ;
        RECT 539.100 3.600 540.900 14.700 ;
        RECT 542.100 3.000 543.900 13.800 ;
        RECT 545.100 3.600 546.900 14.700 ;
        RECT 563.700 9.600 564.900 22.950 ;
        RECT 566.100 21.150 567.900 22.950 ;
        RECT 584.100 15.600 585.300 22.950 ;
        RECT 590.100 21.150 591.900 22.950 ;
        RECT 592.950 18.450 595.050 19.050 ;
        RECT 604.950 18.450 607.050 19.050 ;
        RECT 592.950 17.550 607.050 18.450 ;
        RECT 592.950 16.950 595.050 17.550 ;
        RECT 604.950 16.950 607.050 17.550 ;
        RECT 584.100 14.100 586.500 15.600 ;
        RECT 582.000 11.100 583.800 12.900 ;
        RECT 563.100 3.600 564.900 9.600 ;
        RECT 566.100 3.000 567.900 9.600 ;
        RECT 581.700 3.000 583.500 9.600 ;
        RECT 584.700 3.600 586.500 14.100 ;
        RECT 589.800 3.000 591.600 15.600 ;
        RECT 608.100 9.600 609.300 22.950 ;
        RECT 626.400 21.150 628.200 22.950 ;
        RECT 632.700 22.200 635.100 23.100 ;
        RECT 636.000 22.950 642.900 24.300 ;
        RECT 655.950 22.950 658.050 25.050 ;
        RECT 658.950 22.950 661.050 25.050 ;
        RECT 661.950 22.950 664.050 25.050 ;
        RECT 679.950 22.950 682.050 25.050 ;
        RECT 682.950 22.950 685.050 25.050 ;
        RECT 685.950 22.950 688.050 25.050 ;
        RECT 636.000 22.500 637.800 22.950 ;
        RECT 632.700 22.050 634.200 22.200 ;
        RECT 632.100 19.950 634.200 22.050 ;
        RECT 633.300 18.000 634.200 19.950 ;
        RECT 635.100 19.500 639.000 21.300 ;
        RECT 635.100 19.200 637.200 19.500 ;
        RECT 633.300 16.950 634.800 18.000 ;
        RECT 628.800 15.600 630.900 16.500 ;
        RECT 626.100 14.400 630.900 15.600 ;
        RECT 633.600 15.600 634.800 16.950 ;
        RECT 638.400 15.600 640.500 17.700 ;
        RECT 605.100 3.000 606.900 9.600 ;
        RECT 608.100 3.600 609.900 9.600 ;
        RECT 611.100 3.000 612.900 9.600 ;
        RECT 626.100 3.600 627.900 14.400 ;
        RECT 629.100 3.000 630.900 13.500 ;
        RECT 633.600 3.600 635.400 15.600 ;
        RECT 638.400 14.700 642.900 15.600 ;
        RECT 638.100 3.000 639.900 13.500 ;
        RECT 641.100 3.600 642.900 14.700 ;
        RECT 659.100 9.600 660.300 22.950 ;
        RECT 683.100 9.600 684.300 22.950 ;
        RECT 689.550 17.700 690.450 32.400 ;
        RECT 698.850 31.800 700.650 33.600 ;
        RECT 701.850 33.450 706.800 34.500 ;
        RECT 701.850 32.700 703.650 33.450 ;
        RECT 713.250 33.300 715.650 35.400 ;
        RECT 718.350 32.400 720.150 39.000 ;
        RECT 721.650 32.400 723.450 38.400 ;
        RECT 726.150 34.200 727.950 38.400 ;
        RECT 698.850 30.000 699.900 31.800 ;
        RECT 709.050 30.000 710.850 30.600 ;
        RECT 698.850 28.800 710.850 30.000 ;
        RECT 691.950 27.600 699.900 28.800 ;
        RECT 691.950 25.050 693.750 27.600 ;
        RECT 698.100 27.000 699.900 27.600 ;
        RECT 695.100 25.800 696.900 26.400 ;
        RECT 691.950 22.950 694.050 25.050 ;
        RECT 695.100 24.600 703.200 25.800 ;
        RECT 701.100 22.950 703.200 24.600 ;
        RECT 699.450 17.700 701.250 18.000 ;
        RECT 689.550 17.100 701.250 17.700 ;
        RECT 689.550 16.500 707.850 17.100 ;
        RECT 689.550 15.600 690.450 16.500 ;
        RECT 699.450 16.200 707.850 16.500 ;
        RECT 689.550 13.800 691.950 15.600 ;
        RECT 656.100 3.000 657.900 9.600 ;
        RECT 659.100 3.600 660.900 9.600 ;
        RECT 662.100 3.000 663.900 9.600 ;
        RECT 680.100 3.000 681.900 9.600 ;
        RECT 683.100 3.600 684.900 9.600 ;
        RECT 686.100 3.000 687.900 9.600 ;
        RECT 690.150 3.600 691.950 13.800 ;
        RECT 693.150 3.000 694.950 15.600 ;
        RECT 704.250 14.700 706.050 15.300 ;
        RECT 698.250 13.500 706.050 14.700 ;
        RECT 706.950 14.100 707.850 16.200 ;
        RECT 709.950 16.200 710.850 28.800 ;
        RECT 722.250 25.050 723.450 32.400 ;
        RECT 717.150 23.250 723.450 25.050 ;
        RECT 718.950 22.950 723.450 23.250 ;
        RECT 713.550 20.100 715.650 20.400 ;
        RECT 719.550 20.100 721.350 20.250 ;
        RECT 713.550 18.900 721.350 20.100 ;
        RECT 713.550 18.300 715.650 18.900 ;
        RECT 719.550 18.450 721.350 18.900 ;
        RECT 709.950 15.300 714.750 16.200 ;
        RECT 722.250 15.600 723.450 22.950 ;
        RECT 713.550 14.400 714.750 15.300 ;
        RECT 710.850 14.100 712.650 14.400 ;
        RECT 698.250 12.600 700.350 13.500 ;
        RECT 706.950 13.200 712.650 14.100 ;
        RECT 710.850 12.600 712.650 13.200 ;
        RECT 713.550 12.600 716.550 14.400 ;
        RECT 698.550 3.600 700.350 12.600 ;
        RECT 702.450 11.550 704.250 12.300 ;
        RECT 707.250 11.550 709.050 12.300 ;
        RECT 702.450 10.500 709.050 11.550 ;
        RECT 703.350 3.000 705.150 9.600 ;
        RECT 706.350 3.600 708.150 10.500 ;
        RECT 713.550 9.600 715.650 11.700 ;
        RECT 709.350 3.000 711.150 9.600 ;
        RECT 713.850 3.600 715.650 9.600 ;
        RECT 718.650 3.000 720.450 15.600 ;
        RECT 721.650 3.600 723.450 15.600 ;
        RECT 725.550 32.400 727.950 34.200 ;
        RECT 729.150 32.400 730.950 39.000 ;
        RECT 733.950 36.300 735.750 38.400 ;
        RECT 732.150 35.400 735.750 36.300 ;
        RECT 738.450 35.400 740.250 39.000 ;
        RECT 741.750 35.400 743.550 38.400 ;
        RECT 744.750 35.400 746.550 39.000 ;
        RECT 749.250 35.400 751.050 38.400 ;
        RECT 731.850 34.800 735.750 35.400 ;
        RECT 731.850 33.300 733.950 34.800 ;
        RECT 741.750 34.500 742.800 35.400 ;
        RECT 725.550 17.700 726.450 32.400 ;
        RECT 734.850 31.800 736.650 33.600 ;
        RECT 737.850 33.450 742.800 34.500 ;
        RECT 737.850 32.700 739.650 33.450 ;
        RECT 749.250 33.300 751.650 35.400 ;
        RECT 754.350 32.400 756.150 39.000 ;
        RECT 757.650 32.400 759.450 38.400 ;
        RECT 734.850 30.000 735.900 31.800 ;
        RECT 745.050 30.000 746.850 30.600 ;
        RECT 734.850 28.800 746.850 30.000 ;
        RECT 727.950 27.600 735.900 28.800 ;
        RECT 727.950 25.050 729.750 27.600 ;
        RECT 734.100 27.000 735.900 27.600 ;
        RECT 731.100 25.800 732.900 26.400 ;
        RECT 727.950 22.950 730.050 25.050 ;
        RECT 731.100 24.600 739.200 25.800 ;
        RECT 737.100 22.950 739.200 24.600 ;
        RECT 735.450 17.700 737.250 18.000 ;
        RECT 725.550 17.100 737.250 17.700 ;
        RECT 725.550 16.500 743.850 17.100 ;
        RECT 725.550 15.600 726.450 16.500 ;
        RECT 735.450 16.200 743.850 16.500 ;
        RECT 725.550 13.800 727.950 15.600 ;
        RECT 726.150 3.600 727.950 13.800 ;
        RECT 729.150 3.000 730.950 15.600 ;
        RECT 740.250 14.700 742.050 15.300 ;
        RECT 734.250 13.500 742.050 14.700 ;
        RECT 742.950 14.100 743.850 16.200 ;
        RECT 745.950 16.200 746.850 28.800 ;
        RECT 758.250 25.050 759.450 32.400 ;
        RECT 773.100 35.400 774.900 38.400 ;
        RECT 773.100 31.500 774.300 35.400 ;
        RECT 776.100 32.400 777.900 39.000 ;
        RECT 779.100 32.400 780.900 38.400 ;
        RECT 773.100 30.600 778.800 31.500 ;
        RECT 777.000 29.700 778.800 30.600 ;
        RECT 753.150 23.250 759.450 25.050 ;
        RECT 754.950 22.950 759.450 23.250 ;
        RECT 749.550 20.100 751.650 20.400 ;
        RECT 755.550 20.100 757.350 20.250 ;
        RECT 749.550 18.900 757.350 20.100 ;
        RECT 749.550 18.300 751.650 18.900 ;
        RECT 755.550 18.450 757.350 18.900 ;
        RECT 745.950 15.300 750.750 16.200 ;
        RECT 758.250 15.600 759.450 22.950 ;
        RECT 773.400 22.950 775.500 25.050 ;
        RECT 773.400 21.150 775.200 22.950 ;
        RECT 777.000 18.300 777.900 29.700 ;
        RECT 779.700 25.050 780.900 32.400 ;
        RECT 796.500 30.000 798.300 38.400 ;
        RECT 795.000 28.800 798.300 30.000 ;
        RECT 803.100 29.400 804.900 39.000 ;
        RECT 818.700 31.200 820.500 38.400 ;
        RECT 823.800 32.400 825.600 39.000 ;
        RECT 839.700 31.200 841.500 38.400 ;
        RECT 844.800 32.400 846.600 39.000 ;
        RECT 860.100 35.400 861.900 39.000 ;
        RECT 863.100 35.400 864.900 38.400 ;
        RECT 866.100 35.400 867.900 39.000 ;
        RECT 818.700 30.300 822.900 31.200 ;
        RECT 839.700 30.300 843.900 31.200 ;
        RECT 795.000 25.050 795.900 28.800 ;
        RECT 797.100 25.050 798.900 26.850 ;
        RECT 803.100 25.050 804.900 26.850 ;
        RECT 818.100 25.050 819.900 26.850 ;
        RECT 821.700 25.050 822.900 30.300 ;
        RECT 823.950 25.050 825.750 26.850 ;
        RECT 839.100 25.050 840.900 26.850 ;
        RECT 842.700 25.050 843.900 30.300 ;
        RECT 844.950 25.050 846.750 26.850 ;
        RECT 863.400 25.050 864.300 35.400 ;
        RECT 881.100 32.400 882.900 38.400 ;
        RECT 884.100 32.400 885.900 39.000 ;
        RECT 887.100 35.400 888.900 38.400 ;
        RECT 881.100 25.050 882.300 32.400 ;
        RECT 887.700 31.500 888.900 35.400 ;
        RECT 883.200 30.600 888.900 31.500 ;
        RECT 883.200 29.700 885.000 30.600 ;
        RECT 778.800 22.950 780.900 25.050 ;
        RECT 793.950 22.950 796.050 25.050 ;
        RECT 796.950 22.950 799.050 25.050 ;
        RECT 799.950 22.950 802.050 25.050 ;
        RECT 802.950 22.950 805.050 25.050 ;
        RECT 817.950 22.950 820.050 25.050 ;
        RECT 820.950 22.950 823.050 25.050 ;
        RECT 823.950 22.950 826.050 25.050 ;
        RECT 838.950 22.950 841.050 25.050 ;
        RECT 841.950 22.950 844.050 25.050 ;
        RECT 844.950 22.950 847.050 25.050 ;
        RECT 859.950 22.950 862.050 25.050 ;
        RECT 862.950 22.950 865.050 25.050 ;
        RECT 865.950 22.950 868.050 25.050 ;
        RECT 881.100 22.950 883.200 25.050 ;
        RECT 777.000 17.400 778.800 18.300 ;
        RECT 749.550 14.400 750.750 15.300 ;
        RECT 746.850 14.100 748.650 14.400 ;
        RECT 734.250 12.600 736.350 13.500 ;
        RECT 742.950 13.200 748.650 14.100 ;
        RECT 746.850 12.600 748.650 13.200 ;
        RECT 749.550 12.600 752.550 14.400 ;
        RECT 734.550 3.600 736.350 12.600 ;
        RECT 738.450 11.550 740.250 12.300 ;
        RECT 743.250 11.550 745.050 12.300 ;
        RECT 738.450 10.500 745.050 11.550 ;
        RECT 739.350 3.000 741.150 9.600 ;
        RECT 742.350 3.600 744.150 10.500 ;
        RECT 749.550 9.600 751.650 11.700 ;
        RECT 745.350 3.000 747.150 9.600 ;
        RECT 749.850 3.600 751.650 9.600 ;
        RECT 754.650 3.000 756.450 15.600 ;
        RECT 757.650 3.600 759.450 15.600 ;
        RECT 773.100 16.500 778.800 17.400 ;
        RECT 773.100 9.600 774.300 16.500 ;
        RECT 779.700 15.600 780.900 22.950 ;
        RECT 773.100 3.600 774.900 9.600 ;
        RECT 776.100 3.000 777.900 13.800 ;
        RECT 779.100 3.600 780.900 15.600 ;
        RECT 795.000 10.800 795.900 22.950 ;
        RECT 800.100 21.150 801.900 22.950 ;
        RECT 811.950 15.450 814.050 16.050 ;
        RECT 817.950 15.450 820.050 15.900 ;
        RECT 811.950 14.550 820.050 15.450 ;
        RECT 811.950 13.950 814.050 14.550 ;
        RECT 817.950 13.800 820.050 14.550 ;
        RECT 795.000 9.900 801.600 10.800 ;
        RECT 795.000 9.600 795.900 9.900 ;
        RECT 794.100 3.600 795.900 9.600 ;
        RECT 800.100 9.600 801.600 9.900 ;
        RECT 821.700 9.600 822.900 22.950 ;
        RECT 842.700 9.600 843.900 22.950 ;
        RECT 860.250 21.150 862.050 22.950 ;
        RECT 863.400 15.600 864.300 22.950 ;
        RECT 866.100 21.150 867.900 22.950 ;
        RECT 881.100 15.600 882.300 22.950 ;
        RECT 884.100 18.300 885.000 29.700 ;
        RECT 886.500 22.950 888.600 25.050 ;
        RECT 886.800 21.150 888.600 22.950 ;
        RECT 883.200 17.400 885.000 18.300 ;
        RECT 883.200 16.500 888.900 17.400 ;
        RECT 797.100 3.000 798.900 9.000 ;
        RECT 800.100 3.600 801.900 9.600 ;
        RECT 803.100 3.000 804.900 9.600 ;
        RECT 818.100 3.000 819.900 9.600 ;
        RECT 821.100 3.600 822.900 9.600 ;
        RECT 824.100 3.000 825.900 9.600 ;
        RECT 839.100 3.000 840.900 9.600 ;
        RECT 842.100 3.600 843.900 9.600 ;
        RECT 845.100 3.000 846.900 9.600 ;
        RECT 860.100 3.000 861.900 15.600 ;
        RECT 863.400 14.400 867.000 15.600 ;
        RECT 865.200 3.600 867.000 14.400 ;
        RECT 881.100 3.600 882.900 15.600 ;
        RECT 884.100 3.000 885.900 13.800 ;
        RECT 887.700 9.600 888.900 16.500 ;
        RECT 887.100 3.600 888.900 9.600 ;
      LAYER via1 ;
        RECT 70.950 880.950 73.050 883.050 ;
        RECT 166.950 880.950 169.050 883.050 ;
        RECT 224.550 891.300 226.650 893.400 ;
        RECT 317.550 891.300 319.650 893.400 ;
        RECT 427.950 880.950 430.050 883.050 ;
        RECT 508.950 880.950 511.050 883.050 ;
        RECT 566.550 891.300 568.650 893.400 ;
        RECT 160.950 835.950 163.050 838.050 ;
        RECT 178.800 835.950 180.900 838.050 ;
        RECT 319.950 835.950 322.050 838.050 ;
        RECT 337.800 835.950 339.900 838.050 ;
        RECT 355.950 835.950 358.050 838.050 ;
        RECT 373.800 835.950 375.900 838.050 ;
        RECT 490.950 835.950 493.050 838.050 ;
        RECT 508.800 835.950 510.900 838.050 ;
        RECT 868.950 832.950 871.050 835.050 ;
        RECT 346.800 808.800 348.900 810.900 ;
        RECT 25.950 724.950 28.050 727.050 ;
        RECT 526.950 727.950 529.050 730.050 ;
        RECT 688.950 727.950 691.050 730.050 ;
        RECT 526.950 721.950 529.050 724.050 ;
        RECT 739.950 727.950 742.050 730.050 ;
        RECT 688.950 721.950 691.050 724.050 ;
        RECT 781.950 730.950 784.050 733.050 ;
        RECT 739.950 721.950 742.050 724.050 ;
        RECT 838.950 727.950 841.050 730.050 ;
        RECT 421.800 683.700 423.900 685.800 ;
        RECT 424.800 674.100 426.900 676.200 ;
        RECT 478.950 679.950 481.050 682.050 ;
        RECT 496.800 679.950 498.900 682.050 ;
        RECT 514.950 679.950 517.050 682.050 ;
        RECT 532.800 679.950 534.900 682.050 ;
        RECT 715.800 652.800 717.900 654.900 ;
        RECT 749.100 652.800 751.200 654.900 ;
        RECT 865.950 649.950 868.050 652.050 ;
        RECT 25.950 601.950 28.050 604.050 ;
        RECT 43.800 601.950 45.900 604.050 ;
        RECT 457.950 607.950 460.050 610.050 ;
        RECT 625.950 598.950 628.050 601.050 ;
        RECT 25.950 568.950 28.050 571.050 ;
        RECT 82.950 568.950 85.050 571.050 ;
        RECT 157.950 568.950 160.050 571.050 ;
        RECT 841.950 571.950 844.050 574.050 ;
        RECT 841.950 565.950 844.050 568.050 ;
        RECT 25.950 523.950 28.050 526.050 ;
        RECT 43.800 523.950 45.900 526.050 ;
        RECT 61.950 523.950 64.050 526.050 ;
        RECT 79.800 523.950 81.900 526.050 ;
        RECT 532.950 526.950 535.050 529.050 ;
        RECT 532.950 520.950 535.050 523.050 ;
        RECT 835.950 526.950 838.050 529.050 ;
        RECT 883.950 526.950 886.050 529.050 ;
        RECT 835.950 520.950 838.050 523.050 ;
        RECT 25.950 490.950 28.050 493.050 ;
        RECT 529.950 493.950 532.050 496.050 ;
        RECT 649.950 493.950 652.050 496.050 ;
        RECT 529.950 487.950 532.050 490.050 ;
        RECT 649.950 487.950 652.050 490.050 ;
        RECT 28.950 445.950 31.050 448.050 ;
        RECT 46.800 445.950 48.900 448.050 ;
        RECT 64.950 445.950 67.050 448.050 ;
        RECT 82.800 445.950 84.900 448.050 ;
        RECT 562.950 448.950 565.050 451.050 ;
        RECT 400.950 442.950 403.050 445.050 ;
        RECT 877.950 445.950 880.050 448.050 ;
        RECT 67.950 412.950 70.050 415.050 ;
        RECT 103.950 412.950 106.050 415.050 ;
        RECT 511.950 412.950 514.050 415.050 ;
        RECT 706.950 418.950 709.050 421.050 ;
        RECT 25.950 367.950 28.050 370.050 ;
        RECT 43.800 367.950 45.900 370.050 ;
        RECT 61.950 367.950 64.050 370.050 ;
        RECT 79.800 367.950 81.900 370.050 ;
        RECT 490.500 361.800 492.600 363.900 ;
        RECT 502.800 367.950 504.900 370.050 ;
        RECT 544.500 361.800 546.600 363.900 ;
        RECT 556.800 367.950 558.900 370.050 ;
        RECT 49.950 334.950 52.050 337.050 ;
        RECT 103.950 334.950 106.050 337.050 ;
        RECT 571.950 337.950 574.050 340.050 ;
        RECT 190.950 334.950 193.050 337.050 ;
        RECT 571.950 331.950 574.050 334.050 ;
        RECT 874.950 337.950 877.050 340.050 ;
        RECT 58.950 289.950 61.050 292.050 ;
        RECT 76.800 289.950 78.900 292.050 ;
        RECT 751.950 292.950 754.050 295.050 ;
        RECT 751.950 286.950 754.050 289.050 ;
        RECT 118.950 256.950 121.050 259.050 ;
        RECT 16.500 205.800 18.600 207.900 ;
        RECT 28.800 211.950 30.900 214.050 ;
        RECT 140.100 211.950 142.200 214.050 ;
        RECT 142.500 205.500 144.600 207.600 ;
        RECT 149.100 214.950 151.200 217.050 ;
        RECT 149.100 206.100 151.200 208.200 ;
        RECT 152.400 205.800 154.500 207.900 ;
        RECT 574.950 211.950 577.050 214.050 ;
        RECT 592.800 211.950 594.900 214.050 ;
        RECT 610.950 211.950 613.050 214.050 ;
        RECT 628.800 211.950 630.900 214.050 ;
        RECT 616.800 184.800 618.900 186.900 ;
        RECT 748.950 181.950 751.050 184.050 ;
        RECT 820.950 181.950 823.050 184.050 ;
        RECT 748.950 175.950 751.050 178.050 ;
        RECT 820.950 175.950 823.050 178.050 ;
        RECT 16.500 127.800 18.600 129.900 ;
        RECT 622.800 137.700 624.900 139.800 ;
        RECT 28.800 133.950 30.900 136.050 ;
        RECT 625.800 128.100 627.900 130.200 ;
        RECT 61.950 97.950 64.050 100.050 ;
        RECT 341.550 111.300 343.650 113.400 ;
        RECT 862.950 100.950 865.050 103.050 ;
        RECT 338.100 55.950 340.200 58.050 ;
        RECT 355.950 55.950 358.050 58.050 ;
        RECT 395.100 55.950 397.200 58.050 ;
        RECT 350.550 45.600 352.650 47.700 ;
        RECT 397.500 49.500 399.600 51.600 ;
        RECT 404.100 58.950 406.200 61.050 ;
        RECT 404.100 50.100 406.200 52.200 ;
        RECT 407.400 49.800 409.500 51.900 ;
        RECT 275.550 33.300 277.650 35.400 ;
        RECT 311.550 33.300 313.650 35.400 ;
        RECT 713.550 33.300 715.650 35.400 ;
        RECT 749.550 33.300 751.650 35.400 ;
      LAYER metal2 ;
        RECT 76.350 891.300 78.450 893.400 ;
        RECT 94.050 891.300 96.150 893.400 ;
        RECT 172.350 891.300 174.450 893.400 ;
        RECT 190.050 891.300 192.150 893.400 ;
        RECT 206.850 891.300 208.950 893.400 ;
        RECT 224.550 891.300 226.650 893.400 ;
        RECT 299.850 891.300 301.950 893.400 ;
        RECT 317.550 891.300 319.650 893.400 ;
        RECT 433.350 891.300 435.450 893.400 ;
        RECT 451.050 891.300 453.150 893.400 ;
        RECT 514.350 891.300 516.450 893.400 ;
        RECT 532.050 891.300 534.150 893.400 ;
        RECT 548.850 891.300 550.950 893.400 ;
        RECT 566.550 891.300 568.650 893.400 ;
        RECT 40.950 884.100 43.050 886.200 ;
        RECT 41.400 883.350 42.600 884.100 ;
        RECT 52.950 883.950 55.050 886.050 ;
        RECT 64.950 884.100 67.050 886.200 ;
        RECT 70.950 884.100 73.050 886.200 ;
        RECT 17.100 880.950 19.200 883.050 ;
        RECT 22.500 880.950 24.600 883.050 ;
        RECT 37.950 880.950 40.050 883.050 ;
        RECT 40.950 880.950 43.050 883.050 ;
        RECT 43.950 880.950 46.050 883.050 ;
        RECT 17.400 879.900 18.600 880.650 ;
        RECT 16.950 877.800 19.050 879.900 ;
        RECT 25.950 877.950 28.050 880.050 ;
        RECT 38.400 879.900 39.600 880.650 ;
        RECT 16.950 839.100 19.050 841.200 ;
        RECT 17.400 838.350 18.600 839.100 ;
        RECT 13.950 835.950 16.050 838.050 ;
        RECT 16.950 835.950 19.050 838.050 ;
        RECT 26.400 829.050 27.450 877.950 ;
        RECT 37.950 877.800 40.050 879.900 ;
        RECT 44.400 878.400 45.600 880.650 ;
        RECT 44.400 850.050 45.450 878.400 ;
        RECT 43.950 847.950 46.050 850.050 ;
        RECT 53.400 841.200 54.450 883.950 ;
        RECT 65.400 883.350 66.600 884.100 ;
        RECT 71.400 883.350 72.600 884.100 ;
        RECT 59.100 880.950 61.200 883.050 ;
        RECT 64.500 880.950 66.600 883.050 ;
        RECT 70.950 880.950 73.050 883.050 ;
        RECT 77.250 878.400 78.450 891.300 ;
        RECT 88.800 880.950 90.900 883.050 ;
        RECT 89.400 879.000 90.600 880.650 ;
        RECT 76.350 876.300 78.450 878.400 ;
        RECT 77.250 869.700 78.450 876.300 ;
        RECT 88.950 874.950 91.050 879.000 ;
        RECT 94.650 872.700 95.850 891.300 ;
        RECT 160.950 884.100 163.050 886.200 ;
        RECT 166.950 884.100 169.050 886.200 ;
        RECT 161.400 883.350 162.600 884.100 ;
        RECT 167.400 883.350 168.600 884.100 ;
        RECT 97.950 880.950 100.050 883.050 ;
        RECT 119.100 880.950 121.200 883.050 ;
        RECT 137.100 880.950 139.200 883.050 ;
        RECT 155.100 880.950 157.200 883.050 ;
        RECT 160.500 880.950 162.600 883.050 ;
        RECT 166.950 880.950 169.050 883.050 ;
        RECT 98.400 879.900 99.600 880.650 ;
        RECT 119.400 879.900 120.600 880.650 ;
        RECT 97.950 877.800 100.050 879.900 ;
        RECT 118.950 877.800 121.050 879.900 ;
        RECT 173.250 878.400 174.450 891.300 ;
        RECT 184.800 880.950 186.900 883.050 ;
        RECT 91.650 871.500 95.850 872.700 ;
        RECT 91.650 870.600 93.750 871.500 ;
        RECT 76.350 867.600 78.450 869.700 ;
        RECT 119.400 853.050 120.450 877.800 ;
        RECT 172.350 876.300 174.450 878.400 ;
        RECT 142.950 871.950 145.050 874.050 ;
        RECT 118.950 850.950 121.050 853.050 ;
        RECT 76.950 847.950 79.050 850.050 ;
        RECT 100.950 847.950 103.050 850.050 ;
        RECT 28.950 838.950 31.050 841.050 ;
        RECT 34.950 839.100 37.050 841.200 ;
        RECT 40.950 839.100 43.050 841.200 ;
        RECT 52.950 840.450 55.050 841.200 ;
        RECT 77.400 840.600 78.450 847.950 ;
        RECT 101.400 840.600 102.450 847.950 ;
        RECT 56.400 840.450 57.600 840.600 ;
        RECT 52.950 839.400 57.600 840.450 ;
        RECT 52.950 839.100 55.050 839.400 ;
        RECT 25.950 826.950 28.050 829.050 ;
        RECT 26.400 814.050 27.450 826.950 ;
        RECT 19.950 811.950 22.050 814.050 ;
        RECT 25.950 811.950 28.050 814.050 ;
        RECT 13.950 806.100 16.050 808.200 ;
        RECT 20.400 807.600 21.450 811.950 ;
        RECT 14.400 805.350 15.600 806.100 ;
        RECT 20.400 805.350 21.600 807.600 ;
        RECT 13.950 802.950 16.050 805.050 ;
        RECT 16.950 802.950 19.050 805.050 ;
        RECT 19.950 802.950 22.050 805.050 ;
        RECT 22.950 802.950 25.050 805.050 ;
        RECT 17.400 801.900 18.600 802.650 ;
        RECT 16.950 799.800 19.050 801.900 ;
        RECT 23.400 800.400 24.600 802.650 ;
        RECT 29.400 801.900 30.450 838.950 ;
        RECT 35.400 838.350 36.600 839.100 ;
        RECT 41.400 838.350 42.600 839.100 ;
        RECT 56.400 838.350 57.600 839.400 ;
        RECT 77.400 838.350 78.600 840.600 ;
        RECT 101.400 838.350 102.600 840.600 ;
        RECT 118.950 839.100 121.050 841.200 ;
        RECT 127.950 839.100 130.050 841.200 ;
        RECT 133.950 839.100 136.050 841.200 ;
        RECT 34.950 835.950 37.050 838.050 ;
        RECT 37.950 835.950 40.050 838.050 ;
        RECT 40.950 835.950 43.050 838.050 ;
        RECT 55.950 835.950 58.050 838.050 ;
        RECT 58.950 835.950 61.050 838.050 ;
        RECT 61.950 835.950 64.050 838.050 ;
        RECT 76.950 835.950 79.050 838.050 ;
        RECT 79.950 835.950 82.050 838.050 ;
        RECT 82.950 835.950 85.050 838.050 ;
        RECT 85.950 835.950 88.050 838.050 ;
        RECT 100.950 835.950 103.050 838.050 ;
        RECT 103.950 835.950 106.050 838.050 ;
        RECT 106.950 835.950 109.050 838.050 ;
        RECT 109.950 835.950 112.050 838.050 ;
        RECT 38.400 833.400 39.600 835.650 ;
        RECT 59.400 833.400 60.600 835.650 ;
        RECT 80.400 834.900 81.600 835.650 ;
        RECT 38.400 820.050 39.450 833.400 ;
        RECT 37.950 817.950 40.050 820.050 ;
        RECT 52.950 811.950 55.050 814.050 ;
        RECT 31.950 805.950 34.050 808.050 ;
        RECT 37.950 806.100 40.050 808.200 ;
        RECT 43.950 806.100 46.050 808.200 ;
        RECT 13.950 761.100 16.050 763.200 ;
        RECT 14.400 760.350 15.600 761.100 ;
        RECT 13.950 757.950 16.050 760.050 ;
        RECT 16.950 757.950 19.050 760.050 ;
        RECT 17.400 755.400 18.600 757.650 ;
        RECT 17.400 742.050 18.450 755.400 ;
        RECT 16.950 739.950 19.050 742.050 ;
        RECT 19.950 729.000 22.050 733.050 ;
        RECT 23.400 730.050 24.450 800.400 ;
        RECT 28.950 799.800 31.050 801.900 ;
        RECT 32.400 796.050 33.450 805.950 ;
        RECT 38.400 805.350 39.600 806.100 ;
        RECT 44.400 805.350 45.600 806.100 ;
        RECT 37.950 802.950 40.050 805.050 ;
        RECT 40.950 802.950 43.050 805.050 ;
        RECT 43.950 802.950 46.050 805.050 ;
        RECT 46.950 802.950 49.050 805.050 ;
        RECT 34.950 799.950 37.050 802.050 ;
        RECT 41.400 801.000 42.600 802.650 ;
        RECT 31.950 793.950 34.050 796.050 ;
        RECT 35.400 769.050 36.450 799.950 ;
        RECT 40.950 796.950 43.050 801.000 ;
        RECT 47.400 800.400 48.600 802.650 ;
        RECT 47.400 799.050 48.450 800.400 ;
        RECT 46.950 798.450 49.050 799.050 ;
        RECT 44.400 797.400 49.050 798.450 ;
        RECT 37.950 795.450 40.050 796.050 ;
        RECT 44.400 795.450 45.450 797.400 ;
        RECT 46.950 796.950 49.050 797.400 ;
        RECT 37.950 794.400 45.450 795.450 ;
        RECT 37.950 793.950 40.050 794.400 ;
        RECT 34.950 766.950 37.050 769.050 ;
        RECT 40.950 766.950 43.050 769.050 ;
        RECT 34.950 761.100 37.050 763.200 ;
        RECT 41.400 762.600 42.450 766.950 ;
        RECT 35.400 760.350 36.600 761.100 ;
        RECT 41.400 760.350 42.600 762.600 ;
        RECT 34.950 757.950 37.050 760.050 ;
        RECT 37.950 757.950 40.050 760.050 ;
        RECT 40.950 757.950 43.050 760.050 ;
        RECT 43.950 757.950 46.050 760.050 ;
        RECT 38.400 755.400 39.600 757.650 ;
        RECT 44.400 756.900 45.600 757.650 ;
        RECT 53.400 756.900 54.450 811.950 ;
        RECT 59.400 808.200 60.450 833.400 ;
        RECT 79.950 832.800 82.050 834.900 ;
        RECT 86.400 833.400 87.600 835.650 ;
        RECT 104.400 834.900 105.600 835.650 ;
        RECT 80.400 829.050 81.450 832.800 ;
        RECT 79.950 826.950 82.050 829.050 ;
        RECT 76.950 811.950 79.050 814.050 ;
        RECT 58.950 806.100 61.050 808.200 ;
        RECT 67.950 806.100 70.050 808.200 ;
        RECT 73.950 806.100 76.050 808.200 ;
        RECT 77.400 808.050 78.450 811.950 ;
        RECT 86.400 811.050 87.450 833.400 ;
        RECT 103.950 832.800 106.050 834.900 ;
        RECT 110.400 833.400 111.600 835.650 ;
        RECT 110.400 829.050 111.450 833.400 ;
        RECT 109.950 826.950 112.050 829.050 ;
        RECT 103.950 823.950 106.050 826.050 ;
        RECT 91.950 817.950 94.050 820.050 ;
        RECT 92.400 811.050 93.450 817.950 ;
        RECT 94.950 814.950 97.050 817.050 ;
        RECT 95.400 811.050 96.450 814.950 ;
        RECT 104.400 811.050 105.450 823.950 ;
        RECT 119.400 823.050 120.450 839.100 ;
        RECT 128.400 838.350 129.600 839.100 ;
        RECT 134.400 838.350 135.600 839.100 ;
        RECT 127.950 835.950 130.050 838.050 ;
        RECT 130.950 835.950 133.050 838.050 ;
        RECT 133.950 835.950 136.050 838.050 ;
        RECT 136.950 835.950 139.050 838.050 ;
        RECT 131.400 833.400 132.600 835.650 ;
        RECT 137.400 834.900 138.600 835.650 ;
        RECT 127.950 826.950 130.050 829.050 ;
        RECT 118.950 820.950 121.050 823.050 ;
        RECT 85.950 808.950 88.050 811.050 ;
        RECT 91.950 808.950 94.050 811.050 ;
        RECT 68.400 805.350 69.600 806.100 ;
        RECT 74.400 805.350 75.600 806.100 ;
        RECT 76.950 805.950 79.050 808.050 ;
        RECT 82.950 805.950 85.050 808.050 ;
        RECT 87.000 807.900 90.000 808.050 ;
        RECT 85.950 807.600 90.000 807.900 ;
        RECT 85.950 805.950 90.600 807.600 ;
        RECT 94.950 807.000 97.050 811.050 ;
        RECT 103.950 808.950 106.050 811.050 ;
        RECT 64.950 802.950 67.050 805.050 ;
        RECT 67.950 802.950 70.050 805.050 ;
        RECT 70.950 802.950 73.050 805.050 ;
        RECT 73.950 802.950 76.050 805.050 ;
        RECT 65.400 801.000 66.600 802.650 ;
        RECT 71.400 801.000 72.600 802.650 ;
        RECT 64.950 796.950 67.050 801.000 ;
        RECT 70.950 796.950 73.050 801.000 ;
        RECT 79.950 796.950 82.050 799.050 ;
        RECT 76.950 787.950 79.050 790.050 ;
        RECT 67.950 761.100 70.050 763.200 ;
        RECT 77.400 762.600 78.450 787.950 ;
        RECT 68.400 760.350 69.600 761.100 ;
        RECT 77.400 760.350 78.600 762.600 ;
        RECT 61.800 757.950 63.900 760.050 ;
        RECT 67.950 757.950 70.050 760.050 ;
        RECT 70.950 757.950 73.050 760.050 ;
        RECT 76.500 757.950 78.600 760.050 ;
        RECT 38.400 748.050 39.450 755.400 ;
        RECT 43.950 754.800 46.050 756.900 ;
        RECT 52.950 754.800 55.050 756.900 ;
        RECT 62.400 755.400 63.600 757.650 ;
        RECT 71.400 756.900 72.600 757.650 ;
        RECT 37.950 745.950 40.050 748.050 ;
        RECT 58.950 739.950 61.050 742.050 ;
        RECT 31.350 735.300 33.450 737.400 ;
        RECT 49.050 735.300 51.150 737.400 ;
        RECT 20.400 727.350 21.600 729.000 ;
        RECT 22.950 727.950 25.050 730.050 ;
        RECT 25.950 729.000 28.050 733.050 ;
        RECT 26.400 727.350 27.600 729.000 ;
        RECT 14.100 724.950 16.200 727.050 ;
        RECT 19.500 724.950 21.600 727.050 ;
        RECT 25.950 724.950 28.050 727.050 ;
        RECT 22.950 721.950 25.050 724.050 ;
        RECT 32.250 722.400 33.450 735.300 ;
        RECT 43.800 724.950 45.900 727.050 ;
        RECT 23.400 700.050 24.450 721.950 ;
        RECT 31.350 720.300 33.450 722.400 ;
        RECT 32.250 713.700 33.450 720.300 ;
        RECT 49.650 716.700 50.850 735.300 ;
        RECT 52.950 724.950 55.050 727.050 ;
        RECT 46.650 715.500 50.850 716.700 ;
        RECT 53.400 722.400 54.600 724.650 ;
        RECT 59.400 723.900 60.450 739.950 ;
        RECT 46.650 714.600 48.750 715.500 ;
        RECT 31.350 711.600 33.450 713.700 ;
        RECT 13.950 697.950 16.050 700.050 ;
        RECT 22.950 697.950 25.050 700.050 ;
        RECT 14.400 685.200 15.450 697.950 ;
        RECT 13.950 683.100 16.050 685.200 ;
        RECT 37.950 683.100 40.050 685.200 ;
        RECT 43.950 683.100 46.050 685.200 ;
        RECT 14.400 682.350 15.600 683.100 ;
        RECT 38.400 682.350 39.600 683.100 ;
        RECT 44.400 682.350 45.600 683.100 ;
        RECT 13.950 679.950 16.050 682.050 ;
        RECT 16.950 679.950 19.050 682.050 ;
        RECT 19.950 679.950 22.050 682.050 ;
        RECT 22.950 679.950 25.050 682.050 ;
        RECT 37.950 679.950 40.050 682.050 ;
        RECT 40.950 679.950 43.050 682.050 ;
        RECT 43.950 679.950 46.050 682.050 ;
        RECT 46.950 679.950 49.050 682.050 ;
        RECT 23.400 677.400 24.600 679.650 ;
        RECT 23.400 664.050 24.450 677.400 ;
        RECT 25.950 676.950 28.050 679.050 ;
        RECT 34.950 676.950 37.050 679.050 ;
        RECT 41.400 677.400 42.600 679.650 ;
        RECT 47.400 678.900 48.600 679.650 ;
        RECT 26.400 670.050 27.450 676.950 ;
        RECT 25.950 667.950 28.050 670.050 ;
        RECT 31.950 667.950 34.050 670.050 ;
        RECT 22.950 661.950 25.050 664.050 ;
        RECT 22.950 650.100 25.050 652.200 ;
        RECT 23.400 649.350 24.600 650.100 ;
        RECT 13.950 646.950 16.050 649.050 ;
        RECT 16.950 646.950 19.050 649.050 ;
        RECT 19.950 646.950 22.050 649.050 ;
        RECT 22.950 646.950 25.050 649.050 ;
        RECT 14.400 644.400 15.600 646.650 ;
        RECT 14.400 634.050 15.450 644.400 ;
        RECT 13.950 631.950 16.050 634.050 ;
        RECT 32.400 633.450 33.450 667.950 ;
        RECT 35.400 651.450 36.450 676.950 ;
        RECT 41.400 673.050 42.450 677.400 ;
        RECT 46.950 676.800 49.050 678.900 ;
        RECT 53.400 678.450 54.450 722.400 ;
        RECT 58.950 721.800 61.050 723.900 ;
        RECT 55.950 679.950 58.050 682.050 ;
        RECT 50.400 677.400 54.450 678.450 ;
        RECT 40.950 670.950 43.050 673.050 ;
        RECT 37.950 655.950 40.050 658.050 ;
        RECT 38.400 652.200 39.450 655.950 ;
        RECT 37.950 651.450 40.050 652.200 ;
        RECT 35.400 650.400 40.050 651.450 ;
        RECT 37.950 650.100 40.050 650.400 ;
        RECT 38.400 649.350 39.600 650.100 ;
        RECT 37.950 646.950 40.050 649.050 ;
        RECT 40.950 646.950 43.050 649.050 ;
        RECT 41.400 645.900 42.600 646.650 ;
        RECT 40.950 643.800 43.050 645.900 ;
        RECT 50.400 645.450 51.450 677.400 ;
        RECT 56.400 664.050 57.450 679.950 ;
        RECT 59.400 673.050 60.450 721.800 ;
        RECT 62.400 718.050 63.450 755.400 ;
        RECT 70.950 754.800 73.050 756.900 ;
        RECT 80.400 754.050 81.450 796.950 ;
        RECT 79.950 751.950 82.050 754.050 ;
        RECT 73.950 733.950 76.050 736.050 ;
        RECT 74.400 729.600 75.450 733.950 ;
        RECT 83.400 733.050 84.450 805.950 ;
        RECT 85.950 805.800 88.050 805.950 ;
        RECT 89.400 805.350 90.600 805.950 ;
        RECT 95.400 805.350 96.600 807.000 ;
        RECT 88.950 802.950 91.050 805.050 ;
        RECT 91.950 802.950 94.050 805.050 ;
        RECT 94.950 802.950 97.050 805.050 ;
        RECT 97.950 802.950 100.050 805.050 ;
        RECT 92.400 801.900 93.600 802.650 ;
        RECT 98.400 801.900 99.600 802.650 ;
        RECT 104.400 801.900 105.450 808.950 ;
        RECT 119.400 808.200 120.450 820.950 ;
        RECT 124.950 814.950 127.050 817.050 ;
        RECT 106.950 805.950 109.050 808.050 ;
        RECT 112.950 806.100 115.050 808.200 ;
        RECT 118.950 806.100 121.050 808.200 ;
        RECT 125.400 807.450 126.450 814.950 ;
        RECT 128.400 814.050 129.450 826.950 ;
        RECT 131.400 826.050 132.450 833.400 ;
        RECT 136.950 832.800 139.050 834.900 ;
        RECT 143.400 829.050 144.450 871.950 ;
        RECT 173.250 869.700 174.450 876.300 ;
        RECT 190.650 872.700 191.850 891.300 ;
        RECT 193.950 880.950 196.050 883.050 ;
        RECT 202.950 880.950 205.050 883.050 ;
        RECT 194.400 879.900 195.600 880.650 ;
        RECT 203.400 879.900 204.600 880.650 ;
        RECT 193.950 877.800 196.050 879.900 ;
        RECT 202.950 877.800 205.050 879.900 ;
        RECT 203.400 874.050 204.450 877.800 ;
        RECT 187.650 871.500 191.850 872.700 ;
        RECT 202.950 871.950 205.050 874.050 ;
        RECT 207.150 872.700 208.350 891.300 ;
        RECT 212.100 880.950 214.200 883.050 ;
        RECT 212.400 879.000 213.600 880.650 ;
        RECT 211.950 874.950 214.050 879.000 ;
        RECT 224.550 878.400 225.750 891.300 ;
        RECT 229.950 884.100 232.050 886.200 ;
        RECT 247.950 884.100 250.050 886.200 ;
        RECT 272.400 885.450 273.600 885.600 ;
        RECT 272.400 884.400 279.450 885.450 ;
        RECT 230.400 883.350 231.600 884.100 ;
        RECT 248.400 883.350 249.600 884.100 ;
        RECT 272.400 883.350 273.600 884.400 ;
        RECT 229.950 880.950 232.050 883.050 ;
        RECT 248.400 880.950 250.500 883.050 ;
        RECT 253.800 880.950 255.900 883.050 ;
        RECT 268.950 880.950 271.050 883.050 ;
        RECT 271.950 880.950 274.050 883.050 ;
        RECT 269.400 878.400 270.600 880.650 ;
        RECT 224.550 876.300 226.650 878.400 ;
        RECT 187.650 870.600 189.750 871.500 ;
        RECT 172.350 867.600 174.450 869.700 ;
        RECT 203.400 853.050 204.450 871.950 ;
        RECT 207.150 871.500 211.350 872.700 ;
        RECT 209.250 870.600 211.350 871.500 ;
        RECT 224.550 869.700 225.750 876.300 ;
        RECT 247.950 874.950 250.050 877.050 ;
        RECT 224.550 867.600 226.650 869.700 ;
        RECT 166.350 849.300 168.450 851.400 ;
        RECT 187.950 850.950 190.050 853.050 ;
        RECT 202.950 850.950 205.050 853.050 ;
        RECT 145.950 844.950 148.050 847.050 ;
        RECT 146.400 835.050 147.450 844.950 ;
        RECT 167.250 842.700 168.450 849.300 ;
        RECT 181.650 847.500 183.750 848.400 ;
        RECT 181.650 846.300 185.850 847.500 ;
        RECT 151.950 839.100 154.050 841.200 ;
        RECT 166.350 840.600 168.450 842.700 ;
        RECT 152.400 838.350 153.600 839.100 ;
        RECT 151.950 835.950 154.050 838.050 ;
        RECT 154.950 835.950 157.050 838.050 ;
        RECT 160.950 835.950 163.050 838.050 ;
        RECT 145.950 832.950 148.050 835.050 ;
        RECT 155.400 833.400 156.600 835.650 ;
        RECT 161.400 833.400 162.600 835.650 ;
        RECT 142.950 826.950 145.050 829.050 ;
        RECT 130.950 823.950 133.050 826.050 ;
        RECT 145.950 820.950 148.050 823.050 ;
        RECT 127.950 811.950 130.050 814.050 ;
        RECT 125.400 806.400 129.450 807.450 ;
        RECT 91.950 799.800 94.050 801.900 ;
        RECT 97.950 799.800 100.050 801.900 ;
        RECT 103.950 799.800 106.050 801.900 ;
        RECT 85.950 793.950 88.050 796.050 ;
        RECT 86.400 757.050 87.450 793.950 ;
        RECT 88.950 761.100 91.050 763.200 ;
        RECT 97.950 761.100 100.050 763.200 ;
        RECT 103.950 761.100 106.050 763.200 ;
        RECT 107.400 763.050 108.450 805.950 ;
        RECT 113.400 805.350 114.600 806.100 ;
        RECT 119.400 805.350 120.600 806.100 ;
        RECT 112.950 802.950 115.050 805.050 ;
        RECT 115.950 802.950 118.050 805.050 ;
        RECT 118.950 802.950 121.050 805.050 ;
        RECT 121.950 802.950 124.050 805.050 ;
        RECT 116.400 801.900 117.600 802.650 ;
        RECT 122.400 801.900 123.600 802.650 ;
        RECT 128.400 801.900 129.450 806.400 ;
        RECT 130.950 806.100 133.050 808.200 ;
        RECT 136.950 806.100 139.050 808.200 ;
        RECT 115.950 799.800 118.050 801.900 ;
        RECT 121.950 799.800 124.050 801.900 ;
        RECT 127.950 799.800 130.050 801.900 ;
        RECT 131.400 799.050 132.450 806.100 ;
        RECT 137.400 805.350 138.600 806.100 ;
        RECT 136.950 802.950 139.050 805.050 ;
        RECT 139.950 802.950 142.050 805.050 ;
        RECT 140.400 801.900 141.600 802.650 ;
        RECT 146.400 802.050 147.450 820.950 ;
        RECT 155.400 817.050 156.450 833.400 ;
        RECT 161.400 829.050 162.450 833.400 ;
        RECT 160.950 826.950 163.050 829.050 ;
        RECT 167.250 827.700 168.450 840.600 ;
        RECT 178.950 839.100 181.050 841.200 ;
        RECT 179.400 838.350 180.600 839.100 ;
        RECT 178.800 835.950 180.900 838.050 ;
        RECT 178.950 829.950 181.050 832.050 ;
        RECT 166.350 825.600 168.450 827.700 ;
        RECT 172.950 820.950 175.050 823.050 ;
        RECT 154.950 814.950 157.050 817.050 ;
        RECT 169.950 814.950 172.050 817.050 ;
        RECT 148.950 811.950 151.050 814.050 ;
        RECT 139.950 799.800 142.050 801.900 ;
        RECT 145.800 799.950 147.900 802.050 ;
        RECT 149.400 801.900 150.450 811.950 ;
        RECT 154.950 806.100 157.050 808.200 ;
        RECT 160.950 806.100 163.050 808.200 ;
        RECT 155.400 805.350 156.600 806.100 ;
        RECT 161.400 805.350 162.600 806.100 ;
        RECT 154.950 802.950 157.050 805.050 ;
        RECT 157.950 802.950 160.050 805.050 ;
        RECT 160.950 802.950 163.050 805.050 ;
        RECT 163.950 802.950 166.050 805.050 ;
        RECT 158.400 801.900 159.600 802.650 ;
        RECT 148.950 799.800 151.050 801.900 ;
        RECT 157.950 799.800 160.050 801.900 ;
        RECT 164.400 801.450 165.600 802.650 ;
        RECT 170.400 801.450 171.450 814.950 ;
        RECT 164.400 800.400 171.450 801.450 ;
        RECT 130.950 796.950 133.050 799.050 ;
        RECT 173.400 796.050 174.450 820.950 ;
        RECT 175.950 814.950 178.050 817.050 ;
        RECT 176.400 808.050 177.450 814.950 ;
        RECT 179.400 811.050 180.450 829.950 ;
        RECT 184.650 827.700 185.850 846.300 ;
        RECT 188.400 840.600 189.450 850.950 ;
        RECT 208.950 844.950 211.050 847.050 ;
        RECT 235.950 844.950 238.050 847.050 ;
        RECT 209.400 840.600 210.450 844.950 ;
        RECT 188.400 838.350 189.600 840.600 ;
        RECT 209.400 838.350 210.600 840.600 ;
        RECT 214.950 839.100 217.050 841.200 ;
        RECT 223.950 839.100 226.050 841.200 ;
        RECT 229.950 839.100 232.050 841.200 ;
        RECT 236.400 840.600 237.450 844.950 ;
        RECT 215.400 838.350 216.600 839.100 ;
        RECT 187.950 835.950 190.050 838.050 ;
        RECT 205.950 835.950 208.050 838.050 ;
        RECT 208.950 835.950 211.050 838.050 ;
        RECT 211.950 835.950 214.050 838.050 ;
        RECT 214.950 835.950 217.050 838.050 ;
        RECT 206.400 833.400 207.600 835.650 ;
        RECT 212.400 833.400 213.600 835.650 ;
        RECT 184.050 825.600 186.150 827.700 ;
        RECT 181.950 820.950 184.050 823.050 ;
        RECT 178.950 808.950 181.050 811.050 ;
        RECT 175.950 805.950 178.050 808.050 ;
        RECT 182.400 807.600 183.450 820.950 ;
        RECT 206.400 814.050 207.450 833.400 ;
        RECT 212.400 823.050 213.450 833.400 ;
        RECT 224.400 823.050 225.450 839.100 ;
        RECT 230.400 838.350 231.600 839.100 ;
        RECT 236.400 838.350 237.600 840.600 ;
        RECT 248.400 838.050 249.450 874.950 ;
        RECT 262.950 844.950 265.050 847.050 ;
        RECT 256.950 839.100 259.050 841.200 ;
        RECT 263.400 840.600 264.450 844.950 ;
        RECT 269.400 841.200 270.450 878.400 ;
        RECT 278.400 856.050 279.450 884.400 ;
        RECT 280.950 884.100 283.050 886.200 ;
        RECT 286.950 884.100 289.050 886.200 ;
        RECT 281.400 868.050 282.450 884.100 ;
        RECT 287.400 883.350 288.600 884.100 ;
        RECT 286.950 880.950 289.050 883.050 ;
        RECT 289.950 880.950 292.050 883.050 ;
        RECT 295.950 880.950 298.050 883.050 ;
        RECT 290.400 879.000 291.600 880.650 ;
        RECT 289.950 874.950 292.050 879.000 ;
        RECT 296.400 878.400 297.600 880.650 ;
        RECT 296.400 874.050 297.450 878.400 ;
        RECT 295.950 871.950 298.050 874.050 ;
        RECT 300.150 872.700 301.350 891.300 ;
        RECT 305.100 880.950 307.200 883.050 ;
        RECT 305.400 878.400 306.600 880.650 ;
        RECT 317.550 878.400 318.750 891.300 ;
        RECT 322.950 884.100 325.050 886.200 ;
        RECT 343.950 884.100 346.050 886.200 ;
        RECT 323.400 883.350 324.600 884.100 ;
        RECT 344.400 883.350 345.600 884.100 ;
        RECT 361.950 883.950 364.050 886.050 ;
        RECT 367.950 884.100 370.050 886.200 ;
        RECT 322.950 880.950 325.050 883.050 ;
        RECT 344.400 880.950 346.500 883.050 ;
        RECT 349.800 880.950 351.900 883.050 ;
        RECT 305.400 876.450 306.450 878.400 ;
        RECT 305.400 875.400 309.450 876.450 ;
        RECT 300.150 871.500 304.350 872.700 ;
        RECT 302.250 870.600 304.350 871.500 ;
        RECT 280.950 865.950 283.050 868.050 ;
        RECT 289.950 865.950 292.050 868.050 ;
        RECT 277.950 853.950 280.050 856.050 ;
        RECT 290.400 847.050 291.450 865.950 ;
        RECT 298.950 853.950 301.050 856.050 ;
        RECT 289.950 844.950 292.050 847.050 ;
        RECT 257.400 838.350 258.600 839.100 ;
        RECT 263.400 838.350 264.600 840.600 ;
        RECT 268.950 839.100 271.050 841.200 ;
        RECT 283.950 839.100 286.050 841.200 ;
        RECT 290.400 840.600 291.450 844.950 ;
        RECT 284.400 838.350 285.600 839.100 ;
        RECT 290.400 838.350 291.600 840.600 ;
        RECT 295.950 839.100 298.050 841.200 ;
        RECT 229.950 835.950 232.050 838.050 ;
        RECT 232.950 835.950 235.050 838.050 ;
        RECT 235.950 835.950 238.050 838.050 ;
        RECT 238.950 835.950 241.050 838.050 ;
        RECT 247.950 835.950 250.050 838.050 ;
        RECT 253.950 835.950 256.050 838.050 ;
        RECT 256.950 835.950 259.050 838.050 ;
        RECT 259.950 835.950 262.050 838.050 ;
        RECT 262.950 835.950 265.050 838.050 ;
        RECT 280.950 835.950 283.050 838.050 ;
        RECT 283.950 835.950 286.050 838.050 ;
        RECT 286.950 835.950 289.050 838.050 ;
        RECT 289.950 835.950 292.050 838.050 ;
        RECT 233.400 834.900 234.600 835.650 ;
        RECT 232.950 832.800 235.050 834.900 ;
        RECT 239.400 833.400 240.600 835.650 ;
        RECT 254.400 834.900 255.600 835.650 ;
        RECT 211.950 820.950 214.050 823.050 ;
        RECT 223.950 820.950 226.050 823.050 ;
        RECT 190.950 811.950 193.050 814.050 ;
        RECT 205.950 811.950 208.050 814.050 ;
        RECT 182.400 805.350 183.600 807.600 ;
        RECT 179.100 802.950 181.200 805.050 ;
        RECT 182.400 802.950 184.500 805.050 ;
        RECT 187.800 802.950 189.900 805.050 ;
        RECT 179.400 801.900 180.600 802.650 ;
        RECT 178.950 799.800 181.050 801.900 ;
        RECT 188.400 800.400 189.600 802.650 ;
        RECT 188.400 796.050 189.450 800.400 ;
        RECT 172.950 793.950 175.050 796.050 ;
        RECT 187.950 793.950 190.050 796.050 ;
        RECT 130.950 772.950 133.050 775.050 ;
        RECT 139.950 772.950 142.050 775.050 ;
        RECT 85.950 754.950 88.050 757.050 ;
        RECT 89.400 739.050 90.450 761.100 ;
        RECT 98.400 760.350 99.600 761.100 ;
        RECT 104.400 760.350 105.600 761.100 ;
        RECT 106.950 760.950 109.050 763.050 ;
        RECT 109.950 761.100 112.050 763.200 ;
        RECT 94.950 757.950 97.050 760.050 ;
        RECT 97.950 757.950 100.050 760.050 ;
        RECT 100.950 757.950 103.050 760.050 ;
        RECT 103.950 757.950 106.050 760.050 ;
        RECT 95.400 755.400 96.600 757.650 ;
        RECT 101.400 756.900 102.600 757.650 ;
        RECT 95.400 739.050 96.450 755.400 ;
        RECT 100.950 754.800 103.050 756.900 ;
        RECT 88.950 736.950 91.050 739.050 ;
        RECT 94.950 736.950 97.050 739.050 ;
        RECT 97.950 733.950 100.050 736.050 ;
        RECT 82.950 730.950 85.050 733.050 ;
        RECT 88.950 730.950 91.050 733.050 ;
        RECT 74.400 727.350 75.600 729.600 ;
        RECT 80.400 729.450 81.600 729.600 ;
        RECT 80.400 728.400 87.450 729.450 ;
        RECT 80.400 727.350 81.600 728.400 ;
        RECT 70.950 724.950 73.050 727.050 ;
        RECT 73.950 724.950 76.050 727.050 ;
        RECT 76.950 724.950 79.050 727.050 ;
        RECT 79.950 724.950 82.050 727.050 ;
        RECT 71.400 723.900 72.600 724.650 ;
        RECT 77.400 723.900 78.600 724.650 ;
        RECT 70.950 721.800 73.050 723.900 ;
        RECT 76.950 721.800 79.050 723.900 ;
        RECT 61.950 715.950 64.050 718.050 ;
        RECT 71.400 715.050 72.450 721.800 ;
        RECT 82.950 718.950 85.050 721.050 ;
        RECT 83.400 715.050 84.450 718.950 ;
        RECT 86.400 715.050 87.450 728.400 ;
        RECT 89.400 723.900 90.450 730.950 ;
        RECT 98.400 729.600 99.450 733.950 ;
        RECT 98.400 727.350 99.600 729.600 ;
        RECT 103.950 728.100 106.050 730.200 ;
        RECT 104.400 727.350 105.600 728.100 ;
        RECT 94.950 724.950 97.050 727.050 ;
        RECT 97.950 724.950 100.050 727.050 ;
        RECT 100.950 724.950 103.050 727.050 ;
        RECT 103.950 724.950 106.050 727.050 ;
        RECT 95.400 723.900 96.600 724.650 ;
        RECT 88.950 721.800 91.050 723.900 ;
        RECT 94.950 721.800 97.050 723.900 ;
        RECT 101.400 723.000 102.600 724.650 ;
        RECT 100.950 718.950 103.050 723.000 ;
        RECT 110.400 718.050 111.450 761.100 ;
        RECT 112.950 760.950 115.050 763.050 ;
        RECT 121.950 761.100 124.050 763.200 ;
        RECT 113.400 736.050 114.450 760.950 ;
        RECT 122.400 760.350 123.600 761.100 ;
        RECT 118.950 757.950 121.050 760.050 ;
        RECT 121.950 757.950 124.050 760.050 ;
        RECT 124.950 757.950 127.050 760.050 ;
        RECT 119.400 756.900 120.600 757.650 ;
        RECT 118.950 754.800 121.050 756.900 ;
        RECT 125.400 756.450 126.600 757.650 ;
        RECT 131.400 756.900 132.450 772.950 ;
        RECT 140.400 762.600 141.450 772.950 ;
        RECT 166.950 766.950 169.050 769.050 ;
        RECT 181.950 766.950 184.050 769.050 ;
        RECT 140.400 760.350 141.600 762.600 ;
        RECT 148.950 760.950 151.050 763.050 ;
        RECT 160.950 761.100 163.050 763.200 ;
        RECT 167.400 762.600 168.450 766.950 ;
        RECT 182.400 762.600 183.450 766.950 ;
        RECT 191.400 765.450 192.450 811.950 ;
        RECT 202.950 806.100 205.050 808.200 ;
        RECT 208.950 806.100 211.050 808.200 ;
        RECT 203.400 805.350 204.600 806.100 ;
        RECT 209.400 805.350 210.600 806.100 ;
        RECT 217.950 805.950 220.050 808.050 ;
        RECT 229.950 806.100 232.050 808.200 ;
        RECT 202.950 802.950 205.050 805.050 ;
        RECT 205.950 802.950 208.050 805.050 ;
        RECT 208.950 802.950 211.050 805.050 ;
        RECT 211.950 802.950 214.050 805.050 ;
        RECT 199.950 799.950 202.050 802.050 ;
        RECT 206.400 800.400 207.600 802.650 ;
        RECT 212.400 801.900 213.600 802.650 ;
        RECT 200.400 775.050 201.450 799.950 ;
        RECT 199.950 772.950 202.050 775.050 ;
        RECT 206.400 766.200 207.450 800.400 ;
        RECT 211.950 799.800 214.050 801.900 ;
        RECT 212.400 796.050 213.450 799.800 ;
        RECT 211.950 793.950 214.050 796.050 ;
        RECT 218.400 784.050 219.450 805.950 ;
        RECT 230.400 805.350 231.600 806.100 ;
        RECT 235.950 805.950 238.050 808.050 ;
        RECT 226.950 802.950 229.050 805.050 ;
        RECT 229.950 802.950 232.050 805.050 ;
        RECT 227.400 801.900 228.600 802.650 ;
        RECT 226.950 799.800 229.050 801.900 ;
        RECT 232.950 799.950 235.050 802.050 ;
        RECT 233.400 796.050 234.450 799.950 ;
        RECT 232.950 793.950 235.050 796.050 ;
        RECT 233.400 790.050 234.450 793.950 ;
        RECT 232.950 787.950 235.050 790.050 ;
        RECT 217.950 781.950 220.050 784.050 ;
        RECT 232.950 778.950 235.050 781.050 ;
        RECT 223.950 775.950 226.050 778.050 ;
        RECT 188.400 764.400 192.450 765.450 ;
        RECT 188.400 763.200 189.450 764.400 ;
        RECT 199.950 763.950 202.050 766.050 ;
        RECT 205.950 764.100 208.050 766.200 ;
        RECT 139.950 757.950 142.050 760.050 ;
        RECT 142.950 757.950 145.050 760.050 ;
        RECT 125.400 755.400 129.450 756.450 ;
        RECT 124.950 751.950 127.050 754.050 ;
        RECT 112.950 733.950 115.050 736.050 ;
        RECT 112.950 727.950 115.050 730.050 ;
        RECT 125.400 729.600 126.450 751.950 ;
        RECT 128.400 745.050 129.450 755.400 ;
        RECT 130.950 754.800 133.050 756.900 ;
        RECT 143.400 755.400 144.600 757.650 ;
        RECT 136.950 748.950 139.050 751.050 ;
        RECT 127.950 742.950 130.050 745.050 ;
        RECT 94.950 715.950 97.050 718.050 ;
        RECT 109.950 715.950 112.050 718.050 ;
        RECT 70.950 712.950 73.050 715.050 ;
        RECT 82.800 712.950 84.900 715.050 ;
        RECT 85.950 712.950 88.050 715.050 ;
        RECT 88.950 683.100 91.050 685.200 ;
        RECT 89.400 682.350 90.600 683.100 ;
        RECT 64.950 679.950 67.050 682.050 ;
        RECT 67.950 679.950 70.050 682.050 ;
        RECT 70.950 679.950 73.050 682.050 ;
        RECT 85.950 679.950 88.050 682.050 ;
        RECT 88.950 679.950 91.050 682.050 ;
        RECT 68.400 678.900 69.600 679.650 ;
        RECT 86.400 678.900 87.600 679.650 ;
        RECT 67.950 676.800 70.050 678.900 ;
        RECT 85.950 676.800 88.050 678.900 ;
        RECT 58.950 670.950 61.050 673.050 ;
        RECT 55.950 661.950 58.050 664.050 ;
        RECT 56.400 651.600 57.450 661.950 ;
        RECT 56.400 649.350 57.600 651.600 ;
        RECT 61.950 650.100 64.050 652.200 ;
        RECT 68.400 651.450 69.450 676.800 ;
        RECT 79.950 661.950 82.050 664.050 ;
        RECT 80.400 651.600 81.450 661.950 ;
        RECT 68.400 650.400 72.450 651.450 ;
        RECT 62.400 649.350 63.600 650.100 ;
        RECT 55.950 646.950 58.050 649.050 ;
        RECT 58.950 646.950 61.050 649.050 ;
        RECT 61.950 646.950 64.050 649.050 ;
        RECT 64.950 646.950 67.050 649.050 ;
        RECT 59.400 645.900 60.600 646.650 ;
        RECT 65.400 645.900 66.600 646.650 ;
        RECT 71.400 645.900 72.450 650.400 ;
        RECT 80.400 649.350 81.600 651.600 ;
        RECT 91.950 649.950 94.050 652.050 ;
        RECT 79.950 646.950 82.050 649.050 ;
        RECT 82.950 646.950 85.050 649.050 ;
        RECT 50.400 644.400 54.450 645.450 ;
        RECT 34.950 633.450 37.050 634.050 ;
        RECT 32.400 632.400 37.050 633.450 ;
        RECT 34.950 631.950 37.050 632.400 ;
        RECT 31.350 615.300 33.450 617.400 ;
        RECT 32.250 608.700 33.450 615.300 ;
        RECT 31.350 606.600 33.450 608.700 ;
        RECT 14.100 601.950 16.200 604.050 ;
        RECT 19.500 601.950 21.600 604.050 ;
        RECT 25.950 601.950 28.050 604.050 ;
        RECT 20.400 600.450 21.600 601.650 ;
        RECT 26.400 600.450 27.600 601.650 ;
        RECT 20.400 599.400 27.600 600.450 ;
        RECT 32.250 593.700 33.450 606.600 ;
        RECT 31.350 591.600 33.450 593.700 ;
        RECT 25.950 586.950 28.050 589.050 ;
        RECT 19.950 577.950 22.050 580.050 ;
        RECT 20.400 573.600 21.450 577.950 ;
        RECT 26.400 573.600 27.450 586.950 ;
        RECT 31.350 579.300 33.450 581.400 ;
        RECT 20.400 571.350 21.600 573.600 ;
        RECT 26.400 571.350 27.600 573.600 ;
        RECT 14.100 568.950 16.200 571.050 ;
        RECT 19.500 568.950 21.600 571.050 ;
        RECT 25.950 568.950 28.050 571.050 ;
        RECT 32.250 566.400 33.450 579.300 ;
        RECT 31.350 564.300 33.450 566.400 ;
        RECT 32.250 557.700 33.450 564.300 ;
        RECT 31.350 555.600 33.450 557.700 ;
        RECT 31.350 537.300 33.450 539.400 ;
        RECT 32.250 530.700 33.450 537.300 ;
        RECT 31.350 528.600 33.450 530.700 ;
        RECT 14.100 523.950 16.200 526.050 ;
        RECT 19.500 523.950 21.600 526.050 ;
        RECT 25.950 523.950 28.050 526.050 ;
        RECT 20.400 522.900 21.600 523.650 ;
        RECT 26.400 522.900 27.600 523.650 ;
        RECT 19.950 520.800 22.050 522.900 ;
        RECT 25.950 520.800 28.050 522.900 ;
        RECT 32.250 515.700 33.450 528.600 ;
        RECT 31.350 513.600 33.450 515.700 ;
        RECT 35.400 508.050 36.450 631.950 ;
        RECT 46.650 613.500 48.750 614.400 ;
        RECT 46.650 612.300 50.850 613.500 ;
        RECT 53.400 613.050 54.450 644.400 ;
        RECT 58.950 643.800 61.050 645.900 ;
        RECT 64.950 643.800 67.050 645.900 ;
        RECT 70.950 643.800 73.050 645.900 ;
        RECT 83.400 644.400 84.600 646.650 ;
        RECT 92.400 645.900 93.450 649.950 ;
        RECT 83.400 643.050 84.450 644.400 ;
        RECT 91.950 643.800 94.050 645.900 ;
        RECT 83.400 641.400 88.050 643.050 ;
        RECT 84.000 640.950 88.050 641.400 ;
        RECT 95.400 613.050 96.450 715.950 ;
        RECT 100.950 712.950 103.050 715.050 ;
        RECT 97.950 682.950 100.050 685.050 ;
        RECT 98.400 652.050 99.450 682.950 ;
        RECT 101.400 678.900 102.450 712.950 ;
        RECT 113.400 700.050 114.450 727.950 ;
        RECT 125.400 727.350 126.600 729.600 ;
        RECT 121.950 724.950 124.050 727.050 ;
        RECT 124.950 724.950 127.050 727.050 ;
        RECT 127.950 724.950 130.050 727.050 ;
        RECT 112.950 697.950 115.050 700.050 ;
        RECT 133.950 688.950 136.050 691.050 ;
        RECT 109.950 683.100 112.050 685.200 ;
        RECT 127.950 683.100 130.050 688.050 ;
        RECT 134.400 684.600 135.450 688.950 ;
        RECT 137.400 685.050 138.450 748.950 ;
        RECT 143.400 742.050 144.450 755.400 ;
        RECT 145.950 748.950 148.050 751.050 ;
        RECT 142.950 739.950 145.050 742.050 ;
        RECT 146.400 729.600 147.450 748.950 ;
        RECT 149.400 748.050 150.450 760.950 ;
        RECT 161.400 760.350 162.600 761.100 ;
        RECT 167.400 760.350 168.600 762.600 ;
        RECT 182.400 760.350 183.600 762.600 ;
        RECT 187.950 761.100 190.050 763.200 ;
        RECT 188.400 760.350 189.600 761.100 ;
        RECT 157.950 757.950 160.050 760.050 ;
        RECT 160.950 757.950 163.050 760.050 ;
        RECT 163.950 757.950 166.050 760.050 ;
        RECT 166.950 757.950 169.050 760.050 ;
        RECT 181.950 757.950 184.050 760.050 ;
        RECT 184.950 757.950 187.050 760.050 ;
        RECT 187.950 757.950 190.050 760.050 ;
        RECT 190.950 757.950 193.050 760.050 ;
        RECT 158.400 755.400 159.600 757.650 ;
        RECT 164.400 756.900 165.600 757.650 ;
        RECT 148.950 745.950 151.050 748.050 ;
        RECT 146.400 727.350 147.600 729.600 ;
        RECT 151.950 728.100 154.050 730.200 ;
        RECT 152.400 727.350 153.600 728.100 ;
        RECT 142.950 724.950 145.050 727.050 ;
        RECT 145.950 724.950 148.050 727.050 ;
        RECT 148.950 724.950 151.050 727.050 ;
        RECT 151.950 724.950 154.050 727.050 ;
        RECT 143.400 722.400 144.600 724.650 ;
        RECT 149.400 722.400 150.600 724.650 ;
        RECT 143.400 715.050 144.450 722.400 ;
        RECT 142.950 712.950 145.050 715.050 ;
        RECT 143.400 703.050 144.450 712.950 ;
        RECT 145.950 703.950 148.050 706.050 ;
        RECT 142.950 700.950 145.050 703.050 ;
        RECT 146.400 700.050 147.450 703.950 ;
        RECT 139.950 697.950 142.050 700.050 ;
        RECT 110.400 682.350 111.600 683.100 ;
        RECT 128.400 682.350 129.600 683.100 ;
        RECT 134.400 682.350 135.600 684.600 ;
        RECT 136.950 682.950 139.050 685.050 ;
        RECT 106.950 679.950 109.050 682.050 ;
        RECT 109.950 679.950 112.050 682.050 ;
        RECT 124.950 679.950 127.050 682.050 ;
        RECT 127.950 679.950 130.050 682.050 ;
        RECT 130.950 679.950 133.050 682.050 ;
        RECT 133.950 679.950 136.050 682.050 ;
        RECT 107.400 678.900 108.600 679.650 ;
        RECT 100.950 676.800 103.050 678.900 ;
        RECT 106.950 676.800 109.050 678.900 ;
        RECT 125.400 677.400 126.600 679.650 ;
        RECT 131.400 678.900 132.600 679.650 ;
        RECT 125.400 673.050 126.450 677.400 ;
        RECT 130.950 676.800 133.050 678.900 ;
        RECT 140.400 673.050 141.450 697.950 ;
        RECT 142.950 697.800 145.050 699.900 ;
        RECT 145.950 697.950 148.050 700.050 ;
        RECT 143.400 678.900 144.450 697.800 ;
        RECT 149.400 691.050 150.450 722.400 ;
        RECT 158.400 715.050 159.450 755.400 ;
        RECT 163.950 754.800 166.050 756.900 ;
        RECT 185.400 755.400 186.600 757.650 ;
        RECT 191.400 755.400 192.600 757.650 ;
        RECT 185.400 751.050 186.450 755.400 ;
        RECT 184.950 748.950 187.050 751.050 ;
        RECT 160.950 739.950 163.050 742.050 ;
        RECT 161.400 724.050 162.450 739.950 ;
        RECT 169.950 736.950 172.050 739.050 ;
        RECT 170.400 729.600 171.450 736.950 ;
        RECT 191.400 736.050 192.450 755.400 ;
        RECT 200.400 745.050 201.450 763.950 ;
        RECT 205.950 760.950 208.050 763.050 ;
        RECT 211.950 762.000 214.050 766.050 ;
        RECT 206.400 760.350 207.600 760.950 ;
        RECT 212.400 760.350 213.600 762.000 ;
        RECT 205.950 757.950 208.050 760.050 ;
        RECT 208.950 757.950 211.050 760.050 ;
        RECT 211.950 757.950 214.050 760.050 ;
        RECT 214.950 757.950 217.050 760.050 ;
        RECT 209.400 756.900 210.600 757.650 ;
        RECT 215.400 756.900 216.600 757.650 ;
        RECT 224.400 757.050 225.450 775.950 ;
        RECT 233.400 762.600 234.450 778.950 ;
        RECT 236.400 769.050 237.450 805.950 ;
        RECT 235.950 766.950 238.050 769.050 ;
        RECT 239.400 766.050 240.450 833.400 ;
        RECT 253.950 832.800 256.050 834.900 ;
        RECT 260.400 833.400 261.600 835.650 ;
        RECT 281.400 833.400 282.600 835.650 ;
        RECT 287.400 833.400 288.600 835.650 ;
        RECT 260.400 820.050 261.450 833.400 ;
        RECT 259.950 817.950 262.050 820.050 ;
        RECT 259.950 814.800 262.050 816.900 ;
        RECT 265.950 814.950 268.050 817.050 ;
        RECT 250.950 811.950 253.050 814.050 ;
        RECT 244.950 806.100 247.050 808.200 ;
        RECT 251.400 807.600 252.450 811.950 ;
        RECT 245.400 805.350 246.600 806.100 ;
        RECT 251.400 805.350 252.600 807.600 ;
        RECT 244.950 802.950 247.050 805.050 ;
        RECT 247.950 802.950 250.050 805.050 ;
        RECT 250.950 802.950 253.050 805.050 ;
        RECT 253.950 802.950 256.050 805.050 ;
        RECT 248.400 800.400 249.600 802.650 ;
        RECT 254.400 801.900 255.600 802.650 ;
        RECT 260.400 801.900 261.450 814.800 ;
        RECT 262.950 805.950 265.050 808.050 ;
        RECT 241.950 796.950 244.050 799.050 ;
        RECT 242.400 781.050 243.450 796.950 ;
        RECT 248.400 793.050 249.450 800.400 ;
        RECT 253.950 799.800 256.050 801.900 ;
        RECT 259.950 799.800 262.050 801.900 ;
        RECT 263.400 799.050 264.450 805.950 ;
        RECT 266.400 801.900 267.450 814.950 ;
        RECT 277.950 810.450 280.050 814.050 ;
        RECT 281.400 810.450 282.450 833.400 ;
        RECT 287.400 831.450 288.450 833.400 ;
        RECT 287.400 830.400 291.450 831.450 ;
        RECT 286.950 817.950 289.050 820.050 ;
        RECT 277.950 810.000 282.450 810.450 ;
        RECT 278.400 809.400 282.450 810.000 ;
        RECT 271.950 806.100 274.050 808.200 ;
        RECT 278.400 807.600 279.450 809.400 ;
        RECT 272.400 805.350 273.600 806.100 ;
        RECT 278.400 805.350 279.600 807.600 ;
        RECT 271.950 802.950 274.050 805.050 ;
        RECT 274.950 802.950 277.050 805.050 ;
        RECT 277.950 802.950 280.050 805.050 ;
        RECT 280.950 802.950 283.050 805.050 ;
        RECT 275.400 801.900 276.600 802.650 ;
        RECT 281.400 801.900 282.600 802.650 ;
        RECT 287.400 802.050 288.450 817.950 ;
        RECT 290.400 817.050 291.450 830.400 ;
        RECT 296.400 817.050 297.450 839.100 ;
        RECT 299.400 834.900 300.450 853.950 ;
        RECT 308.400 853.050 309.450 875.400 ;
        RECT 310.950 874.950 313.050 877.050 ;
        RECT 317.550 876.300 319.650 878.400 ;
        RECT 307.950 850.950 310.050 853.050 ;
        RECT 311.400 841.200 312.450 874.950 ;
        RECT 317.550 869.700 318.750 876.300 ;
        RECT 349.950 874.950 352.050 877.050 ;
        RECT 346.950 871.950 349.050 874.050 ;
        RECT 317.550 867.600 319.650 869.700 ;
        RECT 325.350 849.300 327.450 851.400 ;
        RECT 326.250 842.700 327.450 849.300 ;
        RECT 340.650 847.500 342.750 848.400 ;
        RECT 340.650 846.300 344.850 847.500 ;
        RECT 347.400 847.050 348.450 871.950 ;
        RECT 350.400 850.050 351.450 874.950 ;
        RECT 362.400 868.050 363.450 883.950 ;
        RECT 368.400 883.350 369.600 884.100 ;
        RECT 382.950 883.950 385.050 886.050 ;
        RECT 391.950 884.100 394.050 886.200 ;
        RECT 421.950 884.100 424.050 886.200 ;
        RECT 427.950 884.100 430.050 886.200 ;
        RECT 367.950 880.950 370.050 883.050 ;
        RECT 370.950 880.950 373.050 883.050 ;
        RECT 373.950 880.950 376.050 883.050 ;
        RECT 376.950 880.950 379.050 883.050 ;
        RECT 377.400 879.000 378.600 880.650 ;
        RECT 376.950 874.950 379.050 879.000 ;
        RECT 361.950 865.950 364.050 868.050 ;
        RECT 383.400 856.050 384.450 883.950 ;
        RECT 392.400 883.350 393.600 884.100 ;
        RECT 422.400 883.350 423.600 884.100 ;
        RECT 428.400 883.350 429.600 884.100 ;
        RECT 391.950 880.950 394.050 883.050 ;
        RECT 394.950 880.950 397.050 883.050 ;
        RECT 397.950 880.950 400.050 883.050 ;
        RECT 400.950 880.950 403.050 883.050 ;
        RECT 416.100 880.950 418.200 883.050 ;
        RECT 421.500 880.950 423.600 883.050 ;
        RECT 427.950 880.950 430.050 883.050 ;
        RECT 401.400 879.000 402.600 880.650 ;
        RECT 400.950 874.950 403.050 879.000 ;
        RECT 434.250 878.400 435.450 891.300 ;
        RECT 445.800 880.950 447.900 883.050 ;
        RECT 433.350 876.300 435.450 878.400 ;
        RECT 446.400 878.400 447.600 880.650 ;
        RECT 446.400 876.450 447.450 878.400 ;
        RECT 434.250 869.700 435.450 876.300 ;
        RECT 412.950 865.950 415.050 868.050 ;
        RECT 433.350 867.600 435.450 869.700 ;
        RECT 443.400 875.400 447.450 876.450 ;
        RECT 382.950 853.950 385.050 856.050 ;
        RECT 349.950 847.950 352.050 850.050 ;
        RECT 361.350 849.300 363.450 851.400 ;
        RECT 364.950 850.950 367.050 853.050 ;
        RECT 304.950 839.100 307.050 841.200 ;
        RECT 310.950 839.100 313.050 841.200 ;
        RECT 325.350 840.600 327.450 842.700 ;
        RECT 305.400 838.350 306.600 839.100 ;
        RECT 311.400 838.350 312.600 839.100 ;
        RECT 304.950 835.950 307.050 838.050 ;
        RECT 307.950 835.950 310.050 838.050 ;
        RECT 310.950 835.950 313.050 838.050 ;
        RECT 313.950 835.950 316.050 838.050 ;
        RECT 319.950 835.950 322.050 838.050 ;
        RECT 298.950 832.800 301.050 834.900 ;
        RECT 308.400 833.400 309.600 835.650 ;
        RECT 314.400 834.900 315.600 835.650 ;
        RECT 320.400 834.900 321.600 835.650 ;
        RECT 289.950 814.950 292.050 817.050 ;
        RECT 295.950 814.950 298.050 817.050 ;
        RECT 299.400 814.050 300.450 832.800 ;
        RECT 308.400 823.050 309.450 833.400 ;
        RECT 313.950 832.800 316.050 834.900 ;
        RECT 319.950 832.800 322.050 834.900 ;
        RECT 326.250 827.700 327.450 840.600 ;
        RECT 328.800 838.950 330.900 841.050 ;
        RECT 331.950 839.100 334.050 841.200 ;
        RECT 337.950 839.100 340.050 841.200 ;
        RECT 310.950 823.950 313.050 826.050 ;
        RECT 325.350 825.600 327.450 827.700 ;
        RECT 329.400 826.050 330.450 838.950 ;
        RECT 332.400 832.050 333.450 839.100 ;
        RECT 338.400 838.350 339.600 839.100 ;
        RECT 337.800 835.950 339.900 838.050 ;
        RECT 331.950 829.950 334.050 832.050 ;
        RECT 343.650 827.700 344.850 846.300 ;
        RECT 346.950 844.950 349.050 847.050 ;
        RECT 347.400 840.600 348.450 844.950 ;
        RECT 362.250 842.700 363.450 849.300 ;
        RECT 361.350 840.600 363.450 842.700 ;
        RECT 347.400 838.350 348.600 840.600 ;
        RECT 346.950 835.950 349.050 838.050 ;
        RECT 355.950 835.950 358.050 838.050 ;
        RECT 356.400 834.900 357.600 835.650 ;
        RECT 355.950 832.800 358.050 834.900 ;
        RECT 346.950 829.950 349.050 832.050 ;
        RECT 328.950 823.950 331.050 826.050 ;
        RECT 343.050 825.600 345.150 827.700 ;
        RECT 307.950 820.950 310.050 823.050 ;
        RECT 298.950 811.950 301.050 814.050 ;
        RECT 304.950 811.950 307.050 814.050 ;
        RECT 289.950 805.950 292.050 808.050 ;
        RECT 298.950 806.100 301.050 808.200 ;
        RECT 305.400 807.600 306.450 811.950 ;
        RECT 265.950 799.800 268.050 801.900 ;
        RECT 274.950 799.800 277.050 801.900 ;
        RECT 280.950 799.800 283.050 801.900 ;
        RECT 286.950 799.950 289.050 802.050 ;
        RECT 290.400 801.900 291.450 805.950 ;
        RECT 299.400 805.350 300.600 806.100 ;
        RECT 305.400 805.350 306.600 807.600 ;
        RECT 295.950 802.950 298.050 805.050 ;
        RECT 298.950 802.950 301.050 805.050 ;
        RECT 301.950 802.950 304.050 805.050 ;
        RECT 304.950 802.950 307.050 805.050 ;
        RECT 296.400 802.050 297.600 802.650 ;
        RECT 289.950 799.800 292.050 801.900 ;
        RECT 292.950 800.400 297.600 802.050 ;
        RECT 302.400 801.900 303.600 802.650 ;
        RECT 311.400 801.900 312.450 823.950 ;
        RECT 319.950 817.950 322.050 820.050 ;
        RECT 313.950 814.950 316.050 817.050 ;
        RECT 314.400 802.050 315.450 814.950 ;
        RECT 320.400 808.200 321.450 817.950 ;
        RECT 347.400 813.450 348.450 829.950 ;
        RECT 362.250 827.700 363.450 840.600 ;
        RECT 365.400 834.900 366.450 850.950 ;
        RECT 383.400 850.050 384.450 853.950 ;
        RECT 376.650 847.500 378.750 848.400 ;
        RECT 382.950 847.950 385.050 850.050 ;
        RECT 406.950 847.950 409.050 850.050 ;
        RECT 376.650 846.300 380.850 847.500 ;
        RECT 373.950 839.100 376.050 841.200 ;
        RECT 374.400 838.350 375.600 839.100 ;
        RECT 373.800 835.950 375.900 838.050 ;
        RECT 364.950 832.800 367.050 834.900 ;
        RECT 379.650 827.700 380.850 846.300 ;
        RECT 382.950 844.800 385.050 846.900 ;
        RECT 383.400 840.600 384.450 844.800 ;
        RECT 407.400 840.600 408.450 847.950 ;
        RECT 413.400 840.600 414.450 865.950 ;
        RECT 443.400 850.050 444.450 875.400 ;
        RECT 451.650 872.700 452.850 891.300 ;
        RECT 502.950 884.100 505.050 886.200 ;
        RECT 508.950 884.100 511.050 886.200 ;
        RECT 503.400 883.350 504.600 884.100 ;
        RECT 509.400 883.350 510.600 884.100 ;
        RECT 454.950 880.950 457.050 883.050 ;
        RECT 473.100 880.950 475.200 883.050 ;
        RECT 478.500 880.950 480.600 883.050 ;
        RECT 497.100 880.950 499.200 883.050 ;
        RECT 502.500 880.950 504.600 883.050 ;
        RECT 508.950 880.950 511.050 883.050 ;
        RECT 448.650 871.500 452.850 872.700 ;
        RECT 455.400 878.400 456.600 880.650 ;
        RECT 473.400 879.000 474.600 880.650 ;
        RECT 448.650 870.600 450.750 871.500 ;
        RECT 455.400 871.050 456.450 878.400 ;
        RECT 472.950 874.950 475.050 879.000 ;
        RECT 515.250 878.400 516.450 891.300 ;
        RECT 526.800 880.950 528.900 883.050 ;
        RECT 514.350 876.300 516.450 878.400 ;
        RECT 527.400 878.400 528.600 880.650 ;
        RECT 527.400 876.450 528.450 878.400 ;
        RECT 454.950 868.950 457.050 871.050 ;
        RECT 473.400 868.050 474.450 874.950 ;
        RECT 481.950 868.950 484.050 871.050 ;
        RECT 515.250 869.700 516.450 876.300 ;
        RECT 472.950 865.950 475.050 868.050 ;
        RECT 442.950 847.950 445.050 850.050 ;
        RECT 475.950 847.950 478.050 850.050 ;
        RECT 433.800 844.500 435.900 846.600 ;
        RECT 383.400 838.350 384.600 840.600 ;
        RECT 407.400 838.350 408.600 840.600 ;
        RECT 413.400 838.350 414.600 840.600 ;
        RECT 427.950 838.950 430.050 841.050 ;
        RECT 382.950 835.950 385.050 838.050 ;
        RECT 403.950 835.950 406.050 838.050 ;
        RECT 406.950 835.950 409.050 838.050 ;
        RECT 409.950 835.950 412.050 838.050 ;
        RECT 412.950 835.950 415.050 838.050 ;
        RECT 404.400 834.900 405.600 835.650 ;
        RECT 391.950 832.800 394.050 834.900 ;
        RECT 403.950 832.800 406.050 834.900 ;
        RECT 410.400 833.400 411.600 835.650 ;
        RECT 361.350 825.600 363.450 827.700 ;
        RECT 379.050 825.600 381.150 827.700 ;
        RECT 347.400 811.200 348.600 813.450 ;
        RECT 319.950 806.100 322.050 808.200 ;
        RECT 342.900 807.900 345.000 809.700 ;
        RECT 346.800 808.800 348.900 810.900 ;
        RECT 350.100 810.300 352.200 812.400 ;
        RECT 370.950 811.950 373.050 814.050 ;
        RECT 341.400 806.700 350.100 807.900 ;
        RECT 320.400 805.350 321.600 806.100 ;
        RECT 319.950 802.950 322.050 805.050 ;
        RECT 322.950 802.950 325.050 805.050 ;
        RECT 338.100 802.950 340.200 805.050 ;
        RECT 292.950 799.950 297.000 800.400 ;
        RECT 301.950 799.800 304.050 801.900 ;
        RECT 310.800 799.800 312.900 801.900 ;
        RECT 313.950 799.950 316.050 802.050 ;
        RECT 323.400 801.900 324.600 802.650 ;
        RECT 322.950 799.800 325.050 801.900 ;
        RECT 338.400 801.450 339.600 802.650 ;
        RECT 335.400 800.400 339.600 801.450 ;
        RECT 262.950 796.950 265.050 799.050 ;
        RECT 281.400 793.050 282.450 799.800 ;
        RECT 247.950 790.950 250.050 793.050 ;
        RECT 280.950 790.950 283.050 793.050 ;
        RECT 256.950 784.950 259.050 787.050 ;
        RECT 322.950 784.950 325.050 787.050 ;
        RECT 241.950 778.950 244.050 781.050 ;
        RECT 250.950 778.950 253.050 781.050 ;
        RECT 242.400 772.050 243.450 778.950 ;
        RECT 241.950 769.950 244.050 772.050 ;
        RECT 241.950 766.800 244.050 768.900 ;
        RECT 238.950 763.950 241.050 766.050 ;
        RECT 233.400 760.350 234.600 762.600 ;
        RECT 239.400 762.450 240.600 762.600 ;
        RECT 242.400 762.450 243.450 766.800 ;
        RECT 244.950 763.950 247.050 766.050 ;
        RECT 239.400 761.400 243.450 762.450 ;
        RECT 239.400 760.350 240.600 761.400 ;
        RECT 229.950 757.950 232.050 760.050 ;
        RECT 232.950 757.950 235.050 760.050 ;
        RECT 235.950 757.950 238.050 760.050 ;
        RECT 238.950 757.950 241.050 760.050 ;
        RECT 208.950 754.800 211.050 756.900 ;
        RECT 214.950 754.800 217.050 756.900 ;
        RECT 223.950 754.950 226.050 757.050 ;
        RECT 230.400 755.400 231.600 757.650 ;
        RECT 236.400 756.900 237.600 757.650 ;
        RECT 199.950 742.950 202.050 745.050 ;
        RECT 190.950 733.950 193.050 736.050 ;
        RECT 200.400 732.450 201.450 742.950 ;
        RECT 197.400 731.400 201.450 732.450 ;
        RECT 170.400 727.350 171.600 729.600 ;
        RECT 175.950 728.100 178.050 730.200 ;
        RECT 197.400 729.600 198.450 731.400 ;
        RECT 176.400 727.350 177.600 728.100 ;
        RECT 197.400 727.350 198.600 729.600 ;
        RECT 205.950 727.950 208.050 730.050 ;
        RECT 169.950 724.950 172.050 727.050 ;
        RECT 172.950 724.950 175.050 727.050 ;
        RECT 175.950 724.950 178.050 727.050 ;
        RECT 178.950 724.950 181.050 727.050 ;
        RECT 193.950 724.950 196.050 727.050 ;
        RECT 196.950 724.950 199.050 727.050 ;
        RECT 199.950 724.950 202.050 727.050 ;
        RECT 160.950 721.950 163.050 724.050 ;
        RECT 173.400 723.900 174.600 724.650 ;
        RECT 179.400 723.900 180.600 724.650 ;
        RECT 166.950 721.800 169.050 723.900 ;
        RECT 172.950 721.800 175.050 723.900 ;
        RECT 178.950 721.800 181.050 723.900 ;
        RECT 190.950 723.450 193.050 723.900 ;
        RECT 194.400 723.450 195.600 724.650 ;
        RECT 200.400 723.900 201.600 724.650 ;
        RECT 206.400 723.900 207.450 727.950 ;
        RECT 190.950 722.400 195.600 723.450 ;
        RECT 190.950 721.800 193.050 722.400 ;
        RECT 199.950 721.800 202.050 723.900 ;
        RECT 205.950 721.800 208.050 723.900 ;
        RECT 157.950 712.950 160.050 715.050 ;
        RECT 148.950 688.950 151.050 691.050 ;
        RECT 151.950 684.000 154.050 688.050 ;
        RECT 152.400 682.350 153.600 684.000 ;
        RECT 157.950 683.100 160.050 685.200 ;
        RECT 158.400 682.350 159.600 683.100 ;
        RECT 148.950 679.950 151.050 682.050 ;
        RECT 151.950 679.950 154.050 682.050 ;
        RECT 154.950 679.950 157.050 682.050 ;
        RECT 157.950 679.950 160.050 682.050 ;
        RECT 149.400 678.900 150.600 679.650 ;
        RECT 142.950 676.800 145.050 678.900 ;
        RECT 148.950 676.800 151.050 678.900 ;
        RECT 155.400 677.400 156.600 679.650 ;
        RECT 124.950 670.950 127.050 673.050 ;
        RECT 139.950 670.950 142.050 673.050 ;
        RECT 155.400 664.050 156.450 677.400 ;
        RECT 160.950 676.950 163.050 679.050 ;
        RECT 161.400 670.050 162.450 676.950 ;
        RECT 167.400 676.050 168.450 721.800 ;
        RECT 178.950 703.950 181.050 706.050 ;
        RECT 179.400 700.050 180.450 703.950 ;
        RECT 181.950 700.950 184.050 703.050 ;
        RECT 169.950 697.950 172.050 700.050 ;
        RECT 178.950 697.950 181.050 700.050 ;
        RECT 170.400 685.050 171.450 697.950 ;
        RECT 169.950 682.950 172.050 685.050 ;
        RECT 175.950 683.100 178.050 685.200 ;
        RECT 182.400 684.600 183.450 700.950 ;
        RECT 176.400 682.350 177.600 683.100 ;
        RECT 182.400 682.350 183.600 684.600 ;
        RECT 172.950 679.950 175.050 682.050 ;
        RECT 175.950 679.950 178.050 682.050 ;
        RECT 178.950 679.950 181.050 682.050 ;
        RECT 181.950 679.950 184.050 682.050 ;
        RECT 173.400 678.900 174.600 679.650 ;
        RECT 172.950 676.800 175.050 678.900 ;
        RECT 179.400 677.400 180.600 679.650 ;
        RECT 166.950 673.950 169.050 676.050 ;
        RECT 179.400 673.050 180.450 677.400 ;
        RECT 184.950 676.950 187.050 679.050 ;
        RECT 181.950 673.950 184.050 676.050 ;
        RECT 178.950 670.950 181.050 673.050 ;
        RECT 160.950 667.950 163.050 670.050 ;
        RECT 154.950 661.950 157.050 664.050 ;
        RECT 103.950 655.950 106.050 658.050 ;
        RECT 109.950 655.950 112.050 658.050 ;
        RECT 130.950 655.950 133.050 658.050 ;
        RECT 151.950 655.950 154.050 658.050 ;
        RECT 166.950 655.950 169.050 658.050 ;
        RECT 97.950 649.950 100.050 652.050 ;
        RECT 104.400 651.600 105.450 655.950 ;
        RECT 110.400 651.600 111.450 655.950 ;
        RECT 104.400 649.350 105.600 651.600 ;
        RECT 110.400 649.350 111.600 651.600 ;
        RECT 118.950 649.950 121.050 652.050 ;
        RECT 124.950 650.100 127.050 652.200 ;
        RECT 131.400 651.600 132.450 655.950 ;
        RECT 152.400 651.600 153.450 655.950 ;
        RECT 100.950 646.950 103.050 649.050 ;
        RECT 103.950 646.950 106.050 649.050 ;
        RECT 106.950 646.950 109.050 649.050 ;
        RECT 109.950 646.950 112.050 649.050 ;
        RECT 101.400 645.900 102.600 646.650 ;
        RECT 100.950 643.800 103.050 645.900 ;
        RECT 107.400 645.000 108.600 646.650 ;
        RECT 106.950 640.950 109.050 645.000 ;
        RECT 119.400 643.050 120.450 649.950 ;
        RECT 125.400 649.350 126.600 650.100 ;
        RECT 131.400 649.350 132.600 651.600 ;
        RECT 152.400 649.350 153.600 651.600 ;
        RECT 157.950 650.100 160.050 652.200 ;
        RECT 167.400 652.050 168.450 655.950 ;
        RECT 158.400 649.350 159.600 650.100 ;
        RECT 166.800 649.950 168.900 652.050 ;
        RECT 169.950 650.100 172.050 652.200 ;
        RECT 175.950 650.100 178.050 652.200 ;
        RECT 182.400 651.600 183.450 673.950 ;
        RECT 185.400 673.050 186.450 676.950 ;
        RECT 184.950 670.950 187.050 673.050 ;
        RECT 191.400 664.050 192.450 721.800 ;
        RECT 209.400 712.050 210.450 754.800 ;
        RECT 230.400 753.450 231.450 755.400 ;
        RECT 235.950 754.800 238.050 756.900 ;
        RECT 230.400 753.000 234.450 753.450 ;
        RECT 229.950 752.400 234.450 753.000 ;
        RECT 229.950 748.950 232.050 752.400 ;
        RECT 223.950 742.950 226.050 745.050 ;
        RECT 224.400 736.050 225.450 742.950 ;
        RECT 223.950 733.950 226.050 736.050 ;
        RECT 217.950 728.100 220.050 730.200 ;
        RECT 224.400 729.600 225.450 733.950 ;
        RECT 218.400 727.350 219.600 728.100 ;
        RECT 224.400 727.350 225.600 729.600 ;
        RECT 214.950 724.950 217.050 727.050 ;
        RECT 217.950 724.950 220.050 727.050 ;
        RECT 220.950 724.950 223.050 727.050 ;
        RECT 223.950 724.950 226.050 727.050 ;
        RECT 226.950 724.950 229.050 727.050 ;
        RECT 215.400 722.400 216.600 724.650 ;
        RECT 221.400 722.400 222.600 724.650 ;
        RECT 227.400 723.000 228.600 724.650 ;
        RECT 208.950 709.950 211.050 712.050 ;
        RECT 215.400 703.050 216.450 722.400 ;
        RECT 217.950 712.950 220.050 715.050 ;
        RECT 214.950 700.950 217.050 703.050 ;
        RECT 196.950 688.950 199.050 691.050 ;
        RECT 193.950 685.950 196.050 688.050 ;
        RECT 194.400 682.050 195.450 685.950 ;
        RECT 197.400 684.600 198.450 688.950 ;
        RECT 197.400 682.350 198.600 684.600 ;
        RECT 205.950 683.100 208.050 685.200 ;
        RECT 206.400 682.350 207.600 683.100 ;
        RECT 193.950 679.950 196.050 682.050 ;
        RECT 197.100 679.950 199.200 682.050 ;
        RECT 200.400 679.950 202.500 682.050 ;
        RECT 205.800 679.950 207.900 682.050 ;
        RECT 193.950 676.800 196.050 678.900 ;
        RECT 200.400 677.400 201.600 679.650 ;
        RECT 218.400 678.900 219.450 712.950 ;
        RECT 221.400 709.050 222.450 722.400 ;
        RECT 226.950 718.950 229.050 723.000 ;
        RECT 229.950 721.950 232.050 724.050 ;
        RECT 220.950 706.950 223.050 709.050 ;
        RECT 223.950 684.000 226.050 688.050 ;
        RECT 230.400 685.200 231.450 721.950 ;
        RECT 233.400 718.050 234.450 752.400 ;
        RECT 235.950 736.950 238.050 739.050 ;
        RECT 236.400 721.050 237.450 736.950 ;
        RECT 245.400 733.050 246.450 763.950 ;
        RECT 251.400 757.050 252.450 778.950 ;
        RECT 253.950 769.950 256.050 772.050 ;
        RECT 250.950 754.950 253.050 757.050 ;
        RECT 244.950 732.450 247.050 733.050 ;
        RECT 242.400 731.400 247.050 732.450 ;
        RECT 254.400 732.450 255.450 769.950 ;
        RECT 257.400 762.600 258.450 784.950 ;
        RECT 257.400 760.350 258.600 762.600 ;
        RECT 265.950 762.000 268.050 766.050 ;
        RECT 266.400 760.350 267.600 762.000 ;
        RECT 274.950 761.100 277.050 763.200 ;
        RECT 280.950 761.100 283.050 763.200 ;
        RECT 286.950 761.100 289.050 766.050 ;
        RECT 295.950 761.100 298.050 763.200 ;
        RECT 307.950 762.000 310.050 766.050 ;
        RECT 323.400 762.600 324.450 784.950 ;
        RECT 335.400 784.050 336.450 800.400 ;
        RECT 341.400 797.700 342.300 806.700 ;
        RECT 348.000 805.800 350.100 806.700 ;
        RECT 351.000 804.900 351.900 810.300 ;
        RECT 371.400 807.600 372.450 811.950 ;
        RECT 392.400 808.200 393.450 832.800 ;
        RECT 406.950 829.950 409.050 832.050 ;
        RECT 407.400 814.050 408.450 829.950 ;
        RECT 406.950 811.950 409.050 814.050 ;
        RECT 353.400 807.450 354.600 807.600 ;
        RECT 353.400 806.400 357.450 807.450 ;
        RECT 353.400 805.350 354.600 806.400 ;
        RECT 345.000 803.700 351.900 804.900 ;
        RECT 345.000 801.300 345.900 803.700 ;
        RECT 343.800 799.200 345.900 801.300 ;
        RECT 346.800 799.950 348.900 802.050 ;
        RECT 340.500 795.600 342.600 797.700 ;
        RECT 347.400 797.400 348.600 799.650 ;
        RECT 350.700 796.500 351.900 803.700 ;
        RECT 352.800 802.950 354.900 805.050 ;
        RECT 356.400 801.900 357.450 806.400 ;
        RECT 371.400 805.350 372.600 807.600 ;
        RECT 391.950 806.100 394.050 808.200 ;
        RECT 407.400 807.450 408.450 811.950 ;
        RECT 410.400 811.050 411.450 833.400 ;
        RECT 428.400 829.050 429.450 838.950 ;
        RECT 431.100 835.950 433.200 838.050 ;
        RECT 434.100 837.300 435.300 844.500 ;
        RECT 437.400 841.350 438.600 843.600 ;
        RECT 443.400 843.300 445.500 845.400 ;
        RECT 437.100 838.950 439.200 841.050 ;
        RECT 440.100 839.700 442.200 841.800 ;
        RECT 440.100 837.300 441.000 839.700 ;
        RECT 434.100 836.100 441.000 837.300 ;
        RECT 431.400 834.900 432.600 835.650 ;
        RECT 430.950 832.800 433.050 834.900 ;
        RECT 434.100 830.700 435.000 836.100 ;
        RECT 435.900 834.300 438.000 835.200 ;
        RECT 443.700 834.300 444.600 843.300 ;
        RECT 472.950 841.950 475.050 844.050 ;
        RECT 446.400 840.450 447.600 840.600 ;
        RECT 446.400 839.400 450.450 840.450 ;
        RECT 446.400 838.350 447.600 839.400 ;
        RECT 445.800 835.950 447.900 838.050 ;
        RECT 435.900 833.100 444.600 834.300 ;
        RECT 427.950 826.950 430.050 829.050 ;
        RECT 433.800 828.600 435.900 830.700 ;
        RECT 437.100 830.100 439.200 832.200 ;
        RECT 441.000 831.300 443.100 833.100 ;
        RECT 437.400 829.050 438.600 829.800 ;
        RECT 436.950 826.950 439.050 829.050 ;
        RECT 449.400 823.050 450.450 839.400 ;
        RECT 463.800 835.950 465.900 838.050 ;
        RECT 436.950 820.950 439.050 823.050 ;
        RECT 448.950 820.950 451.050 823.050 ;
        RECT 409.950 808.950 412.050 811.050 ;
        RECT 410.400 807.450 411.600 807.600 ;
        RECT 407.400 806.400 411.600 807.450 ;
        RECT 392.400 805.350 393.600 806.100 ;
        RECT 410.400 805.350 411.600 806.400 ;
        RECT 415.950 806.100 418.050 808.200 ;
        RECT 427.950 806.100 430.050 808.200 ;
        RECT 437.400 807.600 438.450 820.950 ;
        RECT 416.400 805.350 417.600 806.100 ;
        RECT 367.950 802.950 370.050 805.050 ;
        RECT 370.950 802.950 373.050 805.050 ;
        RECT 373.950 802.950 376.050 805.050 ;
        RECT 388.950 802.950 391.050 805.050 ;
        RECT 391.950 802.950 394.050 805.050 ;
        RECT 394.950 802.950 397.050 805.050 ;
        RECT 409.950 802.950 412.050 805.050 ;
        RECT 412.950 802.950 415.050 805.050 ;
        RECT 415.950 802.950 418.050 805.050 ;
        RECT 418.950 802.950 421.050 805.050 ;
        RECT 368.400 801.900 369.600 802.650 ;
        RECT 355.950 799.800 358.050 801.900 ;
        RECT 367.950 799.800 370.050 801.900 ;
        RECT 374.400 800.400 375.600 802.650 ;
        RECT 389.400 801.000 390.600 802.650 ;
        RECT 350.100 794.400 352.200 796.500 ;
        RECT 356.400 787.050 357.450 799.800 ;
        RECT 374.400 796.050 375.450 800.400 ;
        RECT 388.950 796.950 391.050 801.000 ;
        RECT 413.400 800.400 414.600 802.650 ;
        RECT 419.400 800.400 420.600 802.650 ;
        RECT 394.950 796.950 397.050 799.050 ;
        RECT 373.950 793.950 376.050 796.050 ;
        RECT 367.950 787.950 370.050 790.050 ;
        RECT 355.950 784.950 358.050 787.050 ;
        RECT 334.950 781.950 337.050 784.050 ;
        RECT 331.950 778.950 334.050 781.050 ;
        RECT 332.400 775.050 333.450 778.950 ;
        RECT 331.950 772.950 334.050 775.050 ;
        RECT 328.950 769.950 331.050 772.050 ;
        RECT 329.400 762.600 330.450 769.950 ;
        RECT 358.950 766.950 361.050 769.050 ;
        RECT 336.000 762.600 340.050 763.050 ;
        RECT 257.100 757.950 259.200 760.050 ;
        RECT 260.400 757.950 262.500 760.050 ;
        RECT 265.800 757.950 267.900 760.050 ;
        RECT 260.400 756.000 261.600 757.650 ;
        RECT 259.950 751.950 262.050 756.000 ;
        RECT 275.400 754.050 276.450 761.100 ;
        RECT 281.400 760.350 282.600 761.100 ;
        RECT 287.400 760.350 288.600 761.100 ;
        RECT 280.950 757.950 283.050 760.050 ;
        RECT 283.950 757.950 286.050 760.050 ;
        RECT 286.950 757.950 289.050 760.050 ;
        RECT 289.950 757.950 292.050 760.050 ;
        RECT 284.400 755.400 285.600 757.650 ;
        RECT 290.400 756.900 291.600 757.650 ;
        RECT 284.400 754.050 285.450 755.400 ;
        RECT 289.950 754.800 292.050 756.900 ;
        RECT 274.950 751.950 277.050 754.050 ;
        RECT 280.800 751.950 282.900 754.050 ;
        RECT 283.950 751.950 286.050 754.050 ;
        RECT 277.950 742.950 280.050 745.050 ;
        RECT 271.950 736.950 274.050 739.050 ;
        RECT 254.400 731.400 258.450 732.450 ;
        RECT 242.400 729.600 243.450 731.400 ;
        RECT 244.950 730.950 247.050 731.400 ;
        RECT 242.400 727.350 243.600 729.600 ;
        RECT 247.950 728.100 250.050 730.200 ;
        RECT 248.400 727.350 249.600 728.100 ;
        RECT 241.950 724.950 244.050 727.050 ;
        RECT 244.950 724.950 247.050 727.050 ;
        RECT 247.950 724.950 250.050 727.050 ;
        RECT 250.950 724.950 253.050 727.050 ;
        RECT 245.400 723.900 246.600 724.650 ;
        RECT 244.950 721.800 247.050 723.900 ;
        RECT 251.400 722.400 252.600 724.650 ;
        RECT 257.400 723.900 258.450 731.400 ;
        RECT 265.950 729.000 268.050 733.050 ;
        RECT 272.400 730.200 273.450 736.950 ;
        RECT 278.400 733.050 279.450 742.950 ;
        RECT 281.400 742.050 282.450 751.950 ;
        RECT 284.400 748.050 285.450 751.950 ;
        RECT 283.950 745.950 286.050 748.050 ;
        RECT 280.950 739.950 283.050 742.050 ;
        RECT 280.950 733.950 283.050 736.050 ;
        RECT 289.950 733.950 292.050 736.050 ;
        RECT 277.950 730.950 280.050 733.050 ;
        RECT 266.400 727.350 267.600 729.000 ;
        RECT 271.950 728.100 274.050 730.200 ;
        RECT 272.400 727.350 273.600 728.100 ;
        RECT 265.950 724.950 268.050 727.050 ;
        RECT 268.950 724.950 271.050 727.050 ;
        RECT 271.950 724.950 274.050 727.050 ;
        RECT 274.950 724.950 277.050 727.050 ;
        RECT 269.400 723.900 270.600 724.650 ;
        RECT 235.950 718.950 238.050 721.050 ;
        RECT 251.400 718.050 252.450 722.400 ;
        RECT 256.950 721.800 259.050 723.900 ;
        RECT 268.950 721.800 271.050 723.900 ;
        RECT 275.400 722.400 276.600 724.650 ;
        RECT 232.950 715.950 235.050 718.050 ;
        RECT 250.950 715.950 253.050 718.050 ;
        RECT 247.950 706.950 250.050 709.050 ;
        RECT 248.400 702.450 249.450 706.950 ;
        RECT 251.400 706.050 252.450 715.950 ;
        RECT 275.400 712.050 276.450 722.400 ;
        RECT 274.950 709.950 277.050 712.050 ;
        RECT 262.950 706.950 265.050 709.050 ;
        RECT 250.950 703.950 253.050 706.050 ;
        RECT 253.950 702.450 256.050 703.050 ;
        RECT 248.400 701.400 256.050 702.450 ;
        RECT 253.950 700.950 256.050 701.400 ;
        RECT 263.400 700.050 264.450 706.950 ;
        RECT 262.950 697.950 265.050 700.050 ;
        RECT 268.950 697.950 271.050 700.050 ;
        RECT 224.400 682.350 225.600 684.000 ;
        RECT 229.950 683.100 232.050 685.200 ;
        RECT 247.950 683.100 250.050 685.200 ;
        RECT 253.950 684.000 256.050 688.050 ;
        RECT 230.400 682.350 231.600 683.100 ;
        RECT 248.400 682.350 249.600 683.100 ;
        RECT 254.400 682.350 255.600 684.000 ;
        RECT 223.950 679.950 226.050 682.050 ;
        RECT 226.950 679.950 229.050 682.050 ;
        RECT 229.950 679.950 232.050 682.050 ;
        RECT 232.950 679.950 235.050 682.050 ;
        RECT 247.950 679.950 250.050 682.050 ;
        RECT 250.950 679.950 253.050 682.050 ;
        RECT 253.950 679.950 256.050 682.050 ;
        RECT 256.950 679.950 259.050 682.050 ;
        RECT 227.400 678.900 228.600 679.650 ;
        RECT 194.400 673.050 195.450 676.800 ;
        RECT 193.950 670.950 196.050 673.050 ;
        RECT 200.400 670.050 201.450 677.400 ;
        RECT 217.950 676.800 220.050 678.900 ;
        RECT 226.950 676.800 229.050 678.900 ;
        RECT 233.400 677.400 234.600 679.650 ;
        RECT 251.400 678.900 252.600 679.650 ;
        RECT 257.400 678.900 258.600 679.650 ;
        RECT 269.400 679.050 270.450 697.950 ;
        RECT 275.400 697.050 276.450 709.950 ;
        RECT 281.400 703.050 282.450 733.950 ;
        RECT 290.400 729.600 291.450 733.950 ;
        RECT 296.400 729.600 297.450 761.100 ;
        RECT 308.400 760.350 309.600 762.000 ;
        RECT 323.400 760.350 324.600 762.600 ;
        RECT 329.400 760.350 330.600 762.600 ;
        RECT 335.400 760.950 340.050 762.600 ;
        RECT 346.950 760.950 349.050 763.200 ;
        RECT 352.950 761.100 355.050 763.200 ;
        RECT 359.400 762.600 360.450 766.950 ;
        RECT 335.400 760.350 336.600 760.950 ;
        RECT 304.950 757.950 307.050 760.050 ;
        RECT 307.950 757.950 310.050 760.050 ;
        RECT 322.950 757.950 325.050 760.050 ;
        RECT 325.950 757.950 328.050 760.050 ;
        RECT 328.950 757.950 331.050 760.050 ;
        RECT 331.950 757.950 334.050 760.050 ;
        RECT 334.950 757.950 337.050 760.050 ;
        RECT 305.400 756.900 306.600 757.650 ;
        RECT 304.950 754.800 307.050 756.900 ;
        RECT 326.400 756.000 327.600 757.650 ;
        RECT 332.400 756.900 333.600 757.650 ;
        RECT 325.950 751.950 328.050 756.000 ;
        RECT 331.950 754.800 334.050 756.900 ;
        RECT 347.400 751.050 348.450 760.950 ;
        RECT 353.400 760.350 354.600 761.100 ;
        RECT 359.400 760.350 360.600 762.600 ;
        RECT 352.950 757.950 355.050 760.050 ;
        RECT 355.950 757.950 358.050 760.050 ;
        RECT 358.950 757.950 361.050 760.050 ;
        RECT 361.950 757.950 364.050 760.050 ;
        RECT 356.400 756.900 357.600 757.650 ;
        RECT 362.400 756.900 363.600 757.650 ;
        RECT 368.400 757.050 369.450 787.950 ;
        RECT 376.950 784.950 379.050 787.050 ;
        RECT 377.400 762.600 378.450 784.950 ;
        RECT 377.400 760.350 378.600 762.600 ;
        RECT 382.950 761.100 385.050 763.200 ;
        RECT 383.400 760.350 384.600 761.100 ;
        RECT 376.950 757.950 379.050 760.050 ;
        RECT 379.950 757.950 382.050 760.050 ;
        RECT 382.950 757.950 385.050 760.050 ;
        RECT 385.950 757.950 388.050 760.050 ;
        RECT 355.950 754.800 358.050 756.900 ;
        RECT 361.950 754.800 364.050 756.900 ;
        RECT 367.950 754.950 370.050 757.050 ;
        RECT 380.400 755.400 381.600 757.650 ;
        RECT 386.400 756.000 387.600 757.650 ;
        RECT 346.950 748.950 349.050 751.050 ;
        RECT 356.400 748.050 357.450 754.800 ;
        RECT 355.950 745.950 358.050 748.050 ;
        RECT 380.400 742.050 381.450 755.400 ;
        RECT 385.950 751.950 388.050 756.000 ;
        RECT 391.950 745.950 394.050 748.050 ;
        RECT 340.950 739.950 343.050 742.050 ;
        RECT 379.950 739.950 382.050 742.050 ;
        RECT 310.950 736.950 313.050 739.050 ;
        RECT 290.400 727.350 291.600 729.600 ;
        RECT 296.400 727.350 297.600 729.600 ;
        RECT 307.950 727.950 310.050 730.050 ;
        RECT 289.950 724.950 292.050 727.050 ;
        RECT 292.950 724.950 295.050 727.050 ;
        RECT 295.950 724.950 298.050 727.050 ;
        RECT 298.950 724.950 301.050 727.050 ;
        RECT 293.400 722.400 294.600 724.650 ;
        RECT 299.400 723.000 300.600 724.650 ;
        RECT 308.400 723.900 309.450 727.950 ;
        RECT 283.950 718.950 286.050 721.050 ;
        RECT 280.950 700.950 283.050 703.050 ;
        RECT 274.950 694.950 277.050 697.050 ;
        RECT 277.950 688.950 280.050 691.050 ;
        RECT 278.400 684.600 279.450 688.950 ;
        RECT 278.400 682.350 279.600 684.600 ;
        RECT 284.400 682.050 285.450 718.950 ;
        RECT 293.400 700.050 294.450 722.400 ;
        RECT 298.950 718.950 301.050 723.000 ;
        RECT 307.950 721.800 310.050 723.900 ;
        RECT 292.950 697.950 295.050 700.050 ;
        RECT 301.950 697.950 304.050 700.050 ;
        RECT 289.950 694.950 292.050 697.050 ;
        RECT 286.950 683.100 289.050 685.200 ;
        RECT 272.400 679.950 274.500 682.050 ;
        RECT 277.800 679.950 279.900 682.050 ;
        RECT 283.950 679.950 286.050 682.050 ;
        RECT 199.950 667.950 202.050 670.050 ;
        RECT 233.400 667.050 234.450 677.400 ;
        RECT 250.950 676.800 253.050 678.900 ;
        RECT 256.950 676.800 259.050 678.900 ;
        RECT 268.950 676.950 271.050 679.050 ;
        RECT 284.400 676.050 285.450 679.950 ;
        RECT 283.950 673.950 286.050 676.050 ;
        RECT 268.950 670.950 271.050 673.050 ;
        RECT 232.950 664.950 235.050 667.050 ;
        RECT 190.950 661.950 193.050 664.050 ;
        RECT 229.950 655.950 232.050 658.050 ;
        RECT 230.400 652.200 231.450 655.950 ;
        RECT 124.950 646.950 127.050 649.050 ;
        RECT 127.950 646.950 130.050 649.050 ;
        RECT 130.950 646.950 133.050 649.050 ;
        RECT 133.950 646.950 136.050 649.050 ;
        RECT 148.950 646.950 151.050 649.050 ;
        RECT 151.950 646.950 154.050 649.050 ;
        RECT 154.950 646.950 157.050 649.050 ;
        RECT 157.950 646.950 160.050 649.050 ;
        RECT 121.950 643.950 124.050 646.050 ;
        RECT 128.400 645.000 129.600 646.650 ;
        RECT 134.400 645.900 135.600 646.650 ;
        RECT 118.950 640.950 121.050 643.050 ;
        RECT 122.400 637.050 123.450 643.950 ;
        RECT 127.950 640.950 130.050 645.000 ;
        RECT 133.950 643.800 136.050 645.900 ;
        RECT 149.400 645.000 150.600 646.650 ;
        RECT 155.400 645.900 156.600 646.650 ;
        RECT 167.400 645.900 168.450 649.950 ;
        RECT 148.950 640.950 151.050 645.000 ;
        RECT 154.950 643.800 157.050 645.900 ;
        RECT 166.950 643.800 169.050 645.900 ;
        RECT 155.400 642.450 156.450 643.800 ;
        RECT 152.400 641.400 156.450 642.450 ;
        RECT 121.950 634.950 124.050 637.050 ;
        RECT 130.950 619.950 133.050 622.050 ;
        RECT 37.950 604.950 40.050 607.050 ;
        RECT 43.950 605.100 46.050 607.200 ;
        RECT 38.400 589.050 39.450 604.950 ;
        RECT 44.400 604.350 45.600 605.100 ;
        RECT 43.800 601.950 45.900 604.050 ;
        RECT 49.650 593.700 50.850 612.300 ;
        RECT 52.950 610.950 55.050 613.050 ;
        RECT 58.950 610.950 61.050 613.050 ;
        RECT 94.950 610.950 97.050 613.050 ;
        RECT 127.950 610.950 130.050 613.050 ;
        RECT 53.400 606.600 54.450 610.950 ;
        RECT 53.400 604.350 54.600 606.600 ;
        RECT 52.950 601.950 55.050 604.050 ;
        RECT 49.050 591.600 51.150 593.700 ;
        RECT 37.950 586.950 40.050 589.050 ;
        RECT 37.950 580.950 40.050 583.050 ;
        RECT 34.950 505.950 37.050 508.050 ;
        RECT 31.350 501.300 33.450 503.400 ;
        RECT 19.950 494.100 22.050 496.200 ;
        RECT 25.950 494.100 28.050 496.200 ;
        RECT 20.400 493.350 21.600 494.100 ;
        RECT 26.400 493.350 27.600 494.100 ;
        RECT 14.100 490.950 16.200 493.050 ;
        RECT 19.500 490.950 21.600 493.050 ;
        RECT 25.950 490.950 28.050 493.050 ;
        RECT 32.250 488.400 33.450 501.300 ;
        RECT 38.400 490.050 39.450 580.950 ;
        RECT 49.050 579.300 51.150 581.400 ;
        RECT 43.800 568.950 45.900 571.050 ;
        RECT 44.400 566.400 45.600 568.650 ;
        RECT 44.400 564.450 45.450 566.400 ;
        RECT 41.400 563.400 45.450 564.450 ;
        RECT 41.400 559.050 42.450 563.400 ;
        RECT 49.650 560.700 50.850 579.300 ;
        RECT 52.950 568.950 55.050 571.050 ;
        RECT 53.400 567.900 54.600 568.650 ;
        RECT 59.400 568.050 60.450 610.950 ;
        RECT 64.950 604.950 67.050 607.050 ;
        RECT 73.950 605.100 76.050 607.200 ;
        RECT 97.950 605.100 100.050 607.200 ;
        RECT 103.950 605.100 106.050 607.200 ;
        RECT 118.950 605.100 121.050 607.200 ;
        RECT 65.400 577.050 66.450 604.950 ;
        RECT 74.400 604.350 75.600 605.100 ;
        RECT 98.400 604.350 99.600 605.100 ;
        RECT 70.950 601.950 73.050 604.050 ;
        RECT 73.950 601.950 76.050 604.050 ;
        RECT 76.950 601.950 79.050 604.050 ;
        RECT 91.950 601.950 94.050 604.050 ;
        RECT 94.950 601.950 97.050 604.050 ;
        RECT 97.950 601.950 100.050 604.050 ;
        RECT 77.400 599.400 78.600 601.650 ;
        RECT 95.400 600.000 96.600 601.650 ;
        RECT 77.400 586.050 78.450 599.400 ;
        RECT 94.950 595.950 97.050 600.000 ;
        RECT 104.400 586.050 105.450 605.100 ;
        RECT 119.400 604.350 120.600 605.100 ;
        RECT 109.950 601.950 112.050 604.050 ;
        RECT 115.950 601.950 118.050 604.050 ;
        RECT 118.950 601.950 121.050 604.050 ;
        RECT 76.950 583.950 79.050 586.050 ;
        RECT 103.950 583.950 106.050 586.050 ;
        RECT 82.950 580.950 85.050 583.050 ;
        RECT 64.950 574.950 67.050 577.050 ;
        RECT 70.950 573.000 73.050 577.050 ;
        RECT 76.950 573.000 79.050 577.050 ;
        RECT 83.400 573.600 84.450 580.950 ;
        RECT 88.350 579.300 90.450 581.400 ;
        RECT 106.050 579.300 108.150 581.400 ;
        RECT 71.400 571.350 72.600 573.000 ;
        RECT 77.400 571.350 78.600 573.000 ;
        RECT 83.400 571.350 84.600 573.600 ;
        RECT 70.950 568.950 73.050 571.050 ;
        RECT 73.950 568.950 76.050 571.050 ;
        RECT 76.950 568.950 79.050 571.050 ;
        RECT 82.950 568.950 85.050 571.050 ;
        RECT 52.950 565.800 55.050 567.900 ;
        RECT 58.950 565.950 61.050 568.050 ;
        RECT 74.400 566.400 75.600 568.650 ;
        RECT 89.250 566.400 90.450 579.300 ;
        RECT 100.800 568.950 102.900 571.050 ;
        RECT 101.400 567.900 102.600 568.650 ;
        RECT 46.650 559.500 50.850 560.700 ;
        RECT 40.950 556.950 43.050 559.050 ;
        RECT 46.650 558.600 48.750 559.500 ;
        RECT 46.650 535.500 48.750 536.400 ;
        RECT 46.650 534.300 50.850 535.500 ;
        RECT 43.950 527.100 46.050 529.200 ;
        RECT 44.400 526.350 45.600 527.100 ;
        RECT 43.800 523.950 45.900 526.050 ;
        RECT 49.650 515.700 50.850 534.300 ;
        RECT 53.400 529.200 54.450 565.800 ;
        RECT 74.400 559.050 75.450 566.400 ;
        RECT 88.350 564.300 90.450 566.400 ;
        RECT 100.950 565.800 103.050 567.900 ;
        RECT 73.950 556.950 76.050 559.050 ;
        RECT 89.250 557.700 90.450 564.300 ;
        RECT 106.650 560.700 107.850 579.300 ;
        RECT 110.400 577.050 111.450 601.950 ;
        RECT 116.400 600.000 117.600 601.650 ;
        RECT 115.950 595.950 118.050 600.000 ;
        RECT 128.400 595.050 129.450 610.950 ;
        RECT 131.400 607.050 132.450 619.950 ;
        RECT 136.950 607.950 139.050 613.050 ;
        RECT 148.950 607.950 151.050 610.050 ;
        RECT 130.950 604.950 133.050 607.050 ;
        RECT 137.400 606.600 138.450 607.950 ;
        RECT 137.400 604.350 138.600 606.600 ;
        RECT 142.950 605.100 145.050 607.200 ;
        RECT 143.400 604.350 144.600 605.100 ;
        RECT 133.950 601.950 136.050 604.050 ;
        RECT 136.950 601.950 139.050 604.050 ;
        RECT 139.950 601.950 142.050 604.050 ;
        RECT 142.950 601.950 145.050 604.050 ;
        RECT 134.400 599.400 135.600 601.650 ;
        RECT 140.400 600.900 141.600 601.650 ;
        RECT 118.950 592.950 121.050 595.050 ;
        RECT 127.950 592.950 130.050 595.050 ;
        RECT 109.950 574.950 112.050 577.050 ;
        RECT 109.950 568.950 112.050 571.050 ;
        RECT 103.650 559.500 107.850 560.700 ;
        RECT 110.400 566.400 111.600 568.650 ;
        RECT 103.650 558.600 105.750 559.500 ;
        RECT 88.350 555.600 90.450 557.700 ;
        RECT 110.400 550.050 111.450 566.400 ;
        RECT 88.950 547.950 91.050 550.050 ;
        RECT 109.950 547.950 112.050 550.050 ;
        RECT 67.350 537.300 69.450 539.400 ;
        RECT 68.250 530.700 69.450 537.300 ;
        RECT 82.650 535.500 84.750 536.400 ;
        RECT 82.650 534.300 86.850 535.500 ;
        RECT 52.950 527.100 55.050 529.200 ;
        RECT 67.350 528.600 69.450 530.700 ;
        RECT 53.400 526.350 54.600 527.100 ;
        RECT 52.950 523.950 55.050 526.050 ;
        RECT 61.950 523.950 64.050 526.050 ;
        RECT 62.400 522.900 63.600 523.650 ;
        RECT 61.950 520.800 64.050 522.900 ;
        RECT 68.250 515.700 69.450 528.600 ;
        RECT 79.950 528.000 82.050 532.050 ;
        RECT 80.400 526.350 81.600 528.000 ;
        RECT 79.800 523.950 81.900 526.050 ;
        RECT 85.650 515.700 86.850 534.300 ;
        RECT 89.400 529.200 90.450 547.950 ;
        RECT 112.950 532.950 115.050 535.050 ;
        RECT 88.950 527.100 91.050 529.200 ;
        RECT 113.400 528.600 114.450 532.950 ;
        RECT 119.400 531.450 120.450 592.950 ;
        RECT 134.400 583.050 135.450 599.400 ;
        RECT 139.950 598.800 142.050 600.900 ;
        RECT 140.400 592.050 141.450 598.800 ;
        RECT 149.400 598.050 150.450 607.950 ;
        RECT 148.950 595.950 151.050 598.050 ;
        RECT 139.950 589.950 142.050 592.050 ;
        RECT 127.950 580.950 130.050 583.050 ;
        RECT 133.950 580.950 136.050 583.050 ;
        RECT 121.950 574.950 124.050 577.050 ;
        RECT 122.400 538.050 123.450 574.950 ;
        RECT 128.400 573.600 129.450 580.950 ;
        RECT 128.400 571.350 129.600 573.600 ;
        RECT 133.950 572.100 136.050 574.200 ;
        RECT 139.950 572.100 142.050 574.200 ;
        RECT 149.400 573.600 150.450 595.950 ;
        RECT 152.400 589.050 153.450 641.400 ;
        RECT 170.400 631.050 171.450 650.100 ;
        RECT 176.400 649.350 177.600 650.100 ;
        RECT 182.400 649.350 183.600 651.600 ;
        RECT 190.950 649.950 193.050 652.050 ;
        RECT 196.950 651.600 201.000 652.050 ;
        RECT 196.950 649.950 201.600 651.600 ;
        RECT 211.950 649.950 214.050 652.050 ;
        RECT 223.950 650.100 226.050 652.200 ;
        RECT 229.950 650.100 232.050 652.200 ;
        RECT 247.950 650.100 250.050 652.200 ;
        RECT 175.950 646.950 178.050 649.050 ;
        RECT 178.950 646.950 181.050 649.050 ;
        RECT 181.950 646.950 184.050 649.050 ;
        RECT 184.950 646.950 187.050 649.050 ;
        RECT 179.400 645.900 180.600 646.650 ;
        RECT 178.950 643.800 181.050 645.900 ;
        RECT 185.400 644.400 186.600 646.650 ;
        RECT 185.400 637.050 186.450 644.400 ;
        RECT 191.400 637.050 192.450 649.950 ;
        RECT 200.400 649.350 201.600 649.950 ;
        RECT 199.950 646.950 202.050 649.050 ;
        RECT 202.950 646.950 205.050 649.050 ;
        RECT 203.400 645.000 204.600 646.650 ;
        RECT 202.950 640.950 205.050 645.000 ;
        RECT 175.950 634.950 178.050 637.050 ;
        RECT 184.950 634.950 187.050 637.050 ;
        RECT 190.950 634.950 193.050 637.050 ;
        RECT 205.950 634.950 208.050 637.050 ;
        RECT 169.950 628.950 172.050 631.050 ;
        RECT 154.950 607.950 157.050 613.050 ;
        RECT 166.950 610.800 169.050 612.900 ;
        RECT 160.950 605.100 163.050 610.050 ;
        RECT 167.400 606.600 168.450 610.800 ;
        RECT 172.950 607.950 175.050 610.050 ;
        RECT 161.400 604.350 162.600 605.100 ;
        RECT 167.400 604.350 168.600 606.600 ;
        RECT 157.950 601.950 160.050 604.050 ;
        RECT 160.950 601.950 163.050 604.050 ;
        RECT 163.950 601.950 166.050 604.050 ;
        RECT 166.950 601.950 169.050 604.050 ;
        RECT 158.400 600.000 159.600 601.650 ;
        RECT 157.950 595.950 160.050 600.000 ;
        RECT 164.400 599.400 165.600 601.650 ;
        RECT 173.400 601.050 174.450 607.950 ;
        RECT 164.400 592.050 165.450 599.400 ;
        RECT 172.950 598.950 175.050 601.050 ;
        RECT 176.400 595.050 177.450 634.950 ;
        RECT 199.950 631.950 202.050 634.050 ;
        RECT 184.950 610.950 187.050 613.050 ;
        RECT 185.400 606.600 186.450 610.950 ;
        RECT 185.400 604.350 186.600 606.600 ;
        RECT 190.950 605.100 193.050 607.200 ;
        RECT 191.400 604.350 192.600 605.100 ;
        RECT 181.950 601.950 184.050 604.050 ;
        RECT 184.950 601.950 187.050 604.050 ;
        RECT 187.950 601.950 190.050 604.050 ;
        RECT 190.950 601.950 193.050 604.050 ;
        RECT 182.400 600.900 183.600 601.650 ;
        RECT 181.950 598.800 184.050 600.900 ;
        RECT 188.400 599.400 189.600 601.650 ;
        RECT 188.400 595.050 189.450 599.400 ;
        RECT 175.950 592.950 178.050 595.050 ;
        RECT 187.950 592.950 190.050 595.050 ;
        RECT 163.950 589.950 166.050 592.050 ;
        RECT 151.950 586.950 154.050 589.050 ;
        RECT 169.950 586.950 172.050 589.050 ;
        RECT 157.950 577.950 160.050 580.050 ;
        RECT 163.350 579.300 165.450 581.400 ;
        RECT 158.400 573.600 159.450 577.950 ;
        RECT 134.400 571.350 135.600 572.100 ;
        RECT 127.950 568.950 130.050 571.050 ;
        RECT 130.950 568.950 133.050 571.050 ;
        RECT 133.950 568.950 136.050 571.050 ;
        RECT 131.400 567.900 132.600 568.650 ;
        RECT 140.400 568.050 141.450 572.100 ;
        RECT 149.400 571.350 150.600 573.600 ;
        RECT 158.400 571.350 159.600 573.600 ;
        RECT 148.950 568.950 151.050 571.050 ;
        RECT 151.950 568.950 154.050 571.050 ;
        RECT 157.950 568.950 160.050 571.050 ;
        RECT 130.950 565.800 133.050 567.900 ;
        RECT 139.950 565.950 142.050 568.050 ;
        RECT 152.400 567.900 153.600 568.650 ;
        RECT 151.950 565.800 154.050 567.900 ;
        RECT 164.250 566.400 165.450 579.300 ;
        RECT 163.350 564.300 165.450 566.400 ;
        RECT 164.250 557.700 165.450 564.300 ;
        RECT 163.350 555.600 165.450 557.700 ;
        RECT 121.950 535.950 124.050 538.050 ;
        RECT 133.950 535.950 136.050 538.050 ;
        RECT 160.950 535.950 163.050 538.050 ;
        RECT 121.950 531.450 124.050 532.050 ;
        RECT 119.400 530.400 124.050 531.450 ;
        RECT 121.950 529.950 124.050 530.400 ;
        RECT 89.400 526.350 90.600 527.100 ;
        RECT 113.400 526.350 114.600 528.600 ;
        RECT 88.950 523.950 91.050 526.050 ;
        RECT 109.950 523.950 112.050 526.050 ;
        RECT 112.950 523.950 115.050 526.050 ;
        RECT 115.950 523.950 118.050 526.050 ;
        RECT 110.400 521.400 111.600 523.650 ;
        RECT 116.400 522.900 117.600 523.650 ;
        RECT 122.400 522.900 123.450 529.950 ;
        RECT 134.400 528.600 135.450 535.950 ;
        RECT 134.400 526.350 135.600 528.600 ;
        RECT 139.950 527.100 142.050 529.200 ;
        RECT 145.950 527.100 148.050 529.200 ;
        RECT 154.950 527.100 157.050 529.200 ;
        RECT 161.400 528.600 162.450 535.950 ;
        RECT 140.400 526.350 141.600 527.100 ;
        RECT 130.950 523.950 133.050 526.050 ;
        RECT 133.950 523.950 136.050 526.050 ;
        RECT 136.950 523.950 139.050 526.050 ;
        RECT 139.950 523.950 142.050 526.050 ;
        RECT 110.400 517.050 111.450 521.400 ;
        RECT 115.950 520.800 118.050 522.900 ;
        RECT 121.950 520.800 124.050 522.900 ;
        RECT 131.400 521.400 132.600 523.650 ;
        RECT 137.400 522.900 138.600 523.650 ;
        RECT 131.400 517.050 132.450 521.400 ;
        RECT 136.950 520.800 139.050 522.900 ;
        RECT 49.050 513.600 51.150 515.700 ;
        RECT 67.350 513.600 69.450 515.700 ;
        RECT 85.050 513.600 87.150 515.700 ;
        RECT 109.950 514.950 112.050 517.050 ;
        RECT 130.950 514.950 133.050 517.050 ;
        RECT 88.950 505.950 91.050 508.050 ;
        RECT 49.050 501.300 51.150 503.400 ;
        RECT 43.800 490.950 45.900 493.050 ;
        RECT 31.350 486.300 33.450 488.400 ;
        RECT 37.950 487.950 40.050 490.050 ;
        RECT 44.400 489.900 45.600 490.650 ;
        RECT 43.950 487.800 46.050 489.900 ;
        RECT 32.250 479.700 33.450 486.300 ;
        RECT 49.650 482.700 50.850 501.300 ;
        RECT 73.950 494.100 76.050 496.200 ;
        RECT 74.400 493.350 75.600 494.100 ;
        RECT 52.950 490.950 55.050 493.050 ;
        RECT 73.950 490.950 76.050 493.050 ;
        RECT 76.950 490.950 79.050 493.050 ;
        RECT 79.950 490.950 82.050 493.050 ;
        RECT 82.950 490.950 85.050 493.050 ;
        RECT 46.650 481.500 50.850 482.700 ;
        RECT 53.400 488.400 54.600 490.650 ;
        RECT 83.400 489.900 84.600 490.650 ;
        RECT 89.400 489.900 90.450 505.950 ;
        RECT 146.400 505.050 147.450 527.100 ;
        RECT 155.400 526.350 156.600 527.100 ;
        RECT 161.400 526.350 162.600 528.600 ;
        RECT 154.950 523.950 157.050 526.050 ;
        RECT 157.950 523.950 160.050 526.050 ;
        RECT 160.950 523.950 163.050 526.050 ;
        RECT 163.950 523.950 166.050 526.050 ;
        RECT 158.400 522.900 159.600 523.650 ;
        RECT 164.400 522.900 165.600 523.650 ;
        RECT 157.950 520.800 160.050 522.900 ;
        RECT 163.950 520.800 166.050 522.900 ;
        RECT 170.400 522.450 171.450 586.950 ;
        RECT 190.950 583.950 193.050 586.050 ;
        RECT 181.050 579.300 183.150 581.400 ;
        RECT 175.800 568.950 177.900 571.050 ;
        RECT 176.400 567.450 177.600 568.650 ;
        RECT 173.400 566.400 177.600 567.450 ;
        RECT 173.400 556.050 174.450 566.400 ;
        RECT 181.650 560.700 182.850 579.300 ;
        RECT 184.950 568.950 187.050 571.050 ;
        RECT 178.650 559.500 182.850 560.700 ;
        RECT 185.400 566.400 186.600 568.650 ;
        RECT 178.650 558.600 180.750 559.500 ;
        RECT 172.950 553.950 175.050 556.050 ;
        RECT 185.400 550.050 186.450 566.400 ;
        RECT 191.400 565.050 192.450 583.950 ;
        RECT 200.400 573.450 201.450 631.950 ;
        RECT 206.400 631.050 207.450 634.950 ;
        RECT 205.950 628.950 208.050 631.050 ;
        RECT 206.400 606.600 207.450 628.950 ;
        RECT 208.950 625.950 211.050 628.050 ;
        RECT 209.400 613.050 210.450 625.950 ;
        RECT 212.400 622.050 213.450 649.950 ;
        RECT 224.400 649.350 225.600 650.100 ;
        RECT 230.400 649.350 231.600 650.100 ;
        RECT 248.400 649.350 249.600 650.100 ;
        RECT 256.950 649.950 259.050 652.050 ;
        RECT 269.400 651.600 270.450 670.950 ;
        RECT 280.950 667.950 283.050 670.050 ;
        RECT 220.950 646.950 223.050 649.050 ;
        RECT 223.950 646.950 226.050 649.050 ;
        RECT 226.950 646.950 229.050 649.050 ;
        RECT 229.950 646.950 232.050 649.050 ;
        RECT 247.950 646.950 250.050 649.050 ;
        RECT 250.950 646.950 253.050 649.050 ;
        RECT 221.400 644.400 222.600 646.650 ;
        RECT 227.400 645.000 228.600 646.650 ;
        RECT 221.400 637.050 222.450 644.400 ;
        RECT 226.950 640.950 229.050 645.000 ;
        RECT 251.400 644.400 252.600 646.650 ;
        RECT 220.950 634.950 223.050 637.050 ;
        RECT 251.400 628.050 252.450 644.400 ;
        RECT 250.950 625.950 253.050 628.050 ;
        RECT 211.950 619.950 214.050 622.050 ;
        RECT 208.950 610.950 211.050 613.050 ;
        RECT 206.400 604.350 207.600 606.600 ;
        RECT 214.950 604.950 217.050 607.050 ;
        RECT 226.950 605.100 229.050 607.200 ;
        RECT 238.950 605.100 241.050 607.200 ;
        RECT 247.950 605.100 250.050 607.200 ;
        RECT 254.400 606.450 255.600 606.600 ;
        RECT 257.400 606.450 258.450 649.950 ;
        RECT 269.400 649.350 270.600 651.600 ;
        RECT 274.950 650.100 277.050 652.200 ;
        RECT 275.400 649.350 276.600 650.100 ;
        RECT 265.950 646.950 268.050 649.050 ;
        RECT 268.950 646.950 271.050 649.050 ;
        RECT 271.950 646.950 274.050 649.050 ;
        RECT 274.950 646.950 277.050 649.050 ;
        RECT 266.400 645.900 267.600 646.650 ;
        RECT 265.950 643.800 268.050 645.900 ;
        RECT 272.400 644.400 273.600 646.650 ;
        RECT 281.400 646.050 282.450 667.950 ;
        RECT 272.400 637.050 273.450 644.400 ;
        RECT 280.950 643.950 283.050 646.050 ;
        RECT 280.950 640.800 283.050 642.900 ;
        RECT 271.950 634.950 274.050 637.050 ;
        RECT 262.950 628.950 265.050 631.050 ;
        RECT 254.400 605.400 258.450 606.450 ;
        RECT 205.950 601.950 208.050 604.050 ;
        RECT 208.950 601.950 211.050 604.050 ;
        RECT 209.400 600.900 210.600 601.650 ;
        RECT 215.400 600.900 216.450 604.950 ;
        RECT 227.400 604.350 228.600 605.100 ;
        RECT 223.950 601.950 226.050 604.050 ;
        RECT 226.950 601.950 229.050 604.050 ;
        RECT 229.950 601.950 232.050 604.050 ;
        RECT 208.950 598.800 211.050 600.900 ;
        RECT 214.950 598.800 217.050 600.900 ;
        RECT 224.400 600.000 225.600 601.650 ;
        RECT 230.400 600.900 231.600 601.650 ;
        RECT 203.400 573.450 204.600 573.600 ;
        RECT 200.400 572.400 204.600 573.450 ;
        RECT 209.400 573.450 210.450 598.800 ;
        RECT 223.950 595.950 226.050 600.000 ;
        RECT 229.950 598.800 232.050 600.900 ;
        RECT 214.950 574.950 217.050 577.050 ;
        RECT 209.400 573.000 213.450 573.450 ;
        RECT 209.400 572.400 214.050 573.000 ;
        RECT 203.400 571.350 204.600 572.400 ;
        RECT 202.950 568.950 205.050 571.050 ;
        RECT 205.950 568.950 208.050 571.050 ;
        RECT 211.950 568.950 214.050 572.400 ;
        RECT 206.400 567.900 207.600 568.650 ;
        RECT 215.400 568.050 216.450 574.950 ;
        RECT 220.950 573.000 223.050 577.050 ;
        RECT 221.400 571.350 222.600 573.000 ;
        RECT 226.950 572.100 229.050 574.200 ;
        RECT 230.400 574.050 231.450 598.800 ;
        RECT 239.400 598.050 240.450 605.100 ;
        RECT 248.400 604.350 249.600 605.100 ;
        RECT 254.400 604.350 255.600 605.400 ;
        RECT 263.400 604.050 264.450 628.950 ;
        RECT 277.950 616.950 280.050 619.050 ;
        RECT 271.950 606.000 274.050 610.050 ;
        RECT 278.400 606.600 279.450 616.950 ;
        RECT 281.400 607.050 282.450 640.800 ;
        RECT 272.400 604.350 273.600 606.000 ;
        RECT 278.400 604.350 279.600 606.600 ;
        RECT 280.950 604.950 283.050 607.050 ;
        RECT 244.950 601.950 247.050 604.050 ;
        RECT 247.950 601.950 250.050 604.050 ;
        RECT 250.950 601.950 253.050 604.050 ;
        RECT 253.950 601.950 256.050 604.050 ;
        RECT 262.950 601.950 265.050 604.050 ;
        RECT 268.950 601.950 271.050 604.050 ;
        RECT 271.950 601.950 274.050 604.050 ;
        RECT 274.950 601.950 277.050 604.050 ;
        RECT 277.950 601.950 280.050 604.050 ;
        RECT 245.400 599.400 246.600 601.650 ;
        RECT 251.400 599.400 252.600 601.650 ;
        RECT 269.400 600.900 270.600 601.650 ;
        RECT 238.950 595.950 241.050 598.050 ;
        RECT 245.400 589.050 246.450 599.400 ;
        RECT 251.400 592.050 252.450 599.400 ;
        RECT 268.950 598.800 271.050 600.900 ;
        RECT 275.400 599.400 276.600 601.650 ;
        RECT 275.400 595.050 276.450 599.400 ;
        RECT 280.950 595.950 283.050 598.050 ;
        RECT 274.950 592.950 277.050 595.050 ;
        RECT 250.950 589.950 253.050 592.050 ;
        RECT 244.950 586.950 247.050 589.050 ;
        RECT 253.950 586.950 256.050 589.050 ;
        RECT 244.950 580.950 247.050 583.050 ;
        RECT 227.400 571.350 228.600 572.100 ;
        RECT 229.950 571.950 232.050 574.050 ;
        RECT 232.950 572.100 235.050 574.200 ;
        RECT 245.400 573.600 246.450 580.950 ;
        RECT 254.400 574.200 255.450 586.950 ;
        RECT 220.950 568.950 223.050 571.050 ;
        RECT 223.950 568.950 226.050 571.050 ;
        RECT 226.950 568.950 229.050 571.050 ;
        RECT 205.950 565.800 208.050 567.900 ;
        RECT 214.950 565.950 217.050 568.050 ;
        RECT 224.400 567.000 225.600 568.650 ;
        RECT 190.950 562.950 193.050 565.050 ;
        RECT 223.950 562.950 226.050 567.000 ;
        RECT 184.950 547.950 187.050 550.050 ;
        RECT 199.950 547.950 202.050 550.050 ;
        RECT 178.950 528.000 181.050 532.050 ;
        RECT 200.400 528.600 201.450 547.950 ;
        RECT 233.400 544.050 234.450 572.100 ;
        RECT 245.400 571.350 246.600 573.600 ;
        RECT 253.950 572.100 256.050 574.200 ;
        RECT 265.950 572.100 268.050 574.200 ;
        RECT 271.950 572.100 274.050 574.200 ;
        RECT 241.950 568.950 244.050 571.050 ;
        RECT 244.950 568.950 247.050 571.050 ;
        RECT 247.950 568.950 250.050 571.050 ;
        RECT 242.400 567.900 243.600 568.650 ;
        RECT 241.950 565.800 244.050 567.900 ;
        RECT 248.400 566.400 249.600 568.650 ;
        RECT 254.400 567.450 255.450 572.100 ;
        RECT 266.400 571.350 267.600 572.100 ;
        RECT 272.400 571.350 273.600 572.100 ;
        RECT 265.950 568.950 268.050 571.050 ;
        RECT 268.950 568.950 271.050 571.050 ;
        RECT 271.950 568.950 274.050 571.050 ;
        RECT 274.950 568.950 277.050 571.050 ;
        RECT 269.400 567.900 270.600 568.650 ;
        RECT 275.400 567.900 276.600 568.650 ;
        RECT 251.400 566.400 255.450 567.450 ;
        RECT 248.400 562.050 249.450 566.400 ;
        RECT 247.950 559.950 250.050 562.050 ;
        RECT 241.950 553.950 244.050 556.050 ;
        RECT 232.950 541.950 235.050 544.050 ;
        RECT 226.950 538.950 229.050 541.050 ;
        RECT 179.400 526.350 180.600 528.000 ;
        RECT 200.400 526.350 201.600 528.600 ;
        RECT 178.950 523.950 181.050 526.050 ;
        RECT 181.950 523.950 184.050 526.050 ;
        RECT 200.100 523.950 202.200 526.050 ;
        RECT 218.100 523.950 220.200 526.050 ;
        RECT 182.400 522.900 183.600 523.650 ;
        RECT 167.400 521.400 171.450 522.450 ;
        RECT 139.950 502.950 142.050 505.050 ;
        RECT 145.950 502.950 148.050 505.050 ;
        RECT 91.950 493.950 94.050 496.050 ;
        RECT 106.950 494.100 109.050 496.200 ;
        RECT 46.650 480.600 48.750 481.500 ;
        RECT 31.350 477.600 33.450 479.700 ;
        RECT 53.400 462.450 54.450 488.400 ;
        RECT 82.950 487.800 85.050 489.900 ;
        RECT 88.950 487.800 91.050 489.900 ;
        RECT 92.400 469.050 93.450 493.950 ;
        RECT 107.400 493.350 108.600 494.100 ;
        RECT 115.950 493.950 118.050 496.050 ;
        RECT 121.950 494.100 124.050 496.200 ;
        RECT 140.400 495.600 141.450 502.950 ;
        RECT 97.950 490.950 100.050 493.050 ;
        RECT 100.950 490.950 103.050 493.050 ;
        RECT 103.950 490.950 106.050 493.050 ;
        RECT 106.950 490.950 109.050 493.050 ;
        RECT 98.400 489.900 99.600 490.650 ;
        RECT 97.950 487.800 100.050 489.900 ;
        RECT 91.950 466.950 94.050 469.050 ;
        RECT 106.950 466.950 109.050 469.050 ;
        RECT 55.950 462.450 58.050 463.050 ;
        RECT 53.400 461.400 58.050 462.450 ;
        RECT 34.350 459.300 36.450 461.400 ;
        RECT 55.950 460.950 58.050 461.400 ;
        RECT 35.250 452.700 36.450 459.300 ;
        RECT 49.650 457.500 51.750 458.400 ;
        RECT 49.650 456.300 53.850 457.500 ;
        RECT 34.350 450.600 36.450 452.700 ;
        RECT 17.100 445.950 19.200 448.050 ;
        RECT 22.500 445.950 24.600 448.050 ;
        RECT 28.950 445.950 31.050 448.050 ;
        RECT 23.400 444.900 24.600 445.650 ;
        RECT 29.400 444.900 30.600 445.650 ;
        RECT 22.950 442.800 25.050 444.900 ;
        RECT 28.950 442.800 31.050 444.900 ;
        RECT 35.250 437.700 36.450 450.600 ;
        RECT 46.800 445.950 48.900 448.050 ;
        RECT 52.650 437.700 53.850 456.300 ;
        RECT 56.400 450.600 57.450 460.950 ;
        RECT 70.350 459.300 72.450 461.400 ;
        RECT 76.950 460.950 79.050 463.050 ;
        RECT 91.950 460.950 94.050 463.050 ;
        RECT 71.250 452.700 72.450 459.300 ;
        RECT 70.350 450.600 72.450 452.700 ;
        RECT 56.400 448.350 57.600 450.600 ;
        RECT 55.950 445.950 58.050 448.050 ;
        RECT 64.950 445.950 67.050 448.050 ;
        RECT 65.400 443.400 66.600 445.650 ;
        RECT 34.350 435.600 36.450 437.700 ;
        RECT 52.050 435.600 54.150 437.700 ;
        RECT 65.400 427.050 66.450 443.400 ;
        RECT 71.250 437.700 72.450 450.600 ;
        RECT 70.350 435.600 72.450 437.700 ;
        RECT 40.950 424.950 43.050 427.050 ;
        RECT 64.950 424.950 67.050 427.050 ;
        RECT 19.950 416.100 22.050 418.200 ;
        RECT 41.400 417.600 42.450 424.950 ;
        RECT 73.350 423.300 75.450 425.400 ;
        RECT 20.400 415.350 21.600 416.100 ;
        RECT 41.400 415.350 42.600 417.600 ;
        RECT 61.950 417.000 64.050 421.050 ;
        RECT 62.400 415.350 63.600 417.000 ;
        RECT 67.950 416.100 70.050 418.200 ;
        RECT 68.400 415.350 69.600 416.100 ;
        RECT 14.100 412.950 16.200 415.050 ;
        RECT 19.500 412.950 21.600 415.050 ;
        RECT 35.100 412.950 37.200 415.050 ;
        RECT 40.500 412.950 42.600 415.050 ;
        RECT 56.100 412.950 58.200 415.050 ;
        RECT 61.500 412.950 63.600 415.050 ;
        RECT 67.950 412.950 70.050 415.050 ;
        RECT 74.250 410.400 75.450 423.300 ;
        RECT 73.350 408.300 75.450 410.400 ;
        RECT 74.250 401.700 75.450 408.300 ;
        RECT 73.350 399.600 75.450 401.700 ;
        RECT 31.350 381.300 33.450 383.400 ;
        RECT 67.350 381.300 69.450 383.400 ;
        RECT 32.250 374.700 33.450 381.300 ;
        RECT 46.650 379.500 48.750 380.400 ;
        RECT 46.650 378.300 50.850 379.500 ;
        RECT 31.350 372.600 33.450 374.700 ;
        RECT 14.100 367.950 16.200 370.050 ;
        RECT 19.500 367.950 21.600 370.050 ;
        RECT 25.950 367.950 28.050 370.050 ;
        RECT 20.400 366.900 21.600 367.650 ;
        RECT 26.400 366.900 27.600 367.650 ;
        RECT 19.950 364.800 22.050 366.900 ;
        RECT 25.950 364.800 28.050 366.900 ;
        RECT 32.250 359.700 33.450 372.600 ;
        RECT 43.950 371.100 46.050 373.200 ;
        RECT 44.400 370.350 45.600 371.100 ;
        RECT 43.800 367.950 45.900 370.050 ;
        RECT 49.650 359.700 50.850 378.300 ;
        RECT 52.950 376.950 55.050 379.050 ;
        RECT 53.400 372.600 54.450 376.950 ;
        RECT 68.250 374.700 69.450 381.300 ;
        RECT 77.400 379.050 78.450 460.950 ;
        RECT 85.650 457.500 87.750 458.400 ;
        RECT 85.650 456.300 89.850 457.500 ;
        RECT 82.800 445.950 84.900 448.050 ;
        RECT 88.650 437.700 89.850 456.300 ;
        RECT 92.400 450.600 93.450 460.950 ;
        RECT 92.400 448.350 93.600 450.600 ;
        RECT 91.950 445.950 94.050 448.050 ;
        RECT 107.400 444.900 108.450 466.950 ;
        RECT 116.400 457.050 117.450 493.950 ;
        RECT 122.400 493.350 123.600 494.100 ;
        RECT 140.400 493.350 141.600 495.600 ;
        RECT 145.950 494.100 148.050 496.200 ;
        RECT 146.400 493.350 147.600 494.100 ;
        RECT 121.950 490.950 124.050 493.050 ;
        RECT 124.950 490.950 127.050 493.050 ;
        RECT 139.950 490.950 142.050 493.050 ;
        RECT 142.950 490.950 145.050 493.050 ;
        RECT 145.950 490.950 148.050 493.050 ;
        RECT 148.950 490.950 151.050 493.050 ;
        RECT 154.950 490.950 157.050 493.050 ;
        RECT 125.400 489.900 126.600 490.650 ;
        RECT 143.400 489.900 144.600 490.650 ;
        RECT 124.950 487.800 127.050 489.900 ;
        RECT 142.950 487.800 145.050 489.900 ;
        RECT 149.400 488.400 150.600 490.650 ;
        RECT 145.950 484.950 148.050 487.050 ;
        RECT 115.950 454.950 118.050 457.050 ;
        RECT 124.950 454.950 127.050 457.050 ;
        RECT 115.950 449.100 118.050 451.200 ;
        RECT 116.400 448.350 117.600 449.100 ;
        RECT 112.950 445.950 115.050 448.050 ;
        RECT 115.950 445.950 118.050 448.050 ;
        RECT 113.400 444.900 114.600 445.650 ;
        RECT 125.400 444.900 126.450 454.950 ;
        RECT 133.950 449.100 136.050 451.200 ;
        RECT 139.950 449.100 142.050 451.200 ;
        RECT 134.400 448.350 135.600 449.100 ;
        RECT 140.400 448.350 141.600 449.100 ;
        RECT 130.950 445.950 133.050 448.050 ;
        RECT 133.950 445.950 136.050 448.050 ;
        RECT 136.950 445.950 139.050 448.050 ;
        RECT 139.950 445.950 142.050 448.050 ;
        RECT 131.400 444.900 132.600 445.650 ;
        RECT 106.950 442.800 109.050 444.900 ;
        RECT 112.950 442.800 115.050 444.900 ;
        RECT 124.950 442.800 127.050 444.900 ;
        RECT 130.950 442.800 133.050 444.900 ;
        RECT 137.400 443.400 138.600 445.650 ;
        RECT 137.400 439.050 138.450 443.400 ;
        RECT 142.950 442.950 145.050 445.050 ;
        RECT 88.050 435.600 90.150 437.700 ;
        RECT 136.950 436.950 139.050 439.050 ;
        RECT 91.050 423.300 93.150 425.400 ;
        RECT 109.350 423.300 111.450 425.400 ;
        RECT 127.050 423.300 129.150 425.400 ;
        RECT 85.800 412.950 87.900 415.050 ;
        RECT 91.650 404.700 92.850 423.300 ;
        RECT 103.950 417.000 106.050 421.050 ;
        RECT 104.400 415.350 105.600 417.000 ;
        RECT 94.950 412.950 97.050 415.050 ;
        RECT 103.950 412.950 106.050 415.050 ;
        RECT 88.650 403.500 92.850 404.700 ;
        RECT 95.400 410.400 96.600 412.650 ;
        RECT 110.250 410.400 111.450 423.300 ;
        RECT 121.800 412.950 123.900 415.050 ;
        RECT 88.650 402.600 90.750 403.500 ;
        RECT 95.400 403.050 96.450 410.400 ;
        RECT 109.350 408.300 111.450 410.400 ;
        RECT 94.950 400.950 97.050 403.050 ;
        RECT 110.250 401.700 111.450 408.300 ;
        RECT 127.650 404.700 128.850 423.300 ;
        RECT 130.950 412.950 133.050 415.050 ;
        RECT 124.650 403.500 128.850 404.700 ;
        RECT 131.400 410.400 132.600 412.650 ;
        RECT 143.400 412.050 144.450 442.950 ;
        RECT 146.400 439.050 147.450 484.950 ;
        RECT 149.400 445.050 150.450 488.400 ;
        RECT 155.400 469.050 156.450 490.950 ;
        RECT 158.400 487.050 159.450 520.800 ;
        RECT 157.950 484.950 160.050 487.050 ;
        RECT 154.950 466.950 157.050 469.050 ;
        RECT 155.400 450.600 156.450 466.950 ;
        RECT 167.400 459.450 168.450 521.400 ;
        RECT 181.950 520.800 184.050 522.900 ;
        RECT 220.950 517.950 223.050 520.050 ;
        RECT 202.950 502.950 205.050 505.050 ;
        RECT 170.100 490.950 172.200 493.050 ;
        RECT 188.100 490.950 190.200 493.050 ;
        RECT 170.400 488.400 171.600 490.650 ;
        RECT 170.400 463.050 171.450 488.400 ;
        RECT 169.950 460.950 172.050 463.050 ;
        RECT 167.400 458.400 171.450 459.450 ;
        RECT 160.950 454.950 163.050 457.050 ;
        RECT 161.400 450.600 162.450 454.950 ;
        RECT 155.400 448.350 156.600 450.600 ;
        RECT 161.400 448.350 162.600 450.600 ;
        RECT 154.950 445.950 157.050 448.050 ;
        RECT 157.950 445.950 160.050 448.050 ;
        RECT 160.950 445.950 163.050 448.050 ;
        RECT 163.950 445.950 166.050 448.050 ;
        RECT 148.950 442.950 151.050 445.050 ;
        RECT 158.400 443.400 159.600 445.650 ;
        RECT 164.400 444.000 165.600 445.650 ;
        RECT 148.950 439.800 151.050 441.900 ;
        RECT 145.950 436.950 148.050 439.050 ;
        RECT 149.400 417.600 150.450 439.800 ;
        RECT 158.400 439.050 159.450 443.400 ;
        RECT 163.950 439.950 166.050 444.000 ;
        RECT 170.400 439.050 171.450 458.400 ;
        RECT 203.400 457.050 204.450 502.950 ;
        RECT 209.100 490.950 211.200 493.050 ;
        RECT 214.500 490.950 216.600 493.050 ;
        RECT 217.800 490.950 219.900 493.050 ;
        RECT 218.400 489.450 219.600 490.650 ;
        RECT 221.400 489.450 222.450 517.950 ;
        RECT 218.400 488.400 222.450 489.450 ;
        RECT 227.400 459.450 228.450 538.950 ;
        RECT 242.400 528.600 243.450 553.950 ;
        RECT 242.400 526.350 243.600 528.600 ;
        RECT 236.400 523.950 238.500 526.050 ;
        RECT 241.800 523.950 243.900 526.050 ;
        RECT 235.950 494.100 238.050 496.200 ;
        RECT 251.400 496.050 252.450 566.400 ;
        RECT 268.950 565.800 271.050 567.900 ;
        RECT 274.950 565.800 277.050 567.900 ;
        RECT 275.400 562.050 276.450 565.800 ;
        RECT 281.400 565.050 282.450 595.950 ;
        RECT 284.400 583.050 285.450 673.950 ;
        RECT 287.400 664.050 288.450 683.100 ;
        RECT 290.400 678.450 291.450 694.950 ;
        RECT 295.950 683.100 298.050 685.200 ;
        RECT 302.400 684.600 303.450 697.950 ;
        RECT 311.400 685.050 312.450 736.950 ;
        RECT 319.950 729.000 322.050 733.050 ;
        RECT 320.400 727.350 321.600 729.000 ;
        RECT 325.950 728.100 328.050 730.200 ;
        RECT 326.400 727.350 327.600 728.100 ;
        RECT 334.950 727.950 337.050 730.050 ;
        RECT 341.400 729.600 342.450 739.950 ;
        RECT 346.950 736.950 349.050 739.050 ;
        RECT 347.400 729.600 348.450 736.950 ;
        RECT 379.950 736.800 382.050 738.900 ;
        RECT 316.950 724.950 319.050 727.050 ;
        RECT 319.950 724.950 322.050 727.050 ;
        RECT 322.950 724.950 325.050 727.050 ;
        RECT 325.950 724.950 328.050 727.050 ;
        RECT 317.400 723.900 318.600 724.650 ;
        RECT 316.950 721.800 319.050 723.900 ;
        RECT 323.400 722.400 324.600 724.650 ;
        RECT 335.400 723.900 336.450 727.950 ;
        RECT 341.400 727.350 342.600 729.600 ;
        RECT 347.400 727.350 348.600 729.600 ;
        RECT 355.950 728.100 358.050 730.200 ;
        RECT 367.950 728.100 370.050 730.200 ;
        RECT 373.950 728.100 376.050 730.200 ;
        RECT 340.950 724.950 343.050 727.050 ;
        RECT 343.950 724.950 346.050 727.050 ;
        RECT 346.950 724.950 349.050 727.050 ;
        RECT 349.950 724.950 352.050 727.050 ;
        RECT 344.400 723.900 345.600 724.650 ;
        RECT 323.400 709.050 324.450 722.400 ;
        RECT 334.950 721.800 337.050 723.900 ;
        RECT 325.950 718.950 328.050 721.050 ;
        RECT 343.950 718.950 346.050 723.900 ;
        RECT 350.400 723.000 351.600 724.650 ;
        RECT 349.950 718.950 352.050 723.000 ;
        RECT 356.400 721.050 357.450 728.100 ;
        RECT 368.400 727.350 369.600 728.100 ;
        RECT 374.400 727.350 375.600 728.100 ;
        RECT 364.950 724.950 367.050 727.050 ;
        RECT 367.950 724.950 370.050 727.050 ;
        RECT 370.950 724.950 373.050 727.050 ;
        RECT 373.950 724.950 376.050 727.050 ;
        RECT 365.400 723.000 366.600 724.650 ;
        RECT 355.950 718.950 358.050 721.050 ;
        RECT 364.950 718.950 367.050 723.000 ;
        RECT 371.400 722.400 372.600 724.650 ;
        RECT 322.950 706.950 325.050 709.050 ;
        RECT 316.950 688.950 319.050 691.050 ;
        RECT 296.400 682.350 297.600 683.100 ;
        RECT 302.400 682.350 303.600 684.600 ;
        RECT 310.950 682.950 313.050 685.050 ;
        RECT 295.950 679.950 298.050 682.050 ;
        RECT 298.950 679.950 301.050 682.050 ;
        RECT 301.950 679.950 304.050 682.050 ;
        RECT 304.950 679.950 307.050 682.050 ;
        RECT 290.400 677.400 294.450 678.450 ;
        RECT 286.950 661.950 289.050 664.050 ;
        RECT 293.400 651.600 294.450 677.400 ;
        RECT 299.400 677.400 300.600 679.650 ;
        RECT 305.400 678.000 306.600 679.650 ;
        RECT 299.400 667.050 300.450 677.400 ;
        RECT 304.950 673.950 307.050 678.000 ;
        RECT 298.950 664.950 301.050 667.050 ;
        RECT 317.400 658.050 318.450 688.950 ;
        RECT 326.400 684.600 327.450 718.950 ;
        RECT 371.400 718.050 372.450 722.400 ;
        RECT 331.950 715.950 334.050 718.050 ;
        RECT 370.950 715.950 373.050 718.050 ;
        RECT 332.400 703.050 333.450 715.950 ;
        RECT 355.950 706.950 358.050 709.050 ;
        RECT 334.950 703.950 337.050 706.050 ;
        RECT 331.950 700.950 334.050 703.050 ;
        RECT 326.400 682.350 327.600 684.600 ;
        RECT 322.950 679.950 325.050 682.050 ;
        RECT 325.950 679.950 328.050 682.050 ;
        RECT 323.400 678.000 324.600 679.650 ;
        RECT 322.950 673.950 325.050 678.000 ;
        RECT 316.950 655.950 319.050 658.050 ;
        RECT 293.400 649.350 294.600 651.600 ;
        RECT 313.950 651.000 316.050 655.050 ;
        RECT 322.950 652.950 325.050 655.050 ;
        RECT 314.400 649.350 315.600 651.000 ;
        RECT 289.950 646.950 292.050 649.050 ;
        RECT 292.950 646.950 295.050 649.050 ;
        RECT 295.950 646.950 298.050 649.050 ;
        RECT 310.950 646.950 313.050 649.050 ;
        RECT 313.950 646.950 316.050 649.050 ;
        RECT 316.950 646.950 319.050 649.050 ;
        RECT 290.400 645.450 291.600 646.650 ;
        RECT 287.400 644.400 291.600 645.450 ;
        RECT 296.400 645.000 297.600 646.650 ;
        RECT 287.400 601.050 288.450 644.400 ;
        RECT 295.950 640.950 298.050 645.000 ;
        RECT 323.400 631.050 324.450 652.950 ;
        RECT 335.400 651.600 336.450 703.950 ;
        RECT 352.950 694.950 355.050 697.050 ;
        RECT 340.950 679.950 343.050 682.050 ;
        RECT 343.950 679.950 346.050 682.050 ;
        RECT 346.950 679.950 349.050 682.050 ;
        RECT 344.400 677.400 345.600 679.650 ;
        RECT 344.400 652.200 345.450 677.400 ;
        RECT 335.400 649.350 336.600 651.600 ;
        RECT 343.950 650.100 346.050 652.200 ;
        RECT 353.400 651.450 354.450 694.950 ;
        RECT 356.400 667.050 357.450 706.950 ;
        RECT 358.950 688.950 361.050 691.050 ;
        RECT 359.400 679.050 360.450 688.950 ;
        RECT 367.950 683.100 370.050 685.200 ;
        RECT 368.400 682.350 369.600 683.100 ;
        RECT 376.950 682.950 379.050 685.050 ;
        RECT 364.950 679.950 367.050 682.050 ;
        RECT 367.950 679.950 370.050 682.050 ;
        RECT 358.950 676.950 361.050 679.050 ;
        RECT 365.400 678.900 366.600 679.650 ;
        RECT 377.400 678.900 378.450 682.950 ;
        RECT 364.950 676.800 367.050 678.900 ;
        RECT 370.950 676.800 373.050 678.900 ;
        RECT 376.950 676.800 379.050 678.900 ;
        RECT 361.950 667.950 364.050 670.050 ;
        RECT 355.950 664.950 358.050 667.050 ;
        RECT 350.400 650.400 354.450 651.450 ;
        RECT 355.950 651.000 358.050 655.050 ;
        RECT 362.400 651.600 363.450 667.950 ;
        RECT 331.950 646.950 334.050 649.050 ;
        RECT 334.950 646.950 337.050 649.050 ;
        RECT 337.950 646.950 340.050 649.050 ;
        RECT 332.400 644.400 333.600 646.650 ;
        RECT 338.400 644.400 339.600 646.650 ;
        RECT 344.400 645.900 345.450 650.100 ;
        RECT 332.400 640.050 333.450 644.400 ;
        RECT 331.950 637.950 334.050 640.050 ;
        RECT 322.950 628.950 325.050 631.050 ;
        RECT 289.950 610.950 292.050 613.050 ;
        RECT 319.950 610.950 322.050 613.050 ;
        RECT 332.400 612.450 333.450 637.950 ;
        RECT 332.400 611.400 336.450 612.450 ;
        RECT 286.950 598.950 289.050 601.050 ;
        RECT 286.950 595.800 289.050 597.900 ;
        RECT 283.950 580.950 286.050 583.050 ;
        RECT 287.400 574.050 288.450 595.800 ;
        RECT 290.400 592.050 291.450 610.950 ;
        RECT 298.950 605.100 301.050 607.200 ;
        RECT 304.950 606.000 307.050 610.050 ;
        RECT 320.400 606.600 321.450 610.950 ;
        RECT 299.400 604.350 300.600 605.100 ;
        RECT 305.400 604.350 306.600 606.000 ;
        RECT 320.400 604.350 321.600 606.600 ;
        RECT 325.950 605.100 328.050 607.200 ;
        RECT 326.400 604.350 327.600 605.100 ;
        RECT 331.950 604.950 334.050 610.050 ;
        RECT 295.950 601.950 298.050 604.050 ;
        RECT 298.950 601.950 301.050 604.050 ;
        RECT 301.950 601.950 304.050 604.050 ;
        RECT 304.950 601.950 307.050 604.050 ;
        RECT 319.950 601.950 322.050 604.050 ;
        RECT 322.950 601.950 325.050 604.050 ;
        RECT 325.950 601.950 328.050 604.050 ;
        RECT 328.950 601.950 331.050 604.050 ;
        RECT 296.400 600.900 297.600 601.650 ;
        RECT 295.950 598.800 298.050 600.900 ;
        RECT 302.400 599.400 303.600 601.650 ;
        RECT 292.950 592.950 295.050 595.050 ;
        RECT 289.950 589.950 292.050 592.050 ;
        RECT 293.400 577.050 294.450 592.950 ;
        RECT 302.400 592.050 303.450 599.400 ;
        RECT 316.950 598.950 319.050 601.050 ;
        RECT 323.400 600.900 324.600 601.650 ;
        RECT 301.950 589.950 304.050 592.050 ;
        RECT 292.950 574.950 295.050 577.050 ;
        RECT 286.950 571.950 289.050 574.050 ;
        RECT 304.950 571.950 307.050 574.050 ;
        RECT 317.400 573.600 318.450 598.950 ;
        RECT 322.950 598.800 325.050 600.900 ;
        RECT 329.400 600.000 330.600 601.650 ;
        RECT 319.950 595.950 322.050 598.050 ;
        RECT 328.950 595.950 331.050 600.000 ;
        RECT 335.400 598.050 336.450 611.400 ;
        RECT 334.950 595.950 337.050 598.050 ;
        RECT 320.400 586.050 321.450 595.950 ;
        RECT 338.400 595.050 339.450 644.400 ;
        RECT 343.950 643.800 346.050 645.900 ;
        RECT 350.400 634.050 351.450 650.400 ;
        RECT 356.400 649.350 357.600 651.000 ;
        RECT 362.400 649.350 363.600 651.600 ;
        RECT 355.950 646.950 358.050 649.050 ;
        RECT 358.950 646.950 361.050 649.050 ;
        RECT 361.950 646.950 364.050 649.050 ;
        RECT 364.950 646.950 367.050 649.050 ;
        RECT 359.400 644.400 360.600 646.650 ;
        RECT 365.400 645.900 366.600 646.650 ;
        RECT 349.950 631.950 352.050 634.050 ;
        RECT 343.950 616.950 346.050 619.050 ;
        RECT 344.400 607.200 345.450 616.950 ;
        RECT 343.950 605.100 346.050 607.200 ;
        RECT 359.400 606.450 360.450 644.400 ;
        RECT 364.950 643.800 367.050 645.900 ;
        RECT 371.400 627.450 372.450 676.800 ;
        RECT 380.400 658.050 381.450 736.800 ;
        RECT 382.950 727.950 385.050 730.050 ;
        RECT 392.400 729.600 393.450 745.950 ;
        RECT 395.400 739.050 396.450 796.950 ;
        RECT 406.950 784.950 409.050 787.050 ;
        RECT 400.950 761.100 403.050 763.200 ;
        RECT 407.400 762.600 408.450 784.950 ;
        RECT 409.950 772.950 412.050 775.050 ;
        RECT 410.400 769.050 411.450 772.950 ;
        RECT 413.400 772.050 414.450 800.400 ;
        RECT 419.400 790.050 420.450 800.400 ;
        RECT 428.400 796.050 429.450 806.100 ;
        RECT 437.400 805.350 438.600 807.600 ;
        RECT 445.950 806.100 448.050 808.200 ;
        RECT 454.950 806.100 457.050 808.200 ;
        RECT 433.950 802.950 436.050 805.050 ;
        RECT 436.950 802.950 439.050 805.050 ;
        RECT 439.950 802.950 442.050 805.050 ;
        RECT 434.400 800.400 435.600 802.650 ;
        RECT 440.400 801.000 441.600 802.650 ;
        RECT 427.950 793.950 430.050 796.050 ;
        RECT 427.950 790.800 430.050 792.900 ;
        RECT 418.950 787.950 421.050 790.050 ;
        RECT 428.400 778.050 429.450 790.800 ;
        RECT 434.400 790.050 435.450 800.400 ;
        RECT 439.950 796.950 442.050 801.000 ;
        RECT 433.950 787.950 436.050 790.050 ;
        RECT 427.950 775.950 430.050 778.050 ;
        RECT 412.950 769.950 415.050 772.050 ;
        RECT 409.950 766.950 412.050 769.050 ;
        RECT 401.400 760.350 402.600 761.100 ;
        RECT 407.400 760.350 408.600 762.600 ;
        RECT 418.950 761.100 421.050 763.200 ;
        RECT 428.400 762.600 429.450 775.950 ;
        RECT 446.400 772.050 447.450 806.100 ;
        RECT 455.400 805.350 456.600 806.100 ;
        RECT 463.950 805.950 466.050 808.050 ;
        RECT 454.950 802.950 457.050 805.050 ;
        RECT 457.950 802.950 460.050 805.050 ;
        RECT 458.400 800.400 459.600 802.650 ;
        RECT 458.400 799.050 459.450 800.400 ;
        RECT 454.950 797.400 459.450 799.050 ;
        RECT 454.950 796.950 459.000 797.400 ;
        RECT 464.400 787.050 465.450 805.950 ;
        RECT 463.950 784.950 466.050 787.050 ;
        RECT 448.950 778.950 451.050 781.050 ;
        RECT 466.950 778.950 469.050 781.050 ;
        RECT 445.950 769.950 448.050 772.050 ;
        RECT 449.400 763.200 450.450 778.950 ;
        RECT 454.950 766.950 457.050 769.050 ;
        RECT 400.950 757.950 403.050 760.050 ;
        RECT 403.950 757.950 406.050 760.050 ;
        RECT 406.950 757.950 409.050 760.050 ;
        RECT 409.950 757.950 412.050 760.050 ;
        RECT 404.400 756.900 405.600 757.650 ;
        RECT 403.950 754.800 406.050 756.900 ;
        RECT 410.400 755.400 411.600 757.650 ;
        RECT 397.950 751.950 400.050 754.050 ;
        RECT 394.950 736.950 397.050 739.050 ;
        RECT 398.400 729.600 399.450 751.950 ;
        RECT 404.400 742.050 405.450 754.800 ;
        RECT 403.950 739.950 406.050 742.050 ;
        RECT 406.950 736.950 409.050 739.050 ;
        RECT 383.400 723.900 384.450 727.950 ;
        RECT 392.400 727.350 393.600 729.600 ;
        RECT 398.400 727.350 399.600 729.600 ;
        RECT 388.950 724.950 391.050 727.050 ;
        RECT 391.950 724.950 394.050 727.050 ;
        RECT 394.950 724.950 397.050 727.050 ;
        RECT 397.950 724.950 400.050 727.050 ;
        RECT 389.400 723.900 390.600 724.650 ;
        RECT 382.950 721.800 385.050 723.900 ;
        RECT 388.950 721.800 391.050 723.900 ;
        RECT 395.400 722.400 396.600 724.650 ;
        RECT 407.400 724.050 408.450 736.950 ;
        RECT 410.400 730.200 411.450 755.400 ;
        RECT 415.950 748.950 418.050 751.050 ;
        RECT 416.400 745.050 417.450 748.950 ;
        RECT 419.400 748.050 420.450 761.100 ;
        RECT 428.400 760.350 429.600 762.600 ;
        RECT 433.950 761.100 436.050 763.200 ;
        RECT 448.950 761.100 451.050 763.200 ;
        RECT 455.400 762.600 456.450 766.950 ;
        RECT 463.950 763.950 466.050 766.050 ;
        RECT 434.400 760.350 435.600 761.100 ;
        RECT 449.400 760.350 450.600 761.100 ;
        RECT 455.400 760.350 456.600 762.600 ;
        RECT 424.950 757.950 427.050 760.050 ;
        RECT 427.950 757.950 430.050 760.050 ;
        RECT 430.950 757.950 433.050 760.050 ;
        RECT 433.950 757.950 436.050 760.050 ;
        RECT 448.950 757.950 451.050 760.050 ;
        RECT 451.950 757.950 454.050 760.050 ;
        RECT 454.950 757.950 457.050 760.050 ;
        RECT 457.950 757.950 460.050 760.050 ;
        RECT 425.400 756.900 426.600 757.650 ;
        RECT 431.400 756.900 432.600 757.650 ;
        RECT 452.400 756.900 453.600 757.650 ;
        RECT 424.950 754.800 427.050 756.900 ;
        RECT 430.950 754.800 433.050 756.900 ;
        RECT 451.950 754.800 454.050 756.900 ;
        RECT 458.400 755.400 459.600 757.650 ;
        RECT 418.950 745.950 421.050 748.050 ;
        RECT 415.950 742.950 418.050 745.050 ;
        RECT 409.950 728.100 412.050 730.200 ;
        RECT 416.400 729.600 417.450 742.950 ;
        RECT 419.400 739.050 420.450 745.950 ;
        RECT 418.950 736.950 421.050 739.050 ;
        RECT 454.950 736.950 457.050 739.050 ;
        RECT 445.950 733.050 448.050 733.200 ;
        RECT 430.950 730.950 433.050 733.050 ;
        RECT 442.950 731.100 448.050 733.050 ;
        RECT 442.950 730.950 447.000 731.100 ;
        RECT 416.400 727.350 417.600 729.600 ;
        RECT 421.950 728.100 424.050 730.200 ;
        RECT 422.400 727.350 423.600 728.100 ;
        RECT 415.950 724.950 418.050 727.050 ;
        RECT 418.950 724.950 421.050 727.050 ;
        RECT 421.950 724.950 424.050 727.050 ;
        RECT 424.950 724.950 427.050 727.050 ;
        RECT 395.400 718.050 396.450 722.400 ;
        RECT 406.950 721.950 409.050 724.050 ;
        RECT 412.950 721.950 415.050 724.050 ;
        RECT 419.400 722.400 420.600 724.650 ;
        RECT 425.400 723.900 426.600 724.650 ;
        RECT 431.400 723.900 432.450 730.950 ;
        RECT 433.950 727.950 436.050 730.050 ;
        RECT 439.950 728.100 442.050 730.200 ;
        RECT 394.950 715.950 397.050 718.050 ;
        RECT 385.800 688.500 387.900 690.600 ;
        RECT 383.100 679.950 385.200 682.050 ;
        RECT 386.100 681.300 387.300 688.500 ;
        RECT 389.400 685.350 390.600 687.600 ;
        RECT 395.400 687.300 397.500 689.400 ;
        RECT 409.950 688.950 412.050 691.050 ;
        RECT 389.100 682.950 391.200 685.050 ;
        RECT 392.100 683.700 394.200 685.800 ;
        RECT 392.100 681.300 393.000 683.700 ;
        RECT 386.100 680.100 393.000 681.300 ;
        RECT 383.400 678.900 384.600 679.650 ;
        RECT 382.950 676.800 385.050 678.900 ;
        RECT 386.100 674.700 387.000 680.100 ;
        RECT 387.900 678.300 390.000 679.200 ;
        RECT 395.700 678.300 396.600 687.300 ;
        RECT 398.400 684.450 399.600 684.600 ;
        RECT 400.950 684.450 403.050 685.200 ;
        RECT 398.400 683.400 403.050 684.450 ;
        RECT 398.400 682.350 399.600 683.400 ;
        RECT 400.950 683.100 403.050 683.400 ;
        RECT 397.800 679.950 399.900 682.050 ;
        RECT 387.900 677.100 396.600 678.300 ;
        RECT 385.800 672.600 387.900 674.700 ;
        RECT 389.100 674.100 391.200 676.200 ;
        RECT 393.000 675.300 395.100 677.100 ;
        RECT 389.400 671.550 390.600 673.800 ;
        RECT 389.400 667.050 390.450 671.550 ;
        RECT 401.400 670.050 402.450 683.100 ;
        RECT 410.400 678.900 411.450 688.950 ;
        RECT 409.950 676.800 412.050 678.900 ;
        RECT 400.950 667.950 403.050 670.050 ;
        RECT 388.950 664.950 391.050 667.050 ;
        RECT 379.950 655.950 382.050 658.050 ;
        RECT 401.400 655.050 402.450 667.950 ;
        RECT 413.400 667.050 414.450 721.950 ;
        RECT 419.400 709.050 420.450 722.400 ;
        RECT 424.950 721.800 427.050 723.900 ;
        RECT 430.950 721.800 433.050 723.900 ;
        RECT 434.400 718.050 435.450 727.950 ;
        RECT 440.400 727.350 441.600 728.100 ;
        RECT 445.950 727.950 448.050 730.050 ;
        RECT 446.400 727.350 447.600 727.950 ;
        RECT 439.950 724.950 442.050 727.050 ;
        RECT 442.950 724.950 445.050 727.050 ;
        RECT 445.950 724.950 448.050 727.050 ;
        RECT 448.950 724.950 451.050 727.050 ;
        RECT 443.400 722.400 444.600 724.650 ;
        RECT 449.400 723.900 450.600 724.650 ;
        RECT 433.950 715.950 436.050 718.050 ;
        RECT 418.950 706.950 421.050 709.050 ;
        RECT 443.400 706.050 444.450 722.400 ;
        RECT 448.950 721.800 451.050 723.900 ;
        RECT 433.950 703.950 436.050 706.050 ;
        RECT 442.950 703.950 445.050 706.050 ;
        RECT 418.500 687.300 420.600 689.400 ;
        RECT 428.100 688.500 430.200 690.600 ;
        RECT 415.950 683.100 418.050 685.200 ;
        RECT 416.400 682.350 417.600 683.100 ;
        RECT 416.100 679.950 418.200 682.050 ;
        RECT 419.400 678.300 420.300 687.300 ;
        RECT 421.800 683.700 423.900 685.800 ;
        RECT 425.400 685.350 426.600 687.600 ;
        RECT 423.000 681.300 423.900 683.700 ;
        RECT 424.800 682.950 426.900 685.050 ;
        RECT 428.700 681.300 429.900 688.500 ;
        RECT 423.000 680.100 429.900 681.300 ;
        RECT 426.000 678.300 428.100 679.200 ;
        RECT 419.400 677.100 428.100 678.300 ;
        RECT 420.900 675.300 423.000 677.100 ;
        RECT 424.800 674.100 426.900 676.200 ;
        RECT 429.000 674.700 429.900 680.100 ;
        RECT 430.800 679.950 432.900 682.050 ;
        RECT 431.400 678.900 432.600 679.650 ;
        RECT 430.950 676.800 433.050 678.900 ;
        RECT 425.400 673.050 426.600 673.800 ;
        RECT 424.950 670.950 427.050 673.050 ;
        RECT 428.100 672.600 430.200 674.700 ;
        RECT 434.400 673.050 435.450 703.950 ;
        RECT 455.400 697.050 456.450 736.950 ;
        RECT 458.400 733.050 459.450 755.400 ;
        RECT 464.400 739.050 465.450 763.950 ;
        RECT 467.400 756.900 468.450 778.950 ;
        RECT 473.400 775.050 474.450 841.950 ;
        RECT 476.400 834.900 477.450 847.950 ;
        RECT 482.400 844.050 483.450 868.950 ;
        RECT 514.350 867.600 516.450 869.700 ;
        RECT 524.400 875.400 528.450 876.450 ;
        RECT 496.350 849.300 498.450 851.400 ;
        RECT 481.950 840.000 484.050 844.050 ;
        RECT 497.250 842.700 498.450 849.300 ;
        RECT 511.650 847.500 513.750 848.400 ;
        RECT 511.650 846.300 515.850 847.500 ;
        RECT 496.350 840.600 498.450 842.700 ;
        RECT 482.400 838.350 483.600 840.000 ;
        RECT 481.800 835.950 483.900 838.050 ;
        RECT 490.950 835.950 493.050 838.050 ;
        RECT 491.400 834.900 492.600 835.650 ;
        RECT 475.950 832.800 478.050 834.900 ;
        RECT 490.950 832.800 493.050 834.900 ;
        RECT 497.250 827.700 498.450 840.600 ;
        RECT 508.950 839.100 511.050 841.200 ;
        RECT 509.400 838.350 510.600 839.100 ;
        RECT 508.800 835.950 510.900 838.050 ;
        RECT 514.650 827.700 515.850 846.300 ;
        RECT 517.950 840.000 520.050 844.050 ;
        RECT 518.400 838.350 519.600 840.000 ;
        RECT 517.950 835.950 520.050 838.050 ;
        RECT 524.400 829.050 525.450 875.400 ;
        RECT 532.650 872.700 533.850 891.300 ;
        RECT 535.950 880.950 538.050 883.050 ;
        RECT 544.950 880.950 547.050 883.050 ;
        RECT 536.400 879.900 537.600 880.650 ;
        RECT 545.400 879.900 546.600 880.650 ;
        RECT 535.950 877.800 538.050 879.900 ;
        RECT 544.950 877.800 547.050 879.900 ;
        RECT 529.650 871.500 533.850 872.700 ;
        RECT 529.650 870.600 531.750 871.500 ;
        RECT 536.400 844.050 537.450 877.800 ;
        RECT 549.150 872.700 550.350 891.300 ;
        RECT 554.100 880.950 556.200 883.050 ;
        RECT 554.400 879.000 555.600 880.650 ;
        RECT 553.950 874.950 556.050 879.000 ;
        RECT 566.550 878.400 567.750 891.300 ;
        RECT 709.950 889.950 712.050 892.050 ;
        RECT 760.950 889.950 763.050 892.050 ;
        RECT 571.950 884.100 574.050 886.200 ;
        RECT 592.950 884.100 595.050 886.200 ;
        RECT 655.950 884.100 658.050 886.200 ;
        RECT 664.950 884.100 667.050 886.200 ;
        RECT 670.950 884.100 673.050 886.200 ;
        RECT 572.400 883.350 573.600 884.100 ;
        RECT 593.400 883.350 594.600 884.100 ;
        RECT 571.950 880.950 574.050 883.050 ;
        RECT 593.400 880.950 595.500 883.050 ;
        RECT 598.800 880.950 600.900 883.050 ;
        RECT 614.100 880.950 616.200 883.050 ;
        RECT 619.500 880.950 621.600 883.050 ;
        RECT 638.400 880.950 640.500 883.050 ;
        RECT 643.800 880.950 645.900 883.050 ;
        RECT 614.400 879.000 615.600 880.650 ;
        RECT 566.550 876.300 568.650 878.400 ;
        RECT 549.150 871.500 553.350 872.700 ;
        RECT 551.250 870.600 553.350 871.500 ;
        RECT 566.550 869.700 567.750 876.300 ;
        RECT 613.950 874.950 616.050 879.000 ;
        RECT 644.400 878.400 645.600 880.650 ;
        RECT 566.550 867.600 568.650 869.700 ;
        RECT 644.400 862.050 645.450 878.400 ;
        RECT 656.400 877.050 657.450 884.100 ;
        RECT 665.400 883.350 666.600 884.100 ;
        RECT 671.400 883.350 672.600 884.100 ;
        RECT 682.950 883.950 685.050 886.050 ;
        RECT 710.400 885.600 711.450 889.950 ;
        RECT 661.950 880.950 664.050 883.050 ;
        RECT 664.950 880.950 667.050 883.050 ;
        RECT 667.950 880.950 670.050 883.050 ;
        RECT 670.950 880.950 673.050 883.050 ;
        RECT 662.400 878.400 663.600 880.650 ;
        RECT 668.400 878.400 669.600 880.650 ;
        RECT 655.950 876.450 658.050 877.050 ;
        RECT 653.400 875.400 658.050 876.450 ;
        RECT 643.950 859.950 646.050 862.050 ;
        RECT 625.950 850.950 628.050 853.050 ;
        RECT 616.950 844.950 619.050 847.050 ;
        RECT 535.950 841.950 538.050 844.050 ;
        RECT 538.950 839.100 541.050 841.200 ;
        RECT 547.950 839.100 550.050 841.200 ;
        RECT 562.950 839.100 565.050 841.200 ;
        RECT 568.950 840.000 571.050 844.050 ;
        RECT 539.400 838.350 540.600 839.100 ;
        RECT 535.950 835.950 538.050 838.050 ;
        RECT 538.950 835.950 541.050 838.050 ;
        RECT 541.950 835.950 544.050 838.050 ;
        RECT 536.400 833.400 537.600 835.650 ;
        RECT 542.400 833.400 543.600 835.650 ;
        RECT 490.950 823.950 493.050 826.050 ;
        RECT 496.350 825.600 498.450 827.700 ;
        RECT 514.050 825.600 516.150 827.700 ;
        RECT 523.950 826.950 526.050 829.050 ;
        RECT 536.400 826.050 537.450 833.400 ;
        RECT 535.950 823.950 538.050 826.050 ;
        RECT 476.100 802.950 478.200 805.050 ;
        RECT 481.500 802.950 483.600 805.050 ;
        RECT 476.400 800.400 477.600 802.650 ;
        RECT 472.950 772.950 475.050 775.050 ;
        RECT 476.400 766.050 477.450 800.400 ;
        RECT 487.950 772.950 490.050 775.050 ;
        RECT 478.950 766.950 481.050 769.050 ;
        RECT 475.950 763.950 478.050 766.050 ;
        RECT 472.950 761.100 475.050 763.200 ;
        RECT 479.400 762.600 480.450 766.950 ;
        RECT 473.400 760.350 474.600 761.100 ;
        RECT 479.400 760.350 480.600 762.600 ;
        RECT 472.950 757.950 475.050 760.050 ;
        RECT 475.950 757.950 478.050 760.050 ;
        RECT 478.950 757.950 481.050 760.050 ;
        RECT 481.950 757.950 484.050 760.050 ;
        RECT 476.400 756.900 477.600 757.650 ;
        RECT 466.950 754.800 469.050 756.900 ;
        RECT 475.950 754.800 478.050 756.900 ;
        RECT 482.400 755.400 483.600 757.650 ;
        RECT 478.950 748.950 481.050 751.050 ;
        RECT 463.950 736.950 466.050 739.050 ;
        RECT 469.950 736.950 472.050 739.050 ;
        RECT 457.950 730.950 460.050 733.050 ;
        RECT 460.950 732.450 465.000 733.050 ;
        RECT 460.950 730.950 465.450 732.450 ;
        RECT 464.400 729.600 465.450 730.950 ;
        RECT 470.400 730.200 471.450 736.950 ;
        RECT 464.400 727.350 465.600 729.600 ;
        RECT 469.950 728.100 472.050 730.200 ;
        RECT 470.400 727.350 471.600 728.100 ;
        RECT 463.950 724.950 466.050 727.050 ;
        RECT 466.950 724.950 469.050 727.050 ;
        RECT 469.950 724.950 472.050 727.050 ;
        RECT 472.950 724.950 475.050 727.050 ;
        RECT 467.400 723.900 468.600 724.650 ;
        RECT 466.950 721.800 469.050 723.900 ;
        RECT 473.400 722.400 474.600 724.650 ;
        RECT 460.950 715.950 463.050 718.050 ;
        RECT 454.950 694.950 457.050 697.050 ;
        RECT 451.950 688.950 454.050 691.050 ;
        RECT 436.950 683.100 439.050 685.200 ;
        RECT 445.950 683.100 448.050 685.200 ;
        RECT 452.400 684.600 453.450 688.950 ;
        RECT 433.950 670.950 436.050 673.050 ;
        RECT 437.400 670.050 438.450 683.100 ;
        RECT 446.400 682.350 447.600 683.100 ;
        RECT 452.400 682.350 453.600 684.600 ;
        RECT 445.950 679.950 448.050 682.050 ;
        RECT 448.950 679.950 451.050 682.050 ;
        RECT 451.950 679.950 454.050 682.050 ;
        RECT 449.400 678.900 450.600 679.650 ;
        RECT 461.400 678.900 462.450 715.950 ;
        RECT 473.400 706.050 474.450 722.400 ;
        RECT 472.950 703.950 475.050 706.050 ;
        RECT 479.400 697.050 480.450 748.950 ;
        RECT 482.400 744.450 483.450 755.400 ;
        RECT 488.400 754.050 489.450 772.950 ;
        RECT 491.400 757.050 492.450 823.950 ;
        RECT 514.950 820.950 517.050 823.050 ;
        RECT 499.950 806.100 502.050 808.200 ;
        RECT 505.950 806.100 508.050 808.200 ;
        RECT 511.950 806.100 514.050 808.200 ;
        RECT 500.400 805.350 501.600 806.100 ;
        RECT 506.400 805.350 507.600 806.100 ;
        RECT 496.950 802.950 499.050 805.050 ;
        RECT 499.950 802.950 502.050 805.050 ;
        RECT 502.950 802.950 505.050 805.050 ;
        RECT 505.950 802.950 508.050 805.050 ;
        RECT 497.400 800.400 498.600 802.650 ;
        RECT 503.400 801.000 504.600 802.650 ;
        RECT 497.400 769.050 498.450 800.400 ;
        RECT 502.950 796.950 505.050 801.000 ;
        RECT 512.400 799.050 513.450 806.100 ;
        RECT 515.400 801.900 516.450 820.950 ;
        RECT 523.950 817.950 526.050 820.050 ;
        RECT 524.400 811.050 525.450 817.950 ;
        RECT 542.400 814.050 543.450 833.400 ;
        RECT 548.400 817.050 549.450 839.100 ;
        RECT 563.400 838.350 564.600 839.100 ;
        RECT 569.400 838.350 570.600 840.000 ;
        RECT 574.950 839.100 577.050 841.200 ;
        RECT 586.950 840.000 589.050 844.050 ;
        RECT 598.950 841.950 601.050 844.050 ;
        RECT 559.950 835.950 562.050 838.050 ;
        RECT 562.950 835.950 565.050 838.050 ;
        RECT 565.950 835.950 568.050 838.050 ;
        RECT 568.950 835.950 571.050 838.050 ;
        RECT 560.400 833.400 561.600 835.650 ;
        RECT 566.400 833.400 567.600 835.650 ;
        RECT 556.950 826.950 559.050 829.050 ;
        RECT 547.950 814.950 550.050 817.050 ;
        RECT 541.950 811.950 544.050 814.050 ;
        RECT 523.950 808.950 526.050 811.050 ;
        RECT 538.950 808.950 541.050 811.050 ;
        RECT 520.950 806.100 523.050 808.200 ;
        RECT 526.950 806.100 529.050 808.200 ;
        RECT 535.950 806.100 538.050 808.200 ;
        RECT 521.400 805.350 522.600 806.100 ;
        RECT 527.400 805.350 528.600 806.100 ;
        RECT 520.950 802.950 523.050 805.050 ;
        RECT 523.950 802.950 526.050 805.050 ;
        RECT 526.950 802.950 529.050 805.050 ;
        RECT 529.950 802.950 532.050 805.050 ;
        RECT 524.400 801.900 525.600 802.650 ;
        RECT 511.950 796.950 514.050 799.050 ;
        RECT 514.950 796.950 517.050 801.900 ;
        RECT 523.950 799.800 526.050 801.900 ;
        RECT 530.400 800.400 531.600 802.650 ;
        RECT 499.950 793.950 502.050 796.050 ;
        RECT 496.950 766.950 499.050 769.050 ;
        RECT 500.400 766.050 501.450 793.950 ;
        RECT 530.400 793.050 531.450 800.400 ;
        RECT 529.950 790.950 532.050 793.050 ;
        RECT 505.950 769.950 508.050 772.050 ;
        RECT 526.950 769.950 529.050 772.050 ;
        RECT 499.950 762.000 502.050 766.050 ;
        RECT 506.400 762.600 507.450 769.950 ;
        RECT 500.400 760.350 501.600 762.000 ;
        RECT 506.400 760.350 507.600 762.600 ;
        RECT 520.950 762.000 523.050 766.050 ;
        RECT 527.400 762.600 528.450 769.950 ;
        RECT 521.400 760.350 522.600 762.000 ;
        RECT 527.400 760.350 528.600 762.600 ;
        RECT 496.950 757.950 499.050 760.050 ;
        RECT 499.950 757.950 502.050 760.050 ;
        RECT 502.950 757.950 505.050 760.050 ;
        RECT 505.950 757.950 508.050 760.050 ;
        RECT 520.950 757.950 523.050 760.050 ;
        RECT 523.950 757.950 526.050 760.050 ;
        RECT 526.950 757.950 529.050 760.050 ;
        RECT 529.950 757.950 532.050 760.050 ;
        RECT 490.950 754.950 493.050 757.050 ;
        RECT 497.400 756.900 498.600 757.650 ;
        RECT 496.950 754.800 499.050 756.900 ;
        RECT 503.400 756.000 504.600 757.650 ;
        RECT 487.950 751.950 490.050 754.050 ;
        RECT 502.950 751.950 505.050 756.000 ;
        RECT 524.400 755.400 525.600 757.650 ;
        RECT 530.400 755.400 531.600 757.650 ;
        RECT 536.400 756.450 537.450 806.100 ;
        RECT 539.400 801.900 540.450 808.950 ;
        RECT 548.400 807.600 549.450 814.950 ;
        RECT 548.400 805.350 549.600 807.600 ;
        RECT 544.950 802.950 547.050 805.050 ;
        RECT 547.950 802.950 550.050 805.050 ;
        RECT 550.950 802.950 553.050 805.050 ;
        RECT 545.400 801.900 546.600 802.650 ;
        RECT 538.950 799.800 541.050 801.900 ;
        RECT 544.950 799.800 547.050 801.900 ;
        RECT 551.400 800.400 552.600 802.650 ;
        RECT 533.400 755.400 537.450 756.450 ;
        RECT 524.400 754.050 525.450 755.400 ;
        RECT 523.950 751.950 526.050 754.050 ;
        RECT 487.950 745.950 490.050 748.050 ;
        RECT 482.400 743.400 486.450 744.450 ;
        RECT 481.950 739.950 484.050 742.050 ;
        RECT 482.400 723.900 483.450 739.950 ;
        RECT 485.400 730.050 486.450 743.400 ;
        RECT 484.950 727.950 487.050 730.050 ;
        RECT 488.400 729.600 489.450 745.950 ;
        RECT 499.950 739.950 502.050 742.050 ;
        RECT 505.950 739.950 508.050 742.050 ;
        RECT 488.400 727.350 489.600 729.600 ;
        RECT 493.950 729.000 496.050 733.050 ;
        RECT 500.400 730.050 501.450 739.950 ;
        RECT 502.950 736.950 505.050 739.050 ;
        RECT 494.400 727.350 495.600 729.000 ;
        RECT 499.950 727.950 502.050 730.050 ;
        RECT 487.950 724.950 490.050 727.050 ;
        RECT 490.950 724.950 493.050 727.050 ;
        RECT 493.950 724.950 496.050 727.050 ;
        RECT 496.950 724.950 499.050 727.050 ;
        RECT 491.400 723.900 492.600 724.650 ;
        RECT 497.400 723.900 498.600 724.650 ;
        RECT 503.400 723.900 504.450 736.950 ;
        RECT 481.950 721.800 484.050 723.900 ;
        RECT 490.950 721.800 493.050 723.900 ;
        RECT 496.950 721.800 499.050 723.900 ;
        RECT 502.950 721.800 505.050 723.900 ;
        RECT 506.400 715.050 507.450 739.950 ;
        RECT 514.950 736.950 517.050 739.050 ;
        RECT 515.400 729.600 516.450 736.950 ;
        RECT 520.950 730.950 523.050 733.050 ;
        RECT 515.400 727.350 516.600 729.600 ;
        RECT 511.950 724.950 514.050 727.050 ;
        RECT 514.950 724.950 517.050 727.050 ;
        RECT 512.400 723.900 513.600 724.650 ;
        RECT 511.950 721.800 514.050 723.900 ;
        RECT 487.950 712.950 490.050 715.050 ;
        RECT 505.950 712.950 508.050 715.050 ;
        RECT 478.950 694.950 481.050 697.050 ;
        RECT 484.350 693.300 486.450 695.400 ;
        RECT 485.250 686.700 486.450 693.300 ;
        RECT 484.350 684.600 486.450 686.700 ;
        RECT 467.100 679.950 469.200 682.050 ;
        RECT 472.500 679.950 474.600 682.050 ;
        RECT 478.950 679.950 481.050 682.050 ;
        RECT 448.950 676.800 451.050 678.900 ;
        RECT 460.950 676.800 463.050 678.900 ;
        RECT 473.400 678.000 474.600 679.650 ;
        RECT 479.400 678.000 480.600 679.650 ;
        RECT 472.950 673.950 475.050 678.000 ;
        RECT 478.950 673.950 481.050 678.000 ;
        RECT 485.250 671.700 486.450 684.600 ;
        RECT 436.950 667.950 439.050 670.050 ;
        RECT 484.350 669.600 486.450 671.700 ;
        RECT 488.400 667.050 489.450 712.950 ;
        RECT 521.400 700.050 522.450 730.950 ;
        RECT 520.950 697.950 523.050 700.050 ;
        RECT 505.950 694.950 508.050 697.050 ;
        RECT 511.950 694.950 514.050 697.050 ;
        RECT 499.650 691.500 501.750 692.400 ;
        RECT 499.650 690.300 503.850 691.500 ;
        RECT 490.950 682.950 493.050 685.050 ;
        RECT 496.950 683.100 499.050 685.200 ;
        RECT 491.400 676.050 492.450 682.950 ;
        RECT 497.400 682.350 498.600 683.100 ;
        RECT 496.800 679.950 498.900 682.050 ;
        RECT 490.950 673.950 493.050 676.050 ;
        RECT 502.650 671.700 503.850 690.300 ;
        RECT 506.400 684.600 507.450 694.950 ;
        RECT 512.400 691.050 513.450 694.950 ;
        RECT 520.350 693.300 522.450 695.400 ;
        RECT 524.400 694.050 525.450 751.950 ;
        RECT 526.950 748.950 529.050 751.050 ;
        RECT 527.400 730.050 528.450 748.950 ;
        RECT 530.400 736.050 531.450 755.400 ;
        RECT 529.950 733.950 532.050 736.050 ;
        RECT 533.400 730.200 534.450 755.400 ;
        RECT 539.400 742.050 540.450 799.800 ;
        RECT 551.400 796.050 552.450 800.400 ;
        RECT 544.950 793.950 547.050 796.050 ;
        RECT 550.950 793.950 553.050 796.050 ;
        RECT 545.400 762.600 546.450 793.950 ;
        RECT 557.400 775.050 558.450 826.950 ;
        RECT 560.400 823.050 561.450 833.400 ;
        RECT 566.400 826.050 567.450 833.400 ;
        RECT 565.950 823.950 568.050 826.050 ;
        RECT 559.950 820.950 562.050 823.050 ;
        RECT 575.400 817.050 576.450 839.100 ;
        RECT 587.400 838.350 588.600 840.000 ;
        RECT 592.950 839.100 595.050 841.200 ;
        RECT 593.400 838.350 594.600 839.100 ;
        RECT 583.950 835.950 586.050 838.050 ;
        RECT 586.950 835.950 589.050 838.050 ;
        RECT 589.950 835.950 592.050 838.050 ;
        RECT 592.950 835.950 595.050 838.050 ;
        RECT 584.400 833.400 585.600 835.650 ;
        RECT 590.400 833.400 591.600 835.650 ;
        RECT 574.950 814.950 577.050 817.050 ;
        RECT 559.950 811.950 562.050 814.050 ;
        RECT 556.950 772.950 559.050 775.050 ;
        RECT 556.950 769.800 559.050 771.900 ;
        RECT 545.400 762.450 546.600 762.600 ;
        RECT 542.400 761.400 546.600 762.450 ;
        RECT 542.400 751.050 543.450 761.400 ;
        RECT 545.400 760.350 546.600 761.400 ;
        RECT 553.950 761.100 556.050 763.200 ;
        RECT 554.400 760.350 555.600 761.100 ;
        RECT 545.100 757.950 547.200 760.050 ;
        RECT 550.500 757.950 552.600 760.050 ;
        RECT 553.800 757.950 555.900 760.050 ;
        RECT 551.400 755.400 552.600 757.650 ;
        RECT 551.400 753.450 552.450 755.400 ;
        RECT 548.400 752.400 552.450 753.450 ;
        RECT 541.950 748.950 544.050 751.050 ;
        RECT 548.400 742.050 549.450 752.400 ;
        RECT 550.950 748.950 553.050 751.050 ;
        RECT 551.400 745.050 552.450 748.950 ;
        RECT 550.950 742.950 553.050 745.050 ;
        RECT 538.950 739.950 541.050 742.050 ;
        RECT 547.950 739.950 550.050 742.050 ;
        RECT 541.950 733.950 544.050 736.050 ;
        RECT 547.950 733.950 550.050 736.050 ;
        RECT 526.950 727.950 529.050 730.050 ;
        RECT 532.950 728.100 535.050 730.200 ;
        RECT 538.950 728.100 541.050 730.200 ;
        RECT 542.400 729.450 543.450 733.950 ;
        RECT 542.400 728.400 546.450 729.450 ;
        RECT 533.400 727.350 534.600 728.100 ;
        RECT 539.400 727.350 540.600 728.100 ;
        RECT 529.950 724.950 532.050 727.050 ;
        RECT 532.950 724.950 535.050 727.050 ;
        RECT 535.950 724.950 538.050 727.050 ;
        RECT 538.950 724.950 541.050 727.050 ;
        RECT 526.950 721.950 529.050 724.050 ;
        RECT 530.400 722.400 531.600 724.650 ;
        RECT 536.400 723.900 537.600 724.650 ;
        RECT 511.950 688.950 514.050 691.050 ;
        RECT 521.250 686.700 522.450 693.300 ;
        RECT 523.950 691.950 526.050 694.050 ;
        RECT 520.350 684.600 522.450 686.700 ;
        RECT 506.400 682.350 507.600 684.600 ;
        RECT 505.950 679.950 508.050 682.050 ;
        RECT 514.950 679.950 517.050 682.050 ;
        RECT 515.400 678.000 516.600 679.650 ;
        RECT 514.950 673.950 517.050 678.000 ;
        RECT 502.050 669.600 504.150 671.700 ;
        RECT 514.950 670.800 517.050 672.900 ;
        RECT 521.250 671.700 522.450 684.600 ;
        RECT 527.400 673.050 528.450 721.950 ;
        RECT 530.400 706.050 531.450 722.400 ;
        RECT 535.950 721.800 538.050 723.900 ;
        RECT 541.950 721.950 544.050 724.050 ;
        RECT 529.950 703.950 532.050 706.050 ;
        RECT 542.400 700.050 543.450 721.950 ;
        RECT 541.950 697.950 544.050 700.050 ;
        RECT 535.650 691.500 537.750 692.400 ;
        RECT 535.650 690.300 539.850 691.500 ;
        RECT 532.950 683.100 535.050 685.200 ;
        RECT 533.400 682.350 534.600 683.100 ;
        RECT 532.800 679.950 534.900 682.050 ;
        RECT 412.950 664.950 415.050 667.050 ;
        RECT 439.950 664.950 442.050 667.050 ;
        RECT 487.950 664.950 490.050 667.050 ;
        RECT 409.950 655.950 412.050 658.050 ;
        RECT 424.950 655.950 427.050 658.050 ;
        RECT 379.950 650.100 382.050 652.200 ;
        RECT 385.950 651.000 388.050 655.050 ;
        RECT 400.950 652.950 403.050 655.050 ;
        RECT 410.400 651.600 411.450 655.950 ;
        RECT 380.400 649.350 381.600 650.100 ;
        RECT 386.400 649.350 387.600 651.000 ;
        RECT 410.400 649.350 411.600 651.600 ;
        RECT 415.950 650.100 418.050 652.200 ;
        RECT 416.400 649.350 417.600 650.100 ;
        RECT 379.950 646.950 382.050 649.050 ;
        RECT 382.950 646.950 385.050 649.050 ;
        RECT 385.950 646.950 388.050 649.050 ;
        RECT 388.950 646.950 391.050 649.050 ;
        RECT 406.950 646.950 409.050 649.050 ;
        RECT 409.950 646.950 412.050 649.050 ;
        RECT 412.950 646.950 415.050 649.050 ;
        RECT 415.950 646.950 418.050 649.050 ;
        RECT 383.400 644.400 384.600 646.650 ;
        RECT 389.400 644.400 390.600 646.650 ;
        RECT 413.400 645.900 414.600 646.650 ;
        RECT 383.400 637.050 384.450 644.400 ;
        RECT 389.400 640.050 390.450 644.400 ;
        RECT 412.950 643.800 415.050 645.900 ;
        RECT 388.950 637.950 391.050 640.050 ;
        RECT 413.400 637.050 414.450 643.800 ;
        RECT 425.400 643.050 426.450 655.950 ;
        RECT 433.950 650.100 436.050 652.200 ;
        RECT 440.400 651.600 441.450 664.950 ;
        RECT 493.950 652.950 496.050 655.050 ;
        RECT 434.400 649.350 435.600 650.100 ;
        RECT 440.400 649.350 441.600 651.600 ;
        RECT 445.950 649.950 448.050 652.050 ;
        RECT 454.950 650.100 457.050 652.200 ;
        RECT 481.950 650.100 484.050 652.200 ;
        RECT 430.950 646.950 433.050 649.050 ;
        RECT 433.950 646.950 436.050 649.050 ;
        RECT 436.950 646.950 439.050 649.050 ;
        RECT 439.950 646.950 442.050 649.050 ;
        RECT 431.400 645.000 432.600 646.650 ;
        RECT 437.400 645.900 438.600 646.650 ;
        RECT 446.400 645.900 447.450 649.950 ;
        RECT 455.400 649.350 456.600 650.100 ;
        RECT 482.400 649.350 483.600 650.100 ;
        RECT 490.950 649.950 493.050 652.050 ;
        RECT 454.950 646.950 457.050 649.050 ;
        RECT 457.950 646.950 460.050 649.050 ;
        RECT 460.950 646.950 463.050 649.050 ;
        RECT 463.950 646.950 466.050 649.050 ;
        RECT 478.950 646.950 481.050 649.050 ;
        RECT 481.950 646.950 484.050 649.050 ;
        RECT 484.950 646.950 487.050 649.050 ;
        RECT 458.400 645.900 459.600 646.650 ;
        RECT 421.950 640.950 424.050 643.050 ;
        RECT 424.950 640.950 427.050 643.050 ;
        RECT 430.950 640.950 433.050 645.000 ;
        RECT 436.950 643.800 439.050 645.900 ;
        RECT 445.950 643.800 448.050 645.900 ;
        RECT 457.950 643.800 460.050 645.900 ;
        RECT 479.400 645.000 480.600 646.650 ;
        RECT 491.400 645.900 492.450 649.950 ;
        RECT 478.950 640.950 481.050 645.000 ;
        RECT 490.950 643.800 493.050 645.900 ;
        RECT 382.950 634.950 385.050 637.050 ;
        RECT 412.950 634.950 415.050 637.050 ;
        RECT 371.400 626.400 375.450 627.450 ;
        RECT 356.400 605.400 360.450 606.450 ;
        RECT 344.400 604.350 345.600 605.100 ;
        RECT 343.950 601.950 346.050 604.050 ;
        RECT 346.950 601.950 349.050 604.050 ;
        RECT 340.950 595.950 343.050 601.050 ;
        RECT 347.400 600.900 348.600 601.650 ;
        RECT 346.950 598.800 349.050 600.900 ;
        RECT 337.950 592.950 340.050 595.050 ;
        RECT 343.950 592.950 346.050 595.050 ;
        RECT 319.950 583.950 322.050 586.050 ;
        RECT 337.950 577.950 340.050 580.050 ;
        RECT 338.400 573.600 339.450 577.950 ;
        RECT 344.400 573.600 345.450 592.950 ;
        RECT 347.400 577.050 348.450 598.800 ;
        RECT 346.950 576.450 349.050 577.050 ;
        RECT 346.950 575.400 351.450 576.450 ;
        RECT 346.950 574.950 349.050 575.400 ;
        RECT 290.100 568.950 292.200 571.050 ;
        RECT 295.500 568.950 297.600 571.050 ;
        RECT 298.800 568.950 300.900 571.050 ;
        RECT 299.400 567.900 300.600 568.650 ;
        RECT 298.950 565.800 301.050 567.900 ;
        RECT 305.400 565.050 306.450 571.950 ;
        RECT 317.400 571.350 318.600 573.600 ;
        RECT 338.400 571.350 339.600 573.600 ;
        RECT 344.400 571.350 345.600 573.600 ;
        RECT 350.400 571.050 351.450 575.400 ;
        RECT 313.950 568.950 316.050 571.050 ;
        RECT 316.950 568.950 319.050 571.050 ;
        RECT 319.950 568.950 322.050 571.050 ;
        RECT 334.950 568.950 337.050 571.050 ;
        RECT 337.950 568.950 340.050 571.050 ;
        RECT 340.950 568.950 343.050 571.050 ;
        RECT 343.950 568.950 346.050 571.050 ;
        RECT 349.950 568.950 352.050 571.050 ;
        RECT 314.400 567.900 315.600 568.650 ;
        RECT 313.950 565.800 316.050 567.900 ;
        RECT 320.400 566.400 321.600 568.650 ;
        RECT 335.400 567.900 336.600 568.650 ;
        RECT 280.950 562.950 283.050 565.050 ;
        RECT 304.950 562.950 307.050 565.050 ;
        RECT 320.400 562.050 321.450 566.400 ;
        RECT 334.950 565.800 337.050 567.900 ;
        RECT 341.400 567.000 342.600 568.650 ;
        RECT 340.950 562.950 343.050 567.000 ;
        RECT 274.950 559.950 277.050 562.050 ;
        RECT 319.950 559.950 322.050 562.050 ;
        RECT 322.950 556.950 325.050 559.050 ;
        RECT 259.950 541.950 262.050 544.050 ;
        RECT 310.950 541.950 313.050 544.050 ;
        RECT 260.400 529.200 261.450 541.950 ;
        RECT 301.950 538.950 304.050 541.050 ;
        RECT 259.950 527.100 262.050 529.200 ;
        RECT 260.400 526.350 261.600 527.100 ;
        RECT 268.950 526.950 271.050 529.050 ;
        RECT 277.950 527.100 280.050 529.200 ;
        RECT 295.950 527.100 298.050 529.200 ;
        RECT 302.400 528.600 303.450 538.950 ;
        RECT 256.950 523.950 259.050 526.050 ;
        RECT 259.950 523.950 262.050 526.050 ;
        RECT 269.400 522.900 270.450 526.950 ;
        RECT 278.400 526.350 279.600 527.100 ;
        RECT 296.400 526.350 297.600 527.100 ;
        RECT 302.400 526.350 303.600 528.600 ;
        RECT 274.950 523.950 277.050 526.050 ;
        RECT 277.950 523.950 280.050 526.050 ;
        RECT 280.950 523.950 283.050 526.050 ;
        RECT 295.950 523.950 298.050 526.050 ;
        RECT 298.950 523.950 301.050 526.050 ;
        RECT 301.950 523.950 304.050 526.050 ;
        RECT 304.950 523.950 307.050 526.050 ;
        RECT 275.400 522.900 276.600 523.650 ;
        RECT 268.950 520.800 271.050 522.900 ;
        RECT 274.950 520.800 277.050 522.900 ;
        RECT 281.400 521.400 282.600 523.650 ;
        RECT 299.400 522.000 300.600 523.650 ;
        RECT 305.400 522.900 306.600 523.650 ;
        RECT 311.400 522.900 312.450 541.950 ;
        RECT 323.400 529.200 324.450 556.950 ;
        RECT 356.400 553.050 357.450 605.400 ;
        RECT 361.950 601.950 364.050 604.050 ;
        RECT 364.950 601.950 367.050 604.050 ;
        RECT 367.950 601.950 370.050 604.050 ;
        RECT 365.400 600.900 366.600 601.650 ;
        RECT 364.950 598.800 367.050 600.900 ;
        RECT 364.950 573.000 367.050 577.050 ;
        RECT 365.400 571.350 366.600 573.000 ;
        RECT 361.950 568.950 364.050 571.050 ;
        RECT 364.950 568.950 367.050 571.050 ;
        RECT 367.950 568.950 370.050 571.050 ;
        RECT 374.400 559.050 375.450 626.400 ;
        RECT 383.400 613.050 384.450 634.950 ;
        RECT 418.950 622.950 421.050 625.050 ;
        RECT 376.950 610.950 379.050 613.050 ;
        RECT 382.950 610.950 385.050 613.050 ;
        RECT 391.950 610.950 394.050 613.050 ;
        RECT 377.400 601.050 378.450 610.950 ;
        RECT 385.950 605.100 388.050 607.200 ;
        RECT 392.400 606.600 393.450 610.950 ;
        RECT 386.400 604.350 387.600 605.100 ;
        RECT 392.400 604.350 393.600 606.600 ;
        RECT 400.950 605.100 403.050 607.200 ;
        RECT 382.950 601.950 385.050 604.050 ;
        RECT 385.950 601.950 388.050 604.050 ;
        RECT 388.950 601.950 391.050 604.050 ;
        RECT 391.950 601.950 394.050 604.050 ;
        RECT 376.950 598.950 379.050 601.050 ;
        RECT 383.400 599.400 384.600 601.650 ;
        RECT 389.400 599.400 390.600 601.650 ;
        RECT 383.400 586.050 384.450 599.400 ;
        RECT 389.400 592.050 390.450 599.400 ;
        RECT 388.950 589.950 391.050 592.050 ;
        RECT 382.950 583.950 385.050 586.050 ;
        RECT 385.950 577.950 388.050 580.050 ;
        RECT 386.400 573.600 387.450 577.950 ;
        RECT 386.400 571.350 387.600 573.600 ;
        RECT 391.950 572.100 394.050 574.200 ;
        RECT 392.400 571.350 393.600 572.100 ;
        RECT 382.950 568.950 385.050 571.050 ;
        RECT 385.950 568.950 388.050 571.050 ;
        RECT 388.950 568.950 391.050 571.050 ;
        RECT 391.950 568.950 394.050 571.050 ;
        RECT 383.400 566.400 384.600 568.650 ;
        RECT 389.400 566.400 390.600 568.650 ;
        RECT 401.400 567.450 402.450 605.100 ;
        RECT 406.950 601.950 409.050 604.050 ;
        RECT 409.950 601.950 412.050 604.050 ;
        RECT 412.950 601.950 415.050 604.050 ;
        RECT 410.400 600.900 411.600 601.650 ;
        RECT 409.950 598.800 412.050 600.900 ;
        RECT 415.950 572.100 418.050 574.200 ;
        RECT 406.950 568.950 409.050 571.050 ;
        RECT 409.950 568.950 412.050 571.050 ;
        RECT 410.400 567.900 411.600 568.650 ;
        RECT 416.400 568.050 417.450 572.100 ;
        RECT 401.400 566.400 405.450 567.450 ;
        RECT 383.400 559.050 384.450 566.400 ;
        RECT 385.950 559.950 388.050 562.050 ;
        RECT 373.950 556.950 376.050 559.050 ;
        RECT 382.950 556.950 385.050 559.050 ;
        RECT 355.950 550.950 358.050 553.050 ;
        RECT 386.400 544.050 387.450 559.950 ;
        RECT 389.400 553.050 390.450 566.400 ;
        RECT 388.950 550.950 391.050 553.050 ;
        RECT 389.400 547.050 390.450 550.950 ;
        RECT 404.400 550.050 405.450 566.400 ;
        RECT 409.950 565.800 412.050 567.900 ;
        RECT 415.950 565.950 418.050 568.050 ;
        RECT 419.400 562.050 420.450 622.950 ;
        RECT 422.400 601.050 423.450 640.950 ;
        RECT 494.400 637.050 495.450 652.950 ;
        RECT 499.950 650.100 502.050 652.200 ;
        RECT 505.950 651.000 508.050 655.050 ;
        RECT 500.400 649.350 501.600 650.100 ;
        RECT 506.400 649.350 507.600 651.000 ;
        RECT 499.950 646.950 502.050 649.050 ;
        RECT 502.950 646.950 505.050 649.050 ;
        RECT 505.950 646.950 508.050 649.050 ;
        RECT 508.950 646.950 511.050 649.050 ;
        RECT 503.400 645.900 504.600 646.650 ;
        RECT 509.400 645.900 510.600 646.650 ;
        RECT 515.400 646.050 516.450 670.800 ;
        RECT 520.350 669.600 522.450 671.700 ;
        RECT 526.950 670.950 529.050 673.050 ;
        RECT 538.650 671.700 539.850 690.300 ;
        RECT 541.950 688.950 544.050 691.050 ;
        RECT 542.400 684.600 543.450 688.950 ;
        RECT 545.400 688.050 546.450 728.400 ;
        RECT 548.400 715.050 549.450 733.950 ;
        RECT 557.400 729.600 558.450 769.800 ;
        RECT 560.400 736.050 561.450 811.950 ;
        RECT 568.950 807.000 571.050 811.050 ;
        RECT 569.400 805.350 570.600 807.000 ;
        RECT 574.950 806.100 577.050 808.200 ;
        RECT 575.400 805.350 576.600 806.100 ;
        RECT 565.950 802.950 568.050 805.050 ;
        RECT 568.950 802.950 571.050 805.050 ;
        RECT 571.950 802.950 574.050 805.050 ;
        RECT 574.950 802.950 577.050 805.050 ;
        RECT 577.950 802.950 580.050 805.050 ;
        RECT 566.400 800.400 567.600 802.650 ;
        RECT 572.400 801.000 573.600 802.650 ;
        RECT 566.400 796.050 567.450 800.400 ;
        RECT 571.950 796.950 574.050 801.000 ;
        RECT 578.400 800.400 579.600 802.650 ;
        RECT 578.400 798.450 579.450 800.400 ;
        RECT 580.950 799.950 583.050 802.050 ;
        RECT 575.400 797.400 579.450 798.450 ;
        RECT 565.950 793.950 568.050 796.050 ;
        RECT 575.400 793.050 576.450 797.400 ;
        RECT 577.950 795.450 580.050 796.050 ;
        RECT 581.400 795.450 582.450 799.950 ;
        RECT 577.950 794.400 582.450 795.450 ;
        RECT 577.950 793.950 580.050 794.400 ;
        RECT 574.950 790.950 577.050 793.050 ;
        RECT 562.950 772.950 565.050 775.050 ;
        RECT 563.400 745.050 564.450 772.950 ;
        RECT 571.950 761.100 574.050 763.200 ;
        RECT 578.400 762.600 579.450 793.950 ;
        RECT 584.400 781.050 585.450 833.400 ;
        RECT 590.400 826.050 591.450 833.400 ;
        RECT 599.400 829.050 600.450 841.950 ;
        RECT 604.950 839.100 607.050 841.200 ;
        RECT 610.950 839.100 613.050 841.200 ;
        RECT 617.400 840.600 618.450 844.950 ;
        RECT 598.950 826.950 601.050 829.050 ;
        RECT 589.950 823.950 592.050 826.050 ;
        RECT 605.400 820.050 606.450 839.100 ;
        RECT 611.400 838.350 612.600 839.100 ;
        RECT 617.400 838.350 618.600 840.600 ;
        RECT 610.950 835.950 613.050 838.050 ;
        RECT 613.950 835.950 616.050 838.050 ;
        RECT 616.950 835.950 619.050 838.050 ;
        RECT 619.950 835.950 622.050 838.050 ;
        RECT 614.400 833.400 615.600 835.650 ;
        RECT 620.400 834.900 621.600 835.650 ;
        RECT 626.400 834.900 627.450 850.950 ;
        RECT 637.950 844.950 640.050 847.050 ;
        RECT 649.950 844.950 652.050 847.050 ;
        RECT 638.400 840.600 639.450 844.950 ;
        RECT 638.400 838.350 639.600 840.600 ;
        RECT 643.950 839.100 646.050 841.200 ;
        RECT 644.400 838.350 645.600 839.100 ;
        RECT 634.950 835.950 637.050 838.050 ;
        RECT 637.950 835.950 640.050 838.050 ;
        RECT 640.950 835.950 643.050 838.050 ;
        RECT 643.950 835.950 646.050 838.050 ;
        RECT 635.400 834.900 636.600 835.650 ;
        RECT 614.400 829.050 615.450 833.400 ;
        RECT 619.950 832.800 622.050 834.900 ;
        RECT 625.950 832.800 628.050 834.900 ;
        RECT 634.950 832.800 637.050 834.900 ;
        RECT 641.400 833.400 642.600 835.650 ;
        RECT 650.400 835.050 651.450 844.950 ;
        RECT 613.950 826.950 616.050 829.050 ;
        RECT 625.950 826.950 628.050 829.050 ;
        RECT 626.400 820.050 627.450 826.950 ;
        RECT 604.950 817.950 607.050 820.050 ;
        RECT 625.950 817.950 628.050 820.050 ;
        RECT 592.950 814.950 595.050 817.050 ;
        RECT 593.400 807.600 594.450 814.950 ;
        RECT 641.400 814.050 642.450 833.400 ;
        RECT 649.950 832.950 652.050 835.050 ;
        RECT 643.950 814.950 646.050 817.050 ;
        RECT 631.950 811.950 634.050 814.050 ;
        RECT 640.950 811.950 643.050 814.050 ;
        RECT 593.400 805.350 594.600 807.600 ;
        RECT 598.950 807.000 601.050 811.050 ;
        RECT 607.950 808.950 610.050 811.050 ;
        RECT 599.400 805.350 600.600 807.000 ;
        RECT 592.950 802.950 595.050 805.050 ;
        RECT 595.950 802.950 598.050 805.050 ;
        RECT 598.950 802.950 601.050 805.050 ;
        RECT 601.950 802.950 604.050 805.050 ;
        RECT 596.400 801.900 597.600 802.650 ;
        RECT 595.950 799.800 598.050 801.900 ;
        RECT 602.400 800.400 603.600 802.650 ;
        RECT 602.400 796.050 603.450 800.400 ;
        RECT 601.950 793.950 604.050 796.050 ;
        RECT 608.400 784.050 609.450 808.950 ;
        RECT 613.950 806.100 616.050 808.200 ;
        RECT 619.950 806.100 622.050 808.200 ;
        RECT 614.400 796.050 615.450 806.100 ;
        RECT 620.400 805.350 621.600 806.100 ;
        RECT 619.950 802.950 622.050 805.050 ;
        RECT 622.950 802.950 625.050 805.050 ;
        RECT 623.400 800.400 624.600 802.650 ;
        RECT 613.950 793.950 616.050 796.050 ;
        RECT 607.950 781.950 610.050 784.050 ;
        RECT 583.950 778.950 586.050 781.050 ;
        RECT 604.950 766.950 607.050 769.050 ;
        RECT 613.950 766.950 616.050 769.050 ;
        RECT 572.400 760.350 573.600 761.100 ;
        RECT 578.400 760.350 579.600 762.600 ;
        RECT 595.950 762.000 598.050 766.050 ;
        RECT 596.400 760.350 597.600 762.000 ;
        RECT 568.950 757.950 571.050 760.050 ;
        RECT 571.950 757.950 574.050 760.050 ;
        RECT 574.950 757.950 577.050 760.050 ;
        RECT 577.950 757.950 580.050 760.050 ;
        RECT 592.950 757.950 595.050 760.050 ;
        RECT 595.950 757.950 598.050 760.050 ;
        RECT 569.400 756.900 570.600 757.650 ;
        RECT 575.400 756.900 576.600 757.650 ;
        RECT 568.950 754.800 571.050 756.900 ;
        RECT 574.950 754.800 577.050 756.900 ;
        RECT 593.400 755.400 594.600 757.650 ;
        RECT 593.400 751.050 594.450 755.400 ;
        RECT 565.950 748.950 568.050 751.050 ;
        RECT 592.950 748.950 595.050 751.050 ;
        RECT 562.950 742.950 565.050 745.050 ;
        RECT 562.950 736.950 565.050 739.050 ;
        RECT 559.950 733.950 562.050 736.050 ;
        RECT 563.400 729.600 564.450 736.950 ;
        RECT 566.400 730.050 567.450 748.950 ;
        RECT 568.950 742.950 571.050 745.050 ;
        RECT 557.400 727.350 558.600 729.600 ;
        RECT 563.400 727.350 564.600 729.600 ;
        RECT 565.950 727.950 568.050 730.050 ;
        RECT 553.950 724.950 556.050 727.050 ;
        RECT 556.950 724.950 559.050 727.050 ;
        RECT 559.950 724.950 562.050 727.050 ;
        RECT 562.950 724.950 565.050 727.050 ;
        RECT 554.400 723.900 555.600 724.650 ;
        RECT 553.950 721.800 556.050 723.900 ;
        RECT 560.400 723.000 561.600 724.650 ;
        RECT 559.950 718.950 562.050 723.000 ;
        RECT 547.950 712.950 550.050 715.050 ;
        RECT 562.950 712.950 565.050 715.050 ;
        RECT 544.950 685.950 547.050 688.050 ;
        RECT 542.400 682.350 543.600 684.600 ;
        RECT 550.950 683.100 553.050 685.200 ;
        RECT 563.400 684.600 564.450 712.950 ;
        RECT 569.400 685.050 570.450 742.950 ;
        RECT 605.400 739.050 606.450 766.950 ;
        RECT 614.400 762.600 615.450 766.950 ;
        RECT 623.400 766.050 624.450 800.400 ;
        RECT 632.400 793.050 633.450 811.950 ;
        RECT 637.950 806.100 640.050 808.200 ;
        RECT 644.400 807.600 645.450 814.950 ;
        RECT 638.400 805.350 639.600 806.100 ;
        RECT 644.400 805.350 645.600 807.600 ;
        RECT 637.950 802.950 640.050 805.050 ;
        RECT 640.950 802.950 643.050 805.050 ;
        RECT 643.950 802.950 646.050 805.050 ;
        RECT 646.950 802.950 649.050 805.050 ;
        RECT 641.400 801.900 642.600 802.650 ;
        RECT 647.400 801.900 648.600 802.650 ;
        RECT 640.950 799.800 643.050 801.900 ;
        RECT 646.950 799.800 649.050 801.900 ;
        RECT 631.950 790.950 634.050 793.050 ;
        RECT 614.400 760.350 615.600 762.600 ;
        RECT 619.950 762.000 622.050 766.050 ;
        RECT 622.950 763.950 625.050 766.050 ;
        RECT 632.400 762.450 633.450 790.950 ;
        RECT 620.400 760.350 621.600 762.000 ;
        RECT 629.400 761.400 633.450 762.450 ;
        RECT 610.950 757.950 613.050 760.050 ;
        RECT 613.950 757.950 616.050 760.050 ;
        RECT 616.950 757.950 619.050 760.050 ;
        RECT 619.950 757.950 622.050 760.050 ;
        RECT 611.400 755.400 612.600 757.650 ;
        RECT 617.400 755.400 618.600 757.650 ;
        RECT 629.400 756.900 630.450 761.400 ;
        RECT 634.950 761.100 637.050 763.200 ;
        RECT 640.950 762.000 643.050 766.050 ;
        RECT 653.400 765.450 654.450 875.400 ;
        RECT 655.950 874.950 658.050 875.400 ;
        RECT 662.400 868.050 663.450 878.400 ;
        RECT 668.400 874.050 669.450 878.400 ;
        RECT 667.950 871.950 670.050 874.050 ;
        RECT 661.950 865.950 664.050 868.050 ;
        RECT 667.950 850.950 670.050 853.050 ;
        RECT 668.400 847.050 669.450 850.950 ;
        RECT 683.400 850.050 684.450 883.950 ;
        RECT 710.400 883.350 711.600 885.600 ;
        RECT 730.950 884.100 733.050 886.200 ;
        RECT 731.400 883.350 732.600 884.100 ;
        RECT 739.800 883.950 741.900 886.050 ;
        RECT 742.950 883.950 745.050 886.050 ;
        RECT 751.950 884.100 754.050 886.200 ;
        RECT 688.950 880.950 691.050 883.050 ;
        RECT 691.950 880.950 694.050 883.050 ;
        RECT 706.950 880.950 709.050 883.050 ;
        RECT 709.950 880.950 712.050 883.050 ;
        RECT 712.950 880.950 715.050 883.050 ;
        RECT 727.950 880.950 730.050 883.050 ;
        RECT 730.950 880.950 733.050 883.050 ;
        RECT 733.950 880.950 736.050 883.050 ;
        RECT 689.400 879.000 690.600 880.650 ;
        RECT 707.400 879.000 708.600 880.650 ;
        RECT 713.400 879.900 714.600 880.650 ;
        RECT 728.400 879.900 729.600 880.650 ;
        RECT 688.950 874.950 691.050 879.000 ;
        RECT 706.950 874.950 709.050 879.000 ;
        RECT 712.950 877.800 715.050 879.900 ;
        RECT 727.950 877.800 730.050 879.900 ;
        RECT 740.400 856.050 741.450 883.950 ;
        RECT 743.400 879.900 744.450 883.950 ;
        RECT 752.400 883.350 753.600 884.100 ;
        RECT 748.950 880.950 751.050 883.050 ;
        RECT 751.950 880.950 754.050 883.050 ;
        RECT 754.950 880.950 757.050 883.050 ;
        RECT 742.950 877.800 745.050 879.900 ;
        RECT 749.400 878.400 750.600 880.650 ;
        RECT 755.400 879.900 756.600 880.650 ;
        RECT 749.400 865.050 750.450 878.400 ;
        RECT 754.950 877.800 757.050 879.900 ;
        RECT 748.950 862.950 751.050 865.050 ;
        RECT 715.950 853.950 718.050 856.050 ;
        RECT 739.950 853.950 742.050 856.050 ;
        RECT 682.950 847.950 685.050 850.050 ;
        RECT 709.950 847.950 712.050 850.050 ;
        RECT 667.950 844.950 670.050 847.050 ;
        RECT 663.000 843.450 667.050 844.050 ;
        RECT 662.400 841.950 667.050 843.450 ;
        RECT 662.400 841.200 663.450 841.950 ;
        RECT 661.950 839.100 664.050 841.200 ;
        RECT 679.950 840.000 682.050 844.050 ;
        RECT 662.400 838.350 663.600 839.100 ;
        RECT 680.400 838.350 681.600 840.000 ;
        RECT 685.950 839.100 688.050 841.200 ;
        RECT 691.800 839.100 693.900 841.200 ;
        RECT 694.950 839.100 697.050 841.200 ;
        RECT 703.950 839.100 706.050 841.200 ;
        RECT 710.400 840.600 711.450 847.950 ;
        RECT 686.400 838.350 687.600 839.100 ;
        RECT 658.950 835.950 661.050 838.050 ;
        RECT 661.950 835.950 664.050 838.050 ;
        RECT 676.950 835.950 679.050 838.050 ;
        RECT 679.950 835.950 682.050 838.050 ;
        RECT 682.950 835.950 685.050 838.050 ;
        RECT 685.950 835.950 688.050 838.050 ;
        RECT 659.400 833.400 660.600 835.650 ;
        RECT 677.400 833.400 678.600 835.650 ;
        RECT 683.400 833.400 684.600 835.650 ;
        RECT 659.400 829.050 660.450 833.400 ;
        RECT 658.950 826.950 661.050 829.050 ;
        RECT 655.950 820.950 658.050 823.050 ;
        RECT 656.400 801.900 657.450 820.950 ;
        RECT 659.400 808.050 660.450 826.950 ;
        RECT 677.400 826.050 678.450 833.400 ;
        RECT 676.950 823.950 679.050 826.050 ;
        RECT 683.400 823.050 684.450 833.400 ;
        RECT 682.950 820.950 685.050 823.050 ;
        RECT 688.950 817.950 691.050 820.050 ;
        RECT 664.950 814.950 667.050 817.050 ;
        RECT 658.950 805.950 661.050 808.050 ;
        RECT 665.400 807.600 666.450 814.950 ;
        RECT 665.400 805.350 666.600 807.600 ;
        RECT 670.950 806.100 673.050 808.200 ;
        RECT 689.400 807.600 690.450 817.950 ;
        RECT 692.400 817.050 693.450 839.100 ;
        RECT 695.400 820.050 696.450 839.100 ;
        RECT 704.400 838.350 705.600 839.100 ;
        RECT 710.400 838.350 711.600 840.600 ;
        RECT 700.950 835.950 703.050 838.050 ;
        RECT 703.950 835.950 706.050 838.050 ;
        RECT 706.950 835.950 709.050 838.050 ;
        RECT 709.950 835.950 712.050 838.050 ;
        RECT 701.400 834.900 702.600 835.650 ;
        RECT 700.950 832.800 703.050 834.900 ;
        RECT 707.400 834.000 708.600 835.650 ;
        RECT 706.950 829.950 709.050 834.000 ;
        RECT 712.950 832.950 715.050 835.050 ;
        RECT 713.400 823.050 714.450 832.950 ;
        RECT 716.400 832.050 717.450 853.950 ;
        RECT 727.950 847.950 730.050 850.050 ;
        RECT 728.400 840.600 729.450 847.950 ;
        RECT 728.400 838.350 729.600 840.600 ;
        RECT 733.950 839.100 736.050 841.200 ;
        RECT 734.400 838.350 735.600 839.100 ;
        RECT 724.950 835.950 727.050 838.050 ;
        RECT 727.950 835.950 730.050 838.050 ;
        RECT 730.950 835.950 733.050 838.050 ;
        RECT 733.950 835.950 736.050 838.050 ;
        RECT 725.400 834.900 726.600 835.650 ;
        RECT 731.400 834.900 732.600 835.650 ;
        RECT 740.400 834.900 741.450 853.950 ;
        RECT 745.950 844.950 748.050 847.050 ;
        RECT 746.400 835.050 747.450 844.950 ;
        RECT 761.400 841.200 762.450 889.950 ;
        RECT 871.950 886.950 874.050 889.050 ;
        RECT 793.950 884.100 796.050 886.200 ;
        RECT 794.400 883.350 795.600 884.100 ;
        RECT 802.950 883.950 805.050 886.050 ;
        RECT 808.950 883.950 811.050 886.050 ;
        RECT 817.950 884.100 820.050 886.200 ;
        RECT 829.950 884.100 832.050 886.200 ;
        RECT 835.950 884.100 838.050 886.200 ;
        RECT 841.950 884.100 844.050 886.200 ;
        RECT 847.950 884.100 850.050 886.200 ;
        RECT 862.950 884.100 865.050 886.200 ;
        RECT 868.950 884.100 871.050 886.200 ;
        RECT 770.400 880.950 772.500 883.050 ;
        RECT 775.800 880.950 777.900 883.050 ;
        RECT 790.950 880.950 793.050 883.050 ;
        RECT 793.950 880.950 796.050 883.050 ;
        RECT 796.950 880.950 799.050 883.050 ;
        RECT 776.400 879.900 777.600 880.650 ;
        RECT 775.950 877.800 778.050 879.900 ;
        RECT 797.400 878.400 798.600 880.650 ;
        RECT 803.400 879.900 804.450 883.950 ;
        RECT 776.400 874.050 777.450 877.800 ;
        RECT 797.400 874.050 798.450 878.400 ;
        RECT 802.950 877.800 805.050 879.900 ;
        RECT 775.950 871.950 778.050 874.050 ;
        RECT 784.950 871.950 787.050 874.050 ;
        RECT 796.950 871.950 799.050 874.050 ;
        RECT 769.950 862.950 772.050 865.050 ;
        RECT 754.950 839.100 757.050 841.200 ;
        RECT 760.950 839.100 763.050 841.200 ;
        RECT 755.400 838.350 756.600 839.100 ;
        RECT 761.400 838.350 762.600 839.100 ;
        RECT 766.950 838.800 769.050 840.900 ;
        RECT 751.950 835.950 754.050 838.050 ;
        RECT 754.950 835.950 757.050 838.050 ;
        RECT 757.950 835.950 760.050 838.050 ;
        RECT 760.950 835.950 763.050 838.050 ;
        RECT 724.950 832.800 727.050 834.900 ;
        RECT 730.950 832.800 733.050 834.900 ;
        RECT 739.950 832.800 742.050 834.900 ;
        RECT 745.950 832.950 748.050 835.050 ;
        RECT 752.400 834.900 753.600 835.650 ;
        RECT 751.950 832.800 754.050 834.900 ;
        RECT 758.400 833.400 759.600 835.650 ;
        RECT 715.950 829.950 718.050 832.050 ;
        RECT 754.950 829.950 757.050 832.050 ;
        RECT 751.950 823.950 754.050 826.050 ;
        RECT 712.950 820.950 715.050 823.050 ;
        RECT 694.950 817.950 697.050 820.050 ;
        RECT 733.950 817.950 736.050 820.050 ;
        RECT 748.950 817.950 751.050 820.050 ;
        RECT 691.950 814.950 694.050 817.050 ;
        RECT 706.950 814.950 709.050 817.050 ;
        RECT 724.950 814.950 727.050 817.050 ;
        RECT 707.400 807.600 708.450 814.950 ;
        RECT 721.950 811.950 724.050 814.050 ;
        RECT 671.400 805.350 672.600 806.100 ;
        RECT 689.400 805.350 690.600 807.600 ;
        RECT 707.400 805.350 708.600 807.600 ;
        RECT 712.950 806.100 715.050 808.200 ;
        RECT 713.400 805.350 714.600 806.100 ;
        RECT 661.950 802.950 664.050 805.050 ;
        RECT 664.950 802.950 667.050 805.050 ;
        RECT 667.950 802.950 670.050 805.050 ;
        RECT 670.950 802.950 673.050 805.050 ;
        RECT 685.950 802.950 688.050 805.050 ;
        RECT 688.950 802.950 691.050 805.050 ;
        RECT 691.950 802.950 694.050 805.050 ;
        RECT 706.950 802.950 709.050 805.050 ;
        RECT 709.950 802.950 712.050 805.050 ;
        RECT 712.950 802.950 715.050 805.050 ;
        RECT 715.950 802.950 718.050 805.050 ;
        RECT 662.400 801.900 663.600 802.650 ;
        RECT 655.950 796.950 658.050 801.900 ;
        RECT 661.950 799.800 664.050 801.900 ;
        RECT 668.400 801.000 669.600 802.650 ;
        RECT 667.950 796.950 670.050 801.000 ;
        RECT 673.950 799.950 676.050 802.050 ;
        RECT 710.400 801.000 711.600 802.650 ;
        RECT 716.400 801.900 717.600 802.650 ;
        RECT 722.400 801.900 723.450 811.950 ;
        RECT 725.400 808.200 726.450 814.950 ;
        RECT 724.950 806.100 727.050 808.200 ;
        RECT 734.400 807.600 735.450 817.950 ;
        RECT 749.400 807.600 750.450 817.950 ;
        RECT 752.400 811.050 753.450 823.950 ;
        RECT 755.400 817.050 756.450 829.950 ;
        RECT 758.400 820.050 759.450 833.400 ;
        RECT 757.950 817.950 760.050 820.050 ;
        RECT 763.950 817.950 766.050 820.050 ;
        RECT 754.950 814.950 757.050 817.050 ;
        RECT 758.400 814.050 759.450 817.950 ;
        RECT 757.950 811.950 760.050 814.050 ;
        RECT 751.950 808.950 754.050 811.050 ;
        RECT 725.400 802.050 726.450 806.100 ;
        RECT 734.400 805.350 735.600 807.600 ;
        RECT 749.400 805.350 750.600 807.600 ;
        RECT 754.950 806.100 757.050 808.200 ;
        RECT 755.400 805.350 756.600 806.100 ;
        RECT 730.950 802.950 733.050 805.050 ;
        RECT 733.950 802.950 736.050 805.050 ;
        RECT 748.950 802.950 751.050 805.050 ;
        RECT 751.950 802.950 754.050 805.050 ;
        RECT 754.950 802.950 757.050 805.050 ;
        RECT 757.950 802.950 760.050 805.050 ;
        RECT 674.400 796.050 675.450 799.950 ;
        RECT 709.950 796.950 712.050 801.000 ;
        RECT 715.950 799.800 718.050 801.900 ;
        RECT 721.800 799.800 723.900 801.900 ;
        RECT 724.950 799.950 727.050 802.050 ;
        RECT 731.400 801.900 732.600 802.650 ;
        RECT 752.400 801.900 753.600 802.650 ;
        RECT 758.400 801.900 759.600 802.650 ;
        RECT 764.400 801.900 765.450 817.950 ;
        RECT 730.950 799.800 733.050 801.900 ;
        RECT 751.950 799.800 754.050 801.900 ;
        RECT 757.950 799.800 760.050 801.900 ;
        RECT 763.950 799.800 766.050 801.900 ;
        RECT 767.400 799.050 768.450 838.800 ;
        RECT 770.400 834.900 771.450 862.950 ;
        RECT 785.400 841.200 786.450 871.950 ;
        RECT 790.950 850.950 793.050 853.050 ;
        RECT 784.950 839.100 787.050 841.200 ;
        RECT 785.400 838.350 786.600 839.100 ;
        RECT 775.950 835.950 778.050 838.050 ;
        RECT 778.950 835.950 781.050 838.050 ;
        RECT 781.950 835.950 784.050 838.050 ;
        RECT 784.950 835.950 787.050 838.050 ;
        RECT 769.950 832.800 772.050 834.900 ;
        RECT 776.400 833.400 777.600 835.650 ;
        RECT 782.400 834.900 783.600 835.650 ;
        RECT 776.400 826.050 777.450 833.400 ;
        RECT 781.950 832.800 784.050 834.900 ;
        RECT 782.400 829.050 783.450 832.800 ;
        RECT 781.950 828.450 784.050 829.050 ;
        RECT 781.950 827.400 786.450 828.450 ;
        RECT 781.950 826.950 784.050 827.400 ;
        RECT 775.950 823.950 778.050 826.050 ;
        RECT 775.950 811.950 778.050 814.050 ;
        RECT 776.400 808.200 777.450 811.950 ;
        RECT 775.950 806.100 778.050 808.200 ;
        RECT 776.400 805.350 777.600 806.100 ;
        RECT 772.950 802.950 775.050 805.050 ;
        RECT 775.950 802.950 778.050 805.050 ;
        RECT 778.950 802.950 781.050 805.050 ;
        RECT 779.400 801.450 780.600 802.650 ;
        RECT 785.400 801.450 786.450 827.400 ;
        RECT 791.400 807.450 792.450 850.950 ;
        RECT 809.400 844.200 810.450 883.950 ;
        RECT 818.400 883.350 819.600 884.100 ;
        RECT 814.950 880.950 817.050 883.050 ;
        RECT 817.950 880.950 820.050 883.050 ;
        RECT 820.950 880.950 823.050 883.050 ;
        RECT 815.400 879.900 816.600 880.650 ;
        RECT 814.950 877.800 817.050 879.900 ;
        RECT 815.400 859.050 816.450 877.800 ;
        RECT 830.400 874.050 831.450 884.100 ;
        RECT 836.400 883.350 837.600 884.100 ;
        RECT 842.400 883.350 843.600 884.100 ;
        RECT 835.950 880.950 838.050 883.050 ;
        RECT 838.950 880.950 841.050 883.050 ;
        RECT 841.950 880.950 844.050 883.050 ;
        RECT 839.400 878.400 840.600 880.650 ;
        RECT 839.400 876.450 840.450 878.400 ;
        RECT 848.400 877.050 849.450 884.100 ;
        RECT 863.400 883.350 864.600 884.100 ;
        RECT 859.950 880.950 862.050 883.050 ;
        RECT 862.950 880.950 865.050 883.050 ;
        RECT 860.400 878.400 861.600 880.650 ;
        RECT 836.400 875.400 840.450 876.450 ;
        RECT 829.950 871.950 832.050 874.050 ;
        RECT 814.950 856.950 817.050 859.050 ;
        RECT 836.400 853.050 837.450 875.400 ;
        RECT 847.950 874.950 850.050 877.050 ;
        RECT 838.950 871.950 841.050 874.050 ;
        RECT 835.950 850.950 838.050 853.050 ;
        RECT 808.950 842.100 811.050 844.200 ;
        RECT 817.950 841.950 820.050 844.050 ;
        RECT 808.950 838.950 811.050 841.050 ;
        RECT 809.400 838.350 810.600 838.950 ;
        RECT 799.950 835.950 802.050 838.050 ;
        RECT 802.950 835.950 805.050 838.050 ;
        RECT 805.950 835.950 808.050 838.050 ;
        RECT 808.950 835.950 811.050 838.050 ;
        RECT 800.400 833.400 801.600 835.650 ;
        RECT 806.400 833.400 807.600 835.650 ;
        RECT 800.400 820.050 801.450 833.400 ;
        RECT 806.400 829.050 807.450 833.400 ;
        RECT 805.950 826.950 808.050 829.050 ;
        RECT 808.950 823.950 811.050 826.050 ;
        RECT 799.950 817.950 802.050 820.050 ;
        RECT 805.950 817.950 808.050 820.050 ;
        RECT 795.000 810.450 799.050 811.050 ;
        RECT 779.400 800.400 786.450 801.450 ;
        RECT 788.400 806.400 792.450 807.450 ;
        RECT 794.400 808.950 799.050 810.450 ;
        RECT 794.400 807.600 795.450 808.950 ;
        RECT 806.400 808.200 807.450 817.950 ;
        RECT 766.950 796.950 769.050 799.050 ;
        RECT 673.950 793.950 676.050 796.050 ;
        RECT 769.950 781.950 772.050 784.050 ;
        RECT 770.400 769.050 771.450 781.950 ;
        RECT 769.950 766.950 772.050 769.050 ;
        RECT 650.400 764.400 654.450 765.450 ;
        RECT 635.400 760.350 636.600 761.100 ;
        RECT 641.400 760.350 642.600 762.000 ;
        RECT 634.950 757.950 637.050 760.050 ;
        RECT 637.950 757.950 640.050 760.050 ;
        RECT 640.950 757.950 643.050 760.050 ;
        RECT 643.950 757.950 646.050 760.050 ;
        RECT 638.400 756.900 639.600 757.650 ;
        RECT 644.400 756.900 645.600 757.650 ;
        RECT 604.950 736.950 607.050 739.050 ;
        RECT 611.400 733.050 612.450 755.400 ;
        RECT 617.400 751.050 618.450 755.400 ;
        RECT 628.950 754.800 631.050 756.900 ;
        RECT 637.950 754.800 640.050 756.900 ;
        RECT 643.950 754.800 646.050 756.900 ;
        RECT 616.950 748.950 619.050 751.050 ;
        RECT 650.400 748.050 651.450 764.400 ;
        RECT 655.950 761.100 658.050 763.200 ;
        RECT 664.950 761.100 667.050 763.200 ;
        RECT 670.950 762.000 673.050 766.050 ;
        RECT 634.950 745.950 637.050 748.050 ;
        RECT 649.950 745.950 652.050 748.050 ;
        RECT 613.950 736.950 616.050 739.050 ;
        RECT 571.950 727.950 574.050 730.050 ;
        RECT 577.950 728.100 580.050 730.200 ;
        RECT 583.950 729.000 586.050 733.050 ;
        RECT 572.400 721.050 573.450 727.950 ;
        RECT 578.400 727.350 579.600 728.100 ;
        RECT 584.400 727.350 585.600 729.000 ;
        RECT 595.950 728.100 598.050 733.050 ;
        RECT 610.950 730.950 613.050 733.050 ;
        RECT 604.950 728.100 607.050 730.200 ;
        RECT 611.400 729.450 612.600 729.600 ;
        RECT 614.400 729.450 615.450 736.950 ;
        RECT 616.950 730.950 619.050 733.050 ;
        RECT 611.400 728.400 615.450 729.450 ;
        RECT 577.950 724.950 580.050 727.050 ;
        RECT 580.950 724.950 583.050 727.050 ;
        RECT 583.950 724.950 586.050 727.050 ;
        RECT 586.950 724.950 589.050 727.050 ;
        RECT 581.400 723.900 582.600 724.650 ;
        RECT 580.950 721.800 583.050 723.900 ;
        RECT 587.400 722.400 588.600 724.650 ;
        RECT 571.950 718.950 574.050 721.050 ;
        RECT 581.400 718.050 582.450 721.800 ;
        RECT 580.950 715.950 583.050 718.050 ;
        RECT 587.400 709.050 588.450 722.400 ;
        RECT 596.400 718.050 597.450 728.100 ;
        RECT 605.400 727.350 606.600 728.100 ;
        RECT 611.400 727.350 612.600 728.400 ;
        RECT 601.950 724.950 604.050 727.050 ;
        RECT 604.950 724.950 607.050 727.050 ;
        RECT 607.950 724.950 610.050 727.050 ;
        RECT 610.950 724.950 613.050 727.050 ;
        RECT 602.400 723.900 603.600 724.650 ;
        RECT 601.950 721.800 604.050 723.900 ;
        RECT 608.400 722.400 609.600 724.650 ;
        RECT 595.950 715.950 598.050 718.050 ;
        RECT 608.400 709.050 609.450 722.400 ;
        RECT 586.950 706.950 589.050 709.050 ;
        RECT 607.950 706.950 610.050 709.050 ;
        RECT 586.950 691.950 589.050 694.050 ;
        RECT 571.950 685.950 574.050 688.050 ;
        RECT 541.950 679.950 544.050 682.050 ;
        RECT 538.050 669.600 540.150 671.700 ;
        RECT 535.950 655.950 538.050 658.050 ;
        RECT 551.400 657.450 552.450 683.100 ;
        RECT 563.400 682.350 564.600 684.600 ;
        RECT 568.950 682.950 571.050 685.050 ;
        RECT 562.950 679.950 565.050 682.050 ;
        RECT 565.950 679.950 568.050 682.050 ;
        RECT 566.400 678.900 567.600 679.650 ;
        RECT 572.400 678.900 573.450 685.950 ;
        RECT 574.950 682.950 577.050 685.050 ;
        RECT 580.950 684.000 583.050 688.050 ;
        RECT 587.400 685.200 588.450 691.950 ;
        RECT 617.400 685.200 618.450 730.950 ;
        RECT 619.950 728.100 622.050 730.200 ;
        RECT 625.950 728.100 628.050 730.200 ;
        RECT 620.400 724.050 621.450 728.100 ;
        RECT 626.400 727.350 627.600 728.100 ;
        RECT 625.950 724.950 628.050 727.050 ;
        RECT 628.950 724.950 631.050 727.050 ;
        RECT 619.950 723.450 622.050 724.050 ;
        RECT 629.400 723.900 630.600 724.650 ;
        RECT 619.950 722.400 624.450 723.450 ;
        RECT 619.950 721.950 622.050 722.400 ;
        RECT 619.950 691.950 622.050 694.050 ;
        RECT 565.950 676.800 568.050 678.900 ;
        RECT 571.950 676.800 574.050 678.900 ;
        RECT 562.950 667.950 565.050 670.050 ;
        RECT 526.950 650.100 529.050 652.200 ;
        RECT 527.400 649.350 528.600 650.100 ;
        RECT 523.950 646.950 526.050 649.050 ;
        RECT 526.950 646.950 529.050 649.050 ;
        RECT 529.950 646.950 532.050 649.050 ;
        RECT 502.950 643.800 505.050 645.900 ;
        RECT 508.950 643.800 511.050 645.900 ;
        RECT 514.950 643.950 517.050 646.050 ;
        RECT 524.400 645.000 525.600 646.650 ;
        RECT 493.950 634.950 496.050 637.050 ;
        RECT 509.400 634.050 510.450 643.800 ;
        RECT 523.950 640.950 526.050 645.000 ;
        RECT 460.950 631.950 463.050 634.050 ;
        RECT 508.950 631.950 511.050 634.050 ;
        RECT 430.950 605.100 433.050 607.200 ;
        RECT 445.950 605.100 448.050 607.200 ;
        RECT 451.950 605.100 454.050 607.200 ;
        RECT 457.950 605.100 460.050 610.050 ;
        RECT 431.400 604.350 432.600 605.100 ;
        RECT 446.400 604.350 447.600 605.100 ;
        RECT 452.400 604.350 453.600 605.100 ;
        RECT 427.950 601.950 430.050 604.050 ;
        RECT 430.950 601.950 433.050 604.050 ;
        RECT 445.950 601.950 448.050 604.050 ;
        RECT 448.950 601.950 451.050 604.050 ;
        RECT 451.950 601.950 454.050 604.050 ;
        RECT 454.950 601.950 457.050 604.050 ;
        RECT 421.950 598.950 424.050 601.050 ;
        RECT 428.400 600.900 429.600 601.650 ;
        RECT 427.950 598.800 430.050 600.900 ;
        RECT 449.400 599.400 450.600 601.650 ;
        RECT 455.400 600.900 456.600 601.650 ;
        RECT 461.400 601.050 462.450 631.950 ;
        RECT 536.400 622.050 537.450 655.950 ;
        RECT 551.400 655.200 552.600 657.450 ;
        RECT 547.500 653.100 549.600 655.200 ;
        RECT 538.950 650.100 541.050 652.200 ;
        RECT 544.950 650.100 547.050 652.200 ;
        RECT 539.400 622.050 540.450 650.100 ;
        RECT 545.400 649.350 546.600 650.100 ;
        RECT 545.100 646.950 547.200 649.050 ;
        RECT 548.100 648.000 549.000 653.100 ;
        RECT 550.800 652.800 552.900 654.900 ;
        RECT 557.400 653.400 559.500 655.500 ;
        RECT 555.000 651.000 557.100 651.900 ;
        RECT 549.900 649.800 557.100 651.000 ;
        RECT 549.900 648.900 552.000 649.800 ;
        RECT 555.000 648.000 557.100 648.900 ;
        RECT 548.100 647.100 557.100 648.000 ;
        RECT 548.100 640.500 549.000 647.100 ;
        RECT 555.000 646.800 557.100 647.100 ;
        RECT 550.800 643.950 552.900 646.050 ;
        RECT 551.400 641.400 552.600 643.650 ;
        RECT 558.000 640.800 558.900 653.400 ;
        RECT 559.800 646.950 561.900 649.050 ;
        RECT 560.400 645.450 561.600 646.650 ;
        RECT 563.400 645.450 564.450 667.950 ;
        RECT 566.400 645.900 567.450 676.800 ;
        RECT 575.400 670.050 576.450 682.950 ;
        RECT 581.400 682.350 582.600 684.000 ;
        RECT 586.950 683.100 589.050 685.200 ;
        RECT 587.400 682.350 588.600 683.100 ;
        RECT 595.950 682.950 598.050 685.050 ;
        RECT 602.400 684.450 603.600 684.600 ;
        RECT 599.400 683.400 603.600 684.450 ;
        RECT 580.950 679.950 583.050 682.050 ;
        RECT 583.950 679.950 586.050 682.050 ;
        RECT 586.950 679.950 589.050 682.050 ;
        RECT 584.400 677.400 585.600 679.650 ;
        RECT 596.400 678.900 597.450 682.950 ;
        RECT 584.400 670.050 585.450 677.400 ;
        RECT 595.950 676.800 598.050 678.900 ;
        RECT 568.950 667.950 571.050 670.050 ;
        RECT 574.950 667.950 577.050 670.050 ;
        RECT 583.950 667.950 586.050 670.050 ;
        RECT 560.400 644.400 564.450 645.450 ;
        RECT 565.950 643.800 568.050 645.900 ;
        RECT 548.100 638.400 550.200 640.500 ;
        RECT 557.100 638.700 559.200 640.800 ;
        RECT 526.950 619.950 529.050 622.050 ;
        RECT 535.800 619.950 537.900 622.050 ;
        RECT 538.950 619.950 541.050 622.050 ;
        RECT 553.950 619.950 556.050 622.050 ;
        RECT 569.400 621.450 570.450 667.950 ;
        RECT 574.950 661.950 577.050 664.050 ;
        RECT 575.400 652.200 576.450 661.950 ;
        RECT 580.950 655.950 583.050 658.050 ;
        RECT 574.950 650.100 577.050 652.200 ;
        RECT 581.400 651.600 582.450 655.950 ;
        RECT 575.400 649.350 576.600 650.100 ;
        RECT 581.400 649.350 582.600 651.600 ;
        RECT 586.950 650.100 589.050 652.200 ;
        RECT 587.400 649.350 588.600 650.100 ;
        RECT 574.950 646.950 577.050 649.050 ;
        RECT 577.950 646.950 580.050 649.050 ;
        RECT 580.950 646.950 583.050 649.050 ;
        RECT 583.950 646.950 586.050 649.050 ;
        RECT 586.950 646.950 589.050 649.050 ;
        RECT 578.400 645.900 579.600 646.650 ;
        RECT 577.950 643.800 580.050 645.900 ;
        RECT 584.400 645.000 585.600 646.650 ;
        RECT 583.950 640.950 586.050 645.000 ;
        RECT 599.400 643.050 600.450 683.400 ;
        RECT 602.400 682.350 603.600 683.400 ;
        RECT 611.400 684.450 612.600 684.600 ;
        RECT 611.400 683.400 615.450 684.450 ;
        RECT 611.400 682.350 612.600 683.400 ;
        RECT 602.100 679.950 604.200 682.050 ;
        RECT 605.400 679.950 607.500 682.050 ;
        RECT 610.800 679.950 612.900 682.050 ;
        RECT 605.400 678.900 606.600 679.650 ;
        RECT 604.950 676.800 607.050 678.900 ;
        RECT 607.950 655.950 610.050 658.050 ;
        RECT 608.400 651.600 609.450 655.950 ;
        RECT 608.400 649.350 609.600 651.600 ;
        RECT 604.950 646.950 607.050 649.050 ;
        RECT 607.950 646.950 610.050 649.050 ;
        RECT 605.400 645.900 606.600 646.650 ;
        RECT 614.400 646.050 615.450 683.400 ;
        RECT 616.950 683.100 619.050 685.200 ;
        RECT 620.400 651.450 621.450 691.950 ;
        RECT 623.400 678.450 624.450 722.400 ;
        RECT 628.950 721.800 631.050 723.900 ;
        RECT 635.400 694.050 636.450 745.950 ;
        RECT 637.950 742.950 640.050 745.050 ;
        RECT 646.950 742.950 649.050 745.050 ;
        RECT 656.400 744.450 657.450 761.100 ;
        RECT 665.400 760.350 666.600 761.100 ;
        RECT 671.400 760.350 672.600 762.000 ;
        RECT 676.950 761.100 679.050 766.050 ;
        RECT 685.950 761.100 688.050 763.200 ;
        RECT 691.950 761.100 694.050 763.200 ;
        RECT 712.950 761.100 715.050 763.200 ;
        RECT 661.950 757.950 664.050 760.050 ;
        RECT 664.950 757.950 667.050 760.050 ;
        RECT 667.950 757.950 670.050 760.050 ;
        RECT 670.950 757.950 673.050 760.050 ;
        RECT 662.400 755.400 663.600 757.650 ;
        RECT 668.400 755.400 669.600 757.650 ;
        RECT 662.400 751.050 663.450 755.400 ;
        RECT 661.950 748.950 664.050 751.050 ;
        RECT 658.950 744.450 661.050 745.050 ;
        RECT 656.400 743.400 661.050 744.450 ;
        RECT 658.950 742.950 661.050 743.400 ;
        RECT 634.950 691.950 637.050 694.050 ;
        RECT 638.400 688.050 639.450 742.950 ;
        RECT 643.950 739.950 646.050 742.050 ;
        RECT 640.950 736.950 643.050 739.050 ;
        RECT 641.400 730.050 642.450 736.950 ;
        RECT 640.950 727.950 643.050 730.050 ;
        RECT 644.400 729.600 645.450 739.950 ;
        RECT 647.400 732.450 648.450 742.950 ;
        RECT 649.950 732.450 652.050 736.050 ;
        RECT 647.400 732.000 652.050 732.450 ;
        RECT 647.400 731.400 651.450 732.000 ;
        RECT 650.400 729.600 651.450 731.400 ;
        RECT 659.400 730.050 660.450 742.950 ;
        RECT 668.400 736.050 669.450 755.400 ;
        RECT 677.400 739.050 678.450 761.100 ;
        RECT 686.400 760.350 687.600 761.100 ;
        RECT 692.400 760.350 693.600 761.100 ;
        RECT 713.400 760.350 714.600 761.100 ;
        RECT 724.950 760.950 727.050 763.050 ;
        RECT 733.950 761.100 736.050 766.050 ;
        RECT 739.950 761.100 742.050 763.200 ;
        RECT 685.950 757.950 688.050 760.050 ;
        RECT 688.950 757.950 691.050 760.050 ;
        RECT 691.950 757.950 694.050 760.050 ;
        RECT 694.950 757.950 697.050 760.050 ;
        RECT 709.950 757.950 712.050 760.050 ;
        RECT 712.950 757.950 715.050 760.050 ;
        RECT 682.950 754.950 685.050 757.050 ;
        RECT 689.400 755.400 690.600 757.650 ;
        RECT 695.400 755.400 696.600 757.650 ;
        RECT 710.400 755.400 711.600 757.650 ;
        RECT 683.400 748.050 684.450 754.950 ;
        RECT 685.950 748.950 688.050 751.050 ;
        RECT 682.950 745.950 685.050 748.050 ;
        RECT 673.950 737.400 678.450 739.050 ;
        RECT 673.950 736.950 678.000 737.400 ;
        RECT 667.950 735.450 670.050 736.050 ;
        RECT 667.950 734.400 672.450 735.450 ;
        RECT 667.950 733.950 670.050 734.400 ;
        RECT 671.400 733.050 672.450 734.400 ;
        RECT 676.950 733.950 679.050 736.050 ;
        RECT 682.950 733.950 685.050 736.050 ;
        RECT 671.400 731.400 676.050 733.050 ;
        RECT 672.000 730.950 676.050 731.400 ;
        RECT 644.400 727.350 645.600 729.600 ;
        RECT 650.400 727.350 651.600 729.600 ;
        RECT 658.950 727.950 661.050 730.050 ;
        RECT 670.950 728.100 673.050 730.200 ;
        RECT 677.400 729.600 678.450 733.950 ;
        RECT 643.950 724.950 646.050 727.050 ;
        RECT 646.950 724.950 649.050 727.050 ;
        RECT 649.950 724.950 652.050 727.050 ;
        RECT 652.950 724.950 655.050 727.050 ;
        RECT 647.400 723.900 648.600 724.650 ;
        RECT 653.400 723.900 654.600 724.650 ;
        RECT 659.400 723.900 660.450 727.950 ;
        RECT 671.400 727.350 672.600 728.100 ;
        RECT 677.400 727.350 678.600 729.600 ;
        RECT 667.950 724.950 670.050 727.050 ;
        RECT 670.950 724.950 673.050 727.050 ;
        RECT 673.950 724.950 676.050 727.050 ;
        RECT 676.950 724.950 679.050 727.050 ;
        RECT 646.950 721.800 649.050 723.900 ;
        RECT 652.950 721.800 655.050 723.900 ;
        RECT 658.950 721.800 661.050 723.900 ;
        RECT 668.400 722.400 669.600 724.650 ;
        RECT 674.400 723.000 675.600 724.650 ;
        RECT 643.950 706.950 646.050 709.050 ;
        RECT 631.950 683.100 634.050 685.200 ;
        RECT 637.950 684.000 640.050 688.050 ;
        RECT 632.400 682.350 633.600 683.100 ;
        RECT 638.400 682.350 639.600 684.000 ;
        RECT 628.950 679.950 631.050 682.050 ;
        RECT 631.950 679.950 634.050 682.050 ;
        RECT 634.950 679.950 637.050 682.050 ;
        RECT 637.950 679.950 640.050 682.050 ;
        RECT 629.400 678.450 630.600 679.650 ;
        RECT 623.400 677.400 630.600 678.450 ;
        RECT 635.400 677.400 636.600 679.650 ;
        RECT 644.400 679.050 645.450 706.950 ;
        RECT 668.400 700.050 669.450 722.400 ;
        RECT 673.950 718.950 676.050 723.000 ;
        RECT 679.950 721.950 682.050 724.050 ;
        RECT 680.400 718.050 681.450 721.950 ;
        RECT 683.400 721.050 684.450 733.950 ;
        RECT 686.400 721.050 687.450 748.950 ;
        RECT 689.400 745.050 690.450 755.400 ;
        RECT 688.950 742.950 691.050 745.050 ;
        RECT 695.400 736.050 696.450 755.400 ;
        RECT 700.950 748.950 703.050 751.050 ;
        RECT 688.950 733.950 691.050 736.050 ;
        RECT 694.950 733.950 697.050 736.050 ;
        RECT 689.400 730.050 690.450 733.950 ;
        RECT 688.950 727.950 691.050 730.050 ;
        RECT 694.950 728.100 697.050 730.200 ;
        RECT 701.400 729.600 702.450 748.950 ;
        RECT 710.400 745.050 711.450 755.400 ;
        RECT 721.950 751.950 724.050 754.050 ;
        RECT 715.950 748.950 721.050 751.050 ;
        RECT 703.950 742.950 706.050 745.050 ;
        RECT 709.950 742.950 712.050 745.050 ;
        RECT 704.400 733.050 705.450 742.950 ;
        RECT 703.950 730.950 706.050 733.050 ;
        RECT 695.400 727.350 696.600 728.100 ;
        RECT 701.400 727.350 702.600 729.600 ;
        RECT 715.950 728.100 718.050 730.200 ;
        RECT 722.400 729.600 723.450 751.950 ;
        RECT 725.400 751.050 726.450 760.950 ;
        RECT 734.400 760.350 735.600 761.100 ;
        RECT 740.400 760.350 741.600 761.100 ;
        RECT 748.950 760.950 751.050 763.050 ;
        RECT 754.950 762.000 757.050 766.050 ;
        RECT 730.950 757.950 733.050 760.050 ;
        RECT 733.950 757.950 736.050 760.050 ;
        RECT 736.950 757.950 739.050 760.050 ;
        RECT 739.950 757.950 742.050 760.050 ;
        RECT 731.400 755.400 732.600 757.650 ;
        RECT 737.400 756.000 738.600 757.650 ;
        RECT 749.400 756.900 750.450 760.950 ;
        RECT 755.400 760.350 756.600 762.000 ;
        RECT 760.950 761.100 763.050 763.200 ;
        RECT 761.400 760.350 762.600 761.100 ;
        RECT 754.950 757.950 757.050 760.050 ;
        RECT 757.950 757.950 760.050 760.050 ;
        RECT 760.950 757.950 763.050 760.050 ;
        RECT 763.950 757.950 766.050 760.050 ;
        RECT 758.400 756.900 759.600 757.650 ;
        RECT 731.400 753.450 732.450 755.400 ;
        RECT 736.950 753.450 739.050 756.000 ;
        RECT 748.950 754.800 751.050 756.900 ;
        RECT 757.950 754.800 760.050 756.900 ;
        RECT 764.400 755.400 765.600 757.650 ;
        RECT 728.400 753.000 732.450 753.450 ;
        RECT 727.950 752.400 732.450 753.000 ;
        RECT 734.400 752.400 739.050 753.450 ;
        RECT 724.950 748.950 727.050 751.050 ;
        RECT 727.950 748.950 730.050 752.400 ;
        RECT 730.950 748.950 733.050 751.050 ;
        RECT 724.950 736.950 727.050 739.050 ;
        RECT 725.400 733.050 726.450 736.950 ;
        RECT 724.950 730.950 727.050 733.050 ;
        RECT 716.400 727.350 717.600 728.100 ;
        RECT 722.400 727.350 723.600 729.600 ;
        RECT 691.950 724.950 694.050 727.050 ;
        RECT 694.950 724.950 697.050 727.050 ;
        RECT 697.950 724.950 700.050 727.050 ;
        RECT 700.950 724.950 703.050 727.050 ;
        RECT 715.950 724.950 718.050 727.050 ;
        RECT 718.950 724.950 721.050 727.050 ;
        RECT 721.950 724.950 724.050 727.050 ;
        RECT 724.950 724.950 727.050 727.050 ;
        RECT 688.950 721.950 691.050 724.050 ;
        RECT 692.400 722.400 693.600 724.650 ;
        RECT 698.400 723.000 699.600 724.650 ;
        RECT 682.950 718.950 685.050 721.050 ;
        RECT 685.950 718.950 688.050 721.050 ;
        RECT 679.950 715.950 682.050 718.050 ;
        RECT 655.950 697.950 658.050 700.050 ;
        RECT 667.950 697.950 670.050 700.050 ;
        RECT 656.400 684.600 657.450 697.950 ;
        RECT 679.950 694.950 682.050 697.050 ;
        RECT 661.950 691.950 664.050 694.050 ;
        RECT 662.400 684.600 663.450 691.950 ;
        RECT 680.400 688.050 681.450 694.950 ;
        RECT 685.950 688.950 688.050 691.050 ;
        RECT 667.950 685.950 670.050 688.050 ;
        RECT 656.400 682.350 657.600 684.600 ;
        RECT 662.400 682.350 663.600 684.600 ;
        RECT 668.400 682.050 669.450 685.950 ;
        RECT 679.950 684.000 682.050 688.050 ;
        RECT 686.400 684.600 687.450 688.950 ;
        RECT 680.400 682.350 681.600 684.000 ;
        RECT 686.400 682.350 687.600 684.600 ;
        RECT 689.400 684.450 690.450 721.950 ;
        RECT 692.400 688.050 693.450 722.400 ;
        RECT 697.950 718.950 700.050 723.000 ;
        RECT 712.950 721.950 715.050 724.050 ;
        RECT 719.400 723.900 720.600 724.650 ;
        RECT 725.400 723.900 726.600 724.650 ;
        RECT 731.400 723.900 732.450 748.950 ;
        RECT 698.400 697.050 699.450 718.950 ;
        RECT 697.950 694.950 700.050 697.050 ;
        RECT 713.400 691.050 714.450 721.950 ;
        RECT 718.950 721.800 721.050 723.900 ;
        RECT 724.950 721.800 727.050 723.900 ;
        RECT 730.950 721.800 733.050 723.900 ;
        RECT 721.950 694.950 724.050 697.050 ;
        RECT 712.950 688.950 715.050 691.050 ;
        RECT 691.950 685.950 694.050 688.050 ;
        RECT 689.400 683.400 693.450 684.450 ;
        RECT 706.950 684.000 709.050 688.050 ;
        RECT 713.400 684.600 714.450 688.950 ;
        RECT 652.950 679.950 655.050 682.050 ;
        RECT 655.950 679.950 658.050 682.050 ;
        RECT 658.950 679.950 661.050 682.050 ;
        RECT 661.950 679.950 664.050 682.050 ;
        RECT 667.950 679.950 670.050 682.050 ;
        RECT 676.950 679.950 679.050 682.050 ;
        RECT 679.950 679.950 682.050 682.050 ;
        RECT 682.950 679.950 685.050 682.050 ;
        RECT 685.950 679.950 688.050 682.050 ;
        RECT 625.950 661.950 628.050 664.050 ;
        RECT 617.400 650.400 621.450 651.450 ;
        RECT 626.400 651.600 627.450 661.950 ;
        RECT 604.950 643.800 607.050 645.900 ;
        RECT 613.950 643.950 616.050 646.050 ;
        RECT 598.950 640.950 601.050 643.050 ;
        RECT 569.400 620.400 573.450 621.450 ;
        RECT 523.950 616.950 526.050 619.050 ;
        RECT 520.950 610.950 523.050 613.050 ;
        RECT 493.950 605.100 496.050 607.200 ;
        RECT 511.950 606.000 514.050 610.050 ;
        RECT 517.950 606.450 520.050 607.200 ;
        RECT 521.400 606.450 522.450 610.950 ;
        RECT 494.400 604.350 495.600 605.100 ;
        RECT 512.400 604.350 513.600 606.000 ;
        RECT 517.950 605.400 522.450 606.450 ;
        RECT 517.950 605.100 520.050 605.400 ;
        RECT 518.400 604.350 519.600 605.100 ;
        RECT 469.950 601.950 472.050 604.050 ;
        RECT 472.950 601.950 475.050 604.050 ;
        RECT 475.950 601.950 478.050 604.050 ;
        RECT 490.950 601.950 493.050 604.050 ;
        RECT 493.950 601.950 496.050 604.050 ;
        RECT 508.950 601.950 511.050 604.050 ;
        RECT 511.950 601.950 514.050 604.050 ;
        RECT 514.950 601.950 517.050 604.050 ;
        RECT 517.950 601.950 520.050 604.050 ;
        RECT 449.400 592.050 450.450 599.400 ;
        RECT 454.950 598.800 457.050 600.900 ;
        RECT 457.950 597.450 460.050 601.050 ;
        RECT 460.950 598.950 463.050 601.050 ;
        RECT 473.400 599.400 474.600 601.650 ;
        RECT 491.400 599.400 492.600 601.650 ;
        RECT 509.400 600.000 510.600 601.650 ;
        RECT 515.400 600.900 516.600 601.650 ;
        RECT 524.400 601.050 525.450 616.950 ;
        RECT 455.400 597.000 460.050 597.450 ;
        RECT 455.400 596.400 459.450 597.000 ;
        RECT 448.950 589.950 451.050 592.050 ;
        RECT 445.950 583.950 448.050 586.050 ;
        RECT 446.400 574.200 447.450 583.950 ;
        RECT 445.950 572.100 448.050 574.200 ;
        RECT 455.400 573.600 456.450 596.400 ;
        RECT 473.400 592.050 474.450 599.400 ;
        RECT 481.950 595.950 484.050 598.050 ;
        RECT 472.950 589.950 475.050 592.050 ;
        RECT 425.100 568.950 427.200 571.050 ;
        RECT 430.500 568.950 432.600 571.050 ;
        RECT 433.800 568.950 435.900 571.050 ;
        RECT 434.400 567.900 435.600 568.650 ;
        RECT 433.950 565.800 436.050 567.900 ;
        RECT 418.950 559.950 421.050 562.050 ;
        RECT 434.400 559.050 435.450 565.800 ;
        RECT 433.950 556.950 436.050 559.050 ;
        RECT 421.950 550.950 424.050 553.050 ;
        RECT 403.950 547.950 406.050 550.050 ;
        RECT 388.950 544.950 391.050 547.050 ;
        RECT 385.950 541.950 388.050 544.050 ;
        RECT 322.950 527.100 325.050 529.200 ;
        RECT 329.400 528.450 330.600 528.600 ;
        RECT 334.950 528.450 337.050 529.200 ;
        RECT 329.400 527.400 337.050 528.450 ;
        RECT 323.400 526.350 324.600 527.100 ;
        RECT 329.400 526.350 330.600 527.400 ;
        RECT 334.950 527.100 337.050 527.400 ;
        RECT 343.950 527.100 346.050 529.200 ;
        RECT 349.950 527.100 352.050 529.200 ;
        RECT 355.950 527.100 358.050 529.200 ;
        RECT 364.950 527.100 367.050 532.050 ;
        RECT 370.950 527.100 373.050 529.200 ;
        RECT 379.800 527.100 381.900 529.200 ;
        RECT 382.950 527.100 385.050 529.200 ;
        RECT 388.950 527.100 391.050 529.200 ;
        RECT 394.950 528.000 397.050 532.050 ;
        RECT 322.950 523.950 325.050 526.050 ;
        RECT 325.950 523.950 328.050 526.050 ;
        RECT 328.950 523.950 331.050 526.050 ;
        RECT 281.400 505.050 282.450 521.400 ;
        RECT 298.950 517.950 301.050 522.000 ;
        RECT 304.950 520.800 307.050 522.900 ;
        RECT 310.950 520.800 313.050 522.900 ;
        RECT 326.400 521.400 327.600 523.650 ;
        RECT 301.950 511.950 304.050 514.050 ;
        RECT 268.950 502.950 271.050 505.050 ;
        RECT 280.950 502.950 283.050 505.050 ;
        RECT 236.400 493.350 237.600 494.100 ;
        RECT 244.950 493.950 247.050 496.050 ;
        RECT 250.950 493.950 253.050 496.050 ;
        RECT 232.950 490.950 235.050 493.050 ;
        RECT 235.950 490.950 238.050 493.050 ;
        RECT 238.950 490.950 241.050 493.050 ;
        RECT 245.400 484.050 246.450 493.950 ;
        RECT 244.950 481.950 247.050 484.050 ;
        RECT 224.400 458.400 228.450 459.450 ;
        RECT 202.950 454.950 205.050 457.050 ;
        RECT 211.950 454.950 214.050 457.050 ;
        RECT 203.400 450.600 204.450 454.950 ;
        RECT 203.400 448.350 204.600 450.600 ;
        RECT 178.950 445.950 181.050 448.050 ;
        RECT 181.950 445.950 184.050 448.050 ;
        RECT 184.950 445.950 187.050 448.050 ;
        RECT 199.950 445.950 202.050 448.050 ;
        RECT 202.950 445.950 205.050 448.050 ;
        RECT 182.400 444.000 183.600 445.650 ;
        RECT 181.950 439.950 184.050 444.000 ;
        RECT 157.950 436.950 160.050 439.050 ;
        RECT 169.950 436.950 172.050 439.050 ;
        RECT 149.400 415.350 150.600 417.600 ;
        RECT 212.400 417.450 213.450 454.950 ;
        RECT 224.400 450.600 225.450 458.400 ;
        RECT 224.400 448.350 225.600 450.600 ;
        RECT 251.400 450.450 252.450 493.950 ;
        RECT 254.400 490.950 256.500 493.050 ;
        RECT 259.800 490.950 261.900 493.050 ;
        RECT 260.400 488.400 261.600 490.650 ;
        RECT 269.400 490.050 270.450 502.950 ;
        RECT 274.950 494.100 277.050 496.200 ;
        RECT 280.950 494.100 283.050 496.200 ;
        RECT 302.400 495.600 303.450 511.950 ;
        RECT 326.400 511.050 327.450 521.400 ;
        RECT 335.400 520.050 336.450 527.100 ;
        RECT 344.400 526.350 345.600 527.100 ;
        RECT 350.400 526.350 351.600 527.100 ;
        RECT 343.950 523.950 346.050 526.050 ;
        RECT 346.950 523.950 349.050 526.050 ;
        RECT 349.950 523.950 352.050 526.050 ;
        RECT 347.400 521.400 348.600 523.650 ;
        RECT 334.950 517.950 337.050 520.050 ;
        RECT 347.400 517.050 348.450 521.400 ;
        RECT 349.950 517.950 352.050 520.050 ;
        RECT 346.950 514.950 349.050 517.050 ;
        RECT 325.950 508.950 328.050 511.050 ;
        RECT 334.950 505.950 337.050 508.050 ;
        RECT 275.400 493.350 276.600 494.100 ;
        RECT 281.400 493.350 282.600 494.100 ;
        RECT 302.400 493.350 303.600 495.600 ;
        RECT 322.950 495.000 325.050 499.050 ;
        RECT 331.950 496.950 334.050 499.050 ;
        RECT 323.400 493.350 324.600 495.000 ;
        RECT 274.950 490.950 277.050 493.050 ;
        RECT 277.950 490.950 280.050 493.050 ;
        RECT 280.950 490.950 283.050 493.050 ;
        RECT 283.950 490.950 286.050 493.050 ;
        RECT 298.950 490.950 301.050 493.050 ;
        RECT 301.950 490.950 304.050 493.050 ;
        RECT 304.950 490.950 307.050 493.050 ;
        RECT 310.950 490.950 313.050 493.050 ;
        RECT 319.950 490.950 322.050 493.050 ;
        RECT 322.950 490.950 325.050 493.050 ;
        RECT 260.400 460.050 261.450 488.400 ;
        RECT 268.950 487.950 271.050 490.050 ;
        RECT 278.400 489.900 279.600 490.650 ;
        RECT 277.950 487.800 280.050 489.900 ;
        RECT 284.400 488.400 285.600 490.650 ;
        RECT 299.400 488.400 300.600 490.650 ;
        RECT 305.400 489.900 306.600 490.650 ;
        RECT 278.400 478.050 279.450 487.800 ;
        RECT 284.400 484.050 285.450 488.400 ;
        RECT 299.400 484.050 300.450 488.400 ;
        RECT 304.950 487.800 307.050 489.900 ;
        RECT 283.950 481.950 286.050 484.050 ;
        RECT 298.950 481.950 301.050 484.050 ;
        RECT 277.950 475.950 280.050 478.050 ;
        RECT 301.950 469.950 304.050 472.050 ;
        RECT 286.950 460.950 289.050 463.050 ;
        RECT 259.950 457.950 262.050 460.050 ;
        RECT 268.950 457.950 271.050 460.050 ;
        RECT 269.400 454.050 270.450 457.950 ;
        RECT 268.950 451.950 271.050 454.050 ;
        RECT 280.950 451.950 283.050 454.050 ;
        RECT 269.400 450.600 270.450 451.950 ;
        RECT 251.400 449.400 255.450 450.450 ;
        RECT 217.950 445.950 220.050 448.050 ;
        RECT 220.950 445.950 223.050 448.050 ;
        RECT 223.950 445.950 226.050 448.050 ;
        RECT 226.950 445.950 229.050 448.050 ;
        RECT 229.950 445.950 232.050 448.050 ;
        RECT 244.950 445.950 247.050 448.050 ;
        RECT 247.950 445.950 250.050 448.050 ;
        RECT 245.400 444.900 246.600 445.650 ;
        RECT 254.400 444.900 255.450 449.400 ;
        RECT 269.400 448.350 270.600 450.600 ;
        RECT 262.950 445.950 265.050 448.050 ;
        RECT 265.950 445.950 268.050 448.050 ;
        RECT 268.950 445.950 271.050 448.050 ;
        RECT 244.950 442.800 247.050 444.900 ;
        RECT 253.950 442.800 256.050 444.900 ;
        RECT 266.400 443.400 267.600 445.650 ;
        RECT 254.400 418.200 255.450 442.800 ;
        RECT 266.400 424.050 267.450 443.400 ;
        RECT 268.950 424.950 271.050 427.050 ;
        RECT 265.950 421.950 268.050 424.050 ;
        RECT 212.400 416.400 216.450 417.450 ;
        RECT 148.950 412.950 151.050 415.050 ;
        RECT 151.950 412.950 154.050 415.050 ;
        RECT 170.100 412.950 172.200 415.050 ;
        RECT 188.100 412.950 190.200 415.050 ;
        RECT 205.950 412.950 208.050 415.050 ;
        RECT 208.950 412.950 211.050 415.050 ;
        RECT 124.650 402.600 126.750 403.500 ;
        RECT 109.350 399.600 111.450 401.700 ;
        RECT 131.400 394.050 132.450 410.400 ;
        RECT 142.950 409.950 145.050 412.050 ;
        RECT 152.400 411.900 153.600 412.650 ;
        RECT 151.950 409.800 154.050 411.900 ;
        RECT 170.400 410.400 171.600 412.650 ;
        RECT 206.400 410.400 207.600 412.650 ;
        RECT 170.400 403.050 171.450 410.400 ;
        RECT 145.950 400.950 148.050 403.050 ;
        RECT 169.950 400.950 172.050 403.050 ;
        RECT 88.950 391.950 91.050 394.050 ;
        RECT 130.950 391.950 133.050 394.050 ;
        RECT 82.650 379.500 84.750 380.400 ;
        RECT 76.950 376.950 79.050 379.050 ;
        RECT 82.650 378.300 86.850 379.500 ;
        RECT 89.400 379.050 90.450 391.950 ;
        RECT 67.350 372.600 69.450 374.700 ;
        RECT 53.400 370.350 54.600 372.600 ;
        RECT 52.950 367.950 55.050 370.050 ;
        RECT 61.950 367.950 64.050 370.050 ;
        RECT 62.400 366.900 63.600 367.650 ;
        RECT 61.950 364.800 64.050 366.900 ;
        RECT 68.250 359.700 69.450 372.600 ;
        RECT 79.950 371.100 82.050 373.200 ;
        RECT 80.400 370.350 81.600 371.100 ;
        RECT 79.800 367.950 81.900 370.050 ;
        RECT 85.650 359.700 86.850 378.300 ;
        RECT 88.950 376.950 91.050 379.050 ;
        RECT 89.400 372.600 90.450 376.950 ;
        RECT 89.400 370.350 90.600 372.600 ;
        RECT 94.950 371.100 97.050 373.200 ;
        RECT 121.950 371.100 124.050 373.200 ;
        RECT 130.950 371.100 133.050 373.200 ;
        RECT 136.950 371.100 139.050 373.200 ;
        RECT 88.950 367.950 91.050 370.050 ;
        RECT 31.350 357.600 33.450 359.700 ;
        RECT 49.050 357.600 51.150 359.700 ;
        RECT 67.350 357.600 69.450 359.700 ;
        RECT 85.050 357.600 87.150 359.700 ;
        RECT 95.400 355.050 96.450 371.100 ;
        RECT 106.950 367.950 109.050 370.050 ;
        RECT 109.950 367.950 112.050 370.050 ;
        RECT 112.950 367.950 115.050 370.050 ;
        RECT 110.400 366.900 111.600 367.650 ;
        RECT 122.400 367.050 123.450 371.100 ;
        RECT 131.400 370.350 132.600 371.100 ;
        RECT 137.400 370.350 138.600 371.100 ;
        RECT 127.950 367.950 130.050 370.050 ;
        RECT 130.950 367.950 133.050 370.050 ;
        RECT 133.950 367.950 136.050 370.050 ;
        RECT 136.950 367.950 139.050 370.050 ;
        RECT 139.950 367.950 142.050 370.050 ;
        RECT 109.950 364.800 112.050 366.900 ;
        RECT 121.950 364.950 124.050 367.050 ;
        RECT 128.400 365.400 129.600 367.650 ;
        RECT 134.400 365.400 135.600 367.650 ;
        RECT 140.400 366.900 141.600 367.650 ;
        RECT 94.950 352.950 97.050 355.050 ;
        RECT 55.350 345.300 57.450 347.400 ;
        RECT 73.050 345.300 75.150 347.400 ;
        RECT 97.950 346.950 100.050 349.050 ;
        RECT 22.950 339.000 25.050 343.050 ;
        RECT 23.400 337.350 24.600 339.000 ;
        RECT 43.950 338.100 46.050 340.200 ;
        RECT 49.950 338.100 52.050 340.200 ;
        RECT 44.400 337.350 45.600 338.100 ;
        RECT 50.400 337.350 51.600 338.100 ;
        RECT 17.100 334.950 19.200 337.050 ;
        RECT 22.500 334.950 24.600 337.050 ;
        RECT 38.100 334.950 40.200 337.050 ;
        RECT 43.500 334.950 45.600 337.050 ;
        RECT 49.950 334.950 52.050 337.050 ;
        RECT 56.250 332.400 57.450 345.300 ;
        RECT 67.800 334.950 69.900 337.050 ;
        RECT 55.350 330.300 57.450 332.400 ;
        RECT 68.400 332.400 69.600 334.650 ;
        RECT 68.400 330.450 69.450 332.400 ;
        RECT 56.250 323.700 57.450 330.300 ;
        RECT 55.350 321.600 57.450 323.700 ;
        RECT 65.400 329.400 69.450 330.450 ;
        RECT 65.400 309.450 66.450 329.400 ;
        RECT 73.650 326.700 74.850 345.300 ;
        RECT 98.400 339.600 99.450 346.950 ;
        RECT 109.350 345.300 111.450 347.400 ;
        RECT 112.950 346.950 115.050 349.050 ;
        RECT 98.400 337.350 99.600 339.600 ;
        RECT 103.950 339.000 106.050 343.050 ;
        RECT 104.400 337.350 105.600 339.000 ;
        RECT 76.950 334.950 79.050 337.050 ;
        RECT 94.950 334.950 97.050 337.050 ;
        RECT 97.950 334.950 100.050 337.050 ;
        RECT 103.950 334.950 106.050 337.050 ;
        RECT 77.400 333.000 78.600 334.650 ;
        RECT 76.950 328.950 79.050 333.000 ;
        RECT 95.400 332.400 96.600 334.650 ;
        RECT 110.250 332.400 111.450 345.300 ;
        RECT 85.950 328.950 88.050 331.050 ;
        RECT 70.650 325.500 74.850 326.700 ;
        RECT 70.650 324.600 72.750 325.500 ;
        RECT 65.400 308.400 69.450 309.450 ;
        RECT 10.950 304.950 13.050 307.050 ;
        RECT 46.950 304.950 49.050 307.050 ;
        RECT 11.400 288.450 12.450 304.950 ;
        RECT 16.800 298.500 18.900 300.600 ;
        RECT 14.100 289.950 16.200 292.050 ;
        RECT 17.100 291.300 18.300 298.500 ;
        RECT 20.400 295.350 21.600 297.600 ;
        RECT 26.400 297.300 28.500 299.400 ;
        RECT 20.100 292.950 22.200 295.050 ;
        RECT 23.100 293.700 25.200 295.800 ;
        RECT 23.100 291.300 24.000 293.700 ;
        RECT 17.100 290.100 24.000 291.300 ;
        RECT 14.400 288.450 15.600 289.650 ;
        RECT 11.400 287.400 15.600 288.450 ;
        RECT 17.100 284.700 18.000 290.100 ;
        RECT 18.900 288.300 21.000 289.200 ;
        RECT 26.700 288.300 27.600 297.300 ;
        RECT 28.950 293.100 31.050 295.200 ;
        RECT 47.400 294.600 48.450 304.950 ;
        RECT 64.350 303.300 66.450 305.400 ;
        RECT 52.950 298.950 55.050 301.050 ;
        RECT 53.400 295.200 54.450 298.950 ;
        RECT 65.250 296.700 66.450 303.300 ;
        RECT 29.400 292.350 30.600 293.100 ;
        RECT 47.400 292.350 48.600 294.600 ;
        RECT 52.950 293.100 55.050 295.200 ;
        RECT 64.350 294.600 66.450 296.700 ;
        RECT 53.400 292.350 54.600 293.100 ;
        RECT 28.800 289.950 30.900 292.050 ;
        RECT 46.950 289.950 49.050 292.050 ;
        RECT 49.950 289.950 52.050 292.050 ;
        RECT 52.950 289.950 55.050 292.050 ;
        RECT 58.950 289.950 61.050 292.050 ;
        RECT 18.900 287.100 27.600 288.300 ;
        RECT 50.400 287.400 51.600 289.650 ;
        RECT 59.400 288.900 60.600 289.650 ;
        RECT 16.800 282.600 18.900 284.700 ;
        RECT 20.100 284.100 22.200 286.200 ;
        RECT 24.000 285.300 26.100 287.100 ;
        RECT 20.400 281.550 21.600 283.800 ;
        RECT 20.400 268.050 21.450 281.550 ;
        RECT 22.950 271.950 25.050 274.050 ;
        RECT 34.950 271.950 37.050 274.050 ;
        RECT 19.950 265.950 22.050 268.050 ;
        RECT 23.400 261.600 24.450 271.950 ;
        RECT 28.950 265.950 31.050 268.050 ;
        RECT 29.400 262.050 30.450 265.950 ;
        RECT 31.950 262.950 34.050 265.050 ;
        RECT 23.400 259.350 24.600 261.600 ;
        RECT 28.950 259.950 31.050 262.050 ;
        RECT 16.950 256.950 19.050 259.050 ;
        RECT 19.950 256.950 22.050 259.050 ;
        RECT 22.950 256.950 25.050 259.050 ;
        RECT 25.950 256.950 28.050 259.050 ;
        RECT 20.400 254.400 21.600 256.650 ;
        RECT 26.400 255.900 27.600 256.650 ;
        RECT 32.400 256.050 33.450 262.950 ;
        RECT 20.400 250.050 21.450 254.400 ;
        RECT 25.950 253.800 28.050 255.900 ;
        RECT 31.950 253.950 34.050 256.050 ;
        RECT 31.950 250.800 34.050 252.900 ;
        RECT 19.950 247.950 22.050 250.050 ;
        RECT 17.100 220.500 19.200 222.600 ;
        RECT 14.100 211.950 16.200 214.050 ;
        RECT 17.100 213.900 18.000 220.500 ;
        RECT 26.100 220.200 28.200 222.300 ;
        RECT 20.400 217.350 21.600 219.600 ;
        RECT 19.800 214.950 21.900 217.050 ;
        RECT 24.000 213.900 26.100 214.200 ;
        RECT 17.100 213.000 26.100 213.900 ;
        RECT 17.100 207.900 18.000 213.000 ;
        RECT 24.000 212.100 26.100 213.000 ;
        RECT 18.900 211.200 21.000 212.100 ;
        RECT 18.900 210.000 26.100 211.200 ;
        RECT 24.000 209.100 26.100 210.000 ;
        RECT 16.500 205.800 18.600 207.900 ;
        RECT 19.800 206.100 21.900 208.200 ;
        RECT 27.000 207.600 27.900 220.200 ;
        RECT 28.950 215.100 31.050 217.200 ;
        RECT 29.400 214.350 30.600 215.100 ;
        RECT 28.800 211.950 30.900 214.050 ;
        RECT 20.400 205.050 21.600 205.800 ;
        RECT 26.400 205.500 28.500 207.600 ;
        RECT 19.950 202.950 22.050 205.050 ;
        RECT 16.950 196.950 19.050 199.050 ;
        RECT 17.400 183.600 18.450 196.950 ;
        RECT 17.400 181.350 18.600 183.600 ;
        RECT 32.400 183.450 33.450 250.800 ;
        RECT 35.400 217.200 36.450 271.950 ;
        RECT 40.950 261.000 43.050 265.050 ;
        RECT 41.400 259.350 42.600 261.000 ;
        RECT 40.950 256.950 43.050 259.050 ;
        RECT 43.950 256.950 46.050 259.050 ;
        RECT 44.400 255.900 45.600 256.650 ;
        RECT 43.950 253.800 46.050 255.900 ;
        RECT 34.800 215.100 36.900 217.200 ;
        RECT 37.950 215.100 40.050 217.200 ;
        RECT 43.950 215.100 46.050 217.200 ;
        RECT 50.400 216.600 51.450 287.400 ;
        RECT 58.950 286.800 61.050 288.900 ;
        RECT 65.250 281.700 66.450 294.600 ;
        RECT 68.400 288.900 69.450 308.400 ;
        RECT 79.650 301.500 81.750 302.400 ;
        RECT 79.650 300.300 83.850 301.500 ;
        RECT 70.950 293.100 73.050 295.200 ;
        RECT 76.950 293.100 79.050 295.200 ;
        RECT 67.950 286.800 70.050 288.900 ;
        RECT 71.400 288.450 72.450 293.100 ;
        RECT 77.400 292.350 78.600 293.100 ;
        RECT 76.800 289.950 78.900 292.050 ;
        RECT 71.400 287.400 75.450 288.450 ;
        RECT 64.350 279.600 66.450 281.700 ;
        RECT 52.950 265.950 55.050 268.050 ;
        RECT 58.950 265.950 61.050 268.050 ;
        RECT 53.400 250.050 54.450 265.950 ;
        RECT 59.400 261.600 60.450 265.950 ;
        RECT 59.400 259.350 60.600 261.600 ;
        RECT 64.950 260.100 67.050 262.200 ;
        RECT 65.400 259.350 66.600 260.100 ;
        RECT 58.950 256.950 61.050 259.050 ;
        RECT 61.950 256.950 64.050 259.050 ;
        RECT 64.950 256.950 67.050 259.050 ;
        RECT 67.950 256.950 70.050 259.050 ;
        RECT 62.400 255.900 63.600 256.650 ;
        RECT 68.400 256.050 69.600 256.650 ;
        RECT 74.400 256.050 75.450 287.400 ;
        RECT 82.650 281.700 83.850 300.300 ;
        RECT 86.400 294.600 87.450 328.950 ;
        RECT 95.400 295.200 96.450 332.400 ;
        RECT 109.350 330.300 111.450 332.400 ;
        RECT 110.250 323.700 111.450 330.300 ;
        RECT 109.350 321.600 111.450 323.700 ;
        RECT 113.400 322.050 114.450 346.950 ;
        RECT 122.400 343.050 123.450 364.950 ;
        RECT 128.400 358.050 129.450 365.400 ;
        RECT 127.950 355.950 130.050 358.050 ;
        RECT 127.050 345.300 129.150 347.400 ;
        RECT 121.950 340.950 124.050 343.050 ;
        RECT 121.800 334.950 123.900 337.050 ;
        RECT 122.400 332.400 123.600 334.650 ;
        RECT 122.400 330.450 123.450 332.400 ;
        RECT 119.400 329.400 123.450 330.450 ;
        RECT 112.950 321.450 115.050 322.050 ;
        RECT 112.950 320.400 117.450 321.450 ;
        RECT 112.950 319.950 115.050 320.400 ;
        RECT 86.400 292.350 87.600 294.600 ;
        RECT 94.950 293.100 97.050 295.200 ;
        RECT 103.950 293.100 106.050 295.200 ;
        RECT 109.950 293.100 112.050 295.200 ;
        RECT 85.950 289.950 88.050 292.050 ;
        RECT 82.050 279.600 84.150 281.700 ;
        RECT 95.400 268.050 96.450 293.100 ;
        RECT 104.400 292.350 105.600 293.100 ;
        RECT 110.400 292.350 111.600 293.100 ;
        RECT 97.950 289.950 100.050 292.050 ;
        RECT 103.950 289.950 106.050 292.050 ;
        RECT 106.950 289.950 109.050 292.050 ;
        RECT 109.950 289.950 112.050 292.050 ;
        RECT 94.950 265.950 97.050 268.050 ;
        RECT 98.400 265.050 99.450 289.950 ;
        RECT 107.400 288.900 108.600 289.650 ;
        RECT 106.950 286.800 109.050 288.900 ;
        RECT 116.400 271.050 117.450 320.400 ;
        RECT 106.950 268.950 109.050 271.050 ;
        RECT 115.950 268.950 118.050 271.050 ;
        RECT 97.950 262.950 100.050 265.050 ;
        RECT 98.400 259.050 99.450 262.950 ;
        RECT 107.400 261.600 108.450 268.950 ;
        RECT 107.400 259.350 108.600 261.600 ;
        RECT 112.950 260.100 115.050 262.200 ;
        RECT 119.400 261.600 120.450 329.400 ;
        RECT 127.650 326.700 128.850 345.300 ;
        RECT 134.400 339.450 135.450 365.400 ;
        RECT 139.950 364.800 142.050 366.900 ;
        RECT 134.400 338.400 138.450 339.450 ;
        RECT 130.950 334.950 133.050 337.050 ;
        RECT 131.400 333.000 132.600 334.650 ;
        RECT 130.950 328.950 133.050 333.000 ;
        RECT 124.650 325.500 128.850 326.700 ;
        RECT 124.650 324.600 126.750 325.500 ;
        RECT 137.400 307.050 138.450 338.400 ;
        RECT 146.400 331.050 147.450 400.950 ;
        RECT 206.400 400.050 207.450 410.400 ;
        RECT 205.950 397.950 208.050 400.050 ;
        RECT 206.400 379.050 207.450 397.950 ;
        RECT 196.950 376.950 199.050 379.050 ;
        RECT 205.950 376.950 208.050 379.050 ;
        RECT 154.950 371.100 157.050 373.200 ;
        RECT 178.950 371.100 181.050 373.200 ;
        RECT 155.400 370.350 156.600 371.100 ;
        RECT 179.400 370.350 180.600 371.100 ;
        RECT 184.800 370.950 186.900 373.050 ;
        RECT 187.950 371.100 190.050 373.200 ;
        RECT 197.400 372.600 198.450 376.950 ;
        RECT 148.950 367.950 151.050 370.050 ;
        RECT 154.950 367.950 157.050 370.050 ;
        RECT 157.950 367.950 160.050 370.050 ;
        RECT 160.950 367.950 163.050 370.050 ;
        RECT 166.950 367.950 169.050 370.050 ;
        RECT 175.950 367.950 178.050 370.050 ;
        RECT 178.950 367.950 181.050 370.050 ;
        RECT 149.400 346.050 150.450 367.950 ;
        RECT 158.400 366.900 159.600 367.650 ;
        RECT 157.950 364.800 160.050 366.900 ;
        RECT 148.950 343.950 151.050 346.050 ;
        RECT 149.400 333.450 150.450 343.950 ;
        RECT 158.400 342.450 159.450 364.800 ;
        RECT 167.400 364.050 168.450 367.950 ;
        RECT 176.400 366.000 177.600 367.650 ;
        RECT 185.400 366.900 186.450 370.950 ;
        RECT 166.950 361.950 169.050 364.050 ;
        RECT 175.950 361.950 178.050 366.000 ;
        RECT 184.950 364.800 187.050 366.900 ;
        RECT 188.400 358.050 189.450 371.100 ;
        RECT 197.400 370.350 198.600 372.600 ;
        RECT 202.950 371.100 205.050 373.200 ;
        RECT 215.400 372.450 216.450 416.400 ;
        RECT 253.950 416.100 256.050 418.200 ;
        RECT 262.950 416.100 265.050 421.050 ;
        RECT 269.400 417.600 270.450 424.950 ;
        RECT 277.950 421.950 280.050 424.050 ;
        RECT 263.400 415.350 264.600 416.100 ;
        RECT 269.400 415.350 270.600 417.600 ;
        RECT 226.800 412.950 228.900 415.050 ;
        RECT 244.800 412.950 246.900 415.050 ;
        RECT 262.950 412.950 265.050 415.050 ;
        RECT 265.950 412.950 268.050 415.050 ;
        RECT 268.950 412.950 271.050 415.050 ;
        RECT 271.950 412.950 274.050 415.050 ;
        RECT 245.400 410.400 246.600 412.650 ;
        RECT 266.400 410.400 267.600 412.650 ;
        RECT 272.400 411.000 273.600 412.650 ;
        RECT 245.400 391.050 246.450 410.400 ;
        RECT 266.400 400.050 267.450 410.400 ;
        RECT 271.950 406.950 274.050 411.000 ;
        RECT 278.400 409.050 279.450 421.950 ;
        RECT 281.400 412.050 282.450 451.950 ;
        RECT 287.400 450.600 288.450 460.950 ;
        RECT 287.400 448.350 288.600 450.600 ;
        RECT 287.100 445.950 289.200 448.050 ;
        RECT 290.400 445.950 292.500 448.050 ;
        RECT 295.800 445.950 297.900 448.050 ;
        RECT 292.950 427.950 295.050 430.050 ;
        RECT 286.950 417.000 289.050 421.050 ;
        RECT 293.400 417.600 294.450 427.950 ;
        RECT 287.400 415.350 288.600 417.000 ;
        RECT 293.400 415.350 294.600 417.600 ;
        RECT 286.950 412.950 289.050 415.050 ;
        RECT 289.950 412.950 292.050 415.050 ;
        RECT 292.950 412.950 295.050 415.050 ;
        RECT 295.950 412.950 298.050 415.050 ;
        RECT 280.950 409.950 283.050 412.050 ;
        RECT 290.400 410.400 291.600 412.650 ;
        RECT 296.400 410.400 297.600 412.650 ;
        RECT 277.950 408.450 280.050 409.050 ;
        RECT 277.950 407.400 282.450 408.450 ;
        RECT 277.950 406.950 280.050 407.400 ;
        RECT 265.950 397.950 268.050 400.050 ;
        RECT 244.950 388.950 247.050 391.050 ;
        RECT 265.950 376.950 268.050 379.050 ;
        RECT 212.400 371.400 216.450 372.450 ;
        RECT 203.400 370.350 204.600 371.100 ;
        RECT 193.950 367.950 196.050 370.050 ;
        RECT 196.950 367.950 199.050 370.050 ;
        RECT 199.950 367.950 202.050 370.050 ;
        RECT 202.950 367.950 205.050 370.050 ;
        RECT 208.950 367.950 211.050 370.050 ;
        RECT 194.400 366.900 195.600 367.650 ;
        RECT 193.950 366.450 196.050 366.900 ;
        RECT 191.400 365.400 196.050 366.450 ;
        RECT 175.950 355.950 178.050 358.050 ;
        RECT 187.950 355.950 190.050 358.050 ;
        RECT 155.400 341.400 159.450 342.450 ;
        RECT 155.400 339.600 156.450 341.400 ;
        RECT 169.950 340.950 172.050 343.050 ;
        RECT 155.400 337.350 156.600 339.600 ;
        RECT 152.100 334.950 154.200 337.050 ;
        RECT 155.400 334.950 157.500 337.050 ;
        RECT 160.800 334.950 162.900 337.050 ;
        RECT 152.400 333.450 153.600 334.650 ;
        RECT 149.400 332.400 153.600 333.450 ;
        RECT 161.400 332.400 162.600 334.650 ;
        RECT 145.950 330.450 148.050 331.050 ;
        RECT 143.400 329.400 148.050 330.450 ;
        RECT 136.950 304.950 139.050 307.050 ;
        RECT 133.950 298.950 136.050 301.050 ;
        RECT 134.400 294.600 135.450 298.950 ;
        RECT 125.400 294.450 126.600 294.600 ;
        RECT 122.400 293.400 126.600 294.450 ;
        RECT 122.400 289.050 123.450 293.400 ;
        RECT 125.400 292.350 126.600 293.400 ;
        RECT 134.400 292.350 135.600 294.600 ;
        RECT 125.100 289.950 127.200 292.050 ;
        RECT 130.500 289.950 132.600 292.050 ;
        RECT 133.800 289.950 135.900 292.050 ;
        RECT 121.950 286.950 124.050 289.050 ;
        RECT 131.400 287.400 132.600 289.650 ;
        RECT 131.400 280.050 132.450 287.400 ;
        RECT 130.950 277.950 133.050 280.050 ;
        RECT 143.400 274.050 144.450 329.400 ;
        RECT 145.950 328.950 148.050 329.400 ;
        RECT 152.400 301.050 153.450 332.400 ;
        RECT 151.950 298.950 154.050 301.050 ;
        RECT 151.950 293.100 154.050 295.200 ;
        RECT 152.400 292.350 153.600 293.100 ;
        RECT 148.950 289.950 151.050 292.050 ;
        RECT 151.950 289.950 154.050 292.050 ;
        RECT 154.950 289.950 157.050 292.050 ;
        RECT 149.400 287.400 150.600 289.650 ;
        RECT 155.400 288.000 156.600 289.650 ;
        RECT 161.400 289.050 162.450 332.400 ;
        RECT 170.400 331.050 171.450 340.950 ;
        RECT 176.400 339.600 177.450 355.950 ;
        RECT 181.950 343.950 184.050 346.050 ;
        RECT 182.400 339.600 183.450 343.950 ;
        RECT 176.400 337.350 177.600 339.600 ;
        RECT 182.400 337.350 183.600 339.600 ;
        RECT 191.400 337.050 192.450 365.400 ;
        RECT 193.950 364.800 196.050 365.400 ;
        RECT 200.400 365.400 201.600 367.650 ;
        RECT 200.400 346.050 201.450 365.400 ;
        RECT 209.400 364.050 210.450 367.950 ;
        RECT 208.950 361.950 211.050 364.050 ;
        RECT 199.950 343.950 202.050 346.050 ;
        RECT 205.950 338.100 208.050 340.200 ;
        RECT 212.400 339.600 213.450 371.400 ;
        RECT 238.950 371.100 241.050 373.200 ;
        RECT 266.400 372.600 267.450 376.950 ;
        RECT 239.400 370.350 240.600 371.100 ;
        RECT 266.400 370.350 267.600 372.600 ;
        RECT 271.950 371.100 274.050 373.200 ;
        RECT 272.400 370.350 273.600 371.100 ;
        RECT 217.950 367.950 220.050 370.050 ;
        RECT 220.950 367.950 223.050 370.050 ;
        RECT 223.950 367.950 226.050 370.050 ;
        RECT 238.950 367.950 241.050 370.050 ;
        RECT 241.950 367.950 244.050 370.050 ;
        RECT 244.950 367.950 247.050 370.050 ;
        RECT 259.950 367.950 262.050 370.050 ;
        RECT 262.950 367.950 265.050 370.050 ;
        RECT 265.950 367.950 268.050 370.050 ;
        RECT 268.950 367.950 271.050 370.050 ;
        RECT 271.950 367.950 274.050 370.050 ;
        RECT 221.400 365.400 222.600 367.650 ;
        RECT 242.400 365.400 243.600 367.650 ;
        RECT 221.400 358.050 222.450 365.400 ;
        RECT 220.950 355.950 223.050 358.050 ;
        RECT 217.800 343.950 219.900 346.050 ;
        RECT 206.400 337.350 207.600 338.100 ;
        RECT 212.400 337.350 213.600 339.600 ;
        RECT 175.950 334.950 178.050 337.050 ;
        RECT 178.950 334.950 181.050 337.050 ;
        RECT 181.950 334.950 184.050 337.050 ;
        RECT 184.950 334.950 187.050 337.050 ;
        RECT 190.950 334.950 193.050 337.050 ;
        RECT 202.950 334.950 205.050 337.050 ;
        RECT 205.950 334.950 208.050 337.050 ;
        RECT 208.950 334.950 211.050 337.050 ;
        RECT 211.950 334.950 214.050 337.050 ;
        RECT 179.400 333.000 180.600 334.650 ;
        RECT 185.400 333.900 186.600 334.650 ;
        RECT 169.950 328.950 172.050 331.050 ;
        RECT 178.950 328.950 181.050 333.000 ;
        RECT 184.950 331.800 187.050 333.900 ;
        RECT 187.950 331.950 190.050 334.050 ;
        RECT 203.400 333.900 204.600 334.650 ;
        RECT 179.400 304.050 180.450 328.950 ;
        RECT 178.950 301.950 181.050 304.050 ;
        RECT 178.950 298.800 181.050 300.900 ;
        RECT 172.950 293.100 175.050 295.200 ;
        RECT 179.400 294.600 180.450 298.800 ;
        RECT 173.400 292.350 174.600 293.100 ;
        RECT 179.400 292.350 180.600 294.600 ;
        RECT 163.950 289.950 166.050 292.050 ;
        RECT 169.950 289.950 172.050 292.050 ;
        RECT 172.950 289.950 175.050 292.050 ;
        RECT 175.950 289.950 178.050 292.050 ;
        RECT 178.950 289.950 181.050 292.050 ;
        RECT 149.400 285.450 150.450 287.400 ;
        RECT 149.400 284.400 153.450 285.450 ;
        RECT 152.400 283.050 153.450 284.400 ;
        RECT 154.950 283.950 157.050 288.000 ;
        RECT 160.950 286.950 163.050 289.050 ;
        RECT 164.400 286.050 165.450 289.950 ;
        RECT 166.950 286.950 169.050 289.050 ;
        RECT 170.400 288.900 171.600 289.650 ;
        RECT 163.950 283.950 166.050 286.050 ;
        RECT 151.950 280.950 154.050 283.050 ;
        RECT 142.950 271.950 145.050 274.050 ;
        RECT 124.350 267.300 126.450 269.400 ;
        RECT 142.050 267.300 144.150 269.400 ;
        RECT 113.400 259.350 114.600 260.100 ;
        RECT 119.400 259.350 120.600 261.600 ;
        RECT 85.950 256.950 88.050 259.050 ;
        RECT 88.950 256.950 91.050 259.050 ;
        RECT 97.950 256.950 100.050 259.050 ;
        RECT 103.950 256.950 106.050 259.050 ;
        RECT 106.950 256.950 109.050 259.050 ;
        RECT 109.950 256.950 112.050 259.050 ;
        RECT 112.950 256.950 115.050 259.050 ;
        RECT 118.950 256.950 121.050 259.050 ;
        RECT 61.950 253.800 64.050 255.900 ;
        RECT 68.400 254.400 73.050 256.050 ;
        RECT 69.000 253.950 73.050 254.400 ;
        RECT 73.950 253.950 76.050 256.050 ;
        RECT 82.950 253.950 85.050 256.050 ;
        RECT 86.400 255.900 87.600 256.650 ;
        RECT 110.400 255.900 111.600 256.650 ;
        RECT 67.950 250.950 70.050 253.050 ;
        RECT 52.950 247.950 55.050 250.050 ;
        RECT 68.400 226.050 69.450 250.950 ;
        RECT 67.950 223.950 70.050 226.050 ;
        RECT 67.800 220.500 69.900 222.600 ;
        RECT 38.400 199.050 39.450 215.100 ;
        RECT 44.400 214.350 45.600 215.100 ;
        RECT 50.400 214.350 51.600 216.600 ;
        RECT 43.950 211.950 46.050 214.050 ;
        RECT 46.950 211.950 49.050 214.050 ;
        RECT 49.950 211.950 52.050 214.050 ;
        RECT 65.100 211.950 67.200 214.050 ;
        RECT 68.100 213.300 69.300 220.500 ;
        RECT 71.400 217.350 72.600 219.600 ;
        RECT 77.400 219.300 79.500 221.400 ;
        RECT 83.400 220.050 84.450 253.950 ;
        RECT 85.950 253.800 88.050 255.900 ;
        RECT 109.950 253.800 112.050 255.900 ;
        RECT 115.950 253.950 118.050 256.050 ;
        RECT 125.250 254.400 126.450 267.300 ;
        RECT 136.800 256.950 138.900 259.050 ;
        RECT 137.400 255.000 138.600 256.650 ;
        RECT 109.950 223.950 112.050 226.050 ;
        RECT 71.100 214.950 73.200 217.050 ;
        RECT 74.100 215.700 76.200 217.800 ;
        RECT 74.100 213.300 75.000 215.700 ;
        RECT 68.100 212.100 75.000 213.300 ;
        RECT 47.400 210.000 48.600 211.650 ;
        RECT 65.400 210.450 66.600 211.650 ;
        RECT 46.950 205.950 49.050 210.000 ;
        RECT 62.400 209.400 66.600 210.450 ;
        RECT 62.400 205.050 63.450 209.400 ;
        RECT 68.100 206.700 69.000 212.100 ;
        RECT 69.900 210.300 72.000 211.200 ;
        RECT 77.700 210.300 78.600 219.300 ;
        RECT 82.950 217.950 85.050 220.050 ;
        RECT 80.400 216.450 81.600 216.600 ;
        RECT 80.400 215.400 84.450 216.450 ;
        RECT 80.400 214.350 81.600 215.400 ;
        RECT 79.800 211.950 81.900 214.050 ;
        RECT 83.400 211.050 84.450 215.400 ;
        RECT 88.950 215.100 91.050 217.200 ;
        RECT 97.950 215.100 100.050 217.200 ;
        RECT 103.950 215.100 106.050 217.200 ;
        RECT 69.900 209.100 78.600 210.300 ;
        RECT 61.950 202.950 64.050 205.050 ;
        RECT 67.800 204.600 69.900 206.700 ;
        RECT 71.100 206.100 73.200 208.200 ;
        RECT 75.000 207.300 77.100 209.100 ;
        RECT 82.950 208.950 85.050 211.050 ;
        RECT 89.400 208.050 90.450 215.100 ;
        RECT 98.400 214.350 99.600 215.100 ;
        RECT 104.400 214.350 105.600 215.100 ;
        RECT 94.950 211.950 97.050 214.050 ;
        RECT 97.950 211.950 100.050 214.050 ;
        RECT 100.950 211.950 103.050 214.050 ;
        RECT 103.950 211.950 106.050 214.050 ;
        RECT 95.400 210.900 96.600 211.650 ;
        RECT 94.950 208.800 97.050 210.900 ;
        RECT 101.400 209.400 102.600 211.650 ;
        RECT 71.400 203.550 72.600 205.800 ;
        RECT 37.950 196.950 40.050 199.050 ;
        RECT 46.950 190.950 49.050 193.050 ;
        RECT 29.400 182.400 33.450 183.450 ;
        RECT 37.950 183.000 40.050 187.050 ;
        RECT 43.950 184.950 46.050 187.050 ;
        RECT 13.950 178.950 16.050 181.050 ;
        RECT 16.950 178.950 19.050 181.050 ;
        RECT 19.950 178.950 22.050 181.050 ;
        RECT 20.400 177.900 21.600 178.650 ;
        RECT 29.400 177.900 30.450 182.400 ;
        RECT 38.400 181.350 39.600 183.000 ;
        RECT 34.950 178.950 37.050 181.050 ;
        RECT 37.950 178.950 40.050 181.050 ;
        RECT 35.400 177.900 36.600 178.650 ;
        RECT 19.950 175.800 22.050 177.900 ;
        RECT 28.950 175.800 31.050 177.900 ;
        RECT 34.950 175.800 37.050 177.900 ;
        RECT 29.400 147.450 30.450 175.800 ;
        RECT 44.400 175.050 45.450 184.950 ;
        RECT 47.400 178.050 48.450 190.950 ;
        RECT 71.400 187.050 72.450 203.550 ;
        RECT 76.950 202.950 79.050 205.050 ;
        RECT 82.950 202.950 85.050 207.900 ;
        RECT 88.950 205.950 91.050 208.050 ;
        RECT 70.950 184.950 73.050 187.050 ;
        RECT 55.950 182.100 58.050 184.200 ;
        RECT 56.400 181.350 57.600 182.100 ;
        RECT 67.950 181.950 70.050 184.050 ;
        RECT 77.400 183.600 78.450 202.950 ;
        RECT 101.400 202.050 102.450 209.400 ;
        RECT 110.400 202.050 111.450 223.950 ;
        RECT 116.400 217.200 117.450 253.950 ;
        RECT 124.350 252.300 126.450 254.400 ;
        RECT 125.250 245.700 126.450 252.300 ;
        RECT 136.950 250.950 139.050 255.000 ;
        RECT 142.650 248.700 143.850 267.300 ;
        RECT 145.950 256.950 148.050 259.050 ;
        RECT 146.400 255.900 147.600 256.650 ;
        RECT 145.950 253.800 148.050 255.900 ;
        RECT 139.650 247.500 143.850 248.700 ;
        RECT 139.650 246.600 141.750 247.500 ;
        RECT 124.350 243.600 126.450 245.700 ;
        RECT 152.400 238.050 153.450 280.950 ;
        RECT 167.400 277.050 168.450 286.950 ;
        RECT 169.950 286.800 172.050 288.900 ;
        RECT 176.400 287.400 177.600 289.650 ;
        RECT 188.400 288.900 189.450 331.950 ;
        RECT 190.950 331.800 193.050 333.900 ;
        RECT 202.950 331.800 205.050 333.900 ;
        RECT 209.400 332.400 210.600 334.650 ;
        RECT 191.400 322.050 192.450 331.800 ;
        RECT 209.400 330.450 210.450 332.400 ;
        RECT 209.400 329.400 213.450 330.450 ;
        RECT 190.950 319.950 193.050 322.050 ;
        RECT 166.950 274.950 169.050 277.050 ;
        RECT 172.950 274.950 175.050 277.050 ;
        RECT 154.950 271.950 157.050 274.050 ;
        RECT 155.400 255.900 156.450 271.950 ;
        RECT 173.400 261.450 174.450 274.950 ;
        RECT 176.400 264.450 177.450 287.400 ;
        RECT 187.950 286.800 190.050 288.900 ;
        RECT 191.400 274.050 192.450 319.950 ;
        RECT 212.400 319.050 213.450 329.400 ;
        RECT 211.950 316.950 214.050 319.050 ;
        RECT 196.950 301.950 199.050 304.050 ;
        RECT 197.400 294.600 198.450 301.950 ;
        RECT 208.950 298.950 211.050 301.050 ;
        RECT 209.400 295.200 210.450 298.950 ;
        RECT 197.400 292.350 198.600 294.600 ;
        RECT 202.950 293.100 205.050 295.200 ;
        RECT 208.950 293.100 211.050 295.200 ;
        RECT 203.400 292.350 204.600 293.100 ;
        RECT 196.950 289.950 199.050 292.050 ;
        RECT 199.950 289.950 202.050 292.050 ;
        RECT 202.950 289.950 205.050 292.050 ;
        RECT 205.950 289.950 208.050 292.050 ;
        RECT 200.400 287.400 201.600 289.650 ;
        RECT 206.400 287.400 207.600 289.650 ;
        RECT 200.400 280.050 201.450 287.400 ;
        RECT 199.950 277.950 202.050 280.050 ;
        RECT 190.950 271.950 193.050 274.050 ;
        RECT 199.950 271.950 202.050 274.050 ;
        RECT 187.950 265.950 190.050 268.050 ;
        RECT 176.400 263.400 180.450 264.450 ;
        RECT 173.400 260.400 177.450 261.450 ;
        RECT 166.950 256.950 169.050 259.050 ;
        RECT 169.950 256.950 172.050 259.050 ;
        RECT 154.950 253.800 157.050 255.900 ;
        RECT 163.950 253.950 166.050 256.050 ;
        RECT 167.400 254.400 168.600 256.650 ;
        RECT 157.950 247.950 160.050 250.050 ;
        RECT 151.950 235.950 154.050 238.050 ;
        RECT 124.950 223.950 127.050 226.050 ;
        RECT 115.950 216.450 118.050 217.200 ;
        RECT 125.400 216.600 126.450 223.950 ;
        RECT 142.800 220.200 144.900 222.300 ;
        RECT 151.800 220.500 153.900 222.600 ;
        RECT 119.400 216.450 120.600 216.600 ;
        RECT 115.950 215.400 120.600 216.450 ;
        RECT 115.950 215.100 118.050 215.400 ;
        RECT 119.400 214.350 120.600 215.400 ;
        RECT 125.400 214.350 126.600 216.600 ;
        RECT 130.950 215.100 133.050 217.200 ;
        RECT 139.950 215.100 142.050 217.200 ;
        RECT 118.950 211.950 121.050 214.050 ;
        RECT 121.950 211.950 124.050 214.050 ;
        RECT 124.950 211.950 127.050 214.050 ;
        RECT 122.400 210.900 123.600 211.650 ;
        RECT 121.950 208.800 124.050 210.900 ;
        RECT 131.400 205.050 132.450 215.100 ;
        RECT 140.400 214.350 141.600 215.100 ;
        RECT 140.100 211.950 142.200 214.050 ;
        RECT 143.100 207.600 144.000 220.200 ;
        RECT 149.400 217.350 150.600 219.600 ;
        RECT 149.100 214.950 151.200 217.050 ;
        RECT 144.900 213.900 147.000 214.200 ;
        RECT 153.000 213.900 153.900 220.500 ;
        RECT 144.900 213.000 153.900 213.900 ;
        RECT 144.900 212.100 147.000 213.000 ;
        RECT 150.000 211.200 152.100 212.100 ;
        RECT 144.900 210.000 152.100 211.200 ;
        RECT 144.900 209.100 147.000 210.000 ;
        RECT 142.500 205.500 144.600 207.600 ;
        RECT 149.100 206.100 151.200 208.200 ;
        RECT 153.000 207.900 153.900 213.000 ;
        RECT 154.800 211.950 156.900 214.050 ;
        RECT 155.400 210.900 156.600 211.650 ;
        RECT 154.950 208.800 157.050 210.900 ;
        RECT 152.400 205.800 154.500 207.900 ;
        RECT 130.950 202.950 133.050 205.050 ;
        RECT 149.400 203.550 150.600 205.800 ;
        RECT 100.950 199.950 103.050 202.050 ;
        RECT 109.950 199.950 112.050 202.050 ;
        RECT 149.400 193.050 150.450 203.550 ;
        RECT 158.400 199.050 159.450 247.950 ;
        RECT 151.950 196.950 154.050 199.050 ;
        RECT 157.950 196.950 160.050 199.050 ;
        RECT 103.950 190.950 106.050 193.050 ;
        RECT 112.950 190.950 115.050 193.050 ;
        RECT 148.950 190.950 151.050 193.050 ;
        RECT 85.950 184.950 88.050 187.050 ;
        RECT 52.950 178.950 55.050 181.050 ;
        RECT 55.950 178.950 58.050 181.050 ;
        RECT 58.950 178.950 61.050 181.050 ;
        RECT 46.950 175.950 49.050 178.050 ;
        RECT 53.400 177.000 54.600 178.650 ;
        RECT 59.400 177.900 60.600 178.650 ;
        RECT 68.400 177.900 69.450 181.950 ;
        RECT 77.400 181.350 78.600 183.600 ;
        RECT 86.400 181.050 87.450 184.950 ;
        RECT 88.950 181.950 91.050 184.050 ;
        RECT 97.950 182.100 100.050 184.200 ;
        RECT 104.400 183.600 105.450 190.950 ;
        RECT 73.950 178.950 76.050 181.050 ;
        RECT 76.950 178.950 79.050 181.050 ;
        RECT 79.950 178.950 82.050 181.050 ;
        RECT 85.950 178.950 88.050 181.050 ;
        RECT 74.400 177.900 75.600 178.650 ;
        RECT 80.400 178.050 81.600 178.650 ;
        RECT 89.400 178.050 90.450 181.950 ;
        RECT 98.400 181.350 99.600 182.100 ;
        RECT 104.400 181.350 105.600 183.600 ;
        RECT 97.950 178.950 100.050 181.050 ;
        RECT 100.950 178.950 103.050 181.050 ;
        RECT 103.950 178.950 106.050 181.050 ;
        RECT 106.950 178.950 109.050 181.050 ;
        RECT 43.950 172.950 46.050 175.050 ;
        RECT 52.950 172.950 55.050 177.000 ;
        RECT 58.950 175.800 61.050 177.900 ;
        RECT 67.950 175.800 70.050 177.900 ;
        RECT 73.950 175.800 76.050 177.900 ;
        RECT 80.400 176.400 85.050 178.050 ;
        RECT 81.000 175.950 85.050 176.400 ;
        RECT 88.950 175.950 91.050 178.050 ;
        RECT 101.400 176.400 102.600 178.650 ;
        RECT 107.400 177.900 108.600 178.650 ;
        RECT 101.400 156.450 102.450 176.400 ;
        RECT 106.950 175.800 109.050 177.900 ;
        RECT 98.400 155.400 102.450 156.450 ;
        RECT 29.400 146.400 33.450 147.450 ;
        RECT 17.100 142.500 19.200 144.600 ;
        RECT 14.100 133.950 16.200 136.050 ;
        RECT 17.100 135.900 18.000 142.500 ;
        RECT 26.100 142.200 28.200 144.300 ;
        RECT 20.400 139.350 21.600 141.600 ;
        RECT 19.800 136.950 21.900 139.050 ;
        RECT 24.000 135.900 26.100 136.200 ;
        RECT 17.100 135.000 26.100 135.900 ;
        RECT 17.100 129.900 18.000 135.000 ;
        RECT 24.000 134.100 26.100 135.000 ;
        RECT 18.900 133.200 21.000 134.100 ;
        RECT 18.900 132.000 26.100 133.200 ;
        RECT 24.000 131.100 26.100 132.000 ;
        RECT 16.500 127.800 18.600 129.900 ;
        RECT 19.800 128.100 21.900 130.200 ;
        RECT 27.000 129.600 27.900 142.200 ;
        RECT 29.400 138.450 30.600 138.600 ;
        RECT 32.400 138.450 33.450 146.400 ;
        RECT 51.000 141.450 55.050 142.050 ;
        RECT 29.400 137.400 33.450 138.450 ;
        RECT 50.400 139.950 55.050 141.450 ;
        RECT 50.400 138.600 51.450 139.950 ;
        RECT 29.400 136.350 30.600 137.400 ;
        RECT 50.400 136.350 51.600 138.600 ;
        RECT 58.950 137.100 61.050 139.200 ;
        RECT 64.950 138.000 67.050 142.050 ;
        RECT 28.800 133.950 30.900 136.050 ;
        RECT 46.950 133.950 49.050 136.050 ;
        RECT 49.950 133.950 52.050 136.050 ;
        RECT 47.400 131.400 48.600 133.650 ;
        RECT 20.400 127.050 21.600 127.800 ;
        RECT 26.400 127.500 28.500 129.600 ;
        RECT 47.400 127.050 48.450 131.400 ;
        RECT 19.950 124.950 22.050 127.050 ;
        RECT 34.950 124.950 37.050 127.050 ;
        RECT 46.950 124.950 49.050 127.050 ;
        RECT 10.950 103.950 13.050 106.050 ;
        RECT 16.950 104.100 19.050 106.200 ;
        RECT 22.950 105.000 25.050 109.050 ;
        RECT 11.400 94.050 12.450 103.950 ;
        RECT 17.400 103.350 18.600 104.100 ;
        RECT 23.400 103.350 24.600 105.000 ;
        RECT 16.950 100.950 19.050 103.050 ;
        RECT 19.950 100.950 22.050 103.050 ;
        RECT 22.950 100.950 25.050 103.050 ;
        RECT 25.950 100.950 28.050 103.050 ;
        RECT 20.400 99.000 21.600 100.650 ;
        RECT 26.400 99.900 27.600 100.650 ;
        RECT 19.950 94.950 22.050 99.000 ;
        RECT 25.950 97.800 28.050 99.900 ;
        RECT 10.950 91.950 13.050 94.050 ;
        RECT 16.950 59.100 19.050 61.200 ;
        RECT 17.400 58.350 18.600 59.100 ;
        RECT 16.950 55.950 19.050 58.050 ;
        RECT 19.950 55.950 22.050 58.050 ;
        RECT 20.400 53.400 21.600 55.650 ;
        RECT 26.400 55.050 27.450 97.800 ;
        RECT 35.400 97.050 36.450 124.950 ;
        RECT 49.950 112.950 52.050 115.050 ;
        RECT 43.950 105.000 46.050 109.050 ;
        RECT 50.400 105.600 51.450 112.950 ;
        RECT 59.400 109.050 60.450 137.100 ;
        RECT 65.400 136.350 66.600 138.000 ;
        RECT 70.950 137.100 73.050 139.200 ;
        RECT 88.950 137.100 91.050 139.200 ;
        RECT 71.400 136.350 72.600 137.100 ;
        RECT 89.400 136.350 90.600 137.100 ;
        RECT 64.950 133.950 67.050 136.050 ;
        RECT 67.950 133.950 70.050 136.050 ;
        RECT 70.950 133.950 73.050 136.050 ;
        RECT 85.950 133.950 88.050 136.050 ;
        RECT 88.950 133.950 91.050 136.050 ;
        RECT 68.400 131.400 69.600 133.650 ;
        RECT 86.400 132.900 87.600 133.650 ;
        RECT 68.400 118.050 69.450 131.400 ;
        RECT 73.950 130.800 76.050 132.900 ;
        RECT 85.950 130.800 88.050 132.900 ;
        RECT 67.950 115.950 70.050 118.050 ;
        RECT 74.400 112.050 75.450 130.800 ;
        RECT 98.400 127.050 99.450 155.400 ;
        RECT 113.400 145.050 114.450 190.950 ;
        RECT 152.400 189.450 153.450 196.950 ;
        RECT 124.950 183.000 127.050 187.050 ;
        RECT 148.800 186.300 150.900 188.400 ;
        RECT 152.400 187.200 153.600 189.450 ;
        RECT 125.400 181.350 126.600 183.000 ;
        RECT 130.950 182.100 133.050 184.200 ;
        RECT 142.950 183.450 145.050 184.200 ;
        RECT 146.400 183.450 147.600 183.600 ;
        RECT 142.950 182.400 147.600 183.450 ;
        RECT 142.950 182.100 145.050 182.400 ;
        RECT 131.400 181.350 132.600 182.100 ;
        RECT 121.950 178.950 124.050 181.050 ;
        RECT 124.950 178.950 127.050 181.050 ;
        RECT 127.950 178.950 130.050 181.050 ;
        RECT 130.950 178.950 133.050 181.050 ;
        RECT 118.950 177.450 121.050 177.900 ;
        RECT 122.400 177.450 123.600 178.650 ;
        RECT 118.950 176.400 123.600 177.450 ;
        RECT 128.400 176.400 129.600 178.650 ;
        RECT 118.950 175.800 121.050 176.400 ;
        RECT 112.950 142.950 115.050 145.050 ;
        RECT 106.950 137.100 109.050 139.200 ;
        RECT 113.400 138.600 114.450 142.950 ;
        RECT 107.400 136.350 108.600 137.100 ;
        RECT 113.400 136.350 114.600 138.600 ;
        RECT 103.950 133.950 106.050 136.050 ;
        RECT 106.950 133.950 109.050 136.050 ;
        RECT 109.950 133.950 112.050 136.050 ;
        RECT 112.950 133.950 115.050 136.050 ;
        RECT 104.400 131.400 105.600 133.650 ;
        RECT 110.400 132.900 111.600 133.650 ;
        RECT 119.400 133.050 120.450 175.800 ;
        RECT 128.400 172.050 129.450 176.400 ;
        RECT 127.950 169.950 130.050 172.050 ;
        RECT 139.950 160.950 142.050 163.050 ;
        RECT 121.950 136.950 124.050 139.050 ;
        RECT 130.950 137.100 133.050 139.200 ;
        RECT 97.950 124.950 100.050 127.050 ;
        RECT 79.950 115.950 82.050 118.050 ;
        RECT 73.950 109.950 76.050 112.050 ;
        RECT 55.950 106.950 58.050 109.050 ;
        RECT 58.950 106.950 61.050 109.050 ;
        RECT 44.400 103.350 45.600 105.000 ;
        RECT 50.400 103.350 51.600 105.600 ;
        RECT 40.950 100.950 43.050 103.050 ;
        RECT 43.950 100.950 46.050 103.050 ;
        RECT 46.950 100.950 49.050 103.050 ;
        RECT 49.950 100.950 52.050 103.050 ;
        RECT 41.400 99.900 42.600 100.650 ;
        RECT 40.950 97.800 43.050 99.900 ;
        RECT 47.400 99.000 48.600 100.650 ;
        RECT 34.950 94.950 37.050 97.050 ;
        RECT 46.950 94.950 49.050 99.000 ;
        RECT 56.400 88.050 57.450 106.950 ;
        RECT 58.950 103.800 61.050 105.900 ;
        RECT 67.950 104.100 70.050 106.200 ;
        RECT 74.400 105.600 75.450 109.950 ;
        RECT 59.400 94.050 60.450 103.800 ;
        RECT 68.400 103.350 69.600 104.100 ;
        RECT 74.400 103.350 75.600 105.600 ;
        RECT 64.950 100.950 67.050 103.050 ;
        RECT 67.950 100.950 70.050 103.050 ;
        RECT 70.950 100.950 73.050 103.050 ;
        RECT 73.950 100.950 76.050 103.050 ;
        RECT 61.950 97.950 64.050 100.050 ;
        RECT 65.400 98.400 66.600 100.650 ;
        RECT 71.400 99.000 72.600 100.650 ;
        RECT 62.400 94.050 63.450 97.950 ;
        RECT 58.950 91.950 61.050 94.050 ;
        RECT 61.950 91.950 64.050 94.050 ;
        RECT 49.950 85.950 52.050 88.050 ;
        RECT 55.950 85.950 58.050 88.050 ;
        RECT 46.950 73.950 49.050 76.050 ;
        RECT 40.950 67.950 43.050 70.050 ;
        RECT 34.950 59.100 37.050 61.200 ;
        RECT 41.400 60.600 42.450 67.950 ;
        RECT 35.400 58.350 36.600 59.100 ;
        RECT 41.400 58.350 42.600 60.600 ;
        RECT 34.950 55.950 37.050 58.050 ;
        RECT 37.950 55.950 40.050 58.050 ;
        RECT 40.950 55.950 43.050 58.050 ;
        RECT 20.400 46.050 21.450 53.400 ;
        RECT 25.950 52.950 28.050 55.050 ;
        RECT 31.950 52.950 34.050 55.050 ;
        RECT 38.400 54.900 39.600 55.650 ;
        RECT 19.950 43.950 22.050 46.050 ;
        RECT 25.950 26.100 28.050 28.200 ;
        RECT 16.950 22.950 19.050 25.050 ;
        RECT 19.950 22.950 22.050 25.050 ;
        RECT 20.400 21.900 21.600 22.650 ;
        RECT 26.400 22.050 27.450 26.100 ;
        RECT 19.950 19.800 22.050 21.900 ;
        RECT 25.950 19.950 28.050 22.050 ;
        RECT 32.400 21.450 33.450 52.950 ;
        RECT 37.950 52.800 40.050 54.900 ;
        RECT 40.950 26.100 43.050 28.200 ;
        RECT 41.400 25.350 42.600 26.100 ;
        RECT 35.100 22.950 37.200 25.050 ;
        RECT 40.500 22.950 42.600 25.050 ;
        RECT 43.800 22.950 45.900 25.050 ;
        RECT 35.400 21.900 36.600 22.650 ;
        RECT 34.950 21.450 37.050 21.900 ;
        RECT 32.400 20.400 37.050 21.450 ;
        RECT 44.400 21.450 45.600 22.650 ;
        RECT 47.400 21.450 48.450 73.950 ;
        RECT 50.400 61.200 51.450 85.950 ;
        RECT 58.950 73.950 61.050 76.050 ;
        RECT 49.950 59.100 52.050 61.200 ;
        RECT 59.400 60.600 60.450 73.950 ;
        RECT 65.400 70.050 66.450 98.400 ;
        RECT 70.950 94.950 73.050 99.000 ;
        RECT 80.400 97.050 81.450 115.950 ;
        RECT 104.400 115.050 105.450 131.400 ;
        RECT 109.950 130.800 112.050 132.900 ;
        RECT 118.950 130.950 121.050 133.050 ;
        RECT 122.400 130.050 123.450 136.950 ;
        RECT 131.400 136.350 132.600 137.100 ;
        RECT 127.950 133.950 130.050 136.050 ;
        RECT 130.950 133.950 133.050 136.050 ;
        RECT 133.950 133.950 136.050 136.050 ;
        RECT 124.950 130.950 127.050 133.050 ;
        RECT 128.400 132.000 129.600 133.650 ;
        RECT 121.950 127.950 124.050 130.050 ;
        RECT 121.950 118.950 124.050 121.050 ;
        RECT 103.950 112.950 106.050 115.050 ;
        RECT 106.950 112.950 109.050 115.050 ;
        RECT 88.950 104.100 91.050 106.200 ;
        RECT 107.400 105.600 108.450 112.950 ;
        RECT 89.400 103.350 90.600 104.100 ;
        RECT 107.400 103.350 108.600 105.600 ;
        RECT 112.950 104.100 115.050 106.200 ;
        RECT 113.400 103.350 114.600 104.100 ;
        RECT 88.950 100.950 91.050 103.050 ;
        RECT 91.950 100.950 94.050 103.050 ;
        RECT 106.950 100.950 109.050 103.050 ;
        RECT 109.950 100.950 112.050 103.050 ;
        RECT 112.950 100.950 115.050 103.050 ;
        RECT 115.950 100.950 118.050 103.050 ;
        RECT 92.400 99.900 93.600 100.650 ;
        RECT 110.400 99.900 111.600 100.650 ;
        RECT 116.400 99.900 117.600 100.650 ;
        RECT 122.400 99.900 123.450 118.950 ;
        RECT 91.950 97.800 94.050 99.900 ;
        RECT 109.950 97.800 112.050 99.900 ;
        RECT 115.950 97.800 118.050 99.900 ;
        RECT 121.950 97.800 124.050 99.900 ;
        RECT 79.950 94.950 82.050 97.050 ;
        RECT 70.950 91.800 73.050 93.900 ;
        RECT 61.800 69.000 63.900 70.050 ;
        RECT 61.800 67.950 64.050 69.000 ;
        RECT 64.950 67.950 67.050 70.050 ;
        RECT 61.950 66.450 64.050 67.950 ;
        RECT 61.950 66.000 69.450 66.450 ;
        RECT 62.400 65.400 70.050 66.000 ;
        RECT 67.950 61.950 70.050 65.400 ;
        RECT 50.400 55.050 51.450 59.100 ;
        RECT 59.400 58.350 60.600 60.600 ;
        RECT 64.950 59.100 67.050 61.200 ;
        RECT 65.400 58.350 66.600 59.100 ;
        RECT 55.950 55.950 58.050 58.050 ;
        RECT 58.950 55.950 61.050 58.050 ;
        RECT 61.950 55.950 64.050 58.050 ;
        RECT 64.950 55.950 67.050 58.050 ;
        RECT 49.950 52.950 52.050 55.050 ;
        RECT 56.400 53.400 57.600 55.650 ;
        RECT 62.400 54.900 63.600 55.650 ;
        RECT 71.400 55.050 72.450 91.800 ;
        RECT 73.950 67.950 76.050 70.050 ;
        RECT 106.950 67.950 109.050 70.050 ;
        RECT 44.400 20.400 48.450 21.450 ;
        RECT 34.950 19.800 37.050 20.400 ;
        RECT 47.400 16.050 48.450 20.400 ;
        RECT 50.400 19.050 51.450 52.950 ;
        RECT 56.400 28.050 57.450 53.400 ;
        RECT 61.950 52.800 64.050 54.900 ;
        RECT 70.950 52.950 73.050 55.050 ;
        RECT 74.400 54.450 75.450 67.950 ;
        RECT 82.950 60.000 85.050 64.050 ;
        RECT 107.400 61.200 108.450 67.950 ;
        RECT 83.400 58.350 84.600 60.000 ;
        RECT 94.950 59.100 97.050 61.200 ;
        RECT 100.950 59.100 103.050 61.200 ;
        RECT 106.950 59.100 109.050 61.200 ;
        RECT 79.950 55.950 82.050 58.050 ;
        RECT 82.950 55.950 85.050 58.050 ;
        RECT 85.950 55.950 88.050 58.050 ;
        RECT 80.400 54.450 81.600 55.650 ;
        RECT 74.400 53.400 81.600 54.450 ;
        RECT 86.400 54.450 87.600 55.650 ;
        RECT 91.950 54.450 94.050 55.050 ;
        RECT 86.400 53.400 94.050 54.450 ;
        RECT 91.950 52.950 94.050 53.400 ;
        RECT 95.400 46.050 96.450 59.100 ;
        RECT 101.400 58.350 102.600 59.100 ;
        RECT 107.400 58.350 108.600 59.100 ;
        RECT 100.950 55.950 103.050 58.050 ;
        RECT 103.950 55.950 106.050 58.050 ;
        RECT 106.950 55.950 109.050 58.050 ;
        RECT 109.950 55.950 112.050 58.050 ;
        RECT 104.400 53.400 105.600 55.650 ;
        RECT 110.400 54.900 111.600 55.650 ;
        RECT 61.950 43.950 64.050 46.050 ;
        RECT 94.950 43.950 97.050 46.050 ;
        RECT 55.950 25.950 58.050 28.050 ;
        RECT 62.400 27.600 63.450 43.950 ;
        RECT 104.400 37.050 105.450 53.400 ;
        RECT 109.950 52.800 112.050 54.900 ;
        RECT 116.400 52.050 117.450 97.800 ;
        RECT 125.400 70.050 126.450 130.950 ;
        RECT 127.950 127.950 130.050 132.000 ;
        RECT 134.400 131.400 135.600 133.650 ;
        RECT 134.400 115.050 135.450 131.400 ;
        RECT 140.400 121.050 141.450 160.950 ;
        RECT 143.400 157.050 144.450 182.100 ;
        RECT 146.400 181.350 147.600 182.400 ;
        RECT 146.100 178.950 148.200 181.050 ;
        RECT 149.100 180.900 150.000 186.300 ;
        RECT 152.100 184.800 154.200 186.900 ;
        RECT 156.000 183.900 158.100 185.700 ;
        RECT 150.900 182.700 159.600 183.900 ;
        RECT 150.900 181.800 153.000 182.700 ;
        RECT 149.100 179.700 156.000 180.900 ;
        RECT 149.100 172.500 150.300 179.700 ;
        RECT 152.100 175.950 154.200 178.050 ;
        RECT 155.100 177.300 156.000 179.700 ;
        RECT 152.400 173.400 153.600 175.650 ;
        RECT 155.100 175.200 157.200 177.300 ;
        RECT 158.700 173.700 159.600 182.700 ;
        RECT 160.800 178.950 162.900 181.050 ;
        RECT 161.400 177.900 162.600 178.650 ;
        RECT 160.950 175.800 163.050 177.900 ;
        RECT 148.800 170.400 150.900 172.500 ;
        RECT 158.400 171.600 160.500 173.700 ;
        RECT 142.950 154.950 145.050 157.050 ;
        RECT 151.950 154.950 154.050 157.050 ;
        RECT 142.950 142.950 145.050 145.050 ;
        RECT 139.950 118.950 142.050 121.050 ;
        RECT 133.950 112.950 136.050 115.050 ;
        RECT 143.400 112.050 144.450 142.950 ;
        RECT 145.950 136.950 148.050 139.050 ;
        RECT 152.400 138.600 153.450 154.950 ;
        RECT 130.950 108.450 133.050 112.050 ;
        RECT 142.950 109.950 145.050 112.050 ;
        RECT 136.950 108.450 139.050 109.050 ;
        RECT 130.950 108.000 139.050 108.450 ;
        RECT 131.400 107.400 139.050 108.000 ;
        RECT 136.950 106.950 139.050 107.400 ;
        RECT 142.950 106.800 145.050 108.900 ;
        RECT 133.950 104.100 136.050 106.200 ;
        RECT 134.400 103.350 135.600 104.100 ;
        RECT 130.950 100.950 133.050 103.050 ;
        RECT 133.950 100.950 136.050 103.050 ;
        RECT 136.950 100.950 139.050 103.050 ;
        RECT 131.400 99.900 132.600 100.650 ;
        RECT 130.950 97.800 133.050 99.900 ;
        RECT 137.400 99.000 138.600 100.650 ;
        RECT 136.950 94.950 139.050 99.000 ;
        RECT 143.400 97.050 144.450 106.800 ;
        RECT 146.400 99.900 147.450 136.950 ;
        RECT 152.400 136.350 153.600 138.600 ;
        RECT 160.950 137.100 163.050 139.200 ;
        RECT 151.950 133.950 154.050 136.050 ;
        RECT 154.950 133.950 157.050 136.050 ;
        RECT 155.400 132.450 156.600 133.650 ;
        RECT 161.400 132.450 162.450 137.100 ;
        RECT 155.400 131.400 162.450 132.450 ;
        RECT 148.950 109.950 151.050 112.050 ;
        RECT 158.400 111.450 159.450 131.400 ;
        RECT 164.400 115.050 165.450 253.950 ;
        RECT 167.400 238.050 168.450 254.400 ;
        RECT 166.950 235.950 169.050 238.050 ;
        RECT 176.400 219.450 177.450 260.400 ;
        RECT 179.400 223.050 180.450 263.400 ;
        RECT 188.400 261.600 189.450 265.950 ;
        RECT 188.400 259.350 189.600 261.600 ;
        RECT 193.950 260.100 196.050 262.200 ;
        RECT 194.400 259.350 195.600 260.100 ;
        RECT 184.950 256.950 187.050 259.050 ;
        RECT 187.950 256.950 190.050 259.050 ;
        RECT 190.950 256.950 193.050 259.050 ;
        RECT 193.950 256.950 196.050 259.050 ;
        RECT 185.400 255.000 186.600 256.650 ;
        RECT 191.400 255.900 192.600 256.650 ;
        RECT 200.400 255.900 201.450 271.950 ;
        RECT 206.400 271.050 207.450 287.400 ;
        RECT 212.400 283.050 213.450 316.950 ;
        RECT 218.400 294.450 219.450 343.950 ;
        RECT 223.950 337.950 226.050 340.050 ;
        RECT 232.950 338.100 235.050 340.200 ;
        RECT 224.400 333.900 225.450 337.950 ;
        RECT 233.400 337.350 234.600 338.100 ;
        RECT 229.950 334.950 232.050 337.050 ;
        RECT 232.950 334.950 235.050 337.050 ;
        RECT 235.950 334.950 238.050 337.050 ;
        RECT 223.950 331.800 226.050 333.900 ;
        RECT 242.400 307.050 243.450 365.400 ;
        RECT 256.950 338.100 259.050 340.200 ;
        RECT 257.400 337.350 258.600 338.100 ;
        RECT 268.950 337.950 271.050 340.050 ;
        RECT 274.950 338.100 277.050 340.200 ;
        RECT 281.400 339.600 282.450 407.400 ;
        RECT 290.400 400.050 291.450 410.400 ;
        RECT 296.400 400.050 297.450 410.400 ;
        RECT 289.950 397.950 292.050 400.050 ;
        RECT 295.950 397.950 298.050 400.050 ;
        RECT 283.950 376.950 286.050 379.050 ;
        RECT 302.400 378.450 303.450 469.950 ;
        RECT 305.400 463.050 306.450 487.800 ;
        RECT 311.400 484.050 312.450 490.950 ;
        RECT 310.950 481.950 313.050 484.050 ;
        RECT 332.400 472.050 333.450 496.950 ;
        RECT 335.400 496.050 336.450 505.950 ;
        RECT 334.950 493.950 337.050 496.050 ;
        RECT 340.950 495.000 343.050 499.050 ;
        RECT 341.400 493.350 342.600 495.000 ;
        RECT 337.950 490.950 340.050 493.050 ;
        RECT 340.950 490.950 343.050 493.050 ;
        RECT 343.950 490.950 346.050 493.050 ;
        RECT 338.400 489.900 339.600 490.650 ;
        RECT 344.400 489.900 345.600 490.650 ;
        RECT 350.400 489.900 351.450 517.950 ;
        RECT 356.400 502.050 357.450 527.100 ;
        RECT 365.400 526.350 366.600 527.100 ;
        RECT 371.400 526.350 372.600 527.100 ;
        RECT 364.950 523.950 367.050 526.050 ;
        RECT 367.950 523.950 370.050 526.050 ;
        RECT 370.950 523.950 373.050 526.050 ;
        RECT 373.950 523.950 376.050 526.050 ;
        RECT 361.950 520.950 364.050 523.050 ;
        RECT 368.400 521.400 369.600 523.650 ;
        RECT 374.400 521.400 375.600 523.650 ;
        RECT 380.400 522.900 381.450 527.100 ;
        RECT 362.400 505.050 363.450 520.950 ;
        RECT 368.400 517.050 369.450 521.400 ;
        RECT 367.950 514.950 370.050 517.050 ;
        RECT 361.950 502.950 364.050 505.050 ;
        RECT 355.950 499.950 358.050 502.050 ;
        RECT 362.400 495.600 363.450 502.950 ;
        RECT 374.400 502.050 375.450 521.400 ;
        RECT 379.950 520.800 382.050 522.900 ;
        RECT 380.400 514.050 381.450 520.800 ;
        RECT 383.400 517.050 384.450 527.100 ;
        RECT 389.400 526.350 390.600 527.100 ;
        RECT 395.400 526.350 396.600 528.000 ;
        RECT 388.950 523.950 391.050 526.050 ;
        RECT 391.950 523.950 394.050 526.050 ;
        RECT 394.950 523.950 397.050 526.050 ;
        RECT 397.950 523.950 400.050 526.050 ;
        RECT 392.400 522.900 393.600 523.650 ;
        RECT 398.400 522.900 399.600 523.650 ;
        RECT 391.950 520.800 394.050 522.900 ;
        RECT 397.950 520.800 400.050 522.900 ;
        RECT 382.950 514.950 385.050 517.050 ;
        RECT 379.950 511.950 382.050 514.050 ;
        RECT 391.950 505.950 394.050 508.050 ;
        RECT 404.400 507.450 405.450 547.950 ;
        RECT 406.950 527.100 409.050 529.200 ;
        RECT 415.950 527.100 418.050 529.200 ;
        RECT 422.400 528.600 423.450 550.950 ;
        RECT 446.400 544.050 447.450 572.100 ;
        RECT 455.400 571.350 456.600 573.600 ;
        RECT 472.950 572.100 475.050 574.200 ;
        RECT 473.400 571.350 474.600 572.100 ;
        RECT 451.950 568.950 454.050 571.050 ;
        RECT 454.950 568.950 457.050 571.050 ;
        RECT 457.950 568.950 460.050 571.050 ;
        RECT 472.950 568.950 475.050 571.050 ;
        RECT 475.950 568.950 478.050 571.050 ;
        RECT 452.400 567.900 453.600 568.650 ;
        RECT 458.400 567.900 459.600 568.650 ;
        RECT 451.950 565.800 454.050 567.900 ;
        RECT 457.950 565.800 460.050 567.900 ;
        RECT 469.950 565.800 472.050 567.900 ;
        RECT 470.400 562.050 471.450 565.800 ;
        RECT 469.950 559.950 472.050 562.050 ;
        RECT 466.950 556.950 469.050 559.050 ;
        RECT 467.400 547.050 468.450 556.950 ;
        RECT 482.400 553.050 483.450 595.950 ;
        RECT 491.400 592.050 492.450 599.400 ;
        RECT 508.950 595.950 511.050 600.000 ;
        RECT 514.950 598.800 517.050 600.900 ;
        RECT 523.950 598.950 526.050 601.050 ;
        RECT 502.950 592.950 505.050 595.050 ;
        RECT 490.950 589.950 493.050 592.050 ;
        RECT 491.400 586.050 492.450 589.950 ;
        RECT 490.950 583.950 493.050 586.050 ;
        RECT 503.400 574.050 504.450 592.950 ;
        RECT 505.950 586.950 508.050 589.050 ;
        RECT 502.950 571.950 505.050 574.050 ;
        RECT 491.100 568.950 493.200 571.050 ;
        RECT 496.500 568.950 498.600 571.050 ;
        RECT 499.800 568.950 501.900 571.050 ;
        RECT 491.400 566.400 492.600 568.650 ;
        RECT 500.400 566.400 501.600 568.650 ;
        RECT 491.400 556.050 492.450 566.400 ;
        RECT 500.400 562.050 501.450 566.400 ;
        RECT 506.400 562.050 507.450 586.950 ;
        RECT 523.950 583.950 526.050 586.050 ;
        RECT 508.950 572.100 511.050 574.200 ;
        RECT 514.950 572.100 517.050 574.200 ;
        RECT 499.950 559.950 502.050 562.050 ;
        RECT 505.950 559.950 508.050 562.050 ;
        RECT 509.400 556.050 510.450 572.100 ;
        RECT 515.400 571.350 516.600 572.100 ;
        RECT 514.950 568.950 517.050 571.050 ;
        RECT 517.950 568.950 520.050 571.050 ;
        RECT 518.400 567.900 519.600 568.650 ;
        RECT 517.950 565.800 520.050 567.900 ;
        RECT 490.950 553.950 493.050 556.050 ;
        RECT 508.950 553.950 511.050 556.050 ;
        RECT 481.950 550.950 484.050 553.050 ;
        RECT 466.950 544.950 469.050 547.050 ;
        RECT 430.950 541.950 433.050 544.050 ;
        RECT 445.950 541.950 448.050 544.050 ;
        RECT 454.950 541.950 457.050 544.050 ;
        RECT 407.400 523.050 408.450 527.100 ;
        RECT 416.400 526.350 417.600 527.100 ;
        RECT 422.400 526.350 423.600 528.600 ;
        RECT 412.950 523.950 415.050 526.050 ;
        RECT 415.950 523.950 418.050 526.050 ;
        RECT 418.950 523.950 421.050 526.050 ;
        RECT 421.950 523.950 424.050 526.050 ;
        RECT 406.950 520.950 409.050 523.050 ;
        RECT 413.400 522.900 414.600 523.650 ;
        RECT 412.950 520.800 415.050 522.900 ;
        RECT 419.400 521.400 420.600 523.650 ;
        RECT 401.400 506.400 405.450 507.450 ;
        RECT 367.950 499.950 370.050 502.050 ;
        RECT 373.950 499.950 376.050 502.050 ;
        RECT 368.400 496.050 369.450 499.950 ;
        RECT 370.950 496.950 373.050 499.050 ;
        RECT 362.400 493.350 363.600 495.600 ;
        RECT 367.950 493.950 370.050 496.050 ;
        RECT 358.950 490.950 361.050 493.050 ;
        RECT 361.950 490.950 364.050 493.050 ;
        RECT 364.950 490.950 367.050 493.050 ;
        RECT 337.950 487.800 340.050 489.900 ;
        RECT 343.950 487.800 346.050 489.900 ;
        RECT 349.950 487.800 352.050 489.900 ;
        RECT 371.400 487.050 372.450 496.950 ;
        RECT 392.400 496.200 393.450 505.950 ;
        RECT 376.950 493.950 379.050 496.050 ;
        RECT 391.950 494.100 394.050 496.200 ;
        RECT 370.950 484.950 373.050 487.050 ;
        RECT 377.400 486.450 378.450 493.950 ;
        RECT 392.400 493.350 393.600 494.100 ;
        RECT 382.950 490.950 385.050 493.050 ;
        RECT 385.950 490.950 388.050 493.050 ;
        RECT 388.950 490.950 391.050 493.050 ;
        RECT 391.950 490.950 394.050 493.050 ;
        RECT 394.950 490.950 397.050 493.050 ;
        RECT 389.400 488.400 390.600 490.650 ;
        RECT 395.400 489.900 396.600 490.650 ;
        RECT 377.400 485.400 381.450 486.450 ;
        RECT 361.950 475.950 364.050 478.050 ;
        RECT 331.950 469.950 334.050 472.050 ;
        RECT 304.950 460.950 307.050 463.050 ;
        RECT 346.950 454.950 349.050 457.050 ;
        RECT 313.950 445.950 316.050 448.050 ;
        RECT 316.950 445.950 319.050 448.050 ;
        RECT 319.950 445.950 322.050 448.050 ;
        RECT 334.950 445.950 337.050 448.050 ;
        RECT 337.950 445.950 340.050 448.050 ;
        RECT 340.950 445.950 343.050 448.050 ;
        RECT 317.400 443.400 318.600 445.650 ;
        RECT 338.400 443.400 339.600 445.650 ;
        RECT 347.400 445.050 348.450 454.950 ;
        RECT 349.950 449.100 352.050 451.200 ;
        RECT 355.950 449.100 358.050 451.200 ;
        RECT 362.400 450.600 363.450 475.950 ;
        RECT 380.400 469.050 381.450 485.400 ;
        RECT 389.400 478.050 390.450 488.400 ;
        RECT 394.950 487.800 397.050 489.900 ;
        RECT 395.400 484.050 396.450 487.800 ;
        RECT 394.950 481.950 397.050 484.050 ;
        RECT 388.950 475.950 391.050 478.050 ;
        RECT 379.950 466.950 382.050 469.050 ;
        RECT 401.400 462.450 402.450 506.400 ;
        RECT 409.950 502.950 412.050 505.050 ;
        RECT 403.950 496.950 406.050 499.050 ;
        RECT 404.400 478.050 405.450 496.950 ;
        RECT 410.400 495.600 411.450 502.950 ;
        RECT 413.400 499.050 414.450 520.800 ;
        RECT 419.400 517.050 420.450 521.400 ;
        RECT 427.950 517.950 430.050 520.050 ;
        RECT 418.950 514.950 421.050 517.050 ;
        RECT 428.400 511.050 429.450 517.950 ;
        RECT 431.400 514.050 432.450 541.950 ;
        RECT 445.950 538.800 448.050 540.900 ;
        RECT 439.950 527.100 442.050 529.200 ;
        RECT 446.400 528.600 447.450 538.800 ;
        RECT 440.400 526.350 441.600 527.100 ;
        RECT 446.400 526.350 447.600 528.600 ;
        RECT 448.950 526.950 451.050 532.050 ;
        RECT 436.950 523.950 439.050 526.050 ;
        RECT 439.950 523.950 442.050 526.050 ;
        RECT 442.950 523.950 445.050 526.050 ;
        RECT 445.950 523.950 448.050 526.050 ;
        RECT 451.950 523.950 454.050 526.050 ;
        RECT 437.400 522.900 438.600 523.650 ;
        RECT 443.400 522.900 444.600 523.650 ;
        RECT 436.950 520.800 439.050 522.900 ;
        RECT 442.950 520.800 445.050 522.900 ;
        RECT 430.950 511.950 433.050 514.050 ;
        RECT 448.950 511.950 451.050 514.050 ;
        RECT 427.950 508.950 430.050 511.050 ;
        RECT 433.950 502.950 436.050 505.050 ;
        RECT 442.950 502.950 445.050 505.050 ;
        RECT 420.000 501.450 424.050 502.050 ;
        RECT 419.400 499.950 424.050 501.450 ;
        RECT 430.950 499.950 433.050 502.050 ;
        RECT 412.950 496.950 415.050 499.050 ;
        RECT 410.400 493.350 411.600 495.600 ;
        RECT 409.950 490.950 412.050 493.050 ;
        RECT 412.950 490.950 415.050 493.050 ;
        RECT 413.400 489.900 414.600 490.650 ;
        RECT 419.400 490.050 420.450 499.950 ;
        RECT 421.950 493.950 424.050 496.050 ;
        RECT 431.400 495.600 432.450 499.950 ;
        RECT 434.400 499.050 435.450 502.950 ;
        RECT 436.950 499.950 439.050 502.050 ;
        RECT 433.950 496.950 436.050 499.050 ;
        RECT 437.400 495.600 438.450 499.950 ;
        RECT 412.950 487.800 415.050 489.900 ;
        RECT 418.800 487.950 420.900 490.050 ;
        RECT 422.400 489.900 423.450 493.950 ;
        RECT 431.400 493.350 432.600 495.600 ;
        RECT 437.400 493.350 438.600 495.600 ;
        RECT 443.400 493.050 444.450 502.950 ;
        RECT 445.950 493.950 448.050 496.050 ;
        RECT 427.950 490.950 430.050 493.050 ;
        RECT 430.950 490.950 433.050 493.050 ;
        RECT 433.950 490.950 436.050 493.050 ;
        RECT 436.950 490.950 439.050 493.050 ;
        RECT 442.950 490.950 445.050 493.050 ;
        RECT 428.400 489.900 429.600 490.650 ;
        RECT 421.950 487.800 424.050 489.900 ;
        RECT 427.950 487.800 430.050 489.900 ;
        RECT 434.400 488.400 435.600 490.650 ;
        RECT 434.400 484.050 435.450 488.400 ;
        RECT 433.950 481.950 436.050 484.050 ;
        RECT 412.950 478.950 415.050 481.050 ;
        RECT 424.950 478.950 427.050 481.050 ;
        RECT 403.950 475.950 406.050 478.050 ;
        RECT 413.400 469.050 414.450 478.950 ;
        RECT 418.950 472.950 421.050 475.050 ;
        RECT 412.950 466.950 415.050 469.050 ;
        RECT 398.400 461.400 402.450 462.450 ;
        RECT 394.950 457.950 397.050 460.050 ;
        RECT 379.950 454.950 382.050 457.050 ;
        RECT 370.950 451.950 373.050 454.050 ;
        RECT 317.400 439.050 318.450 443.400 ;
        RECT 316.950 436.950 319.050 439.050 ;
        RECT 338.400 424.050 339.450 443.400 ;
        RECT 346.950 442.950 349.050 445.050 ;
        RECT 337.950 421.950 340.050 424.050 ;
        RECT 314.100 412.950 316.200 415.050 ;
        RECT 319.500 412.950 321.600 415.050 ;
        RECT 322.800 412.950 324.900 415.050 ;
        RECT 338.100 412.950 340.200 415.050 ;
        RECT 343.500 412.950 345.600 415.050 ;
        RECT 346.800 412.950 348.900 415.050 ;
        RECT 310.950 409.950 313.050 412.050 ;
        RECT 314.400 411.900 315.600 412.650 ;
        RECT 299.400 377.400 303.450 378.450 ;
        RECT 284.400 340.050 285.450 376.950 ;
        RECT 286.950 371.100 289.050 373.200 ;
        RECT 295.950 371.100 298.050 373.200 ;
        RECT 287.400 370.350 288.600 371.100 ;
        RECT 296.400 370.350 297.600 371.100 ;
        RECT 287.100 367.950 289.200 370.050 ;
        RECT 292.500 367.950 294.600 370.050 ;
        RECT 295.800 367.950 297.900 370.050 ;
        RECT 299.400 352.050 300.450 377.400 ;
        RECT 311.400 376.050 312.450 409.950 ;
        RECT 313.950 409.800 316.050 411.900 ;
        RECT 323.400 410.400 324.600 412.650 ;
        RECT 347.400 411.000 348.600 412.650 ;
        RECT 323.400 400.050 324.450 410.400 ;
        RECT 346.950 408.450 349.050 411.000 ;
        RECT 350.400 408.450 351.450 449.100 ;
        RECT 356.400 448.350 357.600 449.100 ;
        RECT 362.400 448.350 363.600 450.600 ;
        RECT 355.950 445.950 358.050 448.050 ;
        RECT 358.950 445.950 361.050 448.050 ;
        RECT 361.950 445.950 364.050 448.050 ;
        RECT 364.950 445.950 367.050 448.050 ;
        RECT 359.400 444.900 360.600 445.650 ;
        RECT 358.950 442.800 361.050 444.900 ;
        RECT 365.400 443.400 366.600 445.650 ;
        RECT 365.400 433.050 366.450 443.400 ;
        RECT 364.950 430.950 367.050 433.050 ;
        RECT 371.400 424.050 372.450 451.950 ;
        RECT 380.400 450.600 381.450 454.950 ;
        RECT 380.400 448.350 381.600 450.600 ;
        RECT 385.950 450.000 388.050 454.050 ;
        RECT 386.400 448.350 387.600 450.000 ;
        RECT 379.950 445.950 382.050 448.050 ;
        RECT 382.950 445.950 385.050 448.050 ;
        RECT 385.950 445.950 388.050 448.050 ;
        RECT 388.950 445.950 391.050 448.050 ;
        RECT 383.400 443.400 384.600 445.650 ;
        RECT 389.400 444.900 390.600 445.650 ;
        RECT 395.400 444.900 396.450 457.950 ;
        RECT 383.400 430.050 384.450 443.400 ;
        RECT 388.950 442.800 391.050 444.900 ;
        RECT 394.950 442.800 397.050 444.900 ;
        RECT 391.950 436.950 394.050 439.050 ;
        RECT 382.950 427.950 385.050 430.050 ;
        RECT 370.950 421.950 373.050 424.050 ;
        RECT 382.950 421.950 385.050 424.050 ;
        RECT 364.950 416.100 367.050 418.200 ;
        RECT 365.400 415.350 366.600 416.100 ;
        RECT 376.950 415.950 379.050 418.050 ;
        RECT 383.400 417.600 384.450 421.950 ;
        RECT 361.950 412.950 364.050 415.050 ;
        RECT 364.950 412.950 367.050 415.050 ;
        RECT 367.950 412.950 370.050 415.050 ;
        RECT 362.400 411.000 363.600 412.650 ;
        RECT 346.950 407.400 351.450 408.450 ;
        RECT 346.950 406.950 349.050 407.400 ;
        RECT 361.950 406.950 364.050 411.000 ;
        RECT 368.400 410.400 369.600 412.650 ;
        RECT 368.400 400.050 369.450 410.400 ;
        RECT 377.400 409.050 378.450 415.950 ;
        RECT 383.400 415.350 384.600 417.600 ;
        RECT 382.950 412.950 385.050 415.050 ;
        RECT 385.950 412.950 388.050 415.050 ;
        RECT 386.400 410.400 387.600 412.650 ;
        RECT 386.400 409.050 387.450 410.400 ;
        RECT 376.950 406.950 379.050 409.050 ;
        RECT 386.400 407.400 391.050 409.050 ;
        RECT 387.000 406.950 391.050 407.400 ;
        RECT 322.950 397.950 325.050 400.050 ;
        RECT 367.950 397.950 370.050 400.050 ;
        RECT 379.950 391.950 382.050 394.050 ;
        RECT 316.950 388.950 319.050 391.050 ;
        RECT 325.950 388.950 328.050 391.050 ;
        RECT 317.400 382.050 318.450 388.950 ;
        RECT 316.950 379.950 319.050 382.050 ;
        RECT 304.950 373.950 307.050 376.050 ;
        RECT 310.950 373.950 313.050 376.050 ;
        RECT 298.950 349.950 301.050 352.050 ;
        RECT 286.950 346.950 289.050 349.050 ;
        RECT 253.950 334.950 256.050 337.050 ;
        RECT 256.950 334.950 259.050 337.050 ;
        RECT 259.950 334.950 262.050 337.050 ;
        RECT 232.950 304.950 235.050 307.050 ;
        RECT 241.950 304.950 244.050 307.050 ;
        RECT 250.950 304.950 253.050 307.050 ;
        RECT 269.400 306.450 270.450 337.950 ;
        RECT 275.400 337.350 276.600 338.100 ;
        RECT 281.400 337.350 282.600 339.600 ;
        RECT 283.950 337.950 286.050 340.050 ;
        RECT 274.950 334.950 277.050 337.050 ;
        RECT 277.950 334.950 280.050 337.050 ;
        RECT 280.950 334.950 283.050 337.050 ;
        RECT 278.400 333.900 279.600 334.650 ;
        RECT 287.400 334.050 288.450 346.950 ;
        RECT 289.950 337.950 292.050 340.050 ;
        RECT 298.950 338.100 301.050 340.200 ;
        RECT 305.400 339.450 306.450 373.950 ;
        RECT 311.400 372.600 312.450 373.950 ;
        RECT 311.400 370.350 312.600 372.600 ;
        RECT 310.950 367.950 313.050 370.050 ;
        RECT 313.950 367.950 316.050 370.050 ;
        RECT 316.950 367.950 319.050 370.050 ;
        RECT 314.400 366.000 315.600 367.650 ;
        RECT 313.950 361.950 316.050 366.000 ;
        RECT 326.400 364.050 327.450 388.950 ;
        RECT 380.400 388.050 381.450 391.950 ;
        RECT 370.950 385.950 373.050 388.050 ;
        RECT 379.950 385.950 382.050 388.050 ;
        RECT 371.400 382.050 372.450 385.950 ;
        RECT 370.950 379.950 373.050 382.050 ;
        RECT 373.950 376.950 376.050 379.050 ;
        RECT 374.400 373.200 375.450 376.950 ;
        RECT 331.950 370.950 334.050 373.050 ;
        RECT 337.950 371.100 340.050 373.200 ;
        RECT 373.950 371.100 376.050 373.200 ;
        RECT 332.400 370.350 333.600 370.950 ;
        RECT 338.400 370.350 339.600 371.100 ;
        RECT 374.400 370.350 375.600 371.100 ;
        RECT 385.950 370.950 388.050 373.050 ;
        RECT 331.950 367.950 334.050 370.050 ;
        RECT 334.950 367.950 337.050 370.050 ;
        RECT 337.950 367.950 340.050 370.050 ;
        RECT 352.950 367.950 355.050 370.050 ;
        RECT 355.950 367.950 358.050 370.050 ;
        RECT 358.950 367.950 361.050 370.050 ;
        RECT 367.950 367.950 370.050 370.050 ;
        RECT 374.100 367.950 376.200 370.050 ;
        RECT 377.400 367.950 379.500 370.050 ;
        RECT 382.800 367.950 384.900 370.050 ;
        RECT 335.400 365.400 336.600 367.650 ;
        RECT 356.400 365.400 357.600 367.650 ;
        RECT 325.950 361.950 328.050 364.050 ;
        RECT 335.400 346.050 336.450 365.400 ;
        RECT 340.950 349.950 343.050 352.050 ;
        RECT 334.950 343.950 337.050 346.050 ;
        RECT 305.400 338.400 309.450 339.450 ;
        RECT 277.950 331.800 280.050 333.900 ;
        RECT 286.950 331.950 289.050 334.050 ;
        RECT 269.400 305.400 273.450 306.450 ;
        RECT 215.400 293.400 219.450 294.450 ;
        RECT 211.950 280.950 214.050 283.050 ;
        RECT 215.400 280.050 216.450 293.400 ;
        RECT 220.950 289.950 223.050 292.050 ;
        RECT 223.950 289.950 226.050 292.050 ;
        RECT 226.950 289.950 229.050 292.050 ;
        RECT 224.400 287.400 225.600 289.650 ;
        RECT 214.950 277.950 217.050 280.050 ;
        RECT 220.950 277.950 223.050 280.050 ;
        RECT 214.950 271.950 217.050 274.050 ;
        RECT 205.950 268.950 208.050 271.050 ;
        RECT 202.950 265.950 205.050 268.050 ;
        RECT 208.950 265.950 211.050 268.050 ;
        RECT 184.950 250.950 187.050 255.000 ;
        RECT 190.950 253.800 193.050 255.900 ;
        RECT 199.950 253.800 202.050 255.900 ;
        RECT 203.400 250.050 204.450 265.950 ;
        RECT 209.400 262.200 210.450 265.950 ;
        RECT 208.950 260.100 211.050 262.200 ;
        RECT 215.400 261.600 216.450 271.950 ;
        RECT 209.400 259.350 210.600 260.100 ;
        RECT 215.400 259.350 216.600 261.600 ;
        RECT 208.950 256.950 211.050 259.050 ;
        RECT 211.950 256.950 214.050 259.050 ;
        RECT 214.950 256.950 217.050 259.050 ;
        RECT 212.400 255.900 213.600 256.650 ;
        RECT 211.950 253.800 214.050 255.900 ;
        RECT 221.400 253.050 222.450 277.950 ;
        RECT 220.950 250.950 223.050 253.050 ;
        RECT 202.950 247.950 205.050 250.050 ;
        RECT 203.400 223.050 204.450 247.950 ;
        RECT 224.400 229.050 225.450 287.400 ;
        RECT 233.400 268.050 234.450 304.950 ;
        RECT 241.950 298.950 244.050 301.050 ;
        RECT 242.400 294.600 243.450 298.950 ;
        RECT 242.400 292.350 243.600 294.600 ;
        RECT 241.950 289.950 244.050 292.050 ;
        RECT 244.950 289.950 247.050 292.050 ;
        RECT 251.400 288.900 252.450 304.950 ;
        RECT 253.950 295.950 256.050 298.050 ;
        RECT 250.950 286.800 253.050 288.900 ;
        RECT 254.400 277.050 255.450 295.950 ;
        RECT 262.950 294.000 265.050 298.050 ;
        RECT 263.400 292.350 264.600 294.000 ;
        RECT 259.950 289.950 262.050 292.050 ;
        RECT 262.950 289.950 265.050 292.050 ;
        RECT 265.950 289.950 268.050 292.050 ;
        RECT 260.400 288.900 261.600 289.650 ;
        RECT 266.400 288.900 267.600 289.650 ;
        RECT 272.400 288.900 273.450 305.400 ;
        RECT 290.400 304.050 291.450 337.950 ;
        RECT 299.400 337.350 300.600 338.100 ;
        RECT 295.950 334.950 298.050 337.050 ;
        RECT 298.950 334.950 301.050 337.050 ;
        RECT 301.950 334.950 304.050 337.050 ;
        RECT 302.400 333.900 303.600 334.650 ;
        RECT 308.400 333.900 309.450 338.400 ;
        RECT 310.950 337.950 313.050 340.050 ;
        RECT 337.950 337.950 340.050 340.050 ;
        RECT 301.950 331.800 304.050 333.900 ;
        RECT 307.950 331.800 310.050 333.900 ;
        RECT 298.950 304.950 301.050 307.050 ;
        RECT 289.950 301.950 292.050 304.050 ;
        RECT 289.950 298.800 292.050 300.900 ;
        RECT 277.950 293.100 280.050 295.200 ;
        RECT 283.950 293.100 286.050 295.200 ;
        RECT 290.400 294.600 291.450 298.800 ;
        RECT 259.950 286.800 262.050 288.900 ;
        RECT 265.950 286.800 268.050 288.900 ;
        RECT 271.950 286.800 274.050 288.900 ;
        RECT 278.400 283.050 279.450 293.100 ;
        RECT 284.400 292.350 285.600 293.100 ;
        RECT 290.400 292.350 291.600 294.600 ;
        RECT 283.950 289.950 286.050 292.050 ;
        RECT 286.950 289.950 289.050 292.050 ;
        RECT 289.950 289.950 292.050 292.050 ;
        RECT 292.950 289.950 295.050 292.050 ;
        RECT 287.400 287.400 288.600 289.650 ;
        RECT 293.400 288.000 294.600 289.650 ;
        RECT 268.950 280.950 271.050 283.050 ;
        RECT 277.950 280.950 280.050 283.050 ;
        RECT 253.950 274.950 256.050 277.050 ;
        RECT 241.950 268.950 244.050 271.050 ;
        RECT 232.950 265.950 235.050 268.050 ;
        RECT 232.950 260.100 235.050 262.200 ;
        RECT 233.400 259.350 234.600 260.100 ;
        RECT 232.950 256.950 235.050 259.050 ;
        RECT 235.950 256.950 238.050 259.050 ;
        RECT 236.400 254.400 237.600 256.650 ;
        RECT 242.400 256.050 243.450 268.950 ;
        RECT 250.950 256.950 253.050 259.050 ;
        RECT 253.950 256.950 256.050 259.050 ;
        RECT 232.950 250.950 235.050 253.050 ;
        RECT 211.950 226.950 214.050 229.050 ;
        RECT 223.950 226.950 226.050 229.050 ;
        RECT 178.950 220.950 181.050 223.050 ;
        RECT 184.950 220.950 187.050 223.050 ;
        RECT 202.950 220.950 205.050 223.050 ;
        RECT 208.950 220.950 211.050 223.050 ;
        RECT 173.400 218.400 177.450 219.450 ;
        RECT 173.400 217.200 174.450 218.400 ;
        RECT 172.950 215.100 175.050 217.200 ;
        RECT 178.950 216.000 181.050 219.900 ;
        RECT 173.400 214.350 174.600 215.100 ;
        RECT 179.400 214.350 180.600 216.000 ;
        RECT 169.950 211.950 172.050 214.050 ;
        RECT 172.950 211.950 175.050 214.050 ;
        RECT 175.950 211.950 178.050 214.050 ;
        RECT 178.950 211.950 181.050 214.050 ;
        RECT 170.400 209.400 171.600 211.650 ;
        RECT 176.400 210.900 177.600 211.650 ;
        RECT 185.400 210.900 186.450 220.950 ;
        RECT 193.950 215.100 196.050 217.200 ;
        RECT 199.950 215.100 202.050 220.050 ;
        RECT 194.400 214.350 195.600 215.100 ;
        RECT 200.400 214.350 201.600 215.100 ;
        RECT 193.950 211.950 196.050 214.050 ;
        RECT 196.950 211.950 199.050 214.050 ;
        RECT 199.950 211.950 202.050 214.050 ;
        RECT 202.950 211.950 205.050 214.050 ;
        RECT 197.400 210.900 198.600 211.650 ;
        RECT 170.400 163.050 171.450 209.400 ;
        RECT 175.950 208.800 178.050 210.900 ;
        RECT 184.950 208.800 187.050 210.900 ;
        RECT 196.950 208.800 199.050 210.900 ;
        RECT 203.400 209.400 204.600 211.650 ;
        RECT 199.950 202.950 202.050 205.050 ;
        RECT 190.950 190.950 193.050 193.050 ;
        RECT 178.950 183.000 181.050 187.050 ;
        RECT 179.400 181.350 180.600 183.000 ;
        RECT 184.950 182.100 187.050 184.200 ;
        RECT 185.400 181.350 186.600 182.100 ;
        RECT 178.950 178.950 181.050 181.050 ;
        RECT 181.950 178.950 184.050 181.050 ;
        RECT 184.950 178.950 187.050 181.050 ;
        RECT 182.400 177.900 183.600 178.650 ;
        RECT 191.400 178.050 192.450 190.950 ;
        RECT 193.950 187.950 196.050 190.050 ;
        RECT 181.950 175.800 184.050 177.900 ;
        RECT 190.950 175.950 193.050 178.050 ;
        RECT 169.950 160.950 172.050 163.050 ;
        RECT 194.400 142.200 195.450 187.950 ;
        RECT 200.400 184.200 201.450 202.950 ;
        RECT 203.400 190.050 204.450 209.400 ;
        RECT 202.950 187.950 205.050 190.050 ;
        RECT 209.400 187.050 210.450 220.950 ;
        RECT 212.400 205.050 213.450 226.950 ;
        RECT 220.950 220.950 223.050 223.050 ;
        RECT 221.400 216.600 222.450 220.950 ;
        RECT 221.400 214.350 222.600 216.600 ;
        RECT 226.950 216.000 229.050 220.050 ;
        RECT 227.400 214.350 228.600 216.000 ;
        RECT 217.950 211.950 220.050 214.050 ;
        RECT 220.950 211.950 223.050 214.050 ;
        RECT 223.950 211.950 226.050 214.050 ;
        RECT 226.950 211.950 229.050 214.050 ;
        RECT 218.400 209.400 219.600 211.650 ;
        RECT 224.400 210.900 225.600 211.650 ;
        RECT 218.400 205.050 219.450 209.400 ;
        RECT 223.950 208.800 226.050 210.900 ;
        RECT 233.400 205.050 234.450 250.950 ;
        RECT 236.400 220.050 237.450 254.400 ;
        RECT 241.950 253.950 244.050 256.050 ;
        RECT 251.400 255.900 252.600 256.650 ;
        RECT 250.950 253.800 253.050 255.900 ;
        RECT 269.400 250.050 270.450 280.950 ;
        RECT 277.950 274.950 280.050 277.050 ;
        RECT 278.400 261.600 279.450 274.950 ;
        RECT 287.400 268.050 288.450 287.400 ;
        RECT 292.950 283.950 295.050 288.000 ;
        RECT 299.400 286.050 300.450 304.950 ;
        RECT 304.950 301.950 307.050 304.050 ;
        RECT 305.400 288.900 306.450 301.950 ;
        RECT 311.400 301.050 312.450 337.950 ;
        RECT 316.950 334.950 319.050 337.050 ;
        RECT 319.950 334.950 322.050 337.050 ;
        RECT 322.950 334.950 325.050 337.050 ;
        RECT 325.950 334.950 328.050 337.050 ;
        RECT 328.950 334.950 331.050 337.050 ;
        RECT 317.400 333.900 318.600 334.650 ;
        RECT 316.950 331.800 319.050 333.900 ;
        RECT 323.400 332.400 324.600 334.650 ;
        RECT 323.400 325.050 324.450 332.400 ;
        RECT 338.400 325.050 339.450 337.950 ;
        RECT 322.950 322.950 325.050 325.050 ;
        RECT 337.950 322.950 340.050 325.050 ;
        RECT 341.400 307.050 342.450 349.950 ;
        RECT 356.400 340.200 357.450 365.400 ;
        RECT 368.400 364.050 369.450 367.950 ;
        RECT 386.400 364.050 387.450 370.950 ;
        RECT 392.400 366.900 393.450 436.950 ;
        RECT 398.400 433.050 399.450 461.400 ;
        RECT 400.950 454.950 403.050 457.050 ;
        RECT 406.950 454.950 412.050 457.050 ;
        RECT 401.400 451.050 402.450 454.950 ;
        RECT 400.950 448.950 403.050 451.050 ;
        RECT 403.950 450.000 406.050 454.050 ;
        RECT 409.950 450.000 412.050 453.900 ;
        RECT 404.400 448.350 405.600 450.000 ;
        RECT 410.400 448.350 411.600 450.000 ;
        RECT 403.950 445.950 406.050 448.050 ;
        RECT 406.950 445.950 409.050 448.050 ;
        RECT 409.950 445.950 412.050 448.050 ;
        RECT 412.950 445.950 415.050 448.050 ;
        RECT 400.950 442.950 403.050 445.050 ;
        RECT 407.400 444.900 408.600 445.650 ;
        RECT 397.950 430.950 400.050 433.050 ;
        RECT 401.400 430.050 402.450 442.950 ;
        RECT 406.950 442.800 409.050 444.900 ;
        RECT 413.400 443.400 414.600 445.650 ;
        RECT 419.400 444.450 420.450 472.950 ;
        RECT 421.950 466.950 424.050 469.050 ;
        RECT 416.400 443.400 420.450 444.450 ;
        RECT 413.400 433.050 414.450 443.400 ;
        RECT 412.950 430.950 415.050 433.050 ;
        RECT 400.950 427.950 403.050 430.050 ;
        RECT 403.950 424.950 406.050 427.050 ;
        RECT 404.400 417.600 405.450 424.950 ;
        RECT 404.400 415.350 405.600 417.600 ;
        RECT 409.950 417.000 412.050 421.050 ;
        RECT 410.400 415.350 411.600 417.000 ;
        RECT 400.950 412.950 403.050 415.050 ;
        RECT 403.950 412.950 406.050 415.050 ;
        RECT 406.950 412.950 409.050 415.050 ;
        RECT 409.950 412.950 412.050 415.050 ;
        RECT 401.400 411.000 402.600 412.650 ;
        RECT 407.400 411.900 408.600 412.650 ;
        RECT 400.950 406.950 403.050 411.000 ;
        RECT 406.950 406.950 409.050 411.900 ;
        RECT 401.400 403.050 402.450 406.950 ;
        RECT 400.950 400.950 403.050 403.050 ;
        RECT 403.950 397.950 406.050 400.050 ;
        RECT 397.950 379.950 400.050 382.050 ;
        RECT 398.400 372.600 399.450 379.950 ;
        RECT 404.400 372.600 405.450 397.950 ;
        RECT 409.950 382.950 412.050 385.050 ;
        RECT 398.400 370.350 399.600 372.600 ;
        RECT 404.400 370.350 405.600 372.600 ;
        RECT 397.950 367.950 400.050 370.050 ;
        RECT 400.950 367.950 403.050 370.050 ;
        RECT 403.950 367.950 406.050 370.050 ;
        RECT 391.950 364.800 394.050 366.900 ;
        RECT 401.400 365.400 402.600 367.650 ;
        RECT 367.950 361.950 370.050 364.050 ;
        RECT 385.950 361.950 388.050 364.050 ;
        RECT 401.400 349.050 402.450 365.400 ;
        RECT 410.400 355.050 411.450 382.950 ;
        RECT 416.400 363.450 417.450 443.400 ;
        RECT 422.400 430.050 423.450 466.950 ;
        RECT 425.400 451.050 426.450 478.950 ;
        RECT 442.950 457.950 445.050 460.050 ;
        RECT 430.950 454.950 433.050 457.050 ;
        RECT 436.950 454.950 439.050 457.050 ;
        RECT 431.400 451.200 432.450 454.950 ;
        RECT 424.950 448.950 427.050 451.050 ;
        RECT 430.950 449.100 433.050 451.200 ;
        RECT 437.400 450.600 438.450 454.950 ;
        RECT 431.400 448.350 432.600 449.100 ;
        RECT 437.400 448.350 438.600 450.600 ;
        RECT 427.950 445.950 430.050 448.050 ;
        RECT 430.950 445.950 433.050 448.050 ;
        RECT 433.950 445.950 436.050 448.050 ;
        RECT 436.950 445.950 439.050 448.050 ;
        RECT 424.800 442.950 426.900 445.050 ;
        RECT 428.400 444.900 429.600 445.650 ;
        RECT 425.400 439.050 426.450 442.950 ;
        RECT 427.950 442.800 430.050 444.900 ;
        RECT 434.400 443.400 435.600 445.650 ;
        RECT 424.950 436.950 427.050 439.050 ;
        RECT 421.950 427.950 424.050 430.050 ;
        RECT 418.950 424.950 421.050 427.050 ;
        RECT 419.400 411.900 420.450 424.950 ;
        RECT 418.950 409.800 421.050 411.900 ;
        RECT 422.400 376.050 423.450 427.950 ;
        RECT 428.400 421.050 429.450 442.800 ;
        RECT 434.400 421.050 435.450 443.400 ;
        RECT 436.950 427.950 439.050 430.050 ;
        RECT 427.950 418.950 430.050 421.050 ;
        RECT 433.950 418.950 436.050 421.050 ;
        RECT 430.950 416.100 433.050 418.200 ;
        RECT 437.400 417.600 438.450 427.950 ;
        RECT 431.400 415.350 432.600 416.100 ;
        RECT 437.400 415.350 438.600 417.600 ;
        RECT 427.950 412.950 430.050 415.050 ;
        RECT 430.950 412.950 433.050 415.050 ;
        RECT 433.950 412.950 436.050 415.050 ;
        RECT 436.950 412.950 439.050 415.050 ;
        RECT 428.400 411.900 429.600 412.650 ;
        RECT 427.950 409.800 430.050 411.900 ;
        RECT 434.400 410.400 435.600 412.650 ;
        RECT 434.400 403.050 435.450 410.400 ;
        RECT 443.400 406.050 444.450 457.950 ;
        RECT 442.950 403.950 445.050 406.050 ;
        RECT 433.950 400.950 436.050 403.050 ;
        RECT 446.400 400.050 447.450 493.950 ;
        RECT 449.400 475.050 450.450 511.950 ;
        RECT 452.400 502.050 453.450 523.950 ;
        RECT 455.400 517.050 456.450 541.950 ;
        RECT 457.950 532.950 460.050 535.050 ;
        RECT 482.400 534.450 483.450 550.950 ;
        RECT 518.400 550.050 519.450 565.800 ;
        RECT 524.400 562.050 525.450 583.950 ;
        RECT 523.950 559.950 526.050 562.050 ;
        RECT 517.950 547.950 520.050 550.050 ;
        RECT 514.950 543.450 517.050 544.050 ;
        RECT 514.950 542.400 522.450 543.450 ;
        RECT 514.950 541.950 517.050 542.400 ;
        RECT 517.950 538.950 520.050 541.050 ;
        RECT 518.400 535.050 519.450 538.950 ;
        RECT 521.400 538.050 522.450 542.400 ;
        RECT 520.950 535.950 523.050 538.050 ;
        RECT 479.400 533.400 483.450 534.450 ;
        RECT 458.400 520.050 459.450 532.950 ;
        RECT 469.950 531.450 472.050 532.200 ;
        RECT 475.950 531.450 478.050 532.050 ;
        RECT 469.950 530.400 478.050 531.450 ;
        RECT 469.950 530.100 472.050 530.400 ;
        RECT 475.950 529.950 478.050 530.400 ;
        RECT 463.950 527.100 466.050 529.200 ;
        RECT 479.400 529.050 480.450 533.400 ;
        RECT 487.950 532.950 490.050 535.050 ;
        RECT 502.950 532.950 505.050 535.050 ;
        RECT 517.950 532.950 520.050 535.050 ;
        RECT 464.400 526.350 465.600 527.100 ;
        RECT 469.950 526.950 472.050 529.050 ;
        RECT 478.950 526.950 481.050 529.050 ;
        RECT 488.400 528.600 489.450 532.950 ;
        RECT 470.400 526.350 471.600 526.950 ;
        RECT 488.400 526.350 489.600 528.600 ;
        RECT 493.950 528.000 496.050 532.050 ;
        RECT 494.400 526.350 495.600 528.000 ;
        RECT 463.950 523.950 466.050 526.050 ;
        RECT 466.950 523.950 469.050 526.050 ;
        RECT 469.950 523.950 472.050 526.050 ;
        RECT 472.950 523.950 475.050 526.050 ;
        RECT 487.950 523.950 490.050 526.050 ;
        RECT 490.950 523.950 493.050 526.050 ;
        RECT 493.950 523.950 496.050 526.050 ;
        RECT 496.950 523.950 499.050 526.050 ;
        RECT 467.400 521.400 468.600 523.650 ;
        RECT 473.400 522.900 474.600 523.650 ;
        RECT 491.400 522.900 492.600 523.650 ;
        RECT 457.950 517.950 460.050 520.050 ;
        RECT 454.950 514.950 457.050 517.050 ;
        RECT 454.950 502.950 457.050 505.050 ;
        RECT 451.950 499.950 454.050 502.050 ;
        RECT 455.400 495.600 456.450 502.950 ;
        RECT 467.400 499.050 468.450 521.400 ;
        RECT 472.950 520.800 475.050 522.900 ;
        RECT 490.950 520.800 493.050 522.900 ;
        RECT 497.400 521.400 498.600 523.650 ;
        RECT 497.400 511.050 498.450 521.400 ;
        RECT 499.950 520.950 502.050 523.050 ;
        RECT 496.950 508.950 499.050 511.050 ;
        RECT 500.400 508.050 501.450 520.950 ;
        RECT 503.400 520.050 504.450 532.950 ;
        RECT 511.950 527.100 514.050 529.200 ;
        RECT 518.400 528.600 519.450 532.950 ;
        RECT 512.400 526.350 513.600 527.100 ;
        RECT 518.400 526.350 519.600 528.600 ;
        RECT 511.950 523.950 514.050 526.050 ;
        RECT 514.950 523.950 517.050 526.050 ;
        RECT 517.950 523.950 520.050 526.050 ;
        RECT 520.950 523.950 523.050 526.050 ;
        RECT 515.400 521.400 516.600 523.650 ;
        RECT 521.400 522.900 522.600 523.650 ;
        RECT 502.950 517.950 505.050 520.050 ;
        RECT 515.400 519.450 516.450 521.400 ;
        RECT 520.950 520.800 523.050 522.900 ;
        RECT 512.400 518.400 516.450 519.450 ;
        RECT 505.950 511.950 508.050 514.050 ;
        RECT 478.950 505.950 481.050 508.050 ;
        RECT 499.950 505.950 502.050 508.050 ;
        RECT 479.400 502.050 480.450 505.950 ;
        RECT 469.950 499.950 472.050 502.050 ;
        RECT 478.800 499.950 480.900 502.050 ;
        RECT 466.950 496.950 469.050 499.050 ;
        RECT 455.400 493.350 456.600 495.600 ;
        RECT 460.950 494.100 463.050 496.200 ;
        RECT 461.400 493.350 462.600 494.100 ;
        RECT 454.950 490.950 457.050 493.050 ;
        RECT 457.950 490.950 460.050 493.050 ;
        RECT 460.950 490.950 463.050 493.050 ;
        RECT 463.950 490.950 466.050 493.050 ;
        RECT 458.400 488.400 459.600 490.650 ;
        RECT 464.400 489.900 465.600 490.650 ;
        RECT 470.400 489.900 471.450 499.950 ;
        RECT 475.950 494.100 478.050 496.200 ;
        RECT 458.400 481.050 459.450 488.400 ;
        RECT 463.950 487.800 466.050 489.900 ;
        RECT 469.950 487.800 472.050 489.900 ;
        RECT 476.400 484.050 477.450 494.100 ;
        RECT 479.400 489.450 480.450 499.950 ;
        RECT 487.950 494.100 490.050 496.200 ;
        RECT 488.400 493.350 489.600 494.100 ;
        RECT 482.100 490.950 484.200 493.050 ;
        RECT 487.500 490.950 489.600 493.050 ;
        RECT 490.800 490.950 492.900 493.050 ;
        RECT 482.400 489.450 483.600 490.650 ;
        RECT 479.400 488.400 483.600 489.450 ;
        RECT 491.400 488.400 492.600 490.650 ;
        RECT 475.950 481.950 478.050 484.050 ;
        RECT 457.950 478.950 460.050 481.050 ;
        RECT 472.950 478.950 475.050 481.050 ;
        RECT 448.950 472.950 451.050 475.050 ;
        RECT 473.400 472.050 474.450 478.950 ;
        RECT 472.950 469.950 475.050 472.050 ;
        RECT 475.950 466.950 478.050 469.050 ;
        RECT 460.950 457.950 463.050 460.050 ;
        RECT 454.950 449.100 457.050 451.200 ;
        RECT 461.400 450.600 462.450 457.950 ;
        RECT 472.950 454.950 475.050 457.050 ;
        RECT 466.950 451.950 469.050 454.050 ;
        RECT 455.400 448.350 456.600 449.100 ;
        RECT 461.400 448.350 462.600 450.600 ;
        RECT 451.950 445.950 454.050 448.050 ;
        RECT 454.950 445.950 457.050 448.050 ;
        RECT 457.950 445.950 460.050 448.050 ;
        RECT 460.950 445.950 463.050 448.050 ;
        RECT 452.400 444.900 453.600 445.650 ;
        RECT 458.400 444.900 459.600 445.650 ;
        RECT 467.400 445.050 468.450 451.950 ;
        RECT 473.400 451.050 474.450 454.950 ;
        RECT 472.950 448.950 475.050 451.050 ;
        RECT 476.400 450.600 477.450 466.950 ;
        RECT 481.950 453.450 484.050 454.200 ;
        RECT 487.950 453.450 490.050 454.050 ;
        RECT 481.950 452.400 490.050 453.450 ;
        RECT 481.950 452.100 484.050 452.400 ;
        RECT 487.950 451.950 490.050 452.400 ;
        RECT 491.400 451.050 492.450 488.400 ;
        RECT 493.950 466.950 496.050 469.050 ;
        RECT 476.400 448.350 477.600 450.600 ;
        RECT 481.950 448.950 484.050 451.050 ;
        RECT 490.950 448.950 493.050 451.050 ;
        RECT 482.400 448.350 483.600 448.950 ;
        RECT 475.950 445.950 478.050 448.050 ;
        RECT 478.950 445.950 481.050 448.050 ;
        RECT 481.950 445.950 484.050 448.050 ;
        RECT 484.950 445.950 487.050 448.050 ;
        RECT 451.950 442.800 454.050 444.900 ;
        RECT 457.950 442.800 460.050 444.900 ;
        RECT 466.950 442.950 469.050 445.050 ;
        RECT 479.400 444.900 480.600 445.650 ;
        RECT 485.400 444.900 486.600 445.650 ;
        RECT 478.950 442.800 481.050 444.900 ;
        RECT 484.950 442.800 487.050 444.900 ;
        RECT 466.950 436.950 469.050 439.050 ;
        RECT 467.400 433.050 468.450 436.950 ;
        RECT 494.400 433.050 495.450 466.950 ;
        RECT 506.400 460.050 507.450 511.950 ;
        RECT 512.400 499.050 513.450 518.400 ;
        RECT 523.950 517.950 526.050 520.050 ;
        RECT 511.950 496.950 514.050 499.050 ;
        RECT 520.950 493.950 523.050 496.050 ;
        RECT 509.100 490.950 511.200 493.050 ;
        RECT 514.500 490.950 516.600 493.050 ;
        RECT 517.800 490.950 519.900 493.050 ;
        RECT 518.400 489.900 519.600 490.650 ;
        RECT 517.950 487.800 520.050 489.900 ;
        RECT 505.950 457.950 508.050 460.050 ;
        RECT 499.950 449.100 502.050 451.200 ;
        RECT 505.950 450.000 508.050 454.050 ;
        RECT 500.400 448.350 501.600 449.100 ;
        RECT 506.400 448.350 507.600 450.000 ;
        RECT 514.950 448.950 517.050 451.050 ;
        RECT 521.400 450.450 522.450 493.950 ;
        RECT 524.400 490.050 525.450 517.950 ;
        RECT 527.400 496.050 528.450 619.950 ;
        RECT 541.950 615.450 544.050 616.050 ;
        RECT 536.400 614.400 544.050 615.450 ;
        RECT 536.400 610.200 537.450 614.400 ;
        RECT 541.950 613.950 544.050 614.400 ;
        RECT 540.000 612.900 543.000 613.050 ;
        RECT 538.950 610.950 544.050 612.900 ;
        RECT 547.950 610.950 553.050 613.050 ;
        RECT 538.950 610.800 541.050 610.950 ;
        RECT 541.950 610.800 544.050 610.950 ;
        RECT 535.950 608.100 538.050 610.200 ;
        RECT 554.400 610.050 555.450 619.950 ;
        RECT 568.950 616.950 571.050 619.050 ;
        RECT 559.950 613.950 562.050 616.050 ;
        RECT 535.950 604.950 538.050 607.050 ;
        RECT 541.950 606.000 544.050 609.900 ;
        RECT 553.950 609.450 556.050 610.050 ;
        RECT 551.400 608.400 556.050 609.450 ;
        RECT 536.400 604.350 537.600 604.950 ;
        RECT 542.400 604.350 543.600 606.000 ;
        RECT 532.950 601.950 535.050 604.050 ;
        RECT 535.950 601.950 538.050 604.050 ;
        RECT 538.950 601.950 541.050 604.050 ;
        RECT 541.950 601.950 544.050 604.050 ;
        RECT 533.400 599.400 534.600 601.650 ;
        RECT 539.400 600.000 540.600 601.650 ;
        RECT 533.400 595.050 534.450 599.400 ;
        RECT 538.950 595.950 541.050 600.000 ;
        RECT 547.800 598.950 549.900 601.050 ;
        RECT 551.400 600.900 552.450 608.400 ;
        RECT 553.950 607.950 556.050 608.400 ;
        RECT 560.400 606.600 561.450 613.950 ;
        RECT 560.400 604.350 561.600 606.600 ;
        RECT 556.950 601.950 559.050 604.050 ;
        RECT 559.950 601.950 562.050 604.050 ;
        RECT 562.950 601.950 565.050 604.050 ;
        RECT 557.400 600.900 558.600 601.650 ;
        RECT 532.950 592.950 535.050 595.050 ;
        RECT 533.400 577.050 534.450 592.950 ;
        RECT 532.950 574.950 535.050 577.050 ;
        RECT 529.950 573.600 534.000 574.050 ;
        RECT 529.950 571.950 534.600 573.600 ;
        RECT 538.950 572.100 541.050 574.200 ;
        RECT 533.400 571.350 534.600 571.950 ;
        RECT 539.400 571.350 540.600 572.100 ;
        RECT 532.950 568.950 535.050 571.050 ;
        RECT 535.950 568.950 538.050 571.050 ;
        RECT 538.950 568.950 541.050 571.050 ;
        RECT 541.950 568.950 544.050 571.050 ;
        RECT 529.950 565.800 532.050 567.900 ;
        RECT 536.400 566.400 537.600 568.650 ;
        RECT 542.400 567.900 543.600 568.650 ;
        RECT 530.400 520.050 531.450 565.800 ;
        RECT 536.400 564.450 537.450 566.400 ;
        RECT 541.950 565.800 544.050 567.900 ;
        RECT 533.400 563.400 537.450 564.450 ;
        RECT 533.400 559.050 534.450 563.400 ;
        RECT 548.400 562.050 549.450 598.950 ;
        RECT 550.950 598.800 553.050 600.900 ;
        RECT 556.950 598.800 559.050 600.900 ;
        RECT 563.400 599.400 564.600 601.650 ;
        RECT 563.400 592.050 564.450 599.400 ;
        RECT 569.400 598.050 570.450 616.950 ;
        RECT 568.950 595.950 571.050 598.050 ;
        RECT 562.950 589.950 565.050 592.050 ;
        RECT 572.400 591.450 573.450 620.400 ;
        RECT 583.950 616.950 586.050 619.050 ;
        RECT 589.950 616.950 592.050 619.050 ;
        RECT 574.950 610.950 577.050 613.050 ;
        RECT 575.400 600.900 576.450 610.950 ;
        RECT 584.400 610.050 585.450 616.950 ;
        RECT 577.950 606.000 580.050 610.050 ;
        RECT 583.950 607.950 586.050 610.050 ;
        RECT 578.400 604.350 579.600 606.000 ;
        RECT 586.950 605.100 589.050 607.200 ;
        RECT 587.400 604.350 588.600 605.100 ;
        RECT 578.100 601.950 580.200 604.050 ;
        RECT 583.500 601.950 585.600 604.050 ;
        RECT 586.800 601.950 588.900 604.050 ;
        RECT 574.950 598.800 577.050 600.900 ;
        RECT 584.400 599.400 585.600 601.650 ;
        RECT 584.400 592.050 585.450 599.400 ;
        RECT 569.400 590.400 573.450 591.450 ;
        RECT 569.400 583.050 570.450 590.400 ;
        RECT 583.950 589.950 586.050 592.050 ;
        RECT 571.950 586.950 574.050 589.050 ;
        RECT 550.950 580.950 553.050 583.050 ;
        RECT 568.950 580.950 571.050 583.050 ;
        RECT 547.950 559.950 550.050 562.050 ;
        RECT 532.950 556.950 535.050 559.050 ;
        RECT 533.400 529.050 534.450 556.950 ;
        RECT 541.950 553.950 544.050 556.050 ;
        RECT 542.400 538.050 543.450 553.950 ;
        RECT 544.950 538.950 547.050 541.050 ;
        RECT 538.800 535.950 540.900 538.050 ;
        RECT 541.950 535.950 544.050 538.050 ;
        RECT 539.400 532.050 540.450 535.950 ;
        RECT 545.400 535.050 546.450 538.950 ;
        RECT 544.950 532.950 547.050 535.050 ;
        RECT 539.400 530.400 544.050 532.050 ;
        RECT 540.000 529.950 544.050 530.400 ;
        RECT 532.950 526.950 535.050 529.050 ;
        RECT 538.950 527.100 541.050 529.200 ;
        RECT 551.400 529.050 552.450 580.950 ;
        RECT 554.400 578.400 567.450 579.450 ;
        RECT 554.400 574.050 555.450 578.400 ;
        RECT 553.950 571.950 556.050 574.050 ;
        RECT 556.950 573.000 559.050 577.050 ;
        RECT 562.950 573.000 565.050 577.050 ;
        RECT 566.400 576.450 567.450 578.400 ;
        RECT 566.400 576.000 570.450 576.450 ;
        RECT 566.400 575.400 571.050 576.000 ;
        RECT 557.400 571.350 558.600 573.000 ;
        RECT 563.400 571.350 564.600 573.000 ;
        RECT 568.950 571.950 571.050 575.400 ;
        RECT 556.950 568.950 559.050 571.050 ;
        RECT 559.950 568.950 562.050 571.050 ;
        RECT 562.950 568.950 565.050 571.050 ;
        RECT 565.950 568.950 568.050 571.050 ;
        RECT 553.950 565.950 556.050 568.050 ;
        RECT 560.400 566.400 561.600 568.650 ;
        RECT 566.400 567.900 567.600 568.650 ;
        RECT 572.400 567.900 573.450 586.950 ;
        RECT 575.400 581.400 582.450 582.450 ;
        RECT 575.400 577.050 576.450 581.400 ;
        RECT 577.950 577.950 580.050 580.050 ;
        RECT 574.950 574.950 577.050 577.050 ;
        RECT 578.400 574.050 579.450 577.950 ;
        RECT 581.400 576.450 582.450 581.400 ;
        RECT 581.400 575.400 585.450 576.450 ;
        RECT 574.950 571.800 577.050 573.900 ;
        RECT 577.950 571.950 580.050 574.050 ;
        RECT 584.400 573.600 585.450 575.400 ;
        RECT 590.400 573.600 591.450 616.950 ;
        RECT 617.400 616.050 618.450 650.400 ;
        RECT 626.400 649.350 627.600 651.600 ;
        RECT 622.950 646.950 625.050 649.050 ;
        RECT 625.950 646.950 628.050 649.050 ;
        RECT 628.950 646.950 631.050 649.050 ;
        RECT 623.400 645.900 624.600 646.650 ;
        RECT 629.400 645.900 630.600 646.650 ;
        RECT 622.950 643.800 625.050 645.900 ;
        RECT 628.950 643.800 631.050 645.900 ;
        RECT 616.950 613.950 619.050 616.050 ;
        RECT 623.400 610.050 624.450 643.800 ;
        RECT 625.950 628.950 628.050 631.050 ;
        RECT 595.950 604.950 598.050 607.050 ;
        RECT 604.950 606.000 607.050 610.050 ;
        RECT 610.950 606.000 613.050 610.050 ;
        RECT 619.950 607.950 622.050 610.050 ;
        RECT 622.950 607.950 625.050 610.050 ;
        RECT 554.400 556.050 555.450 565.950 ;
        RECT 560.400 562.050 561.450 566.400 ;
        RECT 565.950 565.800 568.050 567.900 ;
        RECT 571.950 565.800 574.050 567.900 ;
        RECT 572.400 562.050 573.450 565.800 ;
        RECT 575.400 565.050 576.450 571.800 ;
        RECT 584.400 571.350 585.600 573.600 ;
        RECT 590.400 571.350 591.600 573.600 ;
        RECT 580.950 568.950 583.050 571.050 ;
        RECT 583.950 568.950 586.050 571.050 ;
        RECT 586.950 568.950 589.050 571.050 ;
        RECT 589.950 568.950 592.050 571.050 ;
        RECT 581.400 567.900 582.600 568.650 ;
        RECT 580.950 565.800 583.050 567.900 ;
        RECT 587.400 567.000 588.600 568.650 ;
        RECT 574.950 562.950 577.050 565.050 ;
        RECT 586.950 562.950 589.050 567.000 ;
        RECT 596.400 565.050 597.450 604.950 ;
        RECT 605.400 604.350 606.600 606.000 ;
        RECT 611.400 604.350 612.600 606.000 ;
        RECT 604.950 601.950 607.050 604.050 ;
        RECT 607.950 601.950 610.050 604.050 ;
        RECT 610.950 601.950 613.050 604.050 ;
        RECT 613.950 601.950 616.050 604.050 ;
        RECT 608.400 600.900 609.600 601.650 ;
        RECT 614.400 600.900 615.600 601.650 ;
        RECT 607.950 598.800 610.050 600.900 ;
        RECT 613.950 598.800 616.050 600.900 ;
        RECT 604.950 577.950 607.050 580.050 ;
        RECT 605.400 573.600 606.450 577.950 ;
        RECT 605.400 571.350 606.600 573.600 ;
        RECT 610.950 572.100 613.050 574.200 ;
        RECT 620.400 573.450 621.450 607.950 ;
        RECT 626.400 606.450 627.450 628.950 ;
        RECT 631.950 619.950 634.050 622.050 ;
        RECT 623.400 605.400 627.450 606.450 ;
        RECT 632.400 606.600 633.450 619.950 ;
        RECT 635.400 609.450 636.450 677.400 ;
        RECT 643.950 676.950 646.050 679.050 ;
        RECT 653.400 678.900 654.600 679.650 ;
        RECT 652.950 676.800 655.050 678.900 ;
        RECT 659.400 677.400 660.600 679.650 ;
        RECT 677.400 678.900 678.600 679.650 ;
        RECT 659.400 670.050 660.450 677.400 ;
        RECT 676.950 676.800 679.050 678.900 ;
        RECT 683.400 677.400 684.600 679.650 ;
        RECT 683.400 670.050 684.450 677.400 ;
        RECT 658.950 667.950 661.050 670.050 ;
        RECT 682.950 667.950 685.050 670.050 ;
        RECT 692.400 664.050 693.450 683.400 ;
        RECT 707.400 682.350 708.600 684.000 ;
        RECT 713.400 682.350 714.600 684.600 ;
        RECT 703.950 679.950 706.050 682.050 ;
        RECT 706.950 679.950 709.050 682.050 ;
        RECT 709.950 679.950 712.050 682.050 ;
        RECT 712.950 679.950 715.050 682.050 ;
        RECT 704.400 678.900 705.600 679.650 ;
        RECT 703.950 676.800 706.050 678.900 ;
        RECT 710.400 677.400 711.600 679.650 ;
        RECT 710.400 675.450 711.450 677.400 ;
        RECT 715.950 676.950 718.050 679.050 ;
        RECT 722.400 678.450 723.450 694.950 ;
        RECT 725.400 685.050 726.450 721.800 ;
        RECT 734.400 691.050 735.450 752.400 ;
        RECT 736.950 751.950 739.050 752.400 ;
        RECT 736.950 745.950 739.050 748.050 ;
        RECT 737.400 723.900 738.450 745.950 ;
        RECT 758.400 739.050 759.450 754.800 ;
        RECT 764.400 753.450 765.450 755.400 ;
        RECT 764.400 752.400 768.450 753.450 ;
        RECT 763.950 748.950 766.050 751.050 ;
        RECT 757.950 736.950 760.050 739.050 ;
        RECT 739.950 729.600 744.000 730.050 ;
        RECT 739.950 727.950 744.600 729.600 ;
        RECT 748.950 728.100 751.050 730.200 ;
        RECT 757.950 728.100 760.050 730.200 ;
        RECT 743.400 727.350 744.600 727.950 ;
        RECT 749.400 727.350 750.600 728.100 ;
        RECT 742.950 724.950 745.050 727.050 ;
        RECT 745.950 724.950 748.050 727.050 ;
        RECT 748.950 724.950 751.050 727.050 ;
        RECT 751.950 724.950 754.050 727.050 ;
        RECT 736.950 721.800 739.050 723.900 ;
        RECT 739.950 721.950 742.050 724.050 ;
        RECT 746.400 723.900 747.600 724.650 ;
        RECT 733.950 688.950 736.050 691.050 ;
        RECT 724.950 682.950 727.050 685.050 ;
        RECT 730.950 684.000 733.050 688.050 ;
        RECT 736.950 684.450 739.050 685.200 ;
        RECT 740.400 684.450 741.450 721.950 ;
        RECT 745.950 718.950 748.050 723.900 ;
        RECT 752.400 722.400 753.600 724.650 ;
        RECT 758.400 724.050 759.450 728.100 ;
        RECT 752.400 709.050 753.450 722.400 ;
        RECT 757.950 721.950 760.050 724.050 ;
        RECT 764.400 712.050 765.450 748.950 ;
        RECT 767.400 736.050 768.450 752.400 ;
        RECT 770.400 751.050 771.450 766.950 ;
        RECT 778.950 761.100 781.050 763.200 ;
        RECT 779.400 760.350 780.600 761.100 ;
        RECT 778.950 757.950 781.050 760.050 ;
        RECT 781.950 757.950 784.050 760.050 ;
        RECT 782.400 756.000 783.600 757.650 ;
        RECT 781.950 751.950 784.050 756.000 ;
        RECT 769.950 748.950 772.050 751.050 ;
        RECT 788.400 744.450 789.450 806.400 ;
        RECT 794.400 805.350 795.600 807.600 ;
        RECT 799.950 806.100 802.050 808.200 ;
        RECT 805.950 806.100 808.050 808.200 ;
        RECT 800.400 805.350 801.600 806.100 ;
        RECT 793.950 802.950 796.050 805.050 ;
        RECT 796.950 802.950 799.050 805.050 ;
        RECT 799.950 802.950 802.050 805.050 ;
        RECT 802.950 802.950 805.050 805.050 ;
        RECT 790.950 799.950 793.050 802.050 ;
        RECT 797.400 801.900 798.600 802.650 ;
        RECT 803.400 801.900 804.600 802.650 ;
        RECT 809.400 801.900 810.450 823.950 ;
        RECT 818.400 820.050 819.450 841.950 ;
        RECT 826.950 840.000 829.050 844.050 ;
        RECT 827.400 838.350 828.600 840.000 ;
        RECT 832.950 839.100 835.050 841.200 ;
        RECT 833.400 838.350 834.600 839.100 ;
        RECT 823.950 835.950 826.050 838.050 ;
        RECT 826.950 835.950 829.050 838.050 ;
        RECT 829.950 835.950 832.050 838.050 ;
        RECT 832.950 835.950 835.050 838.050 ;
        RECT 824.400 833.400 825.600 835.650 ;
        RECT 824.400 826.050 825.450 833.400 ;
        RECT 823.950 823.950 826.050 826.050 ;
        RECT 817.950 817.950 820.050 820.050 ;
        RECT 814.950 811.950 817.050 814.050 ;
        RECT 811.950 808.950 814.050 811.050 ;
        RECT 791.400 796.050 792.450 799.950 ;
        RECT 796.950 799.800 799.050 801.900 ;
        RECT 802.950 799.800 805.050 801.900 ;
        RECT 808.950 796.950 811.050 801.900 ;
        RECT 790.950 793.950 793.050 796.050 ;
        RECT 812.400 769.050 813.450 808.950 ;
        RECT 815.400 808.050 816.450 811.950 ;
        RECT 818.400 810.450 819.450 817.950 ;
        RECT 818.400 809.400 822.450 810.450 ;
        RECT 814.950 805.950 817.050 808.050 ;
        RECT 821.400 807.600 822.450 809.400 ;
        RECT 835.950 808.950 838.050 811.050 ;
        RECT 821.400 805.350 822.600 807.600 ;
        RECT 826.950 806.100 829.050 808.200 ;
        RECT 832.950 806.100 835.050 808.200 ;
        RECT 827.400 805.350 828.600 806.100 ;
        RECT 817.950 802.950 820.050 805.050 ;
        RECT 820.950 802.950 823.050 805.050 ;
        RECT 823.950 802.950 826.050 805.050 ;
        RECT 826.950 802.950 829.050 805.050 ;
        RECT 818.400 801.900 819.600 802.650 ;
        RECT 817.950 799.800 820.050 801.900 ;
        RECT 824.400 801.000 825.600 802.650 ;
        RECT 833.400 802.050 834.450 806.100 ;
        RECT 823.950 796.950 826.050 801.000 ;
        RECT 832.950 799.950 835.050 802.050 ;
        RECT 820.950 793.950 823.050 796.050 ;
        RECT 821.400 778.050 822.450 793.950 ;
        RECT 836.400 787.050 837.450 808.950 ;
        RECT 835.950 784.950 838.050 787.050 ;
        RECT 820.950 775.950 823.050 778.050 ;
        RECT 805.950 766.950 808.050 769.050 ;
        RECT 811.950 768.450 814.050 769.050 ;
        RECT 811.950 767.400 816.450 768.450 ;
        RECT 811.950 766.950 814.050 767.400 ;
        RECT 799.950 761.100 802.050 763.200 ;
        RECT 806.400 762.600 807.450 766.950 ;
        RECT 800.400 760.350 801.600 761.100 ;
        RECT 806.400 760.350 807.600 762.600 ;
        RECT 811.950 761.100 814.050 763.200 ;
        RECT 796.950 757.950 799.050 760.050 ;
        RECT 799.950 757.950 802.050 760.050 ;
        RECT 802.950 757.950 805.050 760.050 ;
        RECT 805.950 757.950 808.050 760.050 ;
        RECT 797.400 756.000 798.600 757.650 ;
        RECT 796.950 751.950 799.050 756.000 ;
        RECT 803.400 755.400 804.600 757.650 ;
        RECT 812.400 756.450 813.450 761.100 ;
        RECT 809.400 755.400 813.450 756.450 ;
        RECT 785.400 743.400 789.450 744.450 ;
        RECT 772.950 736.950 775.050 739.050 ;
        RECT 766.950 733.950 769.050 736.050 ;
        RECT 773.400 729.600 774.450 736.950 ;
        RECT 773.400 727.350 774.600 729.600 ;
        RECT 778.950 729.450 781.050 730.200 ;
        RECT 781.950 729.450 784.050 733.050 ;
        RECT 778.950 729.000 784.050 729.450 ;
        RECT 778.950 728.400 783.450 729.000 ;
        RECT 778.950 728.100 781.050 728.400 ;
        RECT 779.400 727.350 780.600 728.100 ;
        RECT 769.950 724.950 772.050 727.050 ;
        RECT 772.950 724.950 775.050 727.050 ;
        RECT 775.950 724.950 778.050 727.050 ;
        RECT 778.950 724.950 781.050 727.050 ;
        RECT 770.400 723.000 771.600 724.650 ;
        RECT 769.950 718.950 772.050 723.000 ;
        RECT 776.400 722.400 777.600 724.650 ;
        RECT 763.950 709.950 766.050 712.050 ;
        RECT 751.950 706.950 754.050 709.050 ;
        RECT 776.400 697.050 777.450 722.400 ;
        RECT 781.950 721.950 784.050 724.050 ;
        RECT 778.950 709.950 781.050 712.050 ;
        RECT 779.400 700.050 780.450 709.950 ;
        RECT 778.950 697.950 781.050 700.050 ;
        RECT 775.950 694.950 778.050 697.050 ;
        RECT 742.950 688.950 745.050 691.050 ;
        RECT 731.400 682.350 732.600 684.000 ;
        RECT 736.950 683.400 741.450 684.450 ;
        RECT 736.950 683.100 739.050 683.400 ;
        RECT 737.400 682.350 738.600 683.100 ;
        RECT 727.950 679.950 730.050 682.050 ;
        RECT 730.950 679.950 733.050 682.050 ;
        RECT 733.950 679.950 736.050 682.050 ;
        RECT 736.950 679.950 739.050 682.050 ;
        RECT 728.400 678.450 729.600 679.650 ;
        RECT 734.400 678.900 735.600 679.650 ;
        RECT 722.400 677.400 729.600 678.450 ;
        RECT 710.400 675.000 714.450 675.450 ;
        RECT 710.400 674.400 715.050 675.000 ;
        RECT 710.400 670.050 711.450 674.400 ;
        RECT 712.950 670.950 715.050 674.400 ;
        RECT 709.950 667.950 712.050 670.050 ;
        RECT 676.950 661.950 679.050 664.050 ;
        RECT 691.950 661.950 694.050 664.050 ;
        RECT 655.950 658.950 658.050 661.050 ;
        RECT 637.950 655.950 640.050 658.050 ;
        RECT 638.400 645.900 639.450 655.950 ;
        RECT 646.950 650.100 649.050 652.200 ;
        RECT 647.400 649.350 648.600 650.100 ;
        RECT 643.950 646.950 646.050 649.050 ;
        RECT 646.950 646.950 649.050 649.050 ;
        RECT 649.950 646.950 652.050 649.050 ;
        RECT 637.950 643.800 640.050 645.900 ;
        RECT 644.400 644.400 645.600 646.650 ;
        RECT 650.400 645.900 651.600 646.650 ;
        RECT 656.400 646.050 657.450 658.950 ;
        RECT 658.950 649.950 661.050 652.050 ;
        RECT 664.950 650.100 667.050 652.200 ;
        RECT 644.400 628.050 645.450 644.400 ;
        RECT 649.950 643.800 652.050 645.900 ;
        RECT 655.950 643.950 658.050 646.050 ;
        RECT 650.400 637.050 651.450 643.800 ;
        RECT 649.950 634.950 652.050 637.050 ;
        RECT 643.950 625.950 646.050 628.050 ;
        RECT 643.950 613.950 646.050 616.050 ;
        RECT 635.400 608.400 639.450 609.450 ;
        RECT 638.400 606.600 639.450 608.400 ;
        RECT 623.400 601.050 624.450 605.400 ;
        RECT 632.400 604.350 633.600 606.600 ;
        RECT 638.400 604.350 639.600 606.600 ;
        RECT 628.950 601.950 631.050 604.050 ;
        RECT 631.950 601.950 634.050 604.050 ;
        RECT 634.950 601.950 637.050 604.050 ;
        RECT 637.950 601.950 640.050 604.050 ;
        RECT 629.400 601.050 630.600 601.650 ;
        RECT 622.950 598.950 625.050 601.050 ;
        RECT 625.950 599.400 630.600 601.050 ;
        RECT 635.400 600.900 636.600 601.650 ;
        RECT 625.950 598.950 630.000 599.400 ;
        RECT 634.950 598.800 637.050 600.900 ;
        RECT 644.400 580.050 645.450 613.950 ;
        RECT 659.400 613.050 660.450 649.950 ;
        RECT 665.400 649.350 666.600 650.100 ;
        RECT 664.950 646.950 667.050 649.050 ;
        RECT 667.950 646.950 670.050 649.050 ;
        RECT 668.400 644.400 669.600 646.650 ;
        RECT 658.950 610.950 661.050 613.050 ;
        RECT 668.400 610.050 669.450 644.400 ;
        RECT 677.400 643.050 678.450 661.950 ;
        RECT 703.950 658.950 706.050 661.050 ;
        RECT 685.950 655.950 688.050 658.050 ;
        RECT 686.400 651.600 687.450 655.950 ;
        RECT 686.400 649.350 687.600 651.600 ;
        RECT 691.950 650.100 694.050 652.200 ;
        RECT 697.950 650.100 700.050 652.200 ;
        RECT 692.400 649.350 693.600 650.100 ;
        RECT 682.950 646.950 685.050 649.050 ;
        RECT 685.950 646.950 688.050 649.050 ;
        RECT 688.950 646.950 691.050 649.050 ;
        RECT 691.950 646.950 694.050 649.050 ;
        RECT 683.400 645.000 684.600 646.650 ;
        RECT 676.950 640.950 679.050 643.050 ;
        RECT 682.950 640.950 685.050 645.000 ;
        RECT 689.400 644.400 690.600 646.650 ;
        RECT 689.400 625.050 690.450 644.400 ;
        RECT 698.400 643.050 699.450 650.100 ;
        RECT 704.400 645.450 705.450 658.950 ;
        RECT 716.400 657.450 717.450 676.950 ;
        RECT 733.950 676.800 736.050 678.900 ;
        RECT 743.400 661.050 744.450 688.950 ;
        RECT 745.950 685.950 748.050 688.050 ;
        RECT 742.950 658.950 745.050 661.050 ;
        RECT 746.400 657.450 747.450 685.950 ;
        RECT 757.950 683.100 760.050 685.200 ;
        RECT 763.950 683.100 766.050 685.200 ;
        RECT 776.400 685.050 777.450 694.950 ;
        RECT 758.400 682.350 759.600 683.100 ;
        RECT 764.400 682.350 765.600 683.100 ;
        RECT 769.950 682.950 772.050 685.050 ;
        RECT 775.950 682.950 778.050 685.050 ;
        RECT 779.400 684.600 780.450 697.950 ;
        RECT 782.400 687.450 783.450 721.950 ;
        RECT 785.400 694.050 786.450 743.400 ;
        RECT 787.950 733.950 790.050 736.050 ;
        RECT 784.950 691.950 787.050 694.050 ;
        RECT 788.400 688.050 789.450 733.950 ;
        RECT 803.400 733.050 804.450 755.400 ;
        RECT 793.950 728.100 796.050 730.200 ;
        RECT 799.950 729.000 802.050 733.050 ;
        RECT 802.950 730.950 805.050 733.050 ;
        RECT 794.400 727.350 795.600 728.100 ;
        RECT 800.400 727.350 801.600 729.000 ;
        RECT 793.950 724.950 796.050 727.050 ;
        RECT 796.950 724.950 799.050 727.050 ;
        RECT 799.950 724.950 802.050 727.050 ;
        RECT 802.950 724.950 805.050 727.050 ;
        RECT 790.950 721.950 793.050 724.050 ;
        RECT 797.400 722.400 798.600 724.650 ;
        RECT 803.400 723.900 804.600 724.650 ;
        RECT 782.400 686.400 786.450 687.450 ;
        RECT 785.400 684.600 786.450 686.400 ;
        RECT 787.950 685.950 790.050 688.050 ;
        RECT 791.400 685.050 792.450 721.950 ;
        RECT 797.400 715.050 798.450 722.400 ;
        RECT 802.950 721.800 805.050 723.900 ;
        RECT 796.950 712.950 799.050 715.050 ;
        RECT 809.400 708.450 810.450 755.400 ;
        RECT 811.950 736.950 814.050 739.050 ;
        RECT 812.400 723.900 813.450 736.950 ;
        RECT 815.400 730.050 816.450 767.400 ;
        RECT 821.400 762.600 822.450 775.950 ;
        RECT 826.950 766.950 829.050 769.050 ;
        RECT 827.400 762.600 828.450 766.950 ;
        RECT 821.400 760.350 822.600 762.600 ;
        RECT 827.400 760.350 828.600 762.600 ;
        RECT 820.950 757.950 823.050 760.050 ;
        RECT 823.950 757.950 826.050 760.050 ;
        RECT 826.950 757.950 829.050 760.050 ;
        RECT 829.950 757.950 832.050 760.050 ;
        RECT 824.400 755.400 825.600 757.650 ;
        RECT 830.400 755.400 831.600 757.650 ;
        RECT 839.400 757.050 840.450 871.950 ;
        RECT 851.400 852.000 858.450 852.450 ;
        RECT 851.400 851.400 859.050 852.000 ;
        RECT 851.400 844.050 852.450 851.400 ;
        RECT 856.950 847.950 859.050 851.400 ;
        RECT 850.950 841.950 853.050 844.050 ;
        RECT 847.950 839.100 850.050 841.200 ;
        RECT 860.400 841.050 861.450 878.400 ;
        RECT 862.950 874.950 865.050 877.050 ;
        RECT 848.400 838.350 849.600 839.100 ;
        RECT 859.950 838.950 862.050 841.050 ;
        RECT 847.950 835.950 850.050 838.050 ;
        RECT 850.950 835.950 853.050 838.050 ;
        RECT 853.950 835.950 856.050 838.050 ;
        RECT 856.950 835.950 859.050 838.050 ;
        RECT 857.400 833.400 858.600 835.650 ;
        RECT 853.950 807.000 856.050 811.050 ;
        RECT 857.400 808.050 858.450 833.400 ;
        RECT 863.400 829.050 864.450 874.950 ;
        RECT 869.400 864.450 870.450 884.100 ;
        RECT 872.400 877.050 873.450 886.950 ;
        RECT 877.950 885.000 880.050 889.050 ;
        RECT 878.400 883.350 879.600 885.000 ;
        RECT 877.950 880.950 880.050 883.050 ;
        RECT 880.950 880.950 883.050 883.050 ;
        RECT 881.400 878.400 882.600 880.650 ;
        RECT 871.950 874.950 874.050 877.050 ;
        RECT 866.400 863.400 870.450 864.450 ;
        RECT 862.950 826.950 865.050 829.050 ;
        RECT 866.400 813.450 867.450 863.400 ;
        RECT 871.950 856.950 874.050 859.050 ;
        RECT 872.400 840.600 873.450 856.950 ;
        RECT 877.950 847.950 880.050 850.050 ;
        RECT 878.400 841.200 879.450 847.950 ;
        RECT 872.400 838.350 873.600 840.600 ;
        RECT 877.950 839.100 880.050 841.200 ;
        RECT 881.400 841.050 882.450 878.400 ;
        RECT 878.400 838.350 879.600 839.100 ;
        RECT 880.950 838.950 883.050 841.050 ;
        RECT 886.950 838.950 889.050 841.050 ;
        RECT 892.950 839.100 895.050 841.200 ;
        RECT 871.950 835.950 874.050 838.050 ;
        RECT 874.950 835.950 877.050 838.050 ;
        RECT 877.950 835.950 880.050 838.050 ;
        RECT 868.950 832.950 871.050 835.050 ;
        RECT 875.400 833.400 876.600 835.650 ;
        RECT 869.400 820.050 870.450 832.950 ;
        RECT 868.950 817.950 871.050 820.050 ;
        RECT 875.400 814.050 876.450 833.400 ;
        RECT 880.950 817.950 883.050 820.050 ;
        RECT 868.950 813.450 871.050 814.050 ;
        RECT 866.400 812.400 871.050 813.450 ;
        RECT 868.950 811.950 871.050 812.400 ;
        RECT 874.950 811.950 877.050 814.050 ;
        RECT 854.400 805.350 855.600 807.000 ;
        RECT 856.950 805.950 859.050 808.050 ;
        RECT 862.950 805.950 865.050 808.050 ;
        RECT 869.400 807.600 870.450 811.950 ;
        RECT 844.950 802.950 847.050 805.050 ;
        RECT 847.950 802.950 850.050 805.050 ;
        RECT 850.950 802.950 853.050 805.050 ;
        RECT 853.950 802.950 856.050 805.050 ;
        RECT 841.950 799.950 844.050 802.050 ;
        RECT 845.400 801.000 846.600 802.650 ;
        RECT 842.400 775.050 843.450 799.950 ;
        RECT 844.950 796.950 847.050 801.000 ;
        RECT 859.950 796.950 862.050 799.050 ;
        RECT 841.950 772.950 844.050 775.050 ;
        RECT 847.950 762.000 850.050 766.050 ;
        RECT 853.950 762.000 856.050 766.050 ;
        RECT 848.400 760.350 849.600 762.000 ;
        RECT 854.400 760.350 855.600 762.000 ;
        RECT 844.950 757.950 847.050 760.050 ;
        RECT 847.950 757.950 850.050 760.050 ;
        RECT 850.950 757.950 853.050 760.050 ;
        RECT 853.950 757.950 856.050 760.050 ;
        RECT 824.400 739.050 825.450 755.400 ;
        RECT 830.400 751.050 831.450 755.400 ;
        RECT 832.950 754.950 835.050 757.050 ;
        RECT 838.950 754.950 841.050 757.050 ;
        RECT 845.400 755.400 846.600 757.650 ;
        RECT 851.400 756.900 852.600 757.650 ;
        RECT 829.950 748.950 832.050 751.050 ;
        RECT 823.950 736.950 826.050 739.050 ;
        RECT 814.950 727.950 817.050 730.050 ;
        RECT 817.950 729.000 820.050 733.050 ;
        RECT 824.400 729.600 825.450 736.950 ;
        RECT 818.400 727.350 819.600 729.000 ;
        RECT 824.400 727.350 825.600 729.600 ;
        RECT 817.950 724.950 820.050 727.050 ;
        RECT 820.950 724.950 823.050 727.050 ;
        RECT 823.950 724.950 826.050 727.050 ;
        RECT 826.950 724.950 829.050 727.050 ;
        RECT 811.800 721.800 813.900 723.900 ;
        RECT 814.950 718.950 817.050 724.050 ;
        RECT 821.400 723.900 822.600 724.650 ;
        RECT 820.950 718.950 823.050 723.900 ;
        RECT 827.400 722.400 828.600 724.650 ;
        RECT 827.400 718.050 828.450 722.400 ;
        RECT 833.400 718.050 834.450 754.950 ;
        RECT 845.400 751.050 846.450 755.400 ;
        RECT 850.950 754.800 853.050 756.900 ;
        RECT 844.950 748.950 847.050 751.050 ;
        RECT 838.950 736.950 841.050 739.050 ;
        RECT 835.950 728.100 838.050 730.200 ;
        RECT 839.400 730.050 840.450 736.950 ;
        RECT 845.400 732.450 846.450 748.950 ;
        RECT 842.400 731.400 846.450 732.450 ;
        RECT 836.400 723.450 837.450 728.100 ;
        RECT 838.950 727.950 841.050 730.050 ;
        RECT 842.400 729.600 843.450 731.400 ;
        RECT 842.400 727.350 843.600 729.600 ;
        RECT 847.950 728.100 850.050 730.200 ;
        RECT 856.950 728.100 859.050 730.200 ;
        RECT 848.400 727.350 849.600 728.100 ;
        RECT 841.950 724.950 844.050 727.050 ;
        RECT 844.950 724.950 847.050 727.050 ;
        RECT 847.950 724.950 850.050 727.050 ;
        RECT 850.950 724.950 853.050 727.050 ;
        RECT 845.400 723.900 846.600 724.650 ;
        RECT 836.400 722.400 840.450 723.450 ;
        RECT 820.950 712.950 823.050 717.900 ;
        RECT 826.950 715.950 829.050 718.050 ;
        RECT 832.950 715.950 835.050 718.050 ;
        RECT 811.950 708.450 814.050 709.050 ;
        RECT 809.400 707.400 814.050 708.450 ;
        RECT 811.950 706.950 814.050 707.400 ;
        RECT 805.950 697.950 808.050 700.050 ;
        RECT 796.950 691.950 799.050 694.050 ;
        RECT 793.950 685.950 796.050 688.050 ;
        RECT 754.950 679.950 757.050 682.050 ;
        RECT 757.950 679.950 760.050 682.050 ;
        RECT 760.950 679.950 763.050 682.050 ;
        RECT 763.950 679.950 766.050 682.050 ;
        RECT 755.400 677.400 756.600 679.650 ;
        RECT 761.400 678.900 762.600 679.650 ;
        RECT 755.400 673.050 756.450 677.400 ;
        RECT 760.950 676.800 763.050 678.900 ;
        RECT 766.950 673.950 769.050 679.050 ;
        RECT 754.950 670.950 757.050 673.050 ;
        RECT 763.950 658.950 766.050 661.050 ;
        RECT 748.950 657.450 751.050 658.050 ;
        RECT 716.400 655.200 717.600 657.450 ;
        RECT 746.400 656.400 751.050 657.450 ;
        RECT 711.900 651.900 714.000 653.700 ;
        RECT 715.800 652.800 717.900 654.900 ;
        RECT 719.100 654.300 721.200 656.400 ;
        RECT 748.950 655.950 751.050 656.400 ;
        RECT 710.400 650.700 719.100 651.900 ;
        RECT 707.100 646.950 709.200 649.050 ;
        RECT 707.400 645.900 708.600 646.650 ;
        RECT 706.950 645.450 709.050 645.900 ;
        RECT 704.400 644.400 709.050 645.450 ;
        RECT 706.950 643.800 709.050 644.400 ;
        RECT 691.950 640.950 694.050 643.050 ;
        RECT 697.950 640.950 700.050 643.050 ;
        RECT 710.400 641.700 711.300 650.700 ;
        RECT 717.000 649.800 719.100 650.700 ;
        RECT 720.000 648.900 720.900 654.300 ;
        RECT 742.500 653.400 744.600 655.500 ;
        RECT 749.400 655.200 750.600 655.950 ;
        RECT 722.400 651.450 723.600 651.600 ;
        RECT 722.400 650.400 726.450 651.450 ;
        RECT 722.400 649.350 723.600 650.400 ;
        RECT 714.000 647.700 720.900 648.900 ;
        RECT 714.000 645.300 714.900 647.700 ;
        RECT 712.800 643.200 714.900 645.300 ;
        RECT 715.800 643.950 717.900 646.050 ;
        RECT 688.950 622.950 691.050 625.050 ;
        RECT 655.950 605.100 658.050 607.200 ;
        RECT 661.950 605.100 664.050 607.200 ;
        RECT 667.950 606.450 670.050 610.050 ;
        RECT 667.950 605.400 672.450 606.450 ;
        RECT 656.400 604.350 657.600 605.100 ;
        RECT 662.400 604.350 663.600 605.100 ;
        RECT 667.950 604.950 670.050 605.400 ;
        RECT 652.950 601.950 655.050 604.050 ;
        RECT 655.950 601.950 658.050 604.050 ;
        RECT 658.950 601.950 661.050 604.050 ;
        RECT 661.950 601.950 664.050 604.050 ;
        RECT 667.950 601.800 670.050 603.900 ;
        RECT 653.400 600.900 654.600 601.650 ;
        RECT 652.950 598.800 655.050 600.900 ;
        RECT 659.400 599.400 660.600 601.650 ;
        RECT 659.400 586.050 660.450 599.400 ;
        RECT 668.400 595.050 669.450 601.800 ;
        RECT 667.950 592.950 670.050 595.050 ;
        RECT 658.950 583.950 661.050 586.050 ;
        RECT 643.950 577.950 646.050 580.050 ;
        RECT 658.950 577.950 661.050 580.050 ;
        RECT 622.950 573.450 625.050 574.200 ;
        RECT 620.400 572.400 625.050 573.450 ;
        RECT 622.950 572.100 625.050 572.400 ;
        RECT 631.950 572.100 634.050 574.200 ;
        RECT 611.400 571.350 612.600 572.100 ;
        RECT 604.950 568.950 607.050 571.050 ;
        RECT 607.950 568.950 610.050 571.050 ;
        RECT 610.950 568.950 613.050 571.050 ;
        RECT 613.950 568.950 616.050 571.050 ;
        RECT 601.950 565.950 604.050 568.050 ;
        RECT 608.400 567.000 609.600 568.650 ;
        RECT 614.400 567.900 615.600 568.650 ;
        RECT 623.400 568.050 624.450 572.100 ;
        RECT 632.400 571.350 633.600 572.100 ;
        RECT 628.950 568.950 631.050 571.050 ;
        RECT 631.950 568.950 634.050 571.050 ;
        RECT 634.950 568.950 637.050 571.050 ;
        RECT 595.950 562.950 598.050 565.050 ;
        RECT 559.950 559.950 562.050 562.050 ;
        RECT 565.950 559.950 568.050 562.050 ;
        RECT 571.950 559.950 574.050 562.050 ;
        RECT 553.950 553.950 556.050 556.050 ;
        RECT 539.400 526.350 540.600 527.100 ;
        RECT 544.950 526.950 547.050 529.050 ;
        RECT 550.950 526.950 553.050 529.050 ;
        RECT 553.950 527.100 556.050 529.200 ;
        RECT 559.950 528.000 562.050 532.050 ;
        RECT 566.400 529.050 567.450 559.950 ;
        RECT 602.400 541.050 603.450 565.950 ;
        RECT 607.950 562.950 610.050 567.000 ;
        RECT 613.950 565.800 616.050 567.900 ;
        RECT 622.950 565.950 625.050 568.050 ;
        RECT 629.400 566.400 630.600 568.650 ;
        RECT 635.400 566.400 636.600 568.650 ;
        RECT 629.400 556.050 630.450 566.400 ;
        RECT 635.400 562.050 636.450 566.400 ;
        RECT 634.950 559.950 637.050 562.050 ;
        RECT 628.950 553.950 631.050 556.050 ;
        RECT 640.950 544.950 643.050 547.050 ;
        RECT 601.950 538.950 604.050 541.050 ;
        RECT 628.950 538.950 631.050 541.050 ;
        RECT 577.950 535.950 580.050 538.050 ;
        RECT 616.950 535.950 619.050 538.050 ;
        RECT 535.950 523.950 538.050 526.050 ;
        RECT 538.950 523.950 541.050 526.050 ;
        RECT 529.950 517.950 532.050 520.050 ;
        RECT 532.950 517.950 535.050 523.050 ;
        RECT 536.400 521.400 537.600 523.650 ;
        RECT 536.400 517.050 537.450 521.400 ;
        RECT 541.950 517.950 544.050 520.050 ;
        RECT 535.950 514.950 538.050 517.050 ;
        RECT 542.400 514.050 543.450 517.950 ;
        RECT 541.950 511.950 544.050 514.050 ;
        RECT 545.400 502.050 546.450 526.950 ;
        RECT 554.400 526.350 555.600 527.100 ;
        RECT 560.400 526.350 561.600 528.000 ;
        RECT 565.950 526.950 568.050 529.050 ;
        RECT 571.950 527.100 574.050 529.200 ;
        RECT 578.400 528.600 579.450 535.950 ;
        RECT 553.950 523.950 556.050 526.050 ;
        RECT 556.950 523.950 559.050 526.050 ;
        RECT 559.950 523.950 562.050 526.050 ;
        RECT 562.950 523.950 565.050 526.050 ;
        RECT 550.950 520.950 553.050 523.050 ;
        RECT 557.400 521.400 558.600 523.650 ;
        RECT 563.400 522.450 564.600 523.650 ;
        RECT 568.950 522.450 571.050 526.050 ;
        RECT 563.400 522.000 571.050 522.450 ;
        RECT 563.400 521.400 570.450 522.000 ;
        RECT 551.400 517.050 552.450 520.950 ;
        RECT 553.950 517.950 556.050 520.050 ;
        RECT 550.950 514.950 553.050 517.050 ;
        RECT 550.950 511.800 553.050 513.900 ;
        RECT 551.400 508.050 552.450 511.800 ;
        RECT 550.950 505.950 553.050 508.050 ;
        RECT 529.950 499.950 532.050 502.050 ;
        RECT 544.950 499.950 547.050 502.050 ;
        RECT 530.400 496.050 531.450 499.950 ;
        RECT 526.950 493.950 529.050 496.050 ;
        RECT 529.950 493.950 532.050 496.050 ;
        RECT 535.950 494.100 538.050 496.200 ;
        RECT 541.950 495.000 544.050 499.050 ;
        RECT 536.400 493.350 537.600 494.100 ;
        RECT 542.400 493.350 543.600 495.000 ;
        RECT 526.950 490.800 529.050 492.900 ;
        RECT 532.950 490.950 535.050 493.050 ;
        RECT 535.950 490.950 538.050 493.050 ;
        RECT 538.950 490.950 541.050 493.050 ;
        RECT 541.950 490.950 544.050 493.050 ;
        RECT 544.950 490.950 547.050 493.050 ;
        RECT 523.950 487.950 526.050 490.050 ;
        RECT 518.400 449.400 522.450 450.450 ;
        RECT 527.400 450.600 528.450 490.800 ;
        RECT 529.950 487.950 532.050 490.050 ;
        RECT 533.400 489.900 534.600 490.650 ;
        RECT 530.400 451.050 531.450 487.950 ;
        RECT 532.950 487.800 535.050 489.900 ;
        RECT 539.400 488.400 540.600 490.650 ;
        RECT 545.400 489.450 546.600 490.650 ;
        RECT 545.400 489.000 549.450 489.450 ;
        RECT 545.400 488.400 550.050 489.000 ;
        RECT 535.950 484.950 538.050 487.050 ;
        RECT 499.950 445.950 502.050 448.050 ;
        RECT 502.950 445.950 505.050 448.050 ;
        RECT 505.950 445.950 508.050 448.050 ;
        RECT 508.950 445.950 511.050 448.050 ;
        RECT 503.400 444.900 504.600 445.650 ;
        RECT 502.950 442.800 505.050 444.900 ;
        RECT 509.400 443.400 510.600 445.650 ;
        RECT 509.400 433.050 510.450 443.400 ;
        RECT 466.950 430.950 469.050 433.050 ;
        RECT 478.950 430.950 481.050 433.050 ;
        RECT 493.950 430.950 496.050 433.050 ;
        RECT 508.950 430.950 511.050 433.050 ;
        RECT 457.950 421.950 460.050 424.050 ;
        RECT 451.950 417.000 454.050 421.050 ;
        RECT 458.400 417.600 459.450 421.950 ;
        RECT 452.400 415.350 453.600 417.000 ;
        RECT 458.400 415.350 459.600 417.600 ;
        RECT 467.400 415.050 468.450 430.950 ;
        RECT 479.400 417.600 480.450 430.950 ;
        RECT 515.400 429.450 516.450 448.950 ;
        RECT 512.400 428.400 516.450 429.450 ;
        RECT 518.400 429.450 519.450 449.400 ;
        RECT 527.400 448.350 528.600 450.600 ;
        RECT 529.950 448.950 532.050 451.050 ;
        RECT 523.950 445.950 526.050 448.050 ;
        RECT 526.950 445.950 529.050 448.050 ;
        RECT 524.400 443.400 525.600 445.650 ;
        RECT 536.400 444.900 537.450 484.950 ;
        RECT 539.400 457.050 540.450 488.400 ;
        RECT 544.950 484.950 547.050 487.050 ;
        RECT 547.950 484.950 550.050 488.400 ;
        RECT 554.400 487.050 555.450 517.950 ;
        RECT 557.400 517.050 558.450 521.400 ;
        RECT 572.400 517.050 573.450 527.100 ;
        RECT 578.400 526.350 579.600 528.600 ;
        RECT 598.950 527.100 601.050 529.200 ;
        RECT 604.950 527.100 607.050 529.200 ;
        RECT 613.950 527.100 616.050 529.200 ;
        RECT 599.400 526.350 600.600 527.100 ;
        RECT 605.400 526.350 606.600 527.100 ;
        RECT 577.950 523.950 580.050 526.050 ;
        RECT 580.950 523.950 583.050 526.050 ;
        RECT 583.950 523.950 586.050 526.050 ;
        RECT 598.950 523.950 601.050 526.050 ;
        RECT 601.950 523.950 604.050 526.050 ;
        RECT 604.950 523.950 607.050 526.050 ;
        RECT 581.400 522.900 582.600 523.650 ;
        RECT 580.950 520.800 583.050 522.900 ;
        RECT 602.400 521.400 603.600 523.650 ;
        RECT 556.950 514.950 559.050 517.050 ;
        RECT 571.950 514.950 574.050 517.050 ;
        RECT 559.950 505.950 562.050 508.050 ;
        RECT 560.400 496.200 561.450 505.950 ;
        RECT 559.950 494.100 562.050 496.200 ;
        RECT 565.950 494.100 568.050 496.200 ;
        RECT 581.400 495.450 582.450 520.800 ;
        RECT 595.950 517.950 598.050 520.050 ;
        RECT 584.400 495.450 585.600 495.600 ;
        RECT 581.400 494.400 585.600 495.450 ;
        RECT 560.400 493.350 561.600 494.100 ;
        RECT 566.400 493.350 567.600 494.100 ;
        RECT 584.400 493.350 585.600 494.400 ;
        RECT 559.950 490.950 562.050 493.050 ;
        RECT 562.950 490.950 565.050 493.050 ;
        RECT 565.950 490.950 568.050 493.050 ;
        RECT 568.950 490.950 571.050 493.050 ;
        RECT 583.950 490.950 586.050 493.050 ;
        RECT 586.950 490.950 589.050 493.050 ;
        RECT 563.400 489.000 564.600 490.650 ;
        RECT 569.400 489.900 570.600 490.650 ;
        RECT 587.400 489.900 588.600 490.650 ;
        RECT 553.950 484.950 556.050 487.050 ;
        RECT 545.400 481.050 546.450 484.950 ;
        RECT 559.950 483.450 562.050 487.050 ;
        RECT 562.950 484.950 565.050 489.000 ;
        RECT 568.950 487.800 571.050 489.900 ;
        RECT 574.950 487.800 577.050 489.900 ;
        RECT 586.950 487.800 589.050 489.900 ;
        RECT 565.950 483.450 568.050 484.050 ;
        RECT 559.950 483.000 568.050 483.450 ;
        RECT 560.400 482.400 568.050 483.000 ;
        RECT 565.950 481.950 568.050 482.400 ;
        RECT 575.400 481.050 576.450 487.800 ;
        RECT 596.400 487.050 597.450 517.950 ;
        RECT 602.400 517.050 603.450 521.400 ;
        RECT 614.400 520.050 615.450 527.100 ;
        RECT 613.950 517.950 616.050 520.050 ;
        RECT 601.950 514.950 604.050 517.050 ;
        RECT 613.950 499.950 616.050 502.050 ;
        RECT 598.950 493.950 601.050 496.050 ;
        RECT 607.950 494.100 610.050 496.200 ;
        RECT 614.400 495.600 615.450 499.950 ;
        RECT 599.400 487.050 600.450 493.950 ;
        RECT 608.400 493.350 609.600 494.100 ;
        RECT 614.400 493.350 615.600 495.600 ;
        RECT 617.400 495.450 618.450 535.950 ;
        RECT 622.950 527.100 625.050 529.200 ;
        RECT 629.400 528.600 630.450 538.950 ;
        RECT 623.400 526.350 624.600 527.100 ;
        RECT 629.400 526.350 630.600 528.600 ;
        RECT 622.950 523.950 625.050 526.050 ;
        RECT 625.950 523.950 628.050 526.050 ;
        RECT 628.950 523.950 631.050 526.050 ;
        RECT 631.950 523.950 634.050 526.050 ;
        RECT 626.400 521.400 627.600 523.650 ;
        RECT 632.400 522.900 633.600 523.650 ;
        RECT 626.400 514.050 627.450 521.400 ;
        RECT 631.950 520.800 634.050 522.900 ;
        RECT 625.950 511.950 628.050 514.050 ;
        RECT 632.400 505.050 633.450 520.800 ;
        RECT 622.950 502.950 625.050 505.050 ;
        RECT 631.950 502.950 634.050 505.050 ;
        RECT 617.400 494.400 621.450 495.450 ;
        RECT 604.950 490.950 607.050 493.050 ;
        RECT 607.950 490.950 610.050 493.050 ;
        RECT 610.950 490.950 613.050 493.050 ;
        RECT 613.950 490.950 616.050 493.050 ;
        RECT 605.400 489.000 606.600 490.650 ;
        RECT 595.950 484.950 598.050 487.050 ;
        RECT 598.950 481.950 601.050 487.050 ;
        RECT 604.950 484.950 607.050 489.000 ;
        RECT 611.400 488.400 612.600 490.650 ;
        RECT 611.400 487.050 612.450 488.400 ;
        RECT 610.950 484.950 613.050 487.050 ;
        RECT 544.950 478.950 547.050 481.050 ;
        RECT 574.950 478.950 577.050 481.050 ;
        RECT 538.950 454.950 541.050 457.050 ;
        RECT 545.400 450.600 546.450 478.950 ;
        RECT 571.950 475.950 574.050 478.050 ;
        RECT 562.950 472.950 565.050 475.050 ;
        RECT 545.400 448.350 546.600 450.600 ;
        RECT 550.950 449.100 553.050 451.200 ;
        RECT 559.950 449.100 562.050 451.200 ;
        RECT 563.400 451.050 564.450 472.950 ;
        RECT 551.400 448.350 552.600 449.100 ;
        RECT 541.950 445.950 544.050 448.050 ;
        RECT 544.950 445.950 547.050 448.050 ;
        RECT 547.950 445.950 550.050 448.050 ;
        RECT 550.950 445.950 553.050 448.050 ;
        RECT 542.400 444.900 543.600 445.650 ;
        RECT 548.400 444.900 549.600 445.650 ;
        RECT 518.400 428.400 522.450 429.450 ;
        RECT 484.950 421.950 487.050 424.050 ;
        RECT 490.950 421.950 493.050 424.050 ;
        RECT 485.400 417.600 486.450 421.950 ;
        RECT 479.400 415.350 480.600 417.600 ;
        RECT 485.400 415.350 486.600 417.600 ;
        RECT 451.950 412.950 454.050 415.050 ;
        RECT 454.950 412.950 457.050 415.050 ;
        RECT 457.950 412.950 460.050 415.050 ;
        RECT 460.950 412.950 463.050 415.050 ;
        RECT 466.950 412.950 469.050 415.050 ;
        RECT 475.950 412.950 478.050 415.050 ;
        RECT 478.950 412.950 481.050 415.050 ;
        RECT 481.950 412.950 484.050 415.050 ;
        RECT 484.950 412.950 487.050 415.050 ;
        RECT 455.400 411.900 456.600 412.650 ;
        RECT 454.950 409.800 457.050 411.900 ;
        RECT 461.400 410.400 462.600 412.650 ;
        RECT 476.400 411.450 477.600 412.650 ;
        RECT 482.400 411.900 483.600 412.650 ;
        RECT 491.400 411.900 492.450 421.950 ;
        RECT 502.950 416.100 505.050 418.200 ;
        RECT 512.400 417.600 513.450 428.400 ;
        RECT 517.350 423.300 519.450 425.400 ;
        RECT 503.400 415.350 504.600 416.100 ;
        RECT 512.400 415.350 513.600 417.600 ;
        RECT 499.950 412.950 502.050 415.050 ;
        RECT 502.950 412.950 505.050 415.050 ;
        RECT 505.950 412.950 508.050 415.050 ;
        RECT 511.950 412.950 514.050 415.050 ;
        RECT 500.400 411.900 501.600 412.650 ;
        RECT 506.400 411.900 507.600 412.650 ;
        RECT 473.400 410.400 477.600 411.450 ;
        RECT 457.950 400.950 460.050 403.050 ;
        RECT 445.950 397.950 448.050 400.050 ;
        RECT 439.950 391.950 442.050 397.050 ;
        RECT 448.950 391.950 451.050 397.050 ;
        RECT 442.950 388.950 445.050 391.050 ;
        RECT 421.950 373.950 424.050 376.050 ;
        RECT 418.950 371.100 421.050 373.200 ;
        RECT 443.400 372.600 444.450 388.950 ;
        RECT 454.950 382.950 457.050 385.050 ;
        RECT 419.400 370.350 420.600 371.100 ;
        RECT 443.400 370.350 444.600 372.600 ;
        RECT 448.950 372.000 451.050 376.050 ;
        RECT 449.400 370.350 450.600 372.000 ;
        RECT 419.100 367.950 421.200 370.050 ;
        RECT 424.500 367.950 426.600 370.050 ;
        RECT 439.950 367.950 442.050 370.050 ;
        RECT 442.950 367.950 445.050 370.050 ;
        RECT 445.950 367.950 448.050 370.050 ;
        RECT 448.950 367.950 451.050 370.050 ;
        RECT 440.400 366.900 441.600 367.650 ;
        RECT 439.950 364.800 442.050 366.900 ;
        RECT 446.400 365.400 447.600 367.650 ;
        RECT 416.400 363.000 420.450 363.450 ;
        RECT 416.400 362.400 421.050 363.000 ;
        RECT 418.950 358.950 421.050 362.400 ;
        RECT 442.950 358.950 445.050 361.050 ;
        RECT 409.950 352.950 412.050 355.050 ;
        RECT 433.950 349.950 436.050 352.050 ;
        RECT 376.950 346.950 379.050 349.050 ;
        RECT 391.950 346.950 394.050 349.050 ;
        RECT 400.950 346.950 403.050 349.050 ;
        RECT 418.950 346.950 421.050 349.050 ;
        RECT 358.950 343.950 361.050 346.050 ;
        RECT 346.950 337.950 349.050 340.050 ;
        RECT 355.950 338.100 358.050 340.200 ;
        RECT 347.400 337.350 348.600 337.950 ;
        RECT 346.950 334.950 349.050 337.050 ;
        RECT 349.950 334.950 352.050 337.050 ;
        RECT 350.400 332.400 351.600 334.650 ;
        RECT 350.400 328.050 351.450 332.400 ;
        RECT 349.950 325.950 352.050 328.050 ;
        RECT 356.400 319.050 357.450 338.100 ;
        RECT 343.950 316.950 346.050 319.050 ;
        RECT 355.950 316.950 358.050 319.050 ;
        RECT 344.400 313.050 345.450 316.950 ;
        RECT 343.950 310.950 346.050 313.050 ;
        RECT 340.950 304.950 343.050 307.050 ;
        RECT 359.400 304.050 360.450 343.950 ;
        RECT 367.950 338.100 370.050 340.200 ;
        RECT 377.400 339.600 378.450 346.950 ;
        RECT 388.950 343.950 391.050 346.050 ;
        RECT 368.400 337.350 369.600 338.100 ;
        RECT 377.400 337.350 378.600 339.600 ;
        RECT 367.800 334.950 369.900 337.050 ;
        RECT 373.950 334.950 376.050 337.050 ;
        RECT 376.950 334.950 379.050 337.050 ;
        RECT 382.500 334.950 384.600 337.050 ;
        RECT 374.400 332.400 375.600 334.650 ;
        RECT 383.400 332.400 384.600 334.650 ;
        RECT 374.400 325.050 375.450 332.400 ;
        RECT 373.950 322.950 376.050 325.050 ;
        RECT 383.400 322.050 384.450 332.400 ;
        RECT 389.400 328.050 390.450 343.950 ;
        RECT 392.400 333.900 393.450 346.950 ;
        RECT 394.950 343.950 400.050 346.050 ;
        RECT 394.950 338.100 397.050 340.200 ;
        RECT 400.950 338.100 403.050 340.200 ;
        RECT 406.950 338.100 409.050 340.200 ;
        RECT 391.950 331.800 394.050 333.900 ;
        RECT 388.950 325.950 391.050 328.050 ;
        RECT 395.400 325.050 396.450 338.100 ;
        RECT 401.400 337.350 402.600 338.100 ;
        RECT 407.400 337.350 408.600 338.100 ;
        RECT 400.950 334.950 403.050 337.050 ;
        RECT 403.950 334.950 406.050 337.050 ;
        RECT 406.950 334.950 409.050 337.050 ;
        RECT 409.950 334.950 412.050 337.050 ;
        RECT 404.400 333.900 405.600 334.650 ;
        RECT 403.950 331.800 406.050 333.900 ;
        RECT 410.400 332.400 411.600 334.650 ;
        RECT 419.400 333.900 420.450 346.950 ;
        RECT 427.950 343.950 430.050 346.050 ;
        RECT 428.400 339.600 429.450 343.950 ;
        RECT 434.400 339.600 435.450 349.950 ;
        RECT 428.400 337.350 429.600 339.600 ;
        RECT 434.400 337.350 435.600 339.600 ;
        RECT 439.950 337.950 442.050 340.050 ;
        RECT 424.950 334.950 427.050 337.050 ;
        RECT 427.950 334.950 430.050 337.050 ;
        RECT 430.950 334.950 433.050 337.050 ;
        RECT 433.950 334.950 436.050 337.050 ;
        RECT 425.400 333.900 426.600 334.650 ;
        RECT 394.950 322.950 397.050 325.050 ;
        RECT 403.950 322.950 406.050 325.050 ;
        RECT 382.950 319.950 385.050 322.050 ;
        RECT 394.950 316.950 397.050 319.050 ;
        RECT 343.950 301.950 346.050 304.050 ;
        RECT 349.950 301.950 352.050 304.050 ;
        RECT 358.950 301.950 361.050 304.050 ;
        RECT 379.950 301.950 382.050 304.050 ;
        RECT 310.950 298.950 313.050 301.050 ;
        RECT 322.950 298.950 325.050 301.050 ;
        RECT 313.950 293.100 316.050 295.200 ;
        RECT 314.400 292.350 315.600 293.100 ;
        RECT 310.950 289.950 313.050 292.050 ;
        RECT 313.950 289.950 316.050 292.050 ;
        RECT 304.950 286.800 307.050 288.900 ;
        RECT 307.950 286.950 310.050 289.050 ;
        RECT 311.400 288.900 312.600 289.650 ;
        RECT 323.400 288.900 324.450 298.950 ;
        RECT 331.950 294.000 334.050 298.050 ;
        RECT 332.400 292.350 333.600 294.000 ;
        RECT 340.950 292.950 343.050 295.050 ;
        RECT 328.950 289.950 331.050 292.050 ;
        RECT 331.950 289.950 334.050 292.050 ;
        RECT 329.400 288.900 330.600 289.650 ;
        RECT 298.950 283.950 301.050 286.050 ;
        RECT 301.950 274.950 304.050 277.050 ;
        RECT 286.950 265.950 289.050 268.050 ;
        RECT 295.950 265.950 298.050 268.050 ;
        RECT 278.400 259.350 279.600 261.600 ;
        RECT 286.950 261.000 289.050 264.900 ;
        RECT 287.400 259.350 288.600 261.000 ;
        RECT 292.950 259.950 295.050 262.050 ;
        RECT 272.400 256.950 274.500 259.050 ;
        RECT 277.950 256.950 280.050 259.050 ;
        RECT 280.950 256.950 283.050 259.050 ;
        RECT 287.100 256.950 289.200 259.050 ;
        RECT 272.400 254.400 273.600 256.650 ;
        RECT 281.400 255.900 282.600 256.650 ;
        RECT 293.400 255.900 294.450 259.950 ;
        RECT 268.950 247.950 271.050 250.050 ;
        RECT 272.400 232.050 273.450 254.400 ;
        RECT 280.950 253.800 283.050 255.900 ;
        RECT 292.950 253.800 295.050 255.900 ;
        RECT 271.950 229.950 274.050 232.050 ;
        RECT 296.400 229.050 297.450 265.950 ;
        RECT 302.400 255.900 303.450 274.950 ;
        RECT 308.400 262.200 309.450 286.950 ;
        RECT 310.950 286.800 313.050 288.900 ;
        RECT 322.950 286.800 325.050 288.900 ;
        RECT 328.950 286.800 331.050 288.900 ;
        RECT 323.400 265.050 324.450 286.800 ;
        RECT 329.400 270.450 330.450 286.800 ;
        RECT 341.400 286.050 342.450 292.950 ;
        RECT 340.950 283.950 343.050 286.050 ;
        RECT 329.400 269.400 333.450 270.450 ;
        RECT 322.950 262.950 325.050 265.050 ;
        RECT 307.950 260.100 310.050 262.200 ;
        RECT 313.950 260.100 316.050 262.200 ;
        RECT 308.400 259.350 309.600 260.100 ;
        RECT 314.400 259.350 315.600 260.100 ;
        RECT 307.950 256.950 310.050 259.050 ;
        RECT 310.950 256.950 313.050 259.050 ;
        RECT 313.950 256.950 316.050 259.050 ;
        RECT 316.950 256.950 319.050 259.050 ;
        RECT 311.400 255.900 312.600 256.650 ;
        RECT 317.400 255.900 318.600 256.650 ;
        RECT 323.400 255.900 324.450 262.950 ;
        RECT 332.400 261.600 333.450 269.400 ;
        RECT 332.400 259.350 333.600 261.600 ;
        RECT 337.950 260.100 340.050 262.200 ;
        RECT 344.400 262.050 345.450 301.950 ;
        RECT 350.400 294.600 351.450 301.950 ;
        RECT 350.400 292.350 351.600 294.600 ;
        RECT 355.950 294.000 358.050 298.050 ;
        RECT 373.950 294.000 376.050 298.050 ;
        RECT 380.400 294.600 381.450 301.950 ;
        RECT 356.400 292.350 357.600 294.000 ;
        RECT 374.400 292.350 375.600 294.000 ;
        RECT 380.400 292.350 381.600 294.600 ;
        RECT 349.950 289.950 352.050 292.050 ;
        RECT 352.950 289.950 355.050 292.050 ;
        RECT 355.950 289.950 358.050 292.050 ;
        RECT 358.950 289.950 361.050 292.050 ;
        RECT 373.950 289.950 376.050 292.050 ;
        RECT 376.950 289.950 379.050 292.050 ;
        RECT 379.950 289.950 382.050 292.050 ;
        RECT 382.950 289.950 385.050 292.050 ;
        RECT 353.400 288.000 354.600 289.650 ;
        RECT 352.950 283.950 355.050 288.000 ;
        RECT 359.400 287.400 360.600 289.650 ;
        RECT 377.400 288.900 378.600 289.650 ;
        RECT 359.400 280.050 360.450 287.400 ;
        RECT 376.950 286.800 379.050 288.900 ;
        RECT 383.400 287.400 384.600 289.650 ;
        RECT 395.400 288.900 396.450 316.950 ;
        RECT 404.400 294.600 405.450 322.950 ;
        RECT 410.400 319.050 411.450 332.400 ;
        RECT 418.950 331.800 421.050 333.900 ;
        RECT 424.950 331.800 427.050 333.900 ;
        RECT 431.400 332.400 432.600 334.650 ;
        RECT 409.950 316.950 412.050 319.050 ;
        RECT 419.400 295.200 420.450 331.800 ;
        RECT 431.400 331.050 432.450 332.400 ;
        RECT 430.950 330.450 433.050 331.050 ;
        RECT 428.400 329.400 433.050 330.450 ;
        RECT 404.400 292.350 405.600 294.600 ;
        RECT 409.950 293.100 412.050 295.200 ;
        RECT 418.950 293.100 421.050 295.200 ;
        RECT 428.400 294.600 429.450 329.400 ;
        RECT 430.950 328.950 433.050 329.400 ;
        RECT 440.400 325.050 441.450 337.950 ;
        RECT 439.950 322.950 442.050 325.050 ;
        RECT 439.950 310.950 442.050 313.050 ;
        RECT 410.400 292.350 411.600 293.100 ;
        RECT 428.400 292.350 429.600 294.600 ;
        RECT 400.950 289.950 403.050 292.050 ;
        RECT 403.950 289.950 406.050 292.050 ;
        RECT 406.950 289.950 409.050 292.050 ;
        RECT 409.950 289.950 412.050 292.050 ;
        RECT 424.950 289.950 427.050 292.050 ;
        RECT 427.950 289.950 430.050 292.050 ;
        RECT 401.400 288.900 402.600 289.650 ;
        RECT 358.950 277.950 361.050 280.050 ;
        RECT 373.950 277.950 376.050 280.050 ;
        RECT 338.400 259.350 339.600 260.100 ;
        RECT 343.950 259.950 346.050 262.050 ;
        RECT 346.950 259.950 349.050 262.050 ;
        RECT 325.950 256.950 328.050 259.050 ;
        RECT 331.950 256.950 334.050 259.050 ;
        RECT 334.950 256.950 337.050 259.050 ;
        RECT 337.950 256.950 340.050 259.050 ;
        RECT 340.950 256.950 343.050 259.050 ;
        RECT 301.950 253.800 304.050 255.900 ;
        RECT 310.950 253.800 313.050 255.900 ;
        RECT 316.950 253.800 319.050 255.900 ;
        RECT 322.950 253.800 325.050 255.900 ;
        RECT 326.400 232.050 327.450 256.950 ;
        RECT 335.400 255.000 336.600 256.650 ;
        RECT 341.400 256.050 342.600 256.650 ;
        RECT 334.950 250.950 337.050 255.000 ;
        RECT 341.400 254.400 346.050 256.050 ;
        RECT 342.000 253.950 346.050 254.400 ;
        RECT 325.950 229.950 328.050 232.050 ;
        RECT 295.950 226.950 298.050 229.050 ;
        RECT 310.950 226.950 313.050 229.050 ;
        RECT 271.950 220.950 274.050 223.050 ;
        RECT 235.950 217.950 238.050 220.050 ;
        RECT 244.950 216.000 247.050 220.050 ;
        RECT 250.950 216.000 253.050 220.050 ;
        RECT 245.400 214.350 246.600 216.000 ;
        RECT 251.400 214.350 252.600 216.000 ;
        RECT 259.950 215.100 262.050 220.050 ;
        RECT 265.950 215.100 268.050 217.200 ;
        RECT 272.400 216.600 273.450 220.950 ;
        RECT 241.950 211.950 244.050 214.050 ;
        RECT 244.950 211.950 247.050 214.050 ;
        RECT 247.950 211.950 250.050 214.050 ;
        RECT 250.950 211.950 253.050 214.050 ;
        RECT 242.400 209.400 243.600 211.650 ;
        RECT 248.400 209.400 249.600 211.650 ;
        RECT 211.950 202.950 214.050 205.050 ;
        RECT 217.950 202.950 220.050 205.050 ;
        RECT 232.950 202.950 235.050 205.050 ;
        RECT 211.950 196.950 214.050 199.050 ;
        RECT 208.950 184.950 211.050 187.050 ;
        RECT 199.950 182.100 202.050 184.200 ;
        RECT 212.400 183.450 213.450 196.950 ;
        RECT 217.950 190.950 220.050 193.050 ;
        RECT 238.950 190.950 241.050 193.050 ;
        RECT 209.400 182.400 213.450 183.450 ;
        RECT 218.400 183.600 219.450 190.950 ;
        RECT 235.950 184.950 238.050 187.050 ;
        RECT 200.400 181.350 201.600 182.100 ;
        RECT 199.950 178.950 202.050 181.050 ;
        RECT 202.950 178.950 205.050 181.050 ;
        RECT 203.400 177.900 204.600 178.650 ;
        RECT 209.400 178.050 210.450 182.400 ;
        RECT 218.400 181.350 219.600 183.600 ;
        RECT 223.950 182.100 226.050 184.200 ;
        RECT 224.400 181.350 225.600 182.100 ;
        RECT 232.950 181.950 235.050 184.050 ;
        RECT 217.950 178.950 220.050 181.050 ;
        RECT 220.950 178.950 223.050 181.050 ;
        RECT 223.950 178.950 226.050 181.050 ;
        RECT 226.950 178.950 229.050 181.050 ;
        RECT 202.950 175.800 205.050 177.900 ;
        RECT 208.950 175.950 211.050 178.050 ;
        RECT 221.400 177.000 222.600 178.650 ;
        RECT 220.950 172.950 223.050 177.000 ;
        RECT 227.400 176.400 228.600 178.650 ;
        RECT 199.950 169.950 202.050 172.050 ;
        RECT 187.950 139.950 190.050 142.050 ;
        RECT 193.950 140.100 196.050 142.200 ;
        RECT 169.950 137.100 172.050 139.200 ;
        RECT 175.950 137.100 178.050 139.200 ;
        RECT 184.950 137.100 187.050 139.200 ;
        RECT 170.400 136.350 171.600 137.100 ;
        RECT 176.400 136.350 177.600 137.100 ;
        RECT 169.950 133.950 172.050 136.050 ;
        RECT 172.950 133.950 175.050 136.050 ;
        RECT 175.950 133.950 178.050 136.050 ;
        RECT 178.950 133.950 181.050 136.050 ;
        RECT 173.400 131.400 174.600 133.650 ;
        RECT 179.400 131.400 180.600 133.650 ;
        RECT 173.400 127.050 174.450 131.400 ;
        RECT 172.950 124.950 175.050 127.050 ;
        RECT 163.950 112.950 166.050 115.050 ;
        RECT 175.950 112.950 178.050 115.050 ;
        RECT 149.400 105.450 150.450 109.950 ;
        RECT 158.400 109.200 159.600 111.450 ;
        RECT 154.500 107.100 156.600 109.200 ;
        RECT 152.400 105.450 153.600 105.600 ;
        RECT 149.400 104.400 153.600 105.450 ;
        RECT 152.400 103.350 153.600 104.400 ;
        RECT 152.100 100.950 154.200 103.050 ;
        RECT 155.100 102.000 156.000 107.100 ;
        RECT 157.800 106.800 159.900 108.900 ;
        RECT 164.400 107.400 166.500 109.500 ;
        RECT 162.000 105.000 164.100 105.900 ;
        RECT 156.900 103.800 164.100 105.000 ;
        RECT 156.900 102.900 159.000 103.800 ;
        RECT 162.000 102.000 164.100 102.900 ;
        RECT 155.100 101.100 164.100 102.000 ;
        RECT 145.950 97.800 148.050 99.900 ;
        RECT 142.950 94.950 145.050 97.050 ;
        RECT 155.100 94.500 156.000 101.100 ;
        RECT 162.000 100.800 164.100 101.100 ;
        RECT 157.800 97.950 159.900 100.050 ;
        RECT 158.400 95.400 159.600 97.650 ;
        RECT 165.000 94.800 165.900 107.400 ;
        RECT 166.800 100.950 168.900 103.050 ;
        RECT 167.400 99.900 168.600 100.650 ;
        RECT 166.950 97.800 169.050 99.900 ;
        RECT 176.400 97.050 177.450 112.950 ;
        RECT 179.400 99.450 180.450 131.400 ;
        RECT 185.400 129.450 186.450 137.100 ;
        RECT 188.400 133.050 189.450 139.950 ;
        RECT 193.950 136.950 196.050 139.050 ;
        RECT 200.400 138.600 201.450 169.950 ;
        RECT 227.400 169.050 228.450 176.400 ;
        RECT 226.950 166.950 229.050 169.050 ;
        RECT 233.400 166.050 234.450 181.950 ;
        RECT 236.400 177.900 237.450 184.950 ;
        RECT 239.400 183.450 240.450 190.950 ;
        RECT 242.400 187.050 243.450 209.400 ;
        RECT 248.400 205.050 249.450 209.400 ;
        RECT 247.950 202.950 250.050 205.050 ;
        RECT 260.400 199.050 261.450 215.100 ;
        RECT 266.400 214.350 267.600 215.100 ;
        RECT 272.400 214.350 273.600 216.600 ;
        RECT 283.950 215.100 286.050 217.200 ;
        RECT 293.400 216.450 294.600 216.600 ;
        RECT 287.400 215.400 294.600 216.450 ;
        RECT 265.950 211.950 268.050 214.050 ;
        RECT 268.950 211.950 271.050 214.050 ;
        RECT 271.950 211.950 274.050 214.050 ;
        RECT 274.950 211.950 277.050 214.050 ;
        RECT 269.400 209.400 270.600 211.650 ;
        RECT 275.400 210.900 276.600 211.650 ;
        RECT 284.400 211.050 285.450 215.100 ;
        RECT 287.400 211.050 288.450 215.400 ;
        RECT 293.400 214.350 294.600 215.400 ;
        RECT 298.950 215.100 301.050 220.050 ;
        RECT 299.400 214.350 300.600 215.100 ;
        RECT 292.950 211.950 295.050 214.050 ;
        RECT 295.950 211.950 298.050 214.050 ;
        RECT 298.950 211.950 301.050 214.050 ;
        RECT 301.950 211.950 304.050 214.050 ;
        RECT 269.400 205.050 270.450 209.400 ;
        RECT 274.950 208.800 277.050 210.900 ;
        RECT 277.950 208.950 280.050 211.050 ;
        RECT 283.950 208.950 286.050 211.050 ;
        RECT 286.950 208.950 289.050 211.050 ;
        RECT 296.400 209.400 297.600 211.650 ;
        RECT 302.400 209.400 303.600 211.650 ;
        RECT 311.400 210.900 312.450 226.950 ;
        RECT 347.400 226.050 348.450 259.950 ;
        RECT 355.950 256.950 358.050 259.050 ;
        RECT 358.950 256.950 361.050 259.050 ;
        RECT 361.950 256.950 364.050 259.050 ;
        RECT 364.950 256.950 367.050 259.050 ;
        RECT 367.950 256.950 370.050 259.050 ;
        RECT 362.400 254.400 363.600 256.650 ;
        RECT 362.400 235.050 363.450 254.400 ;
        RECT 361.950 232.950 364.050 235.050 ;
        RECT 370.950 232.950 373.050 235.050 ;
        RECT 364.950 226.950 367.050 229.050 ;
        RECT 346.950 223.950 349.050 226.050 ;
        RECT 352.950 223.950 355.050 226.050 ;
        RECT 319.950 216.000 322.050 220.050 ;
        RECT 320.400 214.350 321.600 216.000 ;
        RECT 325.950 215.100 328.050 217.200 ;
        RECT 334.950 215.100 337.050 217.200 ;
        RECT 340.950 215.100 343.050 217.200 ;
        RECT 326.400 214.350 327.600 215.100 ;
        RECT 316.950 211.950 319.050 214.050 ;
        RECT 319.950 211.950 322.050 214.050 ;
        RECT 322.950 211.950 325.050 214.050 ;
        RECT 325.950 211.950 328.050 214.050 ;
        RECT 268.950 202.950 271.050 205.050 ;
        RECT 259.950 196.950 262.050 199.050 ;
        RECT 241.950 184.950 244.050 187.050 ;
        RECT 259.950 184.950 262.050 187.050 ;
        RECT 242.400 183.450 243.600 183.600 ;
        RECT 239.400 182.400 243.600 183.450 ;
        RECT 242.400 181.350 243.600 182.400 ;
        RECT 247.950 182.100 250.050 184.200 ;
        RECT 248.400 181.350 249.600 182.100 ;
        RECT 256.950 181.950 259.050 184.050 ;
        RECT 241.950 178.950 244.050 181.050 ;
        RECT 244.950 178.950 247.050 181.050 ;
        RECT 247.950 178.950 250.050 181.050 ;
        RECT 250.950 178.950 253.050 181.050 ;
        RECT 245.400 177.900 246.600 178.650 ;
        RECT 235.950 175.800 238.050 177.900 ;
        RECT 244.950 175.800 247.050 177.900 ;
        RECT 251.400 177.000 252.600 178.650 ;
        RECT 250.950 172.950 253.050 177.000 ;
        RECT 232.950 163.950 235.050 166.050 ;
        RECT 253.950 154.950 256.050 157.050 ;
        RECT 247.950 142.950 250.050 145.050 ;
        RECT 207.000 138.600 211.050 139.050 ;
        RECT 194.400 136.350 195.600 136.950 ;
        RECT 200.400 136.350 201.600 138.600 ;
        RECT 206.400 136.950 211.050 138.600 ;
        RECT 211.950 136.950 214.050 139.050 ;
        RECT 214.950 136.950 217.050 139.050 ;
        RECT 220.950 137.100 223.050 139.200 ;
        RECT 232.950 137.100 235.050 139.200 ;
        RECT 241.950 137.100 244.050 139.200 ;
        RECT 248.400 138.600 249.450 142.950 ;
        RECT 206.400 136.350 207.600 136.950 ;
        RECT 193.950 133.950 196.050 136.050 ;
        RECT 196.950 133.950 199.050 136.050 ;
        RECT 199.950 133.950 202.050 136.050 ;
        RECT 202.950 133.950 205.050 136.050 ;
        RECT 205.950 133.950 208.050 136.050 ;
        RECT 187.950 130.950 190.050 133.050 ;
        RECT 197.400 131.400 198.600 133.650 ;
        RECT 203.400 132.000 204.600 133.650 ;
        RECT 185.400 129.000 189.450 129.450 ;
        RECT 185.400 128.400 190.050 129.000 ;
        RECT 187.950 124.950 190.050 128.400 ;
        RECT 197.400 123.450 198.450 131.400 ;
        RECT 202.950 127.950 205.050 132.000 ;
        RECT 208.950 130.950 211.050 133.050 ;
        RECT 197.400 122.400 201.450 123.450 ;
        RECT 196.950 118.950 199.050 121.050 ;
        RECT 184.950 104.100 187.050 106.200 ;
        RECT 185.400 103.350 186.600 104.100 ;
        RECT 182.100 100.950 184.200 103.050 ;
        RECT 185.400 100.950 187.500 103.050 ;
        RECT 190.800 100.950 192.900 103.050 ;
        RECT 182.400 99.450 183.600 100.650 ;
        RECT 191.400 99.900 192.600 100.650 ;
        RECT 179.400 98.400 183.600 99.450 ;
        RECT 190.950 97.800 193.050 99.900 ;
        RECT 175.950 94.950 178.050 97.050 ;
        RECT 155.100 92.400 157.200 94.500 ;
        RECT 164.100 92.700 166.200 94.800 ;
        RECT 118.950 67.950 121.050 70.050 ;
        RECT 124.950 67.950 127.050 70.050 ;
        RECT 119.400 54.900 120.450 67.950 ;
        RECT 197.400 66.450 198.450 118.950 ;
        RECT 200.400 115.050 201.450 122.400 ;
        RECT 199.950 112.950 202.050 115.050 ;
        RECT 200.400 99.900 201.450 112.950 ;
        RECT 209.400 106.200 210.450 130.950 ;
        RECT 212.400 130.050 213.450 136.950 ;
        RECT 215.400 132.450 216.450 136.950 ;
        RECT 221.400 136.350 222.600 137.100 ;
        RECT 220.950 133.950 223.050 136.050 ;
        RECT 223.950 133.950 226.050 136.050 ;
        RECT 215.400 131.400 219.450 132.450 ;
        RECT 211.950 127.950 214.050 130.050 ;
        RECT 208.950 104.100 211.050 106.200 ;
        RECT 209.400 103.350 210.600 104.100 ;
        RECT 205.950 100.950 208.050 103.050 ;
        RECT 208.950 100.950 211.050 103.050 ;
        RECT 211.950 100.950 214.050 103.050 ;
        RECT 199.950 97.800 202.050 99.900 ;
        RECT 206.400 98.400 207.600 100.650 ;
        RECT 212.400 99.450 213.600 100.650 ;
        RECT 214.950 99.450 217.050 100.050 ;
        RECT 212.400 98.400 217.050 99.450 ;
        RECT 206.400 94.050 207.450 98.400 ;
        RECT 214.950 97.950 217.050 98.400 ;
        RECT 205.950 91.950 208.050 94.050 ;
        RECT 194.400 65.400 198.450 66.450 ;
        RECT 177.000 63.450 181.050 64.050 ;
        RECT 176.400 61.950 181.050 63.450 ;
        RECT 124.950 59.100 127.050 61.200 ;
        RECT 133.950 59.100 136.050 61.200 ;
        RECT 145.950 59.100 148.050 61.200 ;
        RECT 152.400 60.450 153.600 60.600 ;
        RECT 152.400 59.400 159.450 60.450 ;
        RECT 125.400 58.350 126.600 59.100 ;
        RECT 124.950 55.950 127.050 58.050 ;
        RECT 127.950 55.950 130.050 58.050 ;
        RECT 118.950 52.800 121.050 54.900 ;
        RECT 128.400 54.000 129.600 55.650 ;
        RECT 115.950 49.950 118.050 52.050 ;
        RECT 127.950 49.950 130.050 54.000 ;
        RECT 127.950 43.950 130.050 46.050 ;
        RECT 121.950 37.950 124.050 40.050 ;
        RECT 103.950 34.950 106.050 37.050 ;
        RECT 112.950 34.950 115.050 37.050 ;
        RECT 70.950 28.950 73.050 31.050 ;
        RECT 79.950 30.450 84.000 31.050 ;
        RECT 79.950 28.950 84.450 30.450 ;
        RECT 62.400 25.350 63.600 27.600 ;
        RECT 58.950 22.950 61.050 25.050 ;
        RECT 61.950 22.950 64.050 25.050 ;
        RECT 64.950 22.950 67.050 25.050 ;
        RECT 59.400 21.900 60.600 22.650 ;
        RECT 65.400 21.900 66.600 22.650 ;
        RECT 71.400 21.900 72.450 28.950 ;
        RECT 73.950 25.950 76.050 28.050 ;
        RECT 83.400 27.600 84.450 28.950 ;
        RECT 74.400 21.900 75.450 25.950 ;
        RECT 83.400 25.350 84.600 27.600 ;
        RECT 103.950 26.100 106.050 28.200 ;
        RECT 104.400 25.350 105.600 26.100 ;
        RECT 79.950 22.950 82.050 25.050 ;
        RECT 82.950 22.950 85.050 25.050 ;
        RECT 85.950 22.950 88.050 25.050 ;
        RECT 100.950 22.950 103.050 25.050 ;
        RECT 103.950 22.950 106.050 25.050 ;
        RECT 106.950 22.950 109.050 25.050 ;
        RECT 80.400 21.900 81.600 22.650 ;
        RECT 58.950 19.800 61.050 21.900 ;
        RECT 64.950 19.800 67.050 21.900 ;
        RECT 70.800 19.800 72.900 21.900 ;
        RECT 73.950 19.800 76.050 21.900 ;
        RECT 79.950 19.800 82.050 21.900 ;
        RECT 86.400 20.400 87.600 22.650 ;
        RECT 101.400 21.000 102.600 22.650 ;
        RECT 107.400 21.900 108.600 22.650 ;
        RECT 113.400 21.900 114.450 34.950 ;
        RECT 122.400 28.200 123.450 37.950 ;
        RECT 121.950 26.100 124.050 28.200 ;
        RECT 128.400 27.600 129.450 43.950 ;
        RECT 134.400 40.050 135.450 59.100 ;
        RECT 146.400 58.350 147.600 59.100 ;
        RECT 152.400 58.350 153.600 59.400 ;
        RECT 145.950 55.950 148.050 58.050 ;
        RECT 148.950 55.950 151.050 58.050 ;
        RECT 151.950 55.950 154.050 58.050 ;
        RECT 149.400 54.900 150.600 55.650 ;
        RECT 148.950 52.800 151.050 54.900 ;
        RECT 133.950 37.950 136.050 40.050 ;
        RECT 122.400 25.350 123.600 26.100 ;
        RECT 128.400 25.350 129.600 27.600 ;
        RECT 136.950 26.100 139.050 28.200 ;
        RECT 146.400 27.450 147.600 27.600 ;
        RECT 149.400 27.450 150.450 52.800 ;
        RECT 158.400 46.050 159.450 59.400 ;
        RECT 166.950 59.100 169.050 61.200 ;
        RECT 176.400 60.600 177.450 61.950 ;
        RECT 194.400 61.200 195.450 65.400 ;
        RECT 167.400 58.350 168.600 59.100 ;
        RECT 176.400 58.350 177.600 60.600 ;
        RECT 187.950 58.950 190.050 61.050 ;
        RECT 193.950 59.100 196.050 61.200 ;
        RECT 199.950 60.000 202.050 64.050 ;
        RECT 167.100 55.950 169.200 58.050 ;
        RECT 170.400 55.950 172.500 58.050 ;
        RECT 175.800 55.950 177.900 58.050 ;
        RECT 170.400 53.400 171.600 55.650 ;
        RECT 170.400 46.050 171.450 53.400 ;
        RECT 157.950 43.950 160.050 46.050 ;
        RECT 169.950 43.950 172.050 46.050 ;
        RECT 166.950 34.950 169.050 37.050 ;
        RECT 146.400 26.400 150.450 27.450 ;
        RECT 121.950 22.950 124.050 25.050 ;
        RECT 124.950 22.950 127.050 25.050 ;
        RECT 127.950 22.950 130.050 25.050 ;
        RECT 125.400 21.900 126.600 22.650 ;
        RECT 137.400 22.050 138.450 26.100 ;
        RECT 146.400 25.350 147.600 26.400 ;
        RECT 160.950 26.100 163.050 28.200 ;
        RECT 167.400 27.600 168.450 34.950 ;
        RECT 188.400 28.200 189.450 58.950 ;
        RECT 194.400 58.350 195.600 59.100 ;
        RECT 200.400 58.350 201.600 60.000 ;
        RECT 193.950 55.950 196.050 58.050 ;
        RECT 196.950 55.950 199.050 58.050 ;
        RECT 199.950 55.950 202.050 58.050 ;
        RECT 202.950 55.950 205.050 58.050 ;
        RECT 197.400 54.900 198.600 55.650 ;
        RECT 196.950 52.800 199.050 54.900 ;
        RECT 203.400 53.400 204.600 55.650 ;
        RECT 203.400 49.050 204.450 53.400 ;
        RECT 208.950 52.950 211.050 55.050 ;
        RECT 215.400 54.450 216.450 97.950 ;
        RECT 218.400 82.050 219.450 131.400 ;
        RECT 224.400 131.400 225.600 133.650 ;
        RECT 224.400 124.050 225.450 131.400 ;
        RECT 233.400 124.050 234.450 137.100 ;
        RECT 242.400 136.350 243.600 137.100 ;
        RECT 248.400 136.350 249.600 138.600 ;
        RECT 238.950 133.950 241.050 136.050 ;
        RECT 241.950 133.950 244.050 136.050 ;
        RECT 244.950 133.950 247.050 136.050 ;
        RECT 247.950 133.950 250.050 136.050 ;
        RECT 239.400 131.400 240.600 133.650 ;
        RECT 245.400 132.900 246.600 133.650 ;
        RECT 254.400 132.900 255.450 154.950 ;
        RECT 257.400 142.050 258.450 181.950 ;
        RECT 260.400 169.050 261.450 184.950 ;
        RECT 268.950 183.000 271.050 187.050 ;
        RECT 269.400 181.350 270.600 183.000 ;
        RECT 274.950 181.950 277.050 184.050 ;
        RECT 265.950 178.950 268.050 181.050 ;
        RECT 268.950 178.950 271.050 181.050 ;
        RECT 266.400 177.900 267.600 178.650 ;
        RECT 265.950 175.800 268.050 177.900 ;
        RECT 266.400 175.050 267.450 175.800 ;
        RECT 262.950 173.400 267.450 175.050 ;
        RECT 262.950 172.950 267.000 173.400 ;
        RECT 259.950 166.950 262.050 169.050 ;
        RECT 265.950 157.950 268.050 160.050 ;
        RECT 256.950 139.950 259.050 142.050 ;
        RECT 266.400 138.600 267.450 157.950 ;
        RECT 275.400 151.050 276.450 181.950 ;
        RECT 278.400 178.050 279.450 208.950 ;
        RECT 296.400 202.050 297.450 209.400 ;
        RECT 295.950 199.950 298.050 202.050 ;
        RECT 298.950 187.950 301.050 190.050 ;
        RECT 283.950 182.100 286.050 184.200 ;
        RECT 289.950 182.100 292.050 184.200 ;
        RECT 284.400 181.350 285.600 182.100 ;
        RECT 290.400 181.350 291.600 182.100 ;
        RECT 283.950 178.950 286.050 181.050 ;
        RECT 286.950 178.950 289.050 181.050 ;
        RECT 289.950 178.950 292.050 181.050 ;
        RECT 292.950 178.950 295.050 181.050 ;
        RECT 277.950 175.950 280.050 178.050 ;
        RECT 287.400 176.400 288.600 178.650 ;
        RECT 293.400 177.900 294.600 178.650 ;
        RECT 287.400 166.050 288.450 176.400 ;
        RECT 292.950 175.800 295.050 177.900 ;
        RECT 286.950 163.950 289.050 166.050 ;
        RECT 299.400 160.050 300.450 187.950 ;
        RECT 302.400 184.200 303.450 209.400 ;
        RECT 310.950 208.800 313.050 210.900 ;
        RECT 317.400 209.400 318.600 211.650 ;
        RECT 323.400 210.900 324.600 211.650 ;
        RECT 335.400 211.050 336.450 215.100 ;
        RECT 341.400 214.350 342.600 215.100 ;
        RECT 340.950 211.950 343.050 214.050 ;
        RECT 343.950 211.950 346.050 214.050 ;
        RECT 311.400 202.050 312.450 208.800 ;
        RECT 310.950 199.950 313.050 202.050 ;
        RECT 317.400 190.050 318.450 209.400 ;
        RECT 322.950 208.800 325.050 210.900 ;
        RECT 328.950 208.950 331.050 211.050 ;
        RECT 334.950 208.950 337.050 211.050 ;
        RECT 337.950 208.950 340.050 211.050 ;
        RECT 344.400 210.900 345.600 211.650 ;
        RECT 353.400 210.900 354.450 223.950 ;
        RECT 365.400 216.600 366.450 226.950 ;
        RECT 371.400 220.200 372.450 232.950 ;
        RECT 370.950 218.100 373.050 220.200 ;
        RECT 365.400 214.350 366.600 216.600 ;
        RECT 370.950 214.950 373.050 217.050 ;
        RECT 374.400 216.450 375.450 277.950 ;
        RECT 383.400 268.050 384.450 287.400 ;
        RECT 394.950 286.800 397.050 288.900 ;
        RECT 400.950 286.800 403.050 288.900 ;
        RECT 407.400 287.400 408.600 289.650 ;
        RECT 425.400 288.900 426.600 289.650 ;
        RECT 382.950 265.950 385.050 268.050 ;
        RECT 397.950 265.950 400.050 268.050 ;
        RECT 376.950 260.100 379.050 262.200 ;
        RECT 385.950 260.100 388.050 262.200 ;
        RECT 391.950 260.100 394.050 262.200 ;
        RECT 377.400 232.050 378.450 260.100 ;
        RECT 386.400 259.350 387.600 260.100 ;
        RECT 392.400 259.350 393.600 260.100 ;
        RECT 382.950 256.950 385.050 259.050 ;
        RECT 385.950 256.950 388.050 259.050 ;
        RECT 388.950 256.950 391.050 259.050 ;
        RECT 391.950 256.950 394.050 259.050 ;
        RECT 383.400 254.400 384.600 256.650 ;
        RECT 389.400 254.400 390.600 256.650 ;
        RECT 383.400 250.050 384.450 254.400 ;
        RECT 382.950 247.950 385.050 250.050 ;
        RECT 389.400 247.050 390.450 254.400 ;
        RECT 398.400 250.050 399.450 265.950 ;
        RECT 407.400 262.200 408.450 287.400 ;
        RECT 424.950 286.800 427.050 288.900 ;
        RECT 400.950 259.950 403.050 262.050 ;
        RECT 406.950 260.100 409.050 262.200 ;
        RECT 397.950 247.950 400.050 250.050 ;
        RECT 388.950 244.950 391.050 247.050 ;
        RECT 389.400 235.050 390.450 244.950 ;
        RECT 401.400 241.050 402.450 259.950 ;
        RECT 407.400 259.350 408.600 260.100 ;
        RECT 418.950 259.950 421.050 262.050 ;
        RECT 406.950 256.950 409.050 259.050 ;
        RECT 409.950 256.950 412.050 259.050 ;
        RECT 410.400 254.400 411.600 256.650 ;
        RECT 403.950 247.950 406.050 250.050 ;
        RECT 400.950 238.950 403.050 241.050 ;
        RECT 382.950 232.950 385.050 235.050 ;
        RECT 388.950 232.950 391.050 235.050 ;
        RECT 376.950 229.950 379.050 232.050 ;
        RECT 379.950 223.950 382.050 226.050 ;
        RECT 374.400 215.400 378.450 216.450 ;
        RECT 371.400 214.350 372.600 214.950 ;
        RECT 361.950 211.950 364.050 214.050 ;
        RECT 364.950 211.950 367.050 214.050 ;
        RECT 367.950 211.950 370.050 214.050 ;
        RECT 370.950 211.950 373.050 214.050 ;
        RECT 316.950 187.950 319.050 190.050 ;
        RECT 322.950 184.950 325.050 187.050 ;
        RECT 301.950 182.100 304.050 184.200 ;
        RECT 310.950 182.100 313.050 184.200 ;
        RECT 316.950 182.100 319.050 184.200 ;
        RECT 311.400 181.350 312.600 182.100 ;
        RECT 317.400 181.350 318.600 182.100 ;
        RECT 323.400 181.050 324.450 184.950 ;
        RECT 325.950 181.950 328.050 184.050 ;
        RECT 307.950 178.950 310.050 181.050 ;
        RECT 310.950 178.950 313.050 181.050 ;
        RECT 313.950 178.950 316.050 181.050 ;
        RECT 316.950 178.950 319.050 181.050 ;
        RECT 322.950 178.950 325.050 181.050 ;
        RECT 308.400 176.400 309.600 178.650 ;
        RECT 314.400 177.900 315.600 178.650 ;
        RECT 308.400 166.050 309.450 176.400 ;
        RECT 313.950 175.800 316.050 177.900 ;
        RECT 307.950 163.950 310.050 166.050 ;
        RECT 280.950 157.950 283.050 160.050 ;
        RECT 298.950 157.950 301.050 160.050 ;
        RECT 274.950 148.950 277.050 151.050 ;
        RECT 277.950 145.950 280.050 148.050 ;
        RECT 271.950 142.950 277.050 145.050 ;
        RECT 278.400 139.200 279.450 145.950 ;
        RECT 266.400 136.350 267.600 138.600 ;
        RECT 271.950 137.100 274.050 139.200 ;
        RECT 277.950 137.100 280.050 139.200 ;
        RECT 272.400 136.350 273.600 137.100 ;
        RECT 265.950 133.950 268.050 136.050 ;
        RECT 268.950 133.950 271.050 136.050 ;
        RECT 271.950 133.950 274.050 136.050 ;
        RECT 239.400 127.050 240.450 131.400 ;
        RECT 244.950 130.800 247.050 132.900 ;
        RECT 253.950 130.800 256.050 132.900 ;
        RECT 269.400 131.400 270.600 133.650 ;
        RECT 278.400 133.050 279.450 137.100 ;
        RECT 238.950 124.950 241.050 127.050 ;
        RECT 223.950 121.950 226.050 124.050 ;
        RECT 232.950 121.950 235.050 124.050 ;
        RECT 253.950 121.950 256.050 124.050 ;
        RECT 235.950 112.950 238.050 115.050 ;
        RECT 223.950 104.100 226.050 106.200 ;
        RECT 229.950 104.100 232.050 106.200 ;
        RECT 236.400 105.600 237.450 112.950 ;
        RECT 224.400 100.050 225.450 104.100 ;
        RECT 230.400 103.350 231.600 104.100 ;
        RECT 236.400 103.350 237.600 105.600 ;
        RECT 247.950 104.100 250.050 106.200 ;
        RECT 254.400 105.600 255.450 121.950 ;
        RECT 269.400 121.050 270.450 131.400 ;
        RECT 277.950 130.950 280.050 133.050 ;
        RECT 281.400 132.900 282.450 157.950 ;
        RECT 307.950 148.950 310.050 151.050 ;
        RECT 319.950 148.950 322.050 151.050 ;
        RECT 283.950 142.950 289.050 145.050 ;
        RECT 289.950 138.000 292.050 142.050 ;
        RECT 290.400 136.350 291.600 138.000 ;
        RECT 295.950 137.100 298.050 139.200 ;
        RECT 296.400 136.350 297.600 137.100 ;
        RECT 286.950 133.950 289.050 136.050 ;
        RECT 289.950 133.950 292.050 136.050 ;
        RECT 292.950 133.950 295.050 136.050 ;
        RECT 295.950 133.950 298.050 136.050 ;
        RECT 287.400 133.050 288.600 133.650 ;
        RECT 280.950 130.800 283.050 132.900 ;
        RECT 283.950 131.400 288.600 133.050 ;
        RECT 293.400 132.900 294.600 133.650 ;
        RECT 283.950 130.950 288.000 131.400 ;
        RECT 292.950 130.800 295.050 132.900 ;
        RECT 308.400 127.050 309.450 148.950 ;
        RECT 313.950 138.000 316.050 142.050 ;
        RECT 320.400 139.200 321.450 148.950 ;
        RECT 314.400 136.350 315.600 138.000 ;
        RECT 319.950 137.100 322.050 139.200 ;
        RECT 326.400 138.450 327.450 181.950 ;
        RECT 329.400 169.050 330.450 208.950 ;
        RECT 338.400 187.050 339.450 208.950 ;
        RECT 343.950 208.800 346.050 210.900 ;
        RECT 352.950 208.800 355.050 210.900 ;
        RECT 362.400 210.000 363.600 211.650 ;
        RECT 337.950 184.950 340.050 187.050 ;
        RECT 335.100 178.950 337.200 181.050 ;
        RECT 340.500 178.950 342.600 181.050 ;
        RECT 343.800 178.950 345.900 181.050 ;
        RECT 344.400 177.900 345.600 178.650 ;
        RECT 343.950 175.800 346.050 177.900 ;
        RECT 328.950 166.950 331.050 169.050 ;
        RECT 353.400 151.050 354.450 208.800 ;
        RECT 361.950 205.950 364.050 210.000 ;
        RECT 368.400 209.400 369.600 211.650 ;
        RECT 368.400 202.050 369.450 209.400 ;
        RECT 373.950 208.950 376.050 211.050 ;
        RECT 377.400 210.900 378.450 215.400 ;
        RECT 367.950 199.950 370.050 202.050 ;
        RECT 358.950 182.100 361.050 184.200 ;
        RECT 364.950 182.100 367.050 184.200 ;
        RECT 359.400 178.050 360.450 182.100 ;
        RECT 365.400 181.350 366.600 182.100 ;
        RECT 362.100 178.950 364.200 181.050 ;
        RECT 365.400 178.950 367.500 181.050 ;
        RECT 370.800 178.950 372.900 181.050 ;
        RECT 358.950 175.950 361.050 178.050 ;
        RECT 362.400 176.400 363.600 178.650 ;
        RECT 371.400 176.400 372.600 178.650 ;
        RECT 352.950 148.950 355.050 151.050 ;
        RECT 337.950 145.950 340.050 148.050 ;
        RECT 328.950 142.950 334.050 145.050 ;
        RECT 338.400 138.600 339.450 145.950 ;
        RECT 340.950 142.950 346.050 145.050 ;
        RECT 326.400 137.400 330.450 138.450 ;
        RECT 320.400 136.350 321.600 137.100 ;
        RECT 313.950 133.950 316.050 136.050 ;
        RECT 316.950 133.950 319.050 136.050 ;
        RECT 319.950 133.950 322.050 136.050 ;
        RECT 322.950 133.950 325.050 136.050 ;
        RECT 317.400 132.900 318.600 133.650 ;
        RECT 316.950 130.800 319.050 132.900 ;
        RECT 323.400 131.400 324.600 133.650 ;
        RECT 307.950 124.950 310.050 127.050 ;
        RECT 268.950 118.950 271.050 121.050 ;
        RECT 323.400 118.050 324.450 131.400 ;
        RECT 322.950 115.950 325.050 118.050 ;
        RECT 289.950 112.950 292.050 115.050 ;
        RECT 229.950 100.950 232.050 103.050 ;
        RECT 232.950 100.950 235.050 103.050 ;
        RECT 235.950 100.950 238.050 103.050 ;
        RECT 238.950 100.950 241.050 103.050 ;
        RECT 223.950 97.950 226.050 100.050 ;
        RECT 233.400 98.400 234.600 100.650 ;
        RECT 239.400 98.400 240.600 100.650 ;
        RECT 233.400 94.050 234.450 98.400 ;
        RECT 239.400 94.050 240.450 98.400 ;
        RECT 241.950 97.800 244.050 99.900 ;
        RECT 232.950 91.950 235.050 94.050 ;
        RECT 238.950 91.950 241.050 94.050 ;
        RECT 217.950 79.950 220.050 82.050 ;
        RECT 233.400 69.450 234.450 91.950 ;
        RECT 233.400 68.400 237.450 69.450 ;
        RECT 220.800 64.500 222.900 66.600 ;
        RECT 218.100 55.950 220.200 58.050 ;
        RECT 221.100 57.300 222.300 64.500 ;
        RECT 224.400 61.350 225.600 63.600 ;
        RECT 230.400 63.300 232.500 65.400 ;
        RECT 224.100 58.950 226.200 61.050 ;
        RECT 227.100 59.700 229.200 61.800 ;
        RECT 227.100 57.300 228.000 59.700 ;
        RECT 221.100 56.100 228.000 57.300 ;
        RECT 218.400 54.450 219.600 55.650 ;
        RECT 215.400 53.400 219.600 54.450 ;
        RECT 202.950 46.950 205.050 49.050 ;
        RECT 161.400 25.350 162.600 26.100 ;
        RECT 167.400 25.350 168.600 27.600 ;
        RECT 187.950 26.100 190.050 28.200 ;
        RECT 188.400 25.350 189.600 26.100 ;
        RECT 196.950 25.950 199.050 28.050 ;
        RECT 209.400 27.600 210.450 52.950 ;
        RECT 215.400 27.600 216.450 53.400 ;
        RECT 221.100 50.700 222.000 56.100 ;
        RECT 222.900 54.300 225.000 55.200 ;
        RECT 230.700 54.300 231.600 63.300 ;
        RECT 233.400 60.450 234.600 60.600 ;
        RECT 236.400 60.450 237.450 68.400 ;
        RECT 233.400 59.400 237.450 60.450 ;
        RECT 233.400 58.350 234.600 59.400 ;
        RECT 232.800 55.950 234.900 58.050 ;
        RECT 222.900 53.100 231.600 54.300 ;
        RECT 220.800 48.600 222.900 50.700 ;
        RECT 224.100 50.100 226.200 52.200 ;
        RECT 228.000 51.300 230.100 53.100 ;
        RECT 224.400 47.550 225.600 49.800 ;
        RECT 224.400 43.050 225.450 47.550 ;
        RECT 242.400 43.050 243.450 97.800 ;
        RECT 248.400 94.050 249.450 104.100 ;
        RECT 254.400 103.350 255.600 105.600 ;
        RECT 259.950 104.100 262.050 106.200 ;
        RECT 260.400 103.350 261.600 104.100 ;
        RECT 268.950 103.950 271.050 106.050 ;
        RECT 280.950 104.100 283.050 106.200 ;
        RECT 253.950 100.950 256.050 103.050 ;
        RECT 256.950 100.950 259.050 103.050 ;
        RECT 259.950 100.950 262.050 103.050 ;
        RECT 262.950 100.950 265.050 103.050 ;
        RECT 257.400 99.900 258.600 100.650 ;
        RECT 263.400 99.900 264.600 100.650 ;
        RECT 256.950 97.800 259.050 99.900 ;
        RECT 262.950 97.800 265.050 99.900 ;
        RECT 247.950 91.950 250.050 94.050 ;
        RECT 248.400 60.600 249.450 91.950 ;
        RECT 262.950 79.950 265.050 82.050 ;
        RECT 248.400 58.350 249.600 60.600 ;
        RECT 253.950 59.100 256.050 61.200 ;
        RECT 254.400 58.350 255.600 59.100 ;
        RECT 247.950 55.950 250.050 58.050 ;
        RECT 250.950 55.950 253.050 58.050 ;
        RECT 253.950 55.950 256.050 58.050 ;
        RECT 256.950 55.950 259.050 58.050 ;
        RECT 251.400 53.400 252.600 55.650 ;
        RECT 257.400 54.000 258.600 55.650 ;
        RECT 263.400 54.900 264.450 79.950 ;
        RECT 269.400 60.450 270.450 103.950 ;
        RECT 281.400 103.350 282.600 104.100 ;
        RECT 277.950 100.950 280.050 103.050 ;
        RECT 280.950 100.950 283.050 103.050 ;
        RECT 283.950 100.950 286.050 103.050 ;
        RECT 278.400 98.400 279.600 100.650 ;
        RECT 284.400 99.900 285.600 100.650 ;
        RECT 290.400 99.900 291.450 112.950 ;
        RECT 295.950 109.950 298.050 112.050 ;
        RECT 304.950 109.950 307.050 112.050 ;
        RECT 323.850 111.300 325.950 113.400 ;
        RECT 329.400 112.050 330.450 137.400 ;
        RECT 338.400 136.350 339.600 138.600 ;
        RECT 343.950 137.100 346.050 139.200 ;
        RECT 359.400 139.050 360.450 175.950 ;
        RECT 362.400 169.050 363.450 176.400 ;
        RECT 371.400 172.050 372.450 176.400 ;
        RECT 374.400 175.050 375.450 208.950 ;
        RECT 376.950 208.800 379.050 210.900 ;
        RECT 380.400 202.050 381.450 223.950 ;
        RECT 383.400 217.050 384.450 232.950 ;
        RECT 388.950 226.950 391.050 229.050 ;
        RECT 382.950 214.950 385.050 217.050 ;
        RECT 389.400 216.600 390.450 226.950 ;
        RECT 389.400 214.350 390.600 216.600 ;
        RECT 395.400 216.450 396.600 216.600 ;
        RECT 400.950 216.450 403.050 217.200 ;
        RECT 395.400 215.400 403.050 216.450 ;
        RECT 395.400 214.350 396.600 215.400 ;
        RECT 400.950 215.100 403.050 215.400 ;
        RECT 385.950 211.950 388.050 214.050 ;
        RECT 388.950 211.950 391.050 214.050 ;
        RECT 391.950 211.950 394.050 214.050 ;
        RECT 394.950 211.950 397.050 214.050 ;
        RECT 386.400 210.900 387.600 211.650 ;
        RECT 385.950 208.800 388.050 210.900 ;
        RECT 392.400 209.400 393.600 211.650 ;
        RECT 379.950 199.950 382.050 202.050 ;
        RECT 392.400 190.050 393.450 209.400 ;
        RECT 401.400 196.050 402.450 215.100 ;
        RECT 404.400 205.050 405.450 247.950 ;
        RECT 410.400 235.050 411.450 254.400 ;
        RECT 419.400 243.450 420.450 259.950 ;
        RECT 425.100 256.950 427.200 259.050 ;
        RECT 428.400 256.950 430.500 259.050 ;
        RECT 433.800 256.950 435.900 259.050 ;
        RECT 425.400 254.400 426.600 256.650 ;
        RECT 440.400 255.900 441.450 310.950 ;
        RECT 443.400 265.050 444.450 358.950 ;
        RECT 446.400 355.050 447.450 365.400 ;
        RECT 455.400 361.050 456.450 382.950 ;
        RECT 458.400 366.900 459.450 400.950 ;
        RECT 461.400 400.050 462.450 410.400 ;
        RECT 473.400 406.050 474.450 410.400 ;
        RECT 481.950 409.800 484.050 411.900 ;
        RECT 490.950 409.800 493.050 411.900 ;
        RECT 499.950 409.800 502.050 411.900 ;
        RECT 505.950 409.800 508.050 411.900 ;
        RECT 518.250 410.400 519.450 423.300 ;
        RECT 506.400 406.050 507.450 409.800 ;
        RECT 511.950 406.950 514.050 409.050 ;
        RECT 517.350 408.300 519.450 410.400 ;
        RECT 472.950 403.950 475.050 406.050 ;
        RECT 505.950 403.950 508.050 406.050 ;
        RECT 460.950 397.950 463.050 400.050 ;
        RECT 512.400 394.050 513.450 406.950 ;
        RECT 518.250 401.700 519.450 408.300 ;
        RECT 517.350 399.600 519.450 401.700 ;
        RECT 511.950 391.950 514.050 394.050 ;
        RECT 511.950 385.950 514.050 388.050 ;
        RECT 491.100 376.500 493.200 378.600 ;
        RECT 463.950 372.000 466.050 376.050 ;
        RECT 464.400 370.350 465.600 372.000 ;
        RECT 472.950 371.100 475.050 373.200 ;
        RECT 473.400 370.350 474.600 371.100 ;
        RECT 464.100 367.950 466.200 370.050 ;
        RECT 469.500 367.950 471.600 370.050 ;
        RECT 472.800 367.950 474.900 370.050 ;
        RECT 488.100 367.950 490.200 370.050 ;
        RECT 491.100 369.900 492.000 376.500 ;
        RECT 500.100 376.200 502.200 378.300 ;
        RECT 494.400 373.350 495.600 375.600 ;
        RECT 493.800 370.950 495.900 373.050 ;
        RECT 498.000 369.900 500.100 370.200 ;
        RECT 491.100 369.000 500.100 369.900 ;
        RECT 470.400 366.900 471.600 367.650 ;
        RECT 457.950 364.800 460.050 366.900 ;
        RECT 469.950 364.800 472.050 366.900 ;
        RECT 488.400 366.450 489.600 367.650 ;
        RECT 485.400 365.400 489.600 366.450 ;
        RECT 454.950 358.950 457.050 361.050 ;
        RECT 445.950 352.950 448.050 355.050 ;
        RECT 463.950 352.950 466.050 355.050 ;
        RECT 451.950 343.950 454.050 346.050 ;
        RECT 452.400 339.600 453.450 343.950 ;
        RECT 452.400 337.350 453.600 339.600 ;
        RECT 457.950 338.100 460.050 340.200 ;
        RECT 458.400 337.350 459.600 338.100 ;
        RECT 448.950 334.950 451.050 337.050 ;
        RECT 451.950 334.950 454.050 337.050 ;
        RECT 454.950 334.950 457.050 337.050 ;
        RECT 457.950 334.950 460.050 337.050 ;
        RECT 449.400 333.000 450.600 334.650 ;
        RECT 455.400 333.900 456.600 334.650 ;
        RECT 448.950 328.950 451.050 333.000 ;
        RECT 454.950 331.800 457.050 333.900 ;
        RECT 454.950 298.950 457.050 301.050 ;
        RECT 455.400 294.600 456.450 298.950 ;
        RECT 464.400 298.050 465.450 352.950 ;
        RECT 472.950 349.950 475.050 352.050 ;
        RECT 473.400 343.050 474.450 349.950 ;
        RECT 485.400 349.050 486.450 365.400 ;
        RECT 491.100 363.900 492.000 369.000 ;
        RECT 498.000 368.100 500.100 369.000 ;
        RECT 492.900 367.200 495.000 368.100 ;
        RECT 492.900 366.000 500.100 367.200 ;
        RECT 498.000 365.100 500.100 366.000 ;
        RECT 490.500 361.800 492.600 363.900 ;
        RECT 493.800 362.100 495.900 364.200 ;
        RECT 496.950 361.950 499.050 364.050 ;
        RECT 501.000 363.600 501.900 376.200 ;
        RECT 503.400 372.450 504.600 372.600 ;
        RECT 505.950 372.450 508.050 376.050 ;
        RECT 503.400 372.000 508.050 372.450 ;
        RECT 503.400 371.400 507.450 372.000 ;
        RECT 503.400 370.350 504.600 371.400 ;
        RECT 502.800 367.950 504.900 370.050 ;
        RECT 505.950 367.950 508.050 370.050 ;
        RECT 494.400 361.050 495.600 361.800 ;
        RECT 493.950 358.950 496.050 361.050 ;
        RECT 484.950 346.950 487.050 349.050 ;
        RECT 472.950 340.950 475.050 343.050 ;
        RECT 466.950 337.950 469.050 340.050 ;
        RECT 473.400 339.600 474.450 340.950 ;
        RECT 467.400 328.050 468.450 337.950 ;
        RECT 473.400 337.350 474.600 339.600 ;
        RECT 478.950 338.100 481.050 340.200 ;
        RECT 490.950 338.100 493.050 340.200 ;
        RECT 497.400 339.450 498.450 361.950 ;
        RECT 500.400 361.500 502.500 363.600 ;
        RECT 494.400 338.400 498.450 339.450 ;
        RECT 499.950 339.000 502.050 343.050 ;
        RECT 506.400 339.600 507.450 367.950 ;
        RECT 512.400 364.050 513.450 385.950 ;
        RECT 521.400 376.050 522.450 428.400 ;
        RECT 524.400 397.050 525.450 443.400 ;
        RECT 535.950 442.800 538.050 444.900 ;
        RECT 541.950 442.800 544.050 444.900 ;
        RECT 547.950 442.800 550.050 444.900 ;
        RECT 535.050 423.300 537.150 425.400 ;
        RECT 529.800 412.950 531.900 415.050 ;
        RECT 530.400 411.450 531.600 412.650 ;
        RECT 527.400 410.400 531.600 411.450 ;
        RECT 523.950 394.950 526.050 397.050 ;
        RECT 527.400 391.050 528.450 410.400 ;
        RECT 535.650 404.700 536.850 423.300 ;
        RECT 542.400 417.450 543.450 442.800 ;
        RECT 553.950 439.950 556.050 445.050 ;
        RECT 560.400 439.050 561.450 449.100 ;
        RECT 562.950 448.950 565.050 451.050 ;
        RECT 565.950 449.100 568.050 451.200 ;
        RECT 572.400 450.600 573.450 475.950 ;
        RECT 598.950 457.950 601.050 460.050 ;
        RECT 566.400 448.350 567.600 449.100 ;
        RECT 572.400 448.350 573.600 450.600 ;
        RECT 592.950 448.950 595.050 451.050 ;
        RECT 599.400 450.600 600.450 457.950 ;
        RECT 593.400 448.350 594.600 448.950 ;
        RECT 599.400 448.350 600.600 450.600 ;
        RECT 604.950 448.950 607.050 451.050 ;
        RECT 565.950 445.950 568.050 448.050 ;
        RECT 568.950 445.950 571.050 448.050 ;
        RECT 571.950 445.950 574.050 448.050 ;
        RECT 589.950 445.950 592.050 448.050 ;
        RECT 592.950 445.950 595.050 448.050 ;
        RECT 595.950 445.950 598.050 448.050 ;
        RECT 598.950 445.950 601.050 448.050 ;
        RECT 569.400 444.900 570.600 445.650 ;
        RECT 568.950 442.800 571.050 444.900 ;
        RECT 590.400 443.400 591.600 445.650 ;
        RECT 596.400 443.400 597.600 445.650 ;
        RECT 590.400 439.050 591.450 443.400 ;
        RECT 559.950 436.950 562.050 439.050 ;
        RECT 571.950 436.950 574.050 439.050 ;
        RECT 589.950 436.950 592.050 439.050 ;
        RECT 550.950 430.950 553.050 433.050 ;
        RECT 542.400 416.400 546.450 417.450 ;
        RECT 538.950 412.950 541.050 415.050 ;
        RECT 539.400 411.000 540.600 412.650 ;
        RECT 538.950 406.950 541.050 411.000 ;
        RECT 532.650 403.500 536.850 404.700 ;
        RECT 532.650 402.600 534.750 403.500 ;
        RECT 539.400 400.050 540.450 406.950 ;
        RECT 538.950 397.950 541.050 400.050 ;
        RECT 535.950 394.950 538.050 397.050 ;
        RECT 526.950 388.950 529.050 391.050 ;
        RECT 532.950 388.950 535.050 391.050 ;
        RECT 520.950 375.450 523.050 376.050 ;
        RECT 525.000 375.450 529.050 376.050 ;
        RECT 520.950 374.400 529.050 375.450 ;
        RECT 520.950 373.950 523.050 374.400 ;
        RECT 525.000 373.950 529.050 374.400 ;
        RECT 517.950 371.100 520.050 373.200 ;
        RECT 518.400 370.350 519.600 371.100 ;
        RECT 523.950 370.950 526.050 373.050 ;
        RECT 524.400 370.350 525.600 370.950 ;
        RECT 517.950 367.950 520.050 370.050 ;
        RECT 520.950 367.950 523.050 370.050 ;
        RECT 523.950 367.950 526.050 370.050 ;
        RECT 526.950 367.950 529.050 370.050 ;
        RECT 521.400 365.400 522.600 367.650 ;
        RECT 527.400 365.400 528.600 367.650 ;
        RECT 511.950 361.950 514.050 364.050 ;
        RECT 521.400 363.450 522.450 365.400 ;
        RECT 521.400 362.400 525.450 363.450 ;
        RECT 517.950 352.950 520.050 355.050 ;
        RECT 514.950 340.950 517.050 343.050 ;
        RECT 479.400 337.350 480.600 338.100 ;
        RECT 472.950 334.950 475.050 337.050 ;
        RECT 475.950 334.950 478.050 337.050 ;
        RECT 478.950 334.950 481.050 337.050 ;
        RECT 481.950 334.950 484.050 337.050 ;
        RECT 469.950 331.950 472.050 334.050 ;
        RECT 476.400 332.400 477.600 334.650 ;
        RECT 482.400 333.900 483.600 334.650 ;
        RECT 466.950 325.950 469.050 328.050 ;
        RECT 470.400 301.050 471.450 331.950 ;
        RECT 476.400 322.050 477.450 332.400 ;
        RECT 481.950 331.800 484.050 333.900 ;
        RECT 484.950 331.950 487.050 334.050 ;
        RECT 491.400 333.900 492.450 338.100 ;
        RECT 494.400 334.050 495.450 338.400 ;
        RECT 500.400 337.350 501.600 339.000 ;
        RECT 506.400 337.350 507.600 339.600 ;
        RECT 499.950 334.950 502.050 337.050 ;
        RECT 502.950 334.950 505.050 337.050 ;
        RECT 505.950 334.950 508.050 337.050 ;
        RECT 508.950 334.950 511.050 337.050 ;
        RECT 475.950 319.950 478.050 322.050 ;
        RECT 485.400 303.450 486.450 331.950 ;
        RECT 490.950 331.800 493.050 333.900 ;
        RECT 493.950 331.950 496.050 334.050 ;
        RECT 496.950 331.800 499.050 333.900 ;
        RECT 503.400 333.000 504.600 334.650 ;
        RECT 491.400 310.050 492.450 331.800 ;
        RECT 493.950 328.800 496.050 330.900 ;
        RECT 494.400 322.050 495.450 328.800 ;
        RECT 497.400 325.050 498.450 331.800 ;
        RECT 502.950 328.950 505.050 333.000 ;
        RECT 509.400 332.400 510.600 334.650 ;
        RECT 496.950 322.950 499.050 325.050 ;
        RECT 493.950 319.950 496.050 322.050 ;
        RECT 502.950 319.950 505.050 322.050 ;
        RECT 490.950 307.950 493.050 310.050 ;
        RECT 482.400 302.400 486.450 303.450 ;
        RECT 469.950 298.950 472.050 301.050 ;
        RECT 475.950 298.950 478.050 301.050 ;
        RECT 463.950 295.950 466.050 298.050 ;
        RECT 455.400 292.350 456.600 294.600 ;
        RECT 463.950 292.800 466.050 294.900 ;
        RECT 469.950 294.000 472.050 297.900 ;
        RECT 476.400 294.600 477.450 298.950 ;
        RECT 482.400 295.050 483.450 302.400 ;
        RECT 484.950 298.950 487.050 301.050 ;
        RECT 446.100 289.950 448.200 292.050 ;
        RECT 451.500 289.950 453.600 292.050 ;
        RECT 454.800 289.950 456.900 292.050 ;
        RECT 454.950 265.950 457.050 268.050 ;
        RECT 442.950 262.950 445.050 265.050 ;
        RECT 448.950 261.000 451.050 265.050 ;
        RECT 455.400 261.600 456.450 265.950 ;
        RECT 449.400 259.350 450.600 261.000 ;
        RECT 455.400 259.350 456.600 261.600 ;
        RECT 460.950 261.450 463.050 262.200 ;
        RECT 464.400 261.450 465.450 292.800 ;
        RECT 470.400 292.350 471.600 294.000 ;
        RECT 476.400 292.350 477.600 294.600 ;
        RECT 481.950 292.950 484.050 295.050 ;
        RECT 469.950 289.950 472.050 292.050 ;
        RECT 472.950 289.950 475.050 292.050 ;
        RECT 475.950 289.950 478.050 292.050 ;
        RECT 478.950 289.950 481.050 292.050 ;
        RECT 473.400 288.000 474.600 289.650 ;
        RECT 472.950 283.950 475.050 288.000 ;
        RECT 479.400 287.400 480.600 289.650 ;
        RECT 475.950 274.950 478.050 277.050 ;
        RECT 472.950 268.950 475.050 271.050 ;
        RECT 466.950 265.950 469.050 268.050 ;
        RECT 460.950 260.400 465.450 261.450 ;
        RECT 460.950 260.100 463.050 260.400 ;
        RECT 461.400 259.350 462.600 260.100 ;
        RECT 448.950 256.950 451.050 259.050 ;
        RECT 451.950 256.950 454.050 259.050 ;
        RECT 454.950 256.950 457.050 259.050 ;
        RECT 457.950 256.950 460.050 259.050 ;
        RECT 460.950 256.950 463.050 259.050 ;
        RECT 452.400 255.900 453.600 256.650 ;
        RECT 425.400 250.050 426.450 254.400 ;
        RECT 439.950 253.800 442.050 255.900 ;
        RECT 451.950 253.800 454.050 255.900 ;
        RECT 458.400 255.000 459.600 256.650 ;
        RECT 457.950 250.950 460.050 255.000 ;
        RECT 424.950 247.950 427.050 250.050 ;
        RECT 448.950 247.950 451.050 250.050 ;
        RECT 416.400 242.400 420.450 243.450 ;
        RECT 410.400 233.400 415.050 235.050 ;
        RECT 411.000 232.950 415.050 233.400 ;
        RECT 409.950 229.950 412.050 232.050 ;
        RECT 410.400 216.600 411.450 229.950 ;
        RECT 416.400 223.050 417.450 242.400 ;
        RECT 439.950 226.950 442.050 229.050 ;
        RECT 415.950 220.950 418.050 223.050 ;
        RECT 433.950 220.950 436.050 223.050 ;
        RECT 410.400 214.350 411.600 216.600 ;
        RECT 415.950 215.100 418.050 217.200 ;
        RECT 416.400 214.350 417.600 215.100 ;
        RECT 427.950 214.950 430.050 217.050 ;
        RECT 434.400 216.600 435.450 220.950 ;
        RECT 440.400 216.600 441.450 226.950 ;
        RECT 409.950 211.950 412.050 214.050 ;
        RECT 412.950 211.950 415.050 214.050 ;
        RECT 415.950 211.950 418.050 214.050 ;
        RECT 418.950 211.950 421.050 214.050 ;
        RECT 413.400 209.400 414.600 211.650 ;
        RECT 419.400 210.900 420.600 211.650 ;
        RECT 413.400 205.050 414.450 209.400 ;
        RECT 418.950 208.800 421.050 210.900 ;
        RECT 424.950 208.950 427.050 211.050 ;
        RECT 403.950 202.950 406.050 205.050 ;
        RECT 412.950 202.950 415.050 205.050 ;
        RECT 412.950 199.800 415.050 201.900 ;
        RECT 400.950 193.950 403.050 196.050 ;
        RECT 413.400 190.050 414.450 199.800 ;
        RECT 391.950 187.950 394.050 190.050 ;
        RECT 412.950 187.950 415.050 190.050 ;
        RECT 388.950 182.100 391.050 184.200 ;
        RECT 394.950 182.100 397.050 184.200 ;
        RECT 389.400 181.350 390.600 182.100 ;
        RECT 395.400 181.350 396.600 182.100 ;
        RECT 400.800 181.950 402.900 184.050 ;
        RECT 403.950 182.100 406.050 184.200 ;
        RECT 409.950 182.100 412.050 184.200 ;
        RECT 415.950 183.000 418.050 187.050 ;
        RECT 385.950 178.950 388.050 181.050 ;
        RECT 388.950 178.950 391.050 181.050 ;
        RECT 391.950 178.950 394.050 181.050 ;
        RECT 394.950 178.950 397.050 181.050 ;
        RECT 386.400 176.400 387.600 178.650 ;
        RECT 392.400 177.000 393.600 178.650 ;
        RECT 373.950 174.450 376.050 175.050 ;
        RECT 373.950 173.400 378.450 174.450 ;
        RECT 373.950 172.950 376.050 173.400 ;
        RECT 370.950 169.950 373.050 172.050 ;
        RECT 361.950 166.950 364.050 169.050 ;
        RECT 362.400 141.450 363.450 166.950 ;
        RECT 362.400 140.400 366.450 141.450 ;
        RECT 344.400 136.350 345.600 137.100 ;
        RECT 352.950 136.950 355.050 139.050 ;
        RECT 358.950 136.950 361.050 139.050 ;
        RECT 365.400 138.600 366.450 140.400 ;
        RECT 337.950 133.950 340.050 136.050 ;
        RECT 340.950 133.950 343.050 136.050 ;
        RECT 343.950 133.950 346.050 136.050 ;
        RECT 346.950 133.950 349.050 136.050 ;
        RECT 341.400 131.400 342.600 133.650 ;
        RECT 347.400 131.400 348.600 133.650 ;
        RECT 341.400 127.050 342.450 131.400 ;
        RECT 340.950 124.950 343.050 127.050 ;
        RECT 334.950 118.950 337.050 121.050 ;
        RECT 278.400 96.450 279.450 98.400 ;
        RECT 283.950 97.800 286.050 99.900 ;
        RECT 289.950 97.800 292.050 99.900 ;
        RECT 278.400 96.000 282.450 96.450 ;
        RECT 277.950 95.400 282.450 96.000 ;
        RECT 277.950 91.950 280.050 95.400 ;
        RECT 266.400 59.400 270.450 60.450 ;
        RECT 223.950 40.950 226.050 43.050 ;
        RECT 241.950 40.950 244.050 43.050 ;
        RECT 224.400 28.050 225.450 40.950 ;
        RECT 235.800 30.300 237.900 32.400 ;
        RECT 238.950 31.950 241.050 34.050 ;
        RECT 239.400 31.200 240.600 31.950 ;
        RECT 142.950 22.950 145.050 25.050 ;
        RECT 145.950 22.950 148.050 25.050 ;
        RECT 160.950 22.950 163.050 25.050 ;
        RECT 163.950 22.950 166.050 25.050 ;
        RECT 166.950 22.950 169.050 25.050 ;
        RECT 169.950 22.950 172.050 25.050 ;
        RECT 184.950 22.950 187.050 25.050 ;
        RECT 187.950 22.950 190.050 25.050 ;
        RECT 193.950 22.950 196.050 25.050 ;
        RECT 49.950 16.950 52.050 19.050 ;
        RECT 86.400 16.050 87.450 20.400 ;
        RECT 100.950 16.950 103.050 21.000 ;
        RECT 106.950 19.800 109.050 21.900 ;
        RECT 112.950 19.800 115.050 21.900 ;
        RECT 124.950 19.800 127.050 21.900 ;
        RECT 136.950 19.950 139.050 22.050 ;
        RECT 143.400 21.900 144.600 22.650 ;
        RECT 164.400 21.900 165.600 22.650 ;
        RECT 170.400 21.900 171.600 22.650 ;
        RECT 185.400 21.900 186.600 22.650 ;
        RECT 142.950 19.800 145.050 21.900 ;
        RECT 163.950 19.800 166.050 21.900 ;
        RECT 169.950 19.800 172.050 21.900 ;
        RECT 184.950 19.800 187.050 21.900 ;
        RECT 194.400 19.050 195.450 22.950 ;
        RECT 197.400 21.900 198.450 25.950 ;
        RECT 209.400 25.350 210.600 27.600 ;
        RECT 215.400 25.350 216.600 27.600 ;
        RECT 223.950 25.950 226.050 28.050 ;
        RECT 229.950 27.600 234.000 28.050 ;
        RECT 229.950 25.950 234.600 27.600 ;
        RECT 233.400 25.350 234.600 25.950 ;
        RECT 205.950 22.950 208.050 25.050 ;
        RECT 208.950 22.950 211.050 25.050 ;
        RECT 211.950 22.950 214.050 25.050 ;
        RECT 214.950 22.950 217.050 25.050 ;
        RECT 233.100 22.950 235.200 25.050 ;
        RECT 236.100 24.900 237.000 30.300 ;
        RECT 239.100 28.800 241.200 30.900 ;
        RECT 243.000 27.900 245.100 29.700 ;
        RECT 251.400 28.050 252.450 53.400 ;
        RECT 256.950 49.950 259.050 54.000 ;
        RECT 262.950 52.800 265.050 54.900 ;
        RECT 266.400 52.050 267.450 59.400 ;
        RECT 274.950 59.100 277.050 61.200 ;
        RECT 275.400 58.350 276.600 59.100 ;
        RECT 271.950 55.950 274.050 58.050 ;
        RECT 274.950 55.950 277.050 58.050 ;
        RECT 272.400 54.900 273.600 55.650 ;
        RECT 281.400 55.050 282.450 95.400 ;
        RECT 296.400 94.050 297.450 109.950 ;
        RECT 305.400 109.200 306.600 109.950 ;
        RECT 301.500 107.100 303.600 109.200 ;
        RECT 298.950 104.100 301.050 106.200 ;
        RECT 299.400 103.350 300.600 104.100 ;
        RECT 299.100 100.950 301.200 103.050 ;
        RECT 302.100 102.000 303.000 107.100 ;
        RECT 304.800 106.800 306.900 108.900 ;
        RECT 311.400 107.400 313.500 109.500 ;
        RECT 309.000 105.000 311.100 105.900 ;
        RECT 303.900 103.800 311.100 105.000 ;
        RECT 303.900 102.900 306.000 103.800 ;
        RECT 309.000 102.000 311.100 102.900 ;
        RECT 302.100 101.100 311.100 102.000 ;
        RECT 302.100 94.500 303.000 101.100 ;
        RECT 309.000 100.800 311.100 101.100 ;
        RECT 304.800 97.950 306.900 100.050 ;
        RECT 305.400 95.400 306.600 97.650 ;
        RECT 312.000 94.800 312.900 107.400 ;
        RECT 313.800 100.950 315.900 103.050 ;
        RECT 319.950 100.950 322.050 103.050 ;
        RECT 314.400 99.900 315.600 100.650 ;
        RECT 313.950 99.450 316.050 99.900 ;
        RECT 313.950 98.400 318.450 99.450 ;
        RECT 320.400 99.000 321.600 100.650 ;
        RECT 313.950 97.800 316.050 98.400 ;
        RECT 295.950 91.950 298.050 94.050 ;
        RECT 302.100 92.400 304.200 94.500 ;
        RECT 311.100 92.700 313.200 94.800 ;
        RECT 317.400 82.050 318.450 98.400 ;
        RECT 319.950 94.950 322.050 99.000 ;
        RECT 316.950 79.950 319.050 82.050 ;
        RECT 286.950 64.950 289.050 67.050 ;
        RECT 295.950 64.950 298.050 67.050 ;
        RECT 316.950 64.950 319.050 67.050 ;
        RECT 271.950 52.800 274.050 54.900 ;
        RECT 280.950 52.950 283.050 55.050 ;
        RECT 265.950 49.950 268.050 52.050 ;
        RECT 287.400 37.050 288.450 64.950 ;
        RECT 296.400 60.600 297.450 64.950 ;
        RECT 303.000 60.600 307.050 61.050 ;
        RECT 296.400 58.350 297.600 60.600 ;
        RECT 302.400 58.950 307.050 60.600 ;
        RECT 310.950 58.950 313.050 61.050 ;
        RECT 317.400 60.600 318.450 64.950 ;
        RECT 320.400 64.050 321.450 94.950 ;
        RECT 324.150 92.700 325.350 111.300 ;
        RECT 328.950 109.950 331.050 112.050 ;
        RECT 335.400 103.050 336.450 118.950 ;
        RECT 347.400 118.050 348.450 131.400 ;
        RECT 353.400 130.050 354.450 136.950 ;
        RECT 365.400 136.350 366.600 138.600 ;
        RECT 370.950 137.100 373.050 139.200 ;
        RECT 371.400 136.350 372.600 137.100 ;
        RECT 361.950 133.950 364.050 136.050 ;
        RECT 364.950 133.950 367.050 136.050 ;
        RECT 367.950 133.950 370.050 136.050 ;
        RECT 370.950 133.950 373.050 136.050 ;
        RECT 358.950 130.950 361.050 133.050 ;
        RECT 362.400 131.400 363.600 133.650 ;
        RECT 368.400 131.400 369.600 133.650 ;
        RECT 352.950 127.950 355.050 130.050 ;
        RECT 337.950 115.950 340.050 118.050 ;
        RECT 346.950 115.950 349.050 118.050 ;
        RECT 329.100 100.950 331.200 103.050 ;
        RECT 334.950 100.950 337.050 103.050 ;
        RECT 329.400 99.000 330.600 100.650 ;
        RECT 328.950 94.950 331.050 99.000 ;
        RECT 338.400 94.050 339.450 115.950 ;
        RECT 341.550 111.300 343.650 113.400 ;
        RECT 341.550 98.400 342.750 111.300 ;
        RECT 346.950 105.000 349.050 109.050 ;
        RECT 352.950 106.950 355.050 109.050 ;
        RECT 347.400 103.350 348.600 105.000 ;
        RECT 346.950 100.950 349.050 103.050 ;
        RECT 341.550 96.300 343.650 98.400 ;
        RECT 324.150 91.500 328.350 92.700 ;
        RECT 337.950 91.950 340.050 94.050 ;
        RECT 326.250 90.600 328.350 91.500 ;
        RECT 341.550 89.700 342.750 96.300 ;
        RECT 341.550 87.600 343.650 89.700 ;
        RECT 353.400 85.050 354.450 106.950 ;
        RECT 359.400 100.050 360.450 130.950 ;
        RECT 362.400 127.050 363.450 131.400 ;
        RECT 361.950 124.950 364.050 127.050 ;
        RECT 368.400 109.050 369.450 131.400 ;
        RECT 373.950 127.950 376.050 130.050 ;
        RECT 367.950 106.950 370.050 109.050 ;
        RECT 369.000 105.600 373.050 106.050 ;
        RECT 368.400 103.950 373.050 105.600 ;
        RECT 368.400 103.350 369.600 103.950 ;
        RECT 364.950 100.950 367.050 103.050 ;
        RECT 367.950 100.950 370.050 103.050 ;
        RECT 358.950 97.950 361.050 100.050 ;
        RECT 365.400 99.900 366.600 100.650 ;
        RECT 364.950 97.800 367.050 99.900 ;
        RECT 340.950 82.950 343.050 85.050 ;
        RECT 352.950 82.950 355.050 85.050 ;
        RECT 367.950 82.950 370.050 85.050 ;
        RECT 335.250 67.500 337.350 68.400 ;
        RECT 333.150 66.300 337.350 67.500 ;
        RECT 319.950 61.950 322.050 64.050 ;
        RECT 302.400 58.350 303.600 58.950 ;
        RECT 292.950 55.950 295.050 58.050 ;
        RECT 295.950 55.950 298.050 58.050 ;
        RECT 298.950 55.950 301.050 58.050 ;
        RECT 301.950 55.950 304.050 58.050 ;
        RECT 307.950 55.950 310.050 58.050 ;
        RECT 293.400 54.900 294.600 55.650 ;
        RECT 292.950 52.800 295.050 54.900 ;
        RECT 299.400 53.400 300.600 55.650 ;
        RECT 299.400 49.050 300.450 53.400 ;
        RECT 308.400 49.050 309.450 55.950 ;
        RECT 311.400 49.050 312.450 58.950 ;
        RECT 317.400 58.350 318.600 60.600 ;
        RECT 322.950 59.100 325.050 61.200 ;
        RECT 328.950 60.000 331.050 64.050 ;
        RECT 323.400 58.350 324.600 59.100 ;
        RECT 329.400 58.350 330.600 60.000 ;
        RECT 316.950 55.950 319.050 58.050 ;
        RECT 319.950 55.950 322.050 58.050 ;
        RECT 322.950 55.950 325.050 58.050 ;
        RECT 328.950 55.950 331.050 58.050 ;
        RECT 320.400 54.900 321.600 55.650 ;
        RECT 319.950 52.800 322.050 54.900 ;
        RECT 298.950 46.950 301.050 49.050 ;
        RECT 307.800 46.950 309.900 49.050 ;
        RECT 310.950 46.950 313.050 49.050 ;
        RECT 333.150 47.700 334.350 66.300 ;
        RECT 341.400 63.450 342.450 82.950 ;
        RECT 343.950 73.950 346.050 76.050 ;
        RECT 338.400 62.400 342.450 63.450 ;
        RECT 338.400 60.600 339.450 62.400 ;
        RECT 338.400 58.350 339.600 60.600 ;
        RECT 338.100 55.950 340.200 58.050 ;
        RECT 344.400 52.050 345.450 73.950 ;
        RECT 350.550 69.300 352.650 71.400 ;
        RECT 350.550 62.700 351.750 69.300 ;
        RECT 350.550 60.600 352.650 62.700 ;
        RECT 343.950 49.950 346.050 52.050 ;
        RECT 350.550 47.700 351.750 60.600 ;
        RECT 355.950 55.950 358.050 58.050 ;
        RECT 356.400 53.400 357.600 55.650 ;
        RECT 368.400 55.050 369.450 82.950 ;
        RECT 374.400 64.050 375.450 127.950 ;
        RECT 377.400 127.050 378.450 173.400 ;
        RECT 386.400 172.050 387.450 176.400 ;
        RECT 391.950 172.950 394.050 177.000 ;
        RECT 385.950 169.950 388.050 172.050 ;
        RECT 385.950 137.100 388.050 139.200 ;
        RECT 401.400 138.450 402.450 181.950 ;
        RECT 404.400 172.050 405.450 182.100 ;
        RECT 410.400 181.350 411.600 182.100 ;
        RECT 416.400 181.350 417.600 183.000 ;
        RECT 409.950 178.950 412.050 181.050 ;
        RECT 412.950 178.950 415.050 181.050 ;
        RECT 415.950 178.950 418.050 181.050 ;
        RECT 413.400 177.900 414.600 178.650 ;
        RECT 412.950 175.800 415.050 177.900 ;
        RECT 403.950 169.950 406.050 172.050 ;
        RECT 406.950 154.950 409.050 157.050 ;
        RECT 407.400 148.050 408.450 154.950 ;
        RECT 406.950 145.950 409.050 148.050 ;
        RECT 398.400 137.400 402.450 138.450 ;
        RECT 407.400 138.600 408.450 145.950 ;
        RECT 386.400 136.350 387.600 137.100 ;
        RECT 385.950 133.950 388.050 136.050 ;
        RECT 388.950 133.950 391.050 136.050 ;
        RECT 376.950 124.950 379.050 127.050 ;
        RECT 382.950 109.950 385.050 112.050 ;
        RECT 376.950 103.950 379.050 106.050 ;
        RECT 383.400 105.600 384.450 109.950 ;
        RECT 390.000 108.450 394.050 109.050 ;
        RECT 389.400 106.950 394.050 108.450 ;
        RECT 389.400 105.600 390.450 106.950 ;
        RECT 377.400 79.050 378.450 103.950 ;
        RECT 383.400 103.350 384.600 105.600 ;
        RECT 389.400 103.350 390.600 105.600 ;
        RECT 382.950 100.950 385.050 103.050 ;
        RECT 385.950 100.950 388.050 103.050 ;
        RECT 388.950 100.950 391.050 103.050 ;
        RECT 391.950 100.950 394.050 103.050 ;
        RECT 386.400 98.400 387.600 100.650 ;
        RECT 392.400 98.400 393.600 100.650 ;
        RECT 386.400 94.050 387.450 98.400 ;
        RECT 385.950 91.950 388.050 94.050 ;
        RECT 392.400 79.050 393.450 98.400 ;
        RECT 376.950 76.950 379.050 79.050 ;
        RECT 385.950 76.950 388.050 79.050 ;
        RECT 391.950 76.950 394.050 79.050 ;
        RECT 373.950 61.950 376.050 64.050 ;
        RECT 374.400 60.600 375.450 61.950 ;
        RECT 374.400 58.350 375.600 60.600 ;
        RECT 373.950 55.950 376.050 58.050 ;
        RECT 376.950 55.950 379.050 58.050 ;
        RECT 379.950 55.950 382.050 58.050 ;
        RECT 332.850 45.600 334.950 47.700 ;
        RECT 350.550 45.600 352.650 47.700 ;
        RECT 257.850 33.300 259.950 35.400 ;
        RECT 237.900 26.700 246.600 27.900 ;
        RECT 237.900 25.800 240.000 26.700 ;
        RECT 236.100 23.700 243.000 24.900 ;
        RECT 206.400 21.900 207.600 22.650 ;
        RECT 196.950 19.800 199.050 21.900 ;
        RECT 205.950 19.800 208.050 21.900 ;
        RECT 212.400 21.000 213.600 22.650 ;
        RECT 193.950 16.950 196.050 19.050 ;
        RECT 211.950 16.950 214.050 21.000 ;
        RECT 236.100 16.500 237.300 23.700 ;
        RECT 239.100 19.950 241.200 22.050 ;
        RECT 242.100 21.300 243.000 23.700 ;
        RECT 239.400 17.400 240.600 19.650 ;
        RECT 242.100 19.200 244.200 21.300 ;
        RECT 245.700 17.700 246.600 26.700 ;
        RECT 250.950 25.950 253.050 28.050 ;
        RECT 247.800 22.950 249.900 25.050 ;
        RECT 253.950 22.950 256.050 25.050 ;
        RECT 248.400 21.900 249.600 22.650 ;
        RECT 247.950 19.800 250.050 21.900 ;
        RECT 254.400 21.000 255.600 22.650 ;
        RECT 46.950 13.950 49.050 16.050 ;
        RECT 85.950 13.950 88.050 16.050 ;
        RECT 235.800 14.400 237.900 16.500 ;
        RECT 245.400 15.600 247.500 17.700 ;
        RECT 253.950 16.950 256.050 21.000 ;
        RECT 258.150 14.700 259.350 33.300 ;
        RECT 265.950 31.950 268.050 34.050 ;
        RECT 275.550 33.300 277.650 35.400 ;
        RECT 286.950 34.950 289.050 37.050 ;
        RECT 293.850 33.300 295.950 35.400 ;
        RECT 311.550 33.300 313.650 35.400 ;
        RECT 266.400 28.050 267.450 31.950 ;
        RECT 265.950 25.950 268.050 28.050 ;
        RECT 271.950 26.100 274.050 28.200 ;
        RECT 263.100 22.950 265.200 25.050 ;
        RECT 263.400 21.900 264.600 22.650 ;
        RECT 262.950 19.800 265.050 21.900 ;
        RECT 258.150 13.500 262.350 14.700 ;
        RECT 260.250 12.600 262.350 13.500 ;
        RECT 272.400 13.050 273.450 26.100 ;
        RECT 275.550 20.400 276.750 33.300 ;
        RECT 280.950 26.100 283.050 28.200 ;
        RECT 281.400 25.350 282.600 26.100 ;
        RECT 280.950 22.950 283.050 25.050 ;
        RECT 289.950 22.950 292.050 25.050 ;
        RECT 290.400 21.900 291.600 22.650 ;
        RECT 275.550 18.300 277.650 20.400 ;
        RECT 271.950 10.950 274.050 13.050 ;
        RECT 275.550 11.700 276.750 18.300 ;
        RECT 289.950 16.950 292.050 21.900 ;
        RECT 294.150 14.700 295.350 33.300 ;
        RECT 299.100 22.950 301.200 25.050 ;
        RECT 299.400 20.400 300.600 22.650 ;
        RECT 311.550 20.400 312.750 33.300 ;
        RECT 356.400 31.050 357.450 53.400 ;
        RECT 367.950 52.950 370.050 55.050 ;
        RECT 377.400 54.000 378.600 55.650 ;
        RECT 376.950 49.950 379.050 54.000 ;
        RECT 373.950 48.600 376.050 49.050 ;
        RECT 379.950 48.600 382.050 49.050 ;
        RECT 373.950 47.550 382.050 48.600 ;
        RECT 373.950 46.950 376.050 47.550 ;
        RECT 379.950 46.950 382.050 47.550 ;
        RECT 373.950 43.800 376.050 45.900 ;
        RECT 367.950 34.950 370.050 37.050 ;
        RECT 355.950 28.950 358.050 31.050 ;
        RECT 316.950 26.100 319.050 28.200 ;
        RECT 334.950 26.100 337.050 28.200 ;
        RECT 361.950 27.000 364.050 31.050 ;
        RECT 317.400 25.350 318.600 26.100 ;
        RECT 335.400 25.350 336.600 26.100 ;
        RECT 362.400 25.350 363.600 27.000 ;
        RECT 316.950 22.950 319.050 25.050 ;
        RECT 335.400 22.950 337.500 25.050 ;
        RECT 340.800 22.950 342.900 25.050 ;
        RECT 356.100 22.950 358.200 25.050 ;
        RECT 361.500 22.950 363.600 25.050 ;
        RECT 368.400 22.050 369.450 34.950 ;
        RECT 299.400 18.450 300.450 20.400 ;
        RECT 299.400 17.400 303.450 18.450 ;
        RECT 294.150 13.500 298.350 14.700 ;
        RECT 296.250 12.600 298.350 13.500 ;
        RECT 302.400 13.050 303.450 17.400 ;
        RECT 311.550 18.300 313.650 20.400 ;
        RECT 367.950 19.950 370.050 22.050 ;
        RECT 374.400 21.450 375.450 43.800 ;
        RECT 386.400 43.050 387.450 76.950 ;
        RECT 398.400 70.050 399.450 137.400 ;
        RECT 407.400 136.350 408.600 138.600 ;
        RECT 412.950 137.100 415.050 139.200 ;
        RECT 418.950 137.100 421.050 139.200 ;
        RECT 425.400 138.450 426.450 208.950 ;
        RECT 428.400 202.050 429.450 214.950 ;
        RECT 434.400 214.350 435.600 216.600 ;
        RECT 440.400 214.350 441.600 216.600 ;
        RECT 433.950 211.950 436.050 214.050 ;
        RECT 436.950 211.950 439.050 214.050 ;
        RECT 439.950 211.950 442.050 214.050 ;
        RECT 442.950 211.950 445.050 214.050 ;
        RECT 437.400 210.900 438.600 211.650 ;
        RECT 436.950 208.800 439.050 210.900 ;
        RECT 443.400 209.400 444.600 211.650 ;
        RECT 430.950 202.950 433.050 205.050 ;
        RECT 427.950 199.950 430.050 202.050 ;
        RECT 431.400 183.600 432.450 202.950 ;
        RECT 436.950 190.950 439.050 193.050 ;
        RECT 437.400 183.600 438.450 190.950 ;
        RECT 443.400 184.050 444.450 209.400 ;
        RECT 449.400 187.050 450.450 247.950 ;
        RECT 454.950 235.950 457.050 238.050 ;
        RECT 455.400 210.900 456.450 235.950 ;
        RECT 460.950 232.950 463.050 235.050 ;
        RECT 457.950 214.950 460.050 220.050 ;
        RECT 461.400 216.600 462.450 232.950 ;
        RECT 467.400 223.050 468.450 265.950 ;
        RECT 469.950 262.950 472.050 265.050 ;
        RECT 470.400 232.050 471.450 262.950 ;
        RECT 473.400 262.050 474.450 268.950 ;
        RECT 476.400 262.200 477.450 274.950 ;
        RECT 479.400 274.050 480.450 287.400 ;
        RECT 478.950 271.950 481.050 274.050 ;
        RECT 485.400 265.050 486.450 298.950 ;
        RECT 487.950 295.950 490.050 298.050 ;
        RECT 488.400 286.050 489.450 295.950 ;
        RECT 496.950 293.100 499.050 295.200 ;
        RECT 503.400 294.600 504.450 319.950 ;
        RECT 509.400 316.050 510.450 332.400 ;
        RECT 508.950 313.950 511.050 316.050 ;
        RECT 515.400 303.450 516.450 340.950 ;
        RECT 518.400 322.050 519.450 352.950 ;
        RECT 524.400 339.600 525.450 362.400 ;
        RECT 527.400 343.050 528.450 365.400 ;
        RECT 533.400 361.050 534.450 388.950 ;
        RECT 532.950 358.950 535.050 361.050 ;
        RECT 536.400 355.050 537.450 394.950 ;
        RECT 545.400 388.050 546.450 416.400 ;
        RECT 547.950 415.950 550.050 418.050 ;
        RECT 548.400 409.050 549.450 415.950 ;
        RECT 551.400 411.900 552.450 430.950 ;
        RECT 561.000 420.450 565.050 421.050 ;
        RECT 560.400 418.950 565.050 420.450 ;
        RECT 560.400 417.600 561.450 418.950 ;
        RECT 560.400 415.350 561.600 417.600 ;
        RECT 556.950 412.950 559.050 415.050 ;
        RECT 559.950 412.950 562.050 415.050 ;
        RECT 562.950 412.950 565.050 415.050 ;
        RECT 557.400 411.900 558.600 412.650 ;
        RECT 550.950 409.800 553.050 411.900 ;
        RECT 556.950 409.800 559.050 411.900 ;
        RECT 563.400 411.450 564.600 412.650 ;
        RECT 565.950 411.450 568.050 411.900 ;
        RECT 563.400 410.400 568.050 411.450 ;
        RECT 565.950 409.800 568.050 410.400 ;
        RECT 547.950 406.950 550.050 409.050 ;
        RECT 559.950 406.950 565.050 409.050 ;
        RECT 566.400 406.050 567.450 409.800 ;
        RECT 565.950 403.950 568.050 406.050 ;
        RECT 572.400 403.050 573.450 436.950 ;
        RECT 586.950 430.950 589.050 433.050 ;
        RECT 577.950 424.950 580.050 427.050 ;
        RECT 574.950 418.950 577.050 421.050 ;
        RECT 571.950 400.950 574.050 403.050 ;
        RECT 565.950 397.950 568.050 400.050 ;
        RECT 544.950 385.950 547.050 388.050 ;
        RECT 545.100 376.500 547.200 378.600 ;
        RECT 542.100 367.950 544.200 370.050 ;
        RECT 545.100 369.900 546.000 376.500 ;
        RECT 554.100 376.200 556.200 378.300 ;
        RECT 548.400 373.350 549.600 375.600 ;
        RECT 547.800 370.950 549.900 373.050 ;
        RECT 552.000 369.900 554.100 370.200 ;
        RECT 545.100 369.000 554.100 369.900 ;
        RECT 542.400 366.450 543.600 367.650 ;
        RECT 539.400 365.400 543.600 366.450 ;
        RECT 535.950 352.950 538.050 355.050 ;
        RECT 526.950 340.950 529.050 343.050 ;
        RECT 524.400 337.350 525.600 339.600 ;
        RECT 529.950 338.100 532.050 340.200 ;
        RECT 530.400 337.350 531.600 338.100 ;
        RECT 523.950 334.950 526.050 337.050 ;
        RECT 526.950 334.950 529.050 337.050 ;
        RECT 529.950 334.950 532.050 337.050 ;
        RECT 532.950 334.950 535.050 337.050 ;
        RECT 527.400 333.900 528.600 334.650 ;
        RECT 526.950 331.800 529.050 333.900 ;
        RECT 533.400 332.400 534.600 334.650 ;
        RECT 533.400 328.050 534.450 332.400 ;
        RECT 532.950 325.950 535.050 328.050 ;
        RECT 517.950 319.950 520.050 322.050 ;
        RECT 526.950 307.950 529.050 310.050 ;
        RECT 512.400 302.400 516.450 303.450 ;
        RECT 497.400 292.350 498.600 293.100 ;
        RECT 503.400 292.350 504.600 294.600 ;
        RECT 508.950 293.100 511.050 295.200 ;
        RECT 493.950 289.950 496.050 292.050 ;
        RECT 496.950 289.950 499.050 292.050 ;
        RECT 499.950 289.950 502.050 292.050 ;
        RECT 502.950 289.950 505.050 292.050 ;
        RECT 494.400 287.400 495.600 289.650 ;
        RECT 500.400 288.900 501.600 289.650 ;
        RECT 509.400 289.050 510.450 293.100 ;
        RECT 487.950 283.950 490.050 286.050 ;
        RECT 494.400 277.050 495.450 287.400 ;
        RECT 499.950 286.800 502.050 288.900 ;
        RECT 508.950 286.950 511.050 289.050 ;
        RECT 496.950 283.950 499.050 286.050 ;
        RECT 493.950 274.950 496.050 277.050 ;
        RECT 487.950 271.950 490.050 274.050 ;
        RECT 484.950 262.950 487.050 265.050 ;
        RECT 472.950 259.950 475.050 262.050 ;
        RECT 475.950 260.100 478.050 262.200 ;
        RECT 481.950 260.100 484.050 262.200 ;
        RECT 488.400 262.050 489.450 271.950 ;
        RECT 493.950 270.450 496.050 271.050 ;
        RECT 497.400 270.450 498.450 283.950 ;
        RECT 493.950 269.400 498.450 270.450 ;
        RECT 493.950 268.950 496.050 269.400 ;
        RECT 490.950 262.800 493.050 264.900 ;
        RECT 476.400 259.350 477.600 260.100 ;
        RECT 482.400 259.350 483.600 260.100 ;
        RECT 487.950 259.950 490.050 262.050 ;
        RECT 475.950 256.950 478.050 259.050 ;
        RECT 478.950 256.950 481.050 259.050 ;
        RECT 481.950 256.950 484.050 259.050 ;
        RECT 484.950 256.950 487.050 259.050 ;
        RECT 472.950 253.950 475.050 256.050 ;
        RECT 479.400 255.000 480.600 256.650 ;
        RECT 485.400 255.900 486.600 256.650 ;
        RECT 473.400 241.050 474.450 253.950 ;
        RECT 478.950 250.950 481.050 255.000 ;
        RECT 484.950 253.800 487.050 255.900 ;
        RECT 487.950 253.950 490.050 256.050 ;
        RECT 491.400 255.900 492.450 262.800 ;
        RECT 472.950 238.950 475.050 241.050 ;
        RECT 488.400 238.050 489.450 253.950 ;
        RECT 490.950 253.800 493.050 255.900 ;
        RECT 487.950 235.950 490.050 238.050 ;
        RECT 469.950 229.950 472.050 232.050 ;
        RECT 466.950 220.950 469.050 223.050 ;
        RECT 478.950 220.950 481.050 223.050 ;
        RECT 487.950 220.950 490.050 223.050 ;
        RECT 461.400 214.350 462.600 216.600 ;
        RECT 466.950 216.000 469.050 219.900 ;
        RECT 467.400 214.350 468.600 216.000 ;
        RECT 460.950 211.950 463.050 214.050 ;
        RECT 463.950 211.950 466.050 214.050 ;
        RECT 466.950 211.950 469.050 214.050 ;
        RECT 469.950 211.950 472.050 214.050 ;
        RECT 475.950 211.950 478.050 214.050 ;
        RECT 464.400 210.900 465.600 211.650 ;
        RECT 454.950 208.800 457.050 210.900 ;
        RECT 463.950 208.800 466.050 210.900 ;
        RECT 470.400 209.400 471.600 211.650 ;
        RECT 470.400 190.050 471.450 209.400 ;
        RECT 476.400 205.050 477.450 211.950 ;
        RECT 475.950 202.950 478.050 205.050 ;
        RECT 469.950 187.950 472.050 190.050 ;
        RECT 448.950 184.950 451.050 187.050 ;
        RECT 466.950 184.950 469.050 187.050 ;
        RECT 431.400 181.350 432.600 183.600 ;
        RECT 437.400 181.350 438.600 183.600 ;
        RECT 442.950 181.950 445.050 184.050 ;
        RECT 445.950 181.950 448.050 184.050 ;
        RECT 430.950 178.950 433.050 181.050 ;
        RECT 433.950 178.950 436.050 181.050 ;
        RECT 436.950 178.950 439.050 181.050 ;
        RECT 439.950 178.950 442.050 181.050 ;
        RECT 434.400 177.900 435.600 178.650 ;
        RECT 440.400 177.900 441.600 178.650 ;
        RECT 433.950 175.800 436.050 177.900 ;
        RECT 439.950 175.800 442.050 177.900 ;
        RECT 442.950 175.950 445.050 178.050 ;
        RECT 446.400 177.900 447.450 181.950 ;
        RECT 443.400 139.200 444.450 175.950 ;
        RECT 445.950 175.800 448.050 177.900 ;
        RECT 449.400 175.050 450.450 184.950 ;
        RECT 457.950 182.100 460.050 184.200 ;
        RECT 458.400 181.350 459.600 182.100 ;
        RECT 454.950 178.950 457.050 181.050 ;
        RECT 457.950 178.950 460.050 181.050 ;
        RECT 460.950 178.950 463.050 181.050 ;
        RECT 455.400 177.000 456.600 178.650 ;
        RECT 461.400 177.000 462.600 178.650 ;
        RECT 448.950 172.950 451.050 175.050 ;
        RECT 454.950 172.950 457.050 177.000 ;
        RECT 460.950 169.950 463.050 177.000 ;
        RECT 467.400 175.050 468.450 184.950 ;
        RECT 476.400 183.600 477.450 202.950 ;
        RECT 479.400 202.050 480.450 220.950 ;
        RECT 488.400 216.600 489.450 220.950 ;
        RECT 491.400 220.050 492.450 253.800 ;
        RECT 494.400 253.050 495.450 268.950 ;
        RECT 499.950 260.100 502.050 262.200 ;
        RECT 505.950 261.000 508.050 265.050 ;
        RECT 512.400 261.450 513.450 302.400 ;
        RECT 514.950 298.950 517.050 301.050 ;
        RECT 520.950 298.950 523.050 301.050 ;
        RECT 515.400 288.900 516.450 298.950 ;
        RECT 521.400 295.200 522.450 298.950 ;
        RECT 520.950 293.100 523.050 295.200 ;
        RECT 527.400 294.600 528.450 307.950 ;
        RECT 532.950 304.950 535.050 307.050 ;
        RECT 533.400 294.600 534.450 304.950 ;
        RECT 539.400 300.450 540.450 365.400 ;
        RECT 545.100 363.900 546.000 369.000 ;
        RECT 552.000 368.100 554.100 369.000 ;
        RECT 546.900 367.200 549.000 368.100 ;
        RECT 546.900 366.000 554.100 367.200 ;
        RECT 552.000 365.100 554.100 366.000 ;
        RECT 544.500 361.800 546.600 363.900 ;
        RECT 547.800 362.100 549.900 364.200 ;
        RECT 555.000 363.600 555.900 376.200 ;
        RECT 562.950 373.950 565.050 376.050 ;
        RECT 556.950 371.100 559.050 373.200 ;
        RECT 557.400 370.350 558.600 371.100 ;
        RECT 556.800 367.950 558.900 370.050 ;
        RECT 563.400 366.900 564.450 373.950 ;
        RECT 562.950 364.800 565.050 366.900 ;
        RECT 548.400 361.050 549.600 361.800 ;
        RECT 554.400 361.500 556.500 363.600 ;
        RECT 547.950 358.950 550.050 361.050 ;
        RECT 541.950 340.950 544.050 343.050 ;
        RECT 542.400 324.450 543.450 340.950 ;
        RECT 550.950 338.100 553.050 340.200 ;
        RECT 556.950 339.000 559.050 343.050 ;
        RECT 551.400 337.350 552.600 338.100 ;
        RECT 557.400 337.350 558.600 339.000 ;
        RECT 562.950 337.950 565.050 340.050 ;
        RECT 547.950 334.950 550.050 337.050 ;
        RECT 550.950 334.950 553.050 337.050 ;
        RECT 553.950 334.950 556.050 337.050 ;
        RECT 556.950 334.950 559.050 337.050 ;
        RECT 548.400 332.400 549.600 334.650 ;
        RECT 554.400 333.900 555.600 334.650 ;
        RECT 563.400 333.900 564.450 337.950 ;
        RECT 548.400 328.050 549.450 332.400 ;
        RECT 553.950 331.800 556.050 333.900 ;
        RECT 562.950 331.800 565.050 333.900 ;
        RECT 547.950 325.950 550.050 328.050 ;
        RECT 542.400 323.400 546.450 324.450 ;
        RECT 539.400 299.400 543.450 300.450 ;
        RECT 538.950 295.950 541.050 298.050 ;
        RECT 521.400 292.350 522.600 293.100 ;
        RECT 527.400 292.350 528.600 294.600 ;
        RECT 533.400 292.350 534.600 294.600 ;
        RECT 520.950 289.950 523.050 292.050 ;
        RECT 523.950 289.950 526.050 292.050 ;
        RECT 526.950 289.950 529.050 292.050 ;
        RECT 529.950 289.950 532.050 292.050 ;
        RECT 532.950 289.950 535.050 292.050 ;
        RECT 514.950 286.800 517.050 288.900 ;
        RECT 524.400 287.400 525.600 289.650 ;
        RECT 530.400 288.900 531.600 289.650 ;
        RECT 524.400 283.050 525.450 287.400 ;
        RECT 529.950 286.800 532.050 288.900 ;
        RECT 539.400 286.050 540.450 295.950 ;
        RECT 538.950 283.950 541.050 286.050 ;
        RECT 523.950 280.950 526.050 283.050 ;
        RECT 535.950 282.900 540.000 283.050 ;
        RECT 535.950 280.950 541.050 282.900 ;
        RECT 538.950 280.800 541.050 280.950 ;
        RECT 542.400 277.050 543.450 299.400 ;
        RECT 545.400 298.050 546.450 323.400 ;
        RECT 554.400 316.050 555.450 331.800 ;
        RECT 556.950 325.950 559.050 328.050 ;
        RECT 553.950 313.950 556.050 316.050 ;
        RECT 557.400 307.050 558.450 325.950 ;
        RECT 556.950 304.950 559.050 307.050 ;
        RECT 550.950 298.950 556.050 301.050 ;
        RECT 544.950 295.950 547.050 298.050 ;
        RECT 547.950 293.100 550.050 295.200 ;
        RECT 554.400 294.450 555.600 294.600 ;
        RECT 557.400 294.450 558.450 304.950 ;
        RECT 559.950 298.950 562.050 301.050 ;
        RECT 566.400 300.450 567.450 397.950 ;
        RECT 575.400 385.050 576.450 418.950 ;
        RECT 578.400 409.050 579.450 424.950 ;
        RECT 587.400 417.600 588.450 430.950 ;
        RECT 587.400 415.350 588.600 417.600 ;
        RECT 581.100 412.950 583.200 415.050 ;
        RECT 586.500 412.950 588.600 415.050 ;
        RECT 589.800 412.950 591.900 415.050 ;
        RECT 581.400 411.900 582.600 412.650 ;
        RECT 580.950 409.800 583.050 411.900 ;
        RECT 590.400 410.400 591.600 412.650 ;
        RECT 577.950 406.950 580.050 409.050 ;
        RECT 583.950 400.950 586.050 403.050 ;
        RECT 574.950 382.950 577.050 385.050 ;
        RECT 576.000 375.450 580.050 376.050 ;
        RECT 575.400 373.950 580.050 375.450 ;
        RECT 575.400 372.600 576.450 373.950 ;
        RECT 575.400 370.350 576.600 372.600 ;
        RECT 580.950 371.100 583.050 373.200 ;
        RECT 571.950 367.950 574.050 370.050 ;
        RECT 574.950 367.950 577.050 370.050 ;
        RECT 572.400 366.900 573.600 367.650 ;
        RECT 581.400 367.050 582.450 371.100 ;
        RECT 584.400 367.050 585.450 400.950 ;
        RECT 590.400 382.050 591.450 410.400 ;
        RECT 589.950 379.950 592.050 382.050 ;
        RECT 596.400 379.050 597.450 443.400 ;
        RECT 605.400 442.050 606.450 448.950 ;
        RECT 611.400 445.050 612.450 484.950 ;
        RECT 620.400 460.050 621.450 494.400 ;
        RECT 623.400 489.900 624.450 502.950 ;
        RECT 641.400 501.450 642.450 544.950 ;
        RECT 644.400 529.200 645.450 577.950 ;
        RECT 659.400 573.600 660.450 577.950 ;
        RECT 659.400 571.350 660.600 573.600 ;
        RECT 649.950 568.950 652.050 571.050 ;
        RECT 652.950 568.950 655.050 571.050 ;
        RECT 655.950 568.950 658.050 571.050 ;
        RECT 658.950 568.950 661.050 571.050 ;
        RECT 661.950 568.950 664.050 571.050 ;
        RECT 656.400 566.400 657.600 568.650 ;
        RECT 656.400 541.050 657.450 566.400 ;
        RECT 671.400 565.050 672.450 605.400 ;
        RECT 676.950 605.100 679.050 607.200 ;
        RECT 682.950 606.000 685.050 610.050 ;
        RECT 677.400 604.350 678.600 605.100 ;
        RECT 683.400 604.350 684.600 606.000 ;
        RECT 676.950 601.950 679.050 604.050 ;
        RECT 679.950 601.950 682.050 604.050 ;
        RECT 682.950 601.950 685.050 604.050 ;
        RECT 685.950 601.950 688.050 604.050 ;
        RECT 680.400 599.400 681.600 601.650 ;
        RECT 686.400 600.450 687.600 601.650 ;
        RECT 692.400 600.450 693.450 640.950 ;
        RECT 709.500 639.600 711.600 641.700 ;
        RECT 716.400 641.400 717.600 643.650 ;
        RECT 719.700 640.500 720.900 647.700 ;
        RECT 721.800 646.950 723.900 649.050 ;
        RECT 719.100 638.400 721.200 640.500 ;
        RECT 725.400 628.050 726.450 650.400 ;
        RECT 740.100 646.950 742.200 649.050 ;
        RECT 740.400 645.900 741.600 646.650 ;
        RECT 739.950 643.800 742.050 645.900 ;
        RECT 743.100 640.800 744.000 653.400 ;
        RECT 749.100 652.800 751.200 654.900 ;
        RECT 752.400 653.100 754.500 655.200 ;
        RECT 744.900 651.000 747.000 651.900 ;
        RECT 744.900 649.800 752.100 651.000 ;
        RECT 750.000 648.900 752.100 649.800 ;
        RECT 744.900 648.000 747.000 648.900 ;
        RECT 753.000 648.000 753.900 653.100 ;
        RECT 755.400 651.450 756.600 651.600 ;
        RECT 755.400 650.400 759.450 651.450 ;
        RECT 755.400 649.350 756.600 650.400 ;
        RECT 744.900 647.100 753.900 648.000 ;
        RECT 744.900 646.800 747.000 647.100 ;
        RECT 749.100 643.950 751.200 646.050 ;
        RECT 749.400 641.400 750.600 643.650 ;
        RECT 742.800 638.700 744.900 640.800 ;
        RECT 753.000 640.500 753.900 647.100 ;
        RECT 754.800 646.950 756.900 649.050 ;
        RECT 751.800 638.400 753.900 640.500 ;
        RECT 758.400 628.050 759.450 650.400 ;
        RECT 764.400 643.050 765.450 658.950 ;
        RECT 770.400 655.050 771.450 682.950 ;
        RECT 779.400 682.350 780.600 684.600 ;
        RECT 785.400 682.350 786.600 684.600 ;
        RECT 790.950 682.950 793.050 685.050 ;
        RECT 778.950 679.950 781.050 682.050 ;
        RECT 781.950 679.950 784.050 682.050 ;
        RECT 784.950 679.950 787.050 682.050 ;
        RECT 787.950 679.950 790.050 682.050 ;
        RECT 774.000 678.900 778.050 679.050 ;
        RECT 782.400 678.900 783.600 679.650 ;
        RECT 788.400 678.900 789.600 679.650 ;
        RECT 772.950 676.950 778.050 678.900 ;
        RECT 772.950 676.800 775.050 676.950 ;
        RECT 781.950 676.800 784.050 678.900 ;
        RECT 787.950 676.800 790.050 678.900 ;
        RECT 784.950 667.950 787.050 670.050 ;
        RECT 769.950 652.950 772.050 655.050 ;
        RECT 770.400 651.600 771.450 652.950 ;
        RECT 770.400 649.350 771.600 651.600 ;
        RECT 775.950 650.100 778.050 652.200 ;
        RECT 776.400 649.350 777.600 650.100 ;
        RECT 785.400 649.050 786.450 667.950 ;
        RECT 787.950 649.950 790.050 652.050 ;
        RECT 794.400 651.450 795.450 685.950 ;
        RECT 797.400 655.050 798.450 691.950 ;
        RECT 806.400 684.600 807.450 697.950 ;
        RECT 812.400 685.200 813.450 706.950 ;
        RECT 817.950 685.950 820.050 688.050 ;
        RECT 806.400 682.350 807.600 684.600 ;
        RECT 811.950 683.100 814.050 685.200 ;
        RECT 812.400 682.350 813.600 683.100 ;
        RECT 802.950 679.950 805.050 682.050 ;
        RECT 805.950 679.950 808.050 682.050 ;
        RECT 808.950 679.950 811.050 682.050 ;
        RECT 811.950 679.950 814.050 682.050 ;
        RECT 803.400 677.400 804.600 679.650 ;
        RECT 809.400 678.900 810.600 679.650 ;
        RECT 803.400 670.050 804.450 677.400 ;
        RECT 808.950 676.800 811.050 678.900 ;
        RECT 818.400 678.450 819.450 685.950 ;
        RECT 815.400 677.400 819.450 678.450 ;
        RECT 811.950 673.950 814.050 676.050 ;
        RECT 802.950 667.950 805.050 670.050 ;
        RECT 799.950 661.950 802.050 664.050 ;
        RECT 796.950 652.950 799.050 655.050 ;
        RECT 791.400 650.400 795.450 651.450 ;
        RECT 800.400 651.600 801.450 661.950 ;
        RECT 808.950 652.950 811.050 655.050 ;
        RECT 769.950 646.950 772.050 649.050 ;
        RECT 772.950 646.950 775.050 649.050 ;
        RECT 775.950 646.950 778.050 649.050 ;
        RECT 778.950 646.950 781.050 649.050 ;
        RECT 784.950 646.950 787.050 649.050 ;
        RECT 773.400 645.900 774.600 646.650 ;
        RECT 772.950 643.800 775.050 645.900 ;
        RECT 779.400 645.000 780.600 646.650 ;
        RECT 763.950 640.950 766.050 643.050 ;
        RECT 778.950 640.950 781.050 645.000 ;
        RECT 724.950 625.950 727.050 628.050 ;
        RECT 757.950 625.950 760.050 628.050 ;
        RECT 697.950 622.950 700.050 625.050 ;
        RECT 698.400 601.050 699.450 622.950 ;
        RECT 718.950 619.950 721.050 622.050 ;
        RECT 706.950 610.950 709.050 613.050 ;
        RECT 707.400 606.600 708.450 610.950 ;
        RECT 707.400 604.350 708.600 606.600 ;
        RECT 712.950 605.100 715.050 607.200 ;
        RECT 713.400 604.350 714.600 605.100 ;
        RECT 703.950 601.950 706.050 604.050 ;
        RECT 706.950 601.950 709.050 604.050 ;
        RECT 709.950 601.950 712.050 604.050 ;
        RECT 712.950 601.950 715.050 604.050 ;
        RECT 686.400 599.400 693.450 600.450 ;
        RECT 680.400 586.050 681.450 599.400 ;
        RECT 697.950 598.950 700.050 601.050 ;
        RECT 704.400 600.900 705.600 601.650 ;
        RECT 703.950 598.800 706.050 600.900 ;
        RECT 710.400 599.400 711.600 601.650 ;
        RECT 719.400 601.050 720.450 619.950 ;
        RECT 736.950 610.950 739.050 613.050 ;
        RECT 745.950 610.950 748.050 613.050 ;
        RECT 757.950 610.950 760.050 613.050 ;
        RECT 778.950 610.950 781.050 613.050 ;
        RECT 730.950 605.100 733.050 607.200 ;
        RECT 737.400 606.600 738.450 610.950 ;
        RECT 731.400 604.350 732.600 605.100 ;
        RECT 737.400 604.350 738.600 606.600 ;
        RECT 742.950 605.100 745.050 607.200 ;
        RECT 727.950 601.950 730.050 604.050 ;
        RECT 730.950 601.950 733.050 604.050 ;
        RECT 733.950 601.950 736.050 604.050 ;
        RECT 736.950 601.950 739.050 604.050 ;
        RECT 706.950 592.950 709.050 595.050 ;
        RECT 682.950 589.950 685.050 592.050 ;
        RECT 679.950 583.950 682.050 586.050 ;
        RECT 680.400 580.050 681.450 583.950 ;
        RECT 679.950 577.950 682.050 580.050 ;
        RECT 683.400 573.600 684.450 589.950 ;
        RECT 683.400 571.350 684.600 573.600 ;
        RECT 697.950 571.950 700.050 574.050 ;
        RECT 707.400 573.600 708.450 592.950 ;
        RECT 710.400 592.050 711.450 599.400 ;
        RECT 718.950 598.950 721.050 601.050 ;
        RECT 728.400 600.900 729.600 601.650 ;
        RECT 727.950 598.800 730.050 600.900 ;
        RECT 734.400 599.400 735.600 601.650 ;
        RECT 743.400 601.050 744.450 605.100 ;
        RECT 734.400 592.050 735.450 599.400 ;
        RECT 742.950 598.950 745.050 601.050 ;
        RECT 709.950 589.950 712.050 592.050 ;
        RECT 733.950 589.950 736.050 592.050 ;
        RECT 730.950 577.950 733.050 580.050 ;
        RECT 739.950 577.950 742.050 580.050 ;
        RECT 679.950 568.950 682.050 571.050 ;
        RECT 682.950 568.950 685.050 571.050 ;
        RECT 685.950 568.950 688.050 571.050 ;
        RECT 670.950 562.950 673.050 565.050 ;
        RECT 655.950 538.950 658.050 541.050 ;
        RECT 698.400 538.050 699.450 571.950 ;
        RECT 707.400 571.350 708.600 573.600 ;
        RECT 712.950 572.100 715.050 574.200 ;
        RECT 713.400 571.350 714.600 572.100 ;
        RECT 718.950 571.950 721.050 574.050 ;
        RECT 731.400 573.600 732.450 577.950 ;
        RECT 703.950 568.950 706.050 571.050 ;
        RECT 706.950 568.950 709.050 571.050 ;
        RECT 709.950 568.950 712.050 571.050 ;
        RECT 712.950 568.950 715.050 571.050 ;
        RECT 704.400 567.000 705.600 568.650 ;
        RECT 710.400 567.900 711.600 568.650 ;
        RECT 703.950 562.950 706.050 567.000 ;
        RECT 709.950 565.800 712.050 567.900 ;
        RECT 719.400 547.050 720.450 571.950 ;
        RECT 731.400 571.350 732.600 573.600 ;
        RECT 727.950 568.950 730.050 571.050 ;
        RECT 730.950 568.950 733.050 571.050 ;
        RECT 728.400 567.900 729.600 568.650 ;
        RECT 740.400 567.900 741.450 577.950 ;
        RECT 746.400 573.600 747.450 610.950 ;
        RECT 758.400 606.600 759.450 610.950 ;
        RECT 758.400 604.350 759.600 606.600 ;
        RECT 763.950 605.100 766.050 607.200 ;
        RECT 769.950 605.100 772.050 607.200 ;
        RECT 779.400 606.600 780.450 610.950 ;
        RECT 788.400 610.050 789.450 649.950 ;
        RECT 791.400 613.050 792.450 650.400 ;
        RECT 800.400 649.350 801.600 651.600 ;
        RECT 796.950 646.950 799.050 649.050 ;
        RECT 799.950 646.950 802.050 649.050 ;
        RECT 802.950 646.950 805.050 649.050 ;
        RECT 797.400 645.900 798.600 646.650 ;
        RECT 796.950 643.800 799.050 645.900 ;
        RECT 803.400 644.400 804.600 646.650 ;
        RECT 797.400 631.050 798.450 643.800 ;
        RECT 796.950 628.950 799.050 631.050 ;
        RECT 803.400 619.050 804.450 644.400 ;
        RECT 809.400 622.050 810.450 652.950 ;
        RECT 808.950 619.950 811.050 622.050 ;
        RECT 812.400 619.050 813.450 673.950 ;
        RECT 815.400 652.050 816.450 677.400 ;
        RECT 817.950 673.950 820.050 676.050 ;
        RECT 814.950 649.950 817.050 652.050 ;
        RECT 818.400 651.600 819.450 673.950 ;
        RECT 821.400 664.050 822.450 712.950 ;
        RECT 832.950 694.950 835.050 697.050 ;
        RECT 826.950 684.000 829.050 688.050 ;
        RECT 833.400 684.600 834.450 694.950 ;
        RECT 839.400 685.200 840.450 722.400 ;
        RECT 844.950 721.800 847.050 723.900 ;
        RECT 851.400 722.400 852.600 724.650 ;
        RECT 847.950 718.950 850.050 721.050 ;
        RECT 827.400 682.350 828.600 684.000 ;
        RECT 833.400 682.350 834.600 684.600 ;
        RECT 838.950 683.100 841.050 685.200 ;
        RECT 844.950 683.100 847.050 685.200 ;
        RECT 839.400 682.350 840.600 683.100 ;
        RECT 826.950 679.950 829.050 682.050 ;
        RECT 829.950 679.950 832.050 682.050 ;
        RECT 832.950 679.950 835.050 682.050 ;
        RECT 835.950 679.950 838.050 682.050 ;
        RECT 838.950 679.950 841.050 682.050 ;
        RECT 830.400 678.000 831.600 679.650 ;
        RECT 836.400 678.900 837.600 679.650 ;
        RECT 829.950 673.950 832.050 678.000 ;
        RECT 835.950 676.800 838.050 678.900 ;
        RECT 832.950 667.950 835.050 670.050 ;
        RECT 820.950 661.950 823.050 664.050 ;
        RECT 818.400 649.350 819.600 651.600 ;
        RECT 823.950 650.100 826.050 652.200 ;
        RECT 824.400 649.350 825.600 650.100 ;
        RECT 817.950 646.950 820.050 649.050 ;
        RECT 820.950 646.950 823.050 649.050 ;
        RECT 823.950 646.950 826.050 649.050 ;
        RECT 826.950 646.950 829.050 649.050 ;
        RECT 821.400 645.000 822.600 646.650 ;
        RECT 827.400 646.050 828.600 646.650 ;
        RECT 820.950 640.950 823.050 645.000 ;
        RECT 827.400 644.400 832.050 646.050 ;
        RECT 828.000 643.950 832.050 644.400 ;
        RECT 826.950 640.950 829.050 643.050 ;
        RECT 820.950 637.800 823.050 639.900 ;
        RECT 802.950 616.950 805.050 619.050 ;
        RECT 811.950 616.950 814.050 619.050 ;
        RECT 790.950 610.950 793.050 613.050 ;
        RECT 787.950 607.950 790.050 610.050 ;
        RECT 796.950 607.950 799.050 610.050 ;
        RECT 764.400 604.350 765.600 605.100 ;
        RECT 754.950 601.950 757.050 604.050 ;
        RECT 757.950 601.950 760.050 604.050 ;
        RECT 760.950 601.950 763.050 604.050 ;
        RECT 763.950 601.950 766.050 604.050 ;
        RECT 755.400 600.900 756.600 601.650 ;
        RECT 761.400 600.900 762.600 601.650 ;
        RECT 754.950 598.800 757.050 600.900 ;
        RECT 760.950 598.800 763.050 600.900 ;
        RECT 770.400 586.050 771.450 605.100 ;
        RECT 779.400 604.350 780.600 606.600 ;
        RECT 784.950 605.100 787.050 607.200 ;
        RECT 793.950 605.100 796.050 607.200 ;
        RECT 785.400 604.350 786.600 605.100 ;
        RECT 778.950 601.950 781.050 604.050 ;
        RECT 781.950 601.950 784.050 604.050 ;
        RECT 784.950 601.950 787.050 604.050 ;
        RECT 787.950 601.950 790.050 604.050 ;
        RECT 775.950 598.800 778.050 600.900 ;
        RECT 782.400 599.400 783.600 601.650 ;
        RECT 788.400 599.400 789.600 601.650 ;
        RECT 760.950 583.950 763.050 586.050 ;
        RECT 769.950 583.950 772.050 586.050 ;
        RECT 746.400 571.350 747.600 573.600 ;
        RECT 751.950 572.100 754.050 574.200 ;
        RECT 752.400 571.350 753.600 572.100 ;
        RECT 745.950 568.950 748.050 571.050 ;
        RECT 748.950 568.950 751.050 571.050 ;
        RECT 751.950 568.950 754.050 571.050 ;
        RECT 754.950 568.950 757.050 571.050 ;
        RECT 727.950 565.800 730.050 567.900 ;
        RECT 739.950 565.800 742.050 567.900 ;
        RECT 749.400 566.400 750.600 568.650 ;
        RECT 755.400 567.900 756.600 568.650 ;
        RECT 749.400 562.050 750.450 566.400 ;
        RECT 754.950 565.800 757.050 567.900 ;
        RECT 748.950 559.950 751.050 562.050 ;
        RECT 757.950 558.450 760.050 559.050 ;
        RECT 761.400 558.450 762.450 583.950 ;
        RECT 772.950 574.950 775.050 580.050 ;
        RECT 776.400 574.200 777.450 598.800 ;
        RECT 782.400 595.050 783.450 599.400 ;
        RECT 788.400 595.050 789.450 599.400 ;
        RECT 781.950 592.950 784.050 595.050 ;
        RECT 787.950 592.950 790.050 595.050 ;
        RECT 794.400 589.050 795.450 605.100 ;
        RECT 784.950 586.950 787.050 589.050 ;
        RECT 793.950 586.950 796.050 589.050 ;
        RECT 763.950 571.950 766.050 574.050 ;
        RECT 769.950 572.100 772.050 574.200 ;
        RECT 775.950 572.100 778.050 574.200 ;
        RECT 764.400 562.050 765.450 571.950 ;
        RECT 770.400 571.350 771.600 572.100 ;
        RECT 776.400 571.350 777.600 572.100 ;
        RECT 769.950 568.950 772.050 571.050 ;
        RECT 772.950 568.950 775.050 571.050 ;
        RECT 775.950 568.950 778.050 571.050 ;
        RECT 778.950 568.950 781.050 571.050 ;
        RECT 773.400 567.000 774.600 568.650 ;
        RECT 772.950 562.950 775.050 567.000 ;
        RECT 779.400 566.400 780.600 568.650 ;
        RECT 763.950 559.950 766.050 562.050 ;
        RECT 779.400 559.050 780.450 566.400 ;
        RECT 781.950 565.950 784.050 568.050 ;
        RECT 782.400 562.050 783.450 565.950 ;
        RECT 781.950 559.950 784.050 562.050 ;
        RECT 757.950 557.400 762.450 558.450 ;
        RECT 757.950 556.950 760.050 557.400 ;
        RECT 778.950 556.950 781.050 559.050 ;
        RECT 733.950 550.950 736.050 553.050 ;
        RECT 718.950 544.950 721.050 547.050 ;
        RECT 697.950 535.950 700.050 538.050 ;
        RECT 715.950 532.950 718.050 535.050 ;
        RECT 661.950 529.800 664.050 531.900 ;
        RECT 643.950 527.100 646.050 529.200 ;
        RECT 652.950 527.100 655.050 529.200 ;
        RECT 653.400 526.350 654.600 527.100 ;
        RECT 646.950 523.950 649.050 526.050 ;
        RECT 649.950 523.950 652.050 526.050 ;
        RECT 652.950 523.950 655.050 526.050 ;
        RECT 650.400 521.400 651.600 523.650 ;
        RECT 646.950 514.950 649.050 517.050 ;
        RECT 641.400 500.400 645.450 501.450 ;
        RECT 640.950 498.450 643.050 499.050 ;
        RECT 632.400 497.400 643.050 498.450 ;
        RECT 632.400 495.600 633.450 497.400 ;
        RECT 640.950 496.950 643.050 497.400 ;
        RECT 632.400 493.350 633.600 495.600 ;
        RECT 637.950 494.100 640.050 496.200 ;
        RECT 638.400 493.350 639.600 494.100 ;
        RECT 628.950 490.950 631.050 493.050 ;
        RECT 631.950 490.950 634.050 493.050 ;
        RECT 634.950 490.950 637.050 493.050 ;
        RECT 637.950 490.950 640.050 493.050 ;
        RECT 629.400 489.900 630.600 490.650 ;
        RECT 622.950 487.800 625.050 489.900 ;
        RECT 628.950 487.800 631.050 489.900 ;
        RECT 635.400 488.400 636.600 490.650 ;
        RECT 635.400 475.050 636.450 488.400 ;
        RECT 634.950 472.950 637.050 475.050 ;
        RECT 619.950 457.950 622.050 460.050 ;
        RECT 634.950 457.950 637.050 460.050 ;
        RECT 619.950 449.100 622.050 451.200 ;
        RECT 625.950 450.000 628.050 454.050 ;
        RECT 620.400 448.350 621.600 449.100 ;
        RECT 626.400 448.350 627.600 450.000 ;
        RECT 616.950 445.950 619.050 448.050 ;
        RECT 619.950 445.950 622.050 448.050 ;
        RECT 622.950 445.950 625.050 448.050 ;
        RECT 625.950 445.950 628.050 448.050 ;
        RECT 610.950 442.950 613.050 445.050 ;
        RECT 617.400 443.400 618.600 445.650 ;
        RECT 623.400 444.900 624.600 445.650 ;
        RECT 604.950 439.950 607.050 442.050 ;
        RECT 604.950 436.800 607.050 438.900 ;
        RECT 605.400 417.600 606.450 436.800 ;
        RECT 605.400 415.350 606.600 417.600 ;
        RECT 610.950 416.100 613.050 418.200 ;
        RECT 617.400 417.450 618.450 443.400 ;
        RECT 622.950 442.800 625.050 444.900 ;
        RECT 628.950 442.800 631.050 444.900 ;
        RECT 617.400 416.400 621.450 417.450 ;
        RECT 611.400 415.350 612.600 416.100 ;
        RECT 604.950 412.950 607.050 415.050 ;
        RECT 607.950 412.950 610.050 415.050 ;
        RECT 610.950 412.950 613.050 415.050 ;
        RECT 613.950 412.950 616.050 415.050 ;
        RECT 608.400 411.000 609.600 412.650 ;
        RECT 614.400 411.900 615.600 412.650 ;
        RECT 607.950 406.950 610.050 411.000 ;
        RECT 613.950 409.800 616.050 411.900 ;
        RECT 595.950 376.950 598.050 379.050 ;
        RECT 595.950 372.000 598.050 375.900 ;
        RECT 620.400 375.450 621.450 416.400 ;
        RECT 622.950 416.100 625.050 418.200 ;
        RECT 629.400 417.600 630.450 442.800 ;
        RECT 635.400 430.050 636.450 457.950 ;
        RECT 644.400 454.050 645.450 500.400 ;
        RECT 647.400 460.050 648.450 514.950 ;
        RECT 650.400 496.050 651.450 521.400 ;
        RECT 662.400 511.050 663.450 529.800 ;
        RECT 667.950 528.000 670.050 532.050 ;
        RECT 668.400 526.350 669.600 528.000 ;
        RECT 673.950 527.100 676.050 529.200 ;
        RECT 688.950 527.100 691.050 529.200 ;
        RECT 697.950 528.000 700.050 532.050 ;
        RECT 703.950 529.950 706.050 532.050 ;
        RECT 674.400 526.350 675.600 527.100 ;
        RECT 689.400 526.350 690.600 527.100 ;
        RECT 698.400 526.350 699.600 528.000 ;
        RECT 667.950 523.950 670.050 526.050 ;
        RECT 670.950 523.950 673.050 526.050 ;
        RECT 673.950 523.950 676.050 526.050 ;
        RECT 689.100 523.950 691.200 526.050 ;
        RECT 694.500 523.950 696.600 526.050 ;
        RECT 697.800 523.950 699.900 526.050 ;
        RECT 671.400 522.900 672.600 523.650 ;
        RECT 670.950 520.800 673.050 522.900 ;
        RECT 695.400 521.400 696.600 523.650 ;
        RECT 695.400 511.050 696.450 521.400 ;
        RECT 661.950 508.950 664.050 511.050 ;
        RECT 694.950 508.950 697.050 511.050 ;
        RECT 704.400 508.050 705.450 529.950 ;
        RECT 716.400 528.600 717.450 532.950 ;
        RECT 716.400 526.350 717.600 528.600 ;
        RECT 721.950 527.100 724.050 529.200 ;
        RECT 727.950 527.100 730.050 529.200 ;
        RECT 722.400 526.350 723.600 527.100 ;
        RECT 712.950 523.950 715.050 526.050 ;
        RECT 715.950 523.950 718.050 526.050 ;
        RECT 718.950 523.950 721.050 526.050 ;
        RECT 721.950 523.950 724.050 526.050 ;
        RECT 713.400 522.900 714.600 523.650 ;
        RECT 712.950 520.800 715.050 522.900 ;
        RECT 719.400 521.400 720.600 523.650 ;
        RECT 703.950 505.950 706.050 508.050 ;
        RECT 709.950 505.950 712.050 508.050 ;
        RECT 670.950 499.950 673.050 502.050 ;
        RECT 703.950 499.950 706.050 502.050 ;
        RECT 649.950 493.950 652.050 496.050 ;
        RECT 655.950 495.000 658.050 499.050 ;
        RECT 656.400 493.350 657.600 495.000 ;
        RECT 671.400 493.050 672.450 499.950 ;
        RECT 691.950 496.950 694.050 499.050 ;
        RECT 697.950 496.950 703.050 499.050 ;
        RECT 688.950 493.950 691.050 496.050 ;
        RECT 652.950 490.950 655.050 493.050 ;
        RECT 655.950 490.950 658.050 493.050 ;
        RECT 658.950 490.950 661.050 493.050 ;
        RECT 664.950 490.950 667.050 493.050 ;
        RECT 670.950 490.950 673.050 493.050 ;
        RECT 674.100 490.950 676.200 493.050 ;
        RECT 677.400 490.950 679.500 493.050 ;
        RECT 682.800 490.950 684.900 493.050 ;
        RECT 653.400 490.050 654.600 490.650 ;
        RECT 649.950 488.400 654.600 490.050 ;
        RECT 659.400 488.400 660.600 490.650 ;
        RECT 649.950 487.950 654.000 488.400 ;
        RECT 650.400 481.050 651.450 487.950 ;
        RECT 649.950 478.950 652.050 481.050 ;
        RECT 659.400 478.050 660.450 488.400 ;
        RECT 665.400 484.050 666.450 490.950 ;
        RECT 674.400 488.400 675.600 490.650 ;
        RECT 664.950 481.950 667.050 484.050 ;
        RECT 674.400 478.050 675.450 488.400 ;
        RECT 689.400 484.050 690.450 493.950 ;
        RECT 692.400 493.050 693.450 496.950 ;
        RECT 694.950 495.600 699.000 496.050 ;
        RECT 704.400 495.600 705.450 499.950 ;
        RECT 710.400 496.050 711.450 505.950 ;
        RECT 694.950 493.950 699.600 495.600 ;
        RECT 698.400 493.350 699.600 493.950 ;
        RECT 704.400 493.350 705.600 495.600 ;
        RECT 709.950 493.950 712.050 496.050 ;
        RECT 691.950 490.950 694.050 493.050 ;
        RECT 697.950 490.950 700.050 493.050 ;
        RECT 700.950 490.950 703.050 493.050 ;
        RECT 703.950 490.950 706.050 493.050 ;
        RECT 706.950 490.950 709.050 493.050 ;
        RECT 701.400 489.000 702.600 490.650 ;
        RECT 707.400 489.900 708.600 490.650 ;
        RECT 700.950 484.950 703.050 489.000 ;
        RECT 706.950 487.800 709.050 489.900 ;
        RECT 688.950 481.950 691.050 484.050 ;
        RECT 694.950 481.950 697.050 484.050 ;
        RECT 658.950 475.950 661.050 478.050 ;
        RECT 673.950 475.950 676.050 478.050 ;
        RECT 646.950 457.950 649.050 460.050 ;
        RECT 643.800 451.950 645.900 454.050 ;
        RECT 646.950 450.000 649.050 454.050 ;
        RECT 652.950 450.000 655.050 454.050 ;
        RECT 661.950 451.950 664.050 454.050 ;
        RECT 664.950 451.950 670.050 454.050 ;
        RECT 647.400 448.350 648.600 450.000 ;
        RECT 653.400 448.350 654.600 450.000 ;
        RECT 658.950 449.100 661.050 451.200 ;
        RECT 643.950 445.950 646.050 448.050 ;
        RECT 646.950 445.950 649.050 448.050 ;
        RECT 649.950 445.950 652.050 448.050 ;
        RECT 652.950 445.950 655.050 448.050 ;
        RECT 644.400 444.000 645.600 445.650 ;
        RECT 643.950 439.950 646.050 444.000 ;
        RECT 650.400 443.400 651.600 445.650 ;
        RECT 650.400 439.050 651.450 443.400 ;
        RECT 659.400 442.050 660.450 449.100 ;
        RECT 662.400 448.050 663.450 451.950 ;
        RECT 670.950 450.000 673.050 454.050 ;
        RECT 695.400 451.200 696.450 481.950 ;
        RECT 719.400 457.050 720.450 521.400 ;
        RECT 728.400 508.050 729.450 527.100 ;
        RECT 734.400 523.050 735.450 550.950 ;
        RECT 739.950 527.100 742.050 529.200 ;
        RECT 745.950 527.100 748.050 532.050 ;
        RECT 740.400 526.350 741.600 527.100 ;
        RECT 746.400 526.350 747.600 527.100 ;
        RECT 754.950 526.950 757.050 529.050 ;
        RECT 739.950 523.950 742.050 526.050 ;
        RECT 742.950 523.950 745.050 526.050 ;
        RECT 745.950 523.950 748.050 526.050 ;
        RECT 748.950 523.950 751.050 526.050 ;
        RECT 733.950 520.950 736.050 523.050 ;
        RECT 743.400 522.000 744.600 523.650 ;
        RECT 749.400 522.900 750.600 523.650 ;
        RECT 742.950 517.950 745.050 522.000 ;
        RECT 748.950 520.800 751.050 522.900 ;
        RECT 727.950 505.950 730.050 508.050 ;
        RECT 721.950 494.100 724.050 499.050 ;
        RECT 728.400 495.600 729.450 505.950 ;
        RECT 743.400 502.050 744.450 517.950 ;
        RECT 755.400 508.050 756.450 526.950 ;
        RECT 758.400 523.050 759.450 556.950 ;
        RECT 760.950 544.950 763.050 547.050 ;
        RECT 757.800 520.950 759.900 523.050 ;
        RECT 761.400 522.900 762.450 544.950 ;
        RECT 778.950 532.950 781.050 535.050 ;
        RECT 763.950 528.600 768.000 529.050 ;
        RECT 763.950 526.950 768.600 528.600 ;
        RECT 772.950 527.100 775.050 529.200 ;
        RECT 779.400 529.050 780.450 532.950 ;
        RECT 785.400 532.050 786.450 586.950 ;
        RECT 797.400 577.050 798.450 607.950 ;
        RECT 802.950 606.000 805.050 610.050 ;
        RECT 803.400 604.350 804.600 606.000 ;
        RECT 808.950 605.100 811.050 607.200 ;
        RECT 809.400 604.350 810.600 605.100 ;
        RECT 802.950 601.950 805.050 604.050 ;
        RECT 805.950 601.950 808.050 604.050 ;
        RECT 808.950 601.950 811.050 604.050 ;
        RECT 811.950 601.950 814.050 604.050 ;
        RECT 806.400 599.400 807.600 601.650 ;
        RECT 812.400 599.400 813.600 601.650 ;
        RECT 806.400 592.050 807.450 599.400 ;
        RECT 812.400 595.050 813.450 599.400 ;
        RECT 811.950 592.950 814.050 595.050 ;
        RECT 805.950 589.950 808.050 592.050 ;
        RECT 821.400 589.050 822.450 637.800 ;
        RECT 823.950 628.950 826.050 631.050 ;
        RECT 824.400 600.900 825.450 628.950 ;
        RECT 827.400 606.600 828.450 640.950 ;
        RECT 833.400 640.050 834.450 667.950 ;
        RECT 836.400 646.050 837.450 676.800 ;
        RECT 845.400 652.200 846.450 683.100 ;
        RECT 848.400 670.050 849.450 718.950 ;
        RECT 851.400 715.050 852.450 722.400 ;
        RECT 850.950 712.950 853.050 715.050 ;
        RECT 857.400 714.450 858.450 728.100 ;
        RECT 860.400 721.050 861.450 796.950 ;
        RECT 863.400 781.050 864.450 805.950 ;
        RECT 869.400 805.350 870.600 807.600 ;
        RECT 874.950 806.100 877.050 808.200 ;
        RECT 881.400 808.050 882.450 817.950 ;
        RECT 883.950 811.950 886.050 814.050 ;
        RECT 875.400 805.350 876.600 806.100 ;
        RECT 880.950 805.950 883.050 808.050 ;
        RECT 868.950 802.950 871.050 805.050 ;
        RECT 871.950 802.950 874.050 805.050 ;
        RECT 874.950 802.950 877.050 805.050 ;
        RECT 877.950 802.950 880.050 805.050 ;
        RECT 865.950 796.950 868.050 802.050 ;
        RECT 872.400 800.400 873.600 802.650 ;
        RECT 878.400 800.400 879.600 802.650 ;
        RECT 872.400 787.050 873.450 800.400 ;
        RECT 878.400 799.050 879.450 800.400 ;
        RECT 880.950 799.950 883.050 802.050 ;
        RECT 877.950 796.950 880.050 799.050 ;
        RECT 874.950 787.950 877.050 790.050 ;
        RECT 871.950 784.950 874.050 787.050 ;
        RECT 862.950 778.950 865.050 781.050 ;
        RECT 862.950 772.950 865.050 775.050 ;
        RECT 863.400 730.050 864.450 772.950 ;
        RECT 868.950 766.950 871.050 769.050 ;
        RECT 869.400 763.200 870.450 766.950 ;
        RECT 875.400 766.050 876.450 787.950 ;
        RECT 878.400 769.050 879.450 796.950 ;
        RECT 877.950 766.950 880.050 769.050 ;
        RECT 881.400 766.050 882.450 799.950 ;
        RECT 884.400 790.050 885.450 811.950 ;
        RECT 883.950 787.950 886.050 790.050 ;
        RECT 883.950 778.950 886.050 781.050 ;
        RECT 874.950 763.950 877.050 766.050 ;
        RECT 880.950 763.950 883.050 766.050 ;
        RECT 868.950 761.100 871.050 763.200 ;
        RECT 875.400 762.600 876.450 763.950 ;
        RECT 869.400 760.350 870.600 761.100 ;
        RECT 875.400 760.350 876.600 762.600 ;
        RECT 868.950 757.950 871.050 760.050 ;
        RECT 871.950 757.950 874.050 760.050 ;
        RECT 874.950 757.950 877.050 760.050 ;
        RECT 877.950 757.950 880.050 760.050 ;
        RECT 872.400 756.900 873.600 757.650 ;
        RECT 871.950 754.800 874.050 756.900 ;
        RECT 878.400 755.400 879.600 757.650 ;
        RECT 865.950 736.950 868.050 739.050 ;
        RECT 862.950 727.950 865.050 730.050 ;
        RECT 866.400 729.600 867.450 736.950 ;
        RECT 866.400 727.350 867.600 729.600 ;
        RECT 871.950 728.100 874.050 730.200 ;
        RECT 878.400 730.050 879.450 755.400 ;
        RECT 872.400 727.350 873.600 728.100 ;
        RECT 877.950 727.950 880.050 730.050 ;
        RECT 865.950 724.950 868.050 727.050 ;
        RECT 868.950 724.950 871.050 727.050 ;
        RECT 871.950 724.950 874.050 727.050 ;
        RECT 874.950 724.950 877.050 727.050 ;
        RECT 869.400 723.000 870.600 724.650 ;
        RECT 875.400 723.900 876.600 724.650 ;
        RECT 859.950 718.950 862.050 721.050 ;
        RECT 868.950 718.950 871.050 723.000 ;
        RECT 874.950 721.800 877.050 723.900 ;
        RECT 869.400 715.050 870.450 718.950 ;
        RECT 871.950 715.950 874.050 718.050 ;
        RECT 857.400 713.400 861.450 714.450 ;
        RECT 850.950 700.950 853.050 703.050 ;
        RECT 847.950 667.950 850.050 670.050 ;
        RECT 851.400 658.050 852.450 700.950 ;
        RECT 860.400 685.200 861.450 713.400 ;
        RECT 868.950 712.950 871.050 715.050 ;
        RECT 859.950 683.100 862.050 685.200 ;
        RECT 865.950 684.000 868.050 688.050 ;
        RECT 860.400 682.350 861.600 683.100 ;
        RECT 866.400 682.350 867.600 684.000 ;
        RECT 856.950 679.950 859.050 682.050 ;
        RECT 859.950 679.950 862.050 682.050 ;
        RECT 862.950 679.950 865.050 682.050 ;
        RECT 865.950 679.950 868.050 682.050 ;
        RECT 857.400 678.900 858.600 679.650 ;
        RECT 856.950 676.800 859.050 678.900 ;
        RECT 863.400 677.400 864.600 679.650 ;
        RECT 850.950 655.950 853.050 658.050 ;
        RECT 844.950 650.100 847.050 652.200 ;
        RECT 850.950 650.100 853.050 652.200 ;
        RECT 857.400 652.050 858.450 676.800 ;
        RECT 863.400 673.050 864.450 677.400 ;
        RECT 872.400 676.050 873.450 715.950 ;
        RECT 875.400 679.050 876.450 721.800 ;
        RECT 877.950 715.950 880.050 721.050 ;
        RECT 884.400 703.050 885.450 778.950 ;
        RECT 883.950 700.950 886.050 703.050 ;
        RECT 887.400 688.050 888.450 838.950 ;
        RECT 893.400 838.350 894.600 839.100 ;
        RECT 892.950 835.950 895.050 838.050 ;
        RECT 895.950 835.950 898.050 838.050 ;
        RECT 898.950 826.950 901.050 829.050 ;
        RECT 895.950 775.950 898.050 778.050 ;
        RECT 896.400 730.200 897.450 775.950 ;
        RECT 899.400 733.050 900.450 826.950 ;
        RECT 898.950 730.950 901.050 733.050 ;
        RECT 895.950 728.100 898.050 730.200 ;
        RECT 896.400 727.350 897.600 728.100 ;
        RECT 892.950 724.950 895.050 727.050 ;
        RECT 895.950 724.950 898.050 727.050 ;
        RECT 889.950 721.950 892.050 724.050 ;
        RECT 893.400 723.000 894.600 724.650 ;
        RECT 890.400 688.050 891.450 721.950 ;
        RECT 892.950 718.950 895.050 723.000 ;
        RECT 898.950 721.950 901.050 724.050 ;
        RECT 877.950 685.950 880.050 688.050 ;
        RECT 886.950 685.950 889.050 688.050 ;
        RECT 874.950 676.950 877.050 679.050 ;
        RECT 865.950 673.950 868.050 676.050 ;
        RECT 871.950 673.950 874.050 676.050 ;
        RECT 862.950 670.950 865.050 673.050 ;
        RECT 862.950 661.950 865.050 664.050 ;
        RECT 859.950 655.950 862.050 658.050 ;
        RECT 845.400 649.350 846.600 650.100 ;
        RECT 851.400 649.350 852.600 650.100 ;
        RECT 856.950 649.950 859.050 652.050 ;
        RECT 841.950 646.950 844.050 649.050 ;
        RECT 844.950 646.950 847.050 649.050 ;
        RECT 847.950 646.950 850.050 649.050 ;
        RECT 850.950 646.950 853.050 649.050 ;
        RECT 856.950 646.800 859.050 648.900 ;
        RECT 835.950 643.950 838.050 646.050 ;
        RECT 842.400 645.000 843.600 646.650 ;
        RECT 841.950 640.950 844.050 645.000 ;
        RECT 848.400 644.400 849.600 646.650 ;
        RECT 832.950 637.950 835.050 640.050 ;
        RECT 848.400 637.050 849.450 644.400 ;
        RECT 853.950 643.950 856.050 646.050 ;
        RECT 847.950 634.950 850.050 637.050 ;
        RECT 838.950 628.950 841.050 631.050 ;
        RECT 835.950 616.950 838.050 619.050 ;
        RECT 836.400 606.600 837.450 616.950 ;
        RECT 827.400 604.350 828.600 606.600 ;
        RECT 836.400 604.350 837.600 606.600 ;
        RECT 827.100 601.950 829.200 604.050 ;
        RECT 830.400 601.950 832.500 604.050 ;
        RECT 835.800 601.950 837.900 604.050 ;
        RECT 830.400 600.900 831.600 601.650 ;
        RECT 823.950 598.800 826.050 600.900 ;
        RECT 829.950 598.800 832.050 600.900 ;
        RECT 808.950 586.950 811.050 589.050 ;
        RECT 820.950 586.950 823.050 589.050 ;
        RECT 799.950 583.950 802.050 586.050 ;
        RECT 787.950 574.950 790.050 577.050 ;
        RECT 790.950 576.450 795.000 577.050 ;
        RECT 790.950 574.950 795.450 576.450 ;
        RECT 796.950 574.950 799.050 577.050 ;
        RECT 788.400 567.900 789.450 574.950 ;
        RECT 794.400 573.600 795.450 574.950 ;
        RECT 800.400 573.600 801.450 583.950 ;
        RECT 794.400 571.350 795.600 573.600 ;
        RECT 800.400 571.350 801.600 573.600 ;
        RECT 793.950 568.950 796.050 571.050 ;
        RECT 796.950 568.950 799.050 571.050 ;
        RECT 799.950 568.950 802.050 571.050 ;
        RECT 802.950 568.950 805.050 571.050 ;
        RECT 797.400 567.900 798.600 568.650 ;
        RECT 787.950 565.800 790.050 567.900 ;
        RECT 796.950 565.800 799.050 567.900 ;
        RECT 803.400 566.400 804.600 568.650 ;
        RECT 809.400 567.450 810.450 586.950 ;
        RECT 835.950 583.950 838.050 586.050 ;
        RECT 826.950 580.950 829.050 583.050 ;
        RECT 827.400 574.200 828.450 580.950 ;
        RECT 832.950 577.950 835.050 580.050 ;
        RECT 811.950 572.100 814.050 574.200 ;
        RECT 820.950 572.100 823.050 574.200 ;
        RECT 826.950 572.100 829.050 574.200 ;
        RECT 806.400 566.400 810.450 567.450 ;
        RECT 803.400 559.050 804.450 566.400 ;
        RECT 806.400 561.450 807.450 566.400 ;
        RECT 812.400 565.050 813.450 572.100 ;
        RECT 821.400 571.350 822.600 572.100 ;
        RECT 827.400 571.350 828.600 572.100 ;
        RECT 817.950 568.950 820.050 571.050 ;
        RECT 820.950 568.950 823.050 571.050 ;
        RECT 823.950 568.950 826.050 571.050 ;
        RECT 826.950 568.950 829.050 571.050 ;
        RECT 818.400 566.400 819.600 568.650 ;
        RECT 824.400 567.900 825.600 568.650 ;
        RECT 811.950 562.950 814.050 565.050 ;
        RECT 806.400 560.400 810.450 561.450 ;
        RECT 802.950 556.950 805.050 559.050 ;
        RECT 793.950 541.950 796.050 544.050 ;
        RECT 784.950 529.950 787.050 532.050 ;
        RECT 767.400 526.350 768.600 526.950 ;
        RECT 773.400 526.350 774.600 527.100 ;
        RECT 778.950 526.950 781.050 529.050 ;
        RECT 784.950 526.800 787.050 528.900 ;
        RECT 794.400 528.600 795.450 541.950 ;
        RECT 766.950 523.950 769.050 526.050 ;
        RECT 769.950 523.950 772.050 526.050 ;
        RECT 772.950 523.950 775.050 526.050 ;
        RECT 775.950 523.950 778.050 526.050 ;
        RECT 770.400 522.900 771.600 523.650 ;
        RECT 776.400 523.050 777.600 523.650 ;
        RECT 785.400 523.050 786.450 526.800 ;
        RECT 794.400 526.350 795.600 528.600 ;
        RECT 799.950 527.100 802.050 529.200 ;
        RECT 805.950 527.100 808.050 529.200 ;
        RECT 800.400 526.350 801.600 527.100 ;
        RECT 790.950 523.950 793.050 526.050 ;
        RECT 793.950 523.950 796.050 526.050 ;
        RECT 796.950 523.950 799.050 526.050 ;
        RECT 799.950 523.950 802.050 526.050 ;
        RECT 760.950 520.800 763.050 522.900 ;
        RECT 769.950 520.800 772.050 522.900 ;
        RECT 776.400 521.400 781.050 523.050 ;
        RECT 777.000 520.950 781.050 521.400 ;
        RECT 784.950 520.950 787.050 523.050 ;
        RECT 791.400 522.900 792.600 523.650 ;
        RECT 797.400 522.900 798.600 523.650 ;
        RECT 790.950 520.800 793.050 522.900 ;
        RECT 796.950 520.800 799.050 522.900 ;
        RECT 806.400 520.050 807.450 527.100 ;
        RECT 775.950 517.950 778.050 520.050 ;
        RECT 805.950 517.950 808.050 520.050 ;
        RECT 754.950 505.950 757.050 508.050 ;
        RECT 742.950 499.950 745.050 502.050 ;
        RECT 760.950 496.950 763.050 499.050 ;
        RECT 728.400 493.350 729.600 495.600 ;
        RECT 745.950 494.100 748.050 496.200 ;
        RECT 746.400 493.350 747.600 494.100 ;
        RECT 724.950 490.950 727.050 493.050 ;
        RECT 727.950 490.950 730.050 493.050 ;
        RECT 743.100 490.950 745.200 493.050 ;
        RECT 746.400 490.950 748.500 493.050 ;
        RECT 751.800 490.950 753.900 493.050 ;
        RECT 725.400 488.400 726.600 490.650 ;
        RECT 743.400 489.900 744.600 490.650 ;
        RECT 725.400 487.050 726.450 488.400 ;
        RECT 742.950 487.800 745.050 489.900 ;
        RECT 752.400 488.400 753.600 490.650 ;
        RECT 721.950 485.400 726.450 487.050 ;
        RECT 721.950 484.950 726.000 485.400 ;
        RECT 743.400 457.050 744.450 487.800 ;
        RECT 752.400 484.050 753.450 488.400 ;
        RECT 751.950 481.950 754.050 484.050 ;
        RECT 761.400 478.050 762.450 496.950 ;
        RECT 769.950 495.000 772.050 499.050 ;
        RECT 776.400 495.600 777.450 517.950 ;
        RECT 809.400 516.450 810.450 560.400 ;
        RECT 818.400 529.200 819.450 566.400 ;
        RECT 823.950 565.800 826.050 567.900 ;
        RECT 823.950 562.650 826.050 564.750 ;
        RECT 824.400 529.200 825.450 562.650 ;
        RECT 833.400 559.050 834.450 577.950 ;
        RECT 836.400 567.900 837.450 583.950 ;
        RECT 835.950 565.800 838.050 567.900 ;
        RECT 836.400 562.050 837.450 565.800 ;
        RECT 835.950 559.950 838.050 562.050 ;
        RECT 832.950 556.950 835.050 559.050 ;
        RECT 839.400 558.450 840.450 628.950 ;
        RECT 854.400 613.050 855.450 643.950 ;
        RECT 857.400 631.050 858.450 646.800 ;
        RECT 856.950 628.950 859.050 631.050 ;
        RECT 844.950 610.950 847.050 613.050 ;
        RECT 853.950 610.950 856.050 613.050 ;
        RECT 841.950 607.950 844.050 610.050 ;
        RECT 842.400 574.050 843.450 607.950 ;
        RECT 845.400 586.050 846.450 610.950 ;
        RECT 860.400 610.050 861.450 655.950 ;
        RECT 863.400 640.050 864.450 661.950 ;
        RECT 866.400 652.050 867.450 673.950 ;
        RECT 875.400 673.050 876.450 676.950 ;
        RECT 874.950 670.950 877.050 673.050 ;
        RECT 865.950 649.950 868.050 652.050 ;
        RECT 868.950 650.100 871.050 652.200 ;
        RECT 869.400 649.350 870.600 650.100 ;
        RECT 868.950 646.950 871.050 649.050 ;
        RECT 871.950 646.950 874.050 649.050 ;
        RECT 872.400 644.400 873.600 646.650 ;
        RECT 862.950 637.950 865.050 640.050 ;
        RECT 872.400 637.050 873.450 644.400 ;
        RECT 871.950 634.950 874.050 637.050 ;
        RECT 865.950 619.950 868.050 622.050 ;
        RECT 859.950 607.950 862.050 610.050 ;
        RECT 853.950 605.100 856.050 607.200 ;
        RECT 861.000 606.600 865.050 607.050 ;
        RECT 854.400 604.350 855.600 605.100 ;
        RECT 860.400 604.950 865.050 606.600 ;
        RECT 860.400 604.350 861.600 604.950 ;
        RECT 850.950 601.950 853.050 604.050 ;
        RECT 853.950 601.950 856.050 604.050 ;
        RECT 856.950 601.950 859.050 604.050 ;
        RECT 859.950 601.950 862.050 604.050 ;
        RECT 847.950 598.950 850.050 601.050 ;
        RECT 851.400 599.400 852.600 601.650 ;
        RECT 857.400 599.400 858.600 601.650 ;
        RECT 844.950 583.950 847.050 586.050 ;
        RECT 844.950 577.950 847.050 580.050 ;
        RECT 841.950 571.950 844.050 574.050 ;
        RECT 845.400 573.600 846.450 577.950 ;
        RECT 848.400 577.050 849.450 598.950 ;
        RECT 851.400 595.050 852.450 599.400 ;
        RECT 850.950 592.950 853.050 595.050 ;
        RECT 857.400 592.050 858.450 599.400 ;
        RECT 856.950 589.950 859.050 592.050 ;
        RECT 857.400 580.050 858.450 589.950 ;
        RECT 850.950 577.950 853.050 580.050 ;
        RECT 856.950 577.950 859.050 580.050 ;
        RECT 847.950 574.950 850.050 577.050 ;
        RECT 851.400 573.600 852.450 577.950 ;
        RECT 866.400 574.050 867.450 619.950 ;
        RECT 878.400 613.050 879.450 685.950 ;
        RECT 883.950 683.100 886.050 685.200 ;
        RECT 889.950 684.000 892.050 688.050 ;
        RECT 884.400 682.350 885.600 683.100 ;
        RECT 890.400 682.350 891.600 684.000 ;
        RECT 883.950 679.950 886.050 682.050 ;
        RECT 886.950 679.950 889.050 682.050 ;
        RECT 889.950 679.950 892.050 682.050 ;
        RECT 892.950 679.950 895.050 682.050 ;
        RECT 887.400 678.900 888.600 679.650 ;
        RECT 886.950 676.800 889.050 678.900 ;
        RECT 893.400 677.400 894.600 679.650 ;
        RECT 893.400 654.450 894.450 677.400 ;
        RECT 893.400 653.400 897.450 654.450 ;
        RECT 880.950 649.950 883.050 652.050 ;
        RECT 889.950 650.100 892.050 652.200 ;
        RECT 896.400 651.600 897.450 653.400 ;
        RECT 899.400 652.050 900.450 721.950 ;
        RECT 877.950 610.950 880.050 613.050 ;
        RECT 881.400 609.450 882.450 649.950 ;
        RECT 890.400 649.350 891.600 650.100 ;
        RECT 896.400 649.350 897.600 651.600 ;
        RECT 898.950 649.950 901.050 652.050 ;
        RECT 886.950 646.950 889.050 649.050 ;
        RECT 889.950 646.950 892.050 649.050 ;
        RECT 892.950 646.950 895.050 649.050 ;
        RECT 895.950 646.950 898.050 649.050 ;
        RECT 887.400 645.900 888.600 646.650 ;
        RECT 886.950 643.800 889.050 645.900 ;
        RECT 893.400 644.400 894.600 646.650 ;
        RECT 893.400 640.050 894.450 644.400 ;
        RECT 898.950 643.950 901.050 646.050 ;
        RECT 892.950 637.950 895.050 640.050 ;
        RECT 889.950 610.950 892.050 613.050 ;
        RECT 881.400 608.400 885.450 609.450 ;
        RECT 884.400 607.200 885.450 608.400 ;
        RECT 868.950 604.950 871.050 607.050 ;
        RECT 877.950 605.100 880.050 607.200 ;
        RECT 883.950 605.100 886.050 607.200 ;
        RECT 869.400 583.050 870.450 604.950 ;
        RECT 878.400 604.350 879.600 605.100 ;
        RECT 884.400 604.350 885.600 605.100 ;
        RECT 874.950 601.950 877.050 604.050 ;
        RECT 877.950 601.950 880.050 604.050 ;
        RECT 880.950 601.950 883.050 604.050 ;
        RECT 883.950 601.950 886.050 604.050 ;
        RECT 875.400 599.400 876.600 601.650 ;
        RECT 881.400 599.400 882.600 601.650 ;
        RECT 875.400 583.050 876.450 599.400 ;
        RECT 877.950 595.950 880.050 598.050 ;
        RECT 868.950 580.950 871.050 583.050 ;
        RECT 874.950 580.950 877.050 583.050 ;
        RECT 878.400 574.200 879.450 595.950 ;
        RECT 881.400 592.050 882.450 599.400 ;
        RECT 883.950 595.950 886.050 598.050 ;
        RECT 880.950 589.950 883.050 592.050 ;
        RECT 845.400 571.350 846.600 573.600 ;
        RECT 851.400 571.350 852.600 573.600 ;
        RECT 859.950 571.950 862.050 574.050 ;
        RECT 862.950 571.950 865.050 574.050 ;
        RECT 865.950 571.950 868.050 574.050 ;
        RECT 871.950 572.100 874.050 574.200 ;
        RECT 877.950 572.100 880.050 574.200 ;
        RECT 844.950 568.950 847.050 571.050 ;
        RECT 847.950 568.950 850.050 571.050 ;
        RECT 850.950 568.950 853.050 571.050 ;
        RECT 853.950 568.950 856.050 571.050 ;
        RECT 841.950 565.950 844.050 568.050 ;
        RECT 848.400 567.900 849.600 568.650 ;
        RECT 854.400 567.900 855.600 568.650 ;
        RECT 836.400 557.400 840.450 558.450 ;
        RECT 832.950 541.950 835.050 544.050 ;
        RECT 817.950 527.100 820.050 529.200 ;
        RECT 823.950 527.100 826.050 529.200 ;
        RECT 829.950 527.100 832.050 529.200 ;
        RECT 818.400 526.350 819.600 527.100 ;
        RECT 824.400 526.350 825.600 527.100 ;
        RECT 814.950 523.950 817.050 526.050 ;
        RECT 817.950 523.950 820.050 526.050 ;
        RECT 820.950 523.950 823.050 526.050 ;
        RECT 823.950 523.950 826.050 526.050 ;
        RECT 806.400 515.400 810.450 516.450 ;
        RECT 815.400 521.400 816.600 523.650 ;
        RECT 821.400 522.000 822.600 523.650 ;
        RECT 796.950 502.950 799.050 505.050 ;
        RECT 797.400 496.200 798.450 502.950 ;
        RECT 770.400 493.350 771.600 495.000 ;
        RECT 776.400 493.350 777.600 495.600 ;
        RECT 784.800 493.950 786.900 496.050 ;
        RECT 787.950 493.950 790.050 496.050 ;
        RECT 796.950 494.100 799.050 496.200 ;
        RECT 766.950 490.950 769.050 493.050 ;
        RECT 769.950 490.950 772.050 493.050 ;
        RECT 772.950 490.950 775.050 493.050 ;
        RECT 775.950 490.950 778.050 493.050 ;
        RECT 767.400 488.400 768.600 490.650 ;
        RECT 773.400 489.900 774.600 490.650 ;
        RECT 785.400 489.900 786.450 493.950 ;
        RECT 754.950 475.950 757.050 478.050 ;
        RECT 760.950 475.950 763.050 478.050 ;
        RECT 706.950 454.950 709.050 457.050 ;
        RECT 718.950 454.950 721.050 457.050 ;
        RECT 742.950 454.950 745.050 457.050 ;
        RECT 748.950 454.950 751.050 457.050 ;
        RECT 671.400 448.350 672.600 450.000 ;
        RECT 676.950 449.100 679.050 451.200 ;
        RECT 677.400 448.350 678.600 449.100 ;
        RECT 682.950 448.950 685.050 451.050 ;
        RECT 694.950 449.100 697.050 451.200 ;
        RECT 700.950 449.100 703.050 451.200 ;
        RECT 661.950 445.950 664.050 448.050 ;
        RECT 667.950 445.950 670.050 448.050 ;
        RECT 670.950 445.950 673.050 448.050 ;
        RECT 673.950 445.950 676.050 448.050 ;
        RECT 676.950 445.950 679.050 448.050 ;
        RECT 658.950 439.950 661.050 442.050 ;
        RECT 649.950 436.950 652.050 439.050 ;
        RECT 634.950 427.950 637.050 430.050 ;
        RECT 652.950 427.950 655.050 430.050 ;
        RECT 646.950 424.950 649.050 427.050 ;
        RECT 623.400 400.050 624.450 416.100 ;
        RECT 629.400 415.350 630.600 417.600 ;
        RECT 634.950 416.100 637.050 418.200 ;
        RECT 635.400 415.350 636.600 416.100 ;
        RECT 628.950 412.950 631.050 415.050 ;
        RECT 631.950 412.950 634.050 415.050 ;
        RECT 634.950 412.950 637.050 415.050 ;
        RECT 637.950 412.950 640.050 415.050 ;
        RECT 632.400 411.900 633.600 412.650 ;
        RECT 638.400 411.900 639.600 412.650 ;
        RECT 631.950 409.800 634.050 411.900 ;
        RECT 622.950 397.950 625.050 400.050 ;
        RECT 632.400 394.050 633.450 409.800 ;
        RECT 637.950 406.950 640.050 411.900 ;
        RECT 638.400 403.050 639.450 406.950 ;
        RECT 637.950 400.950 640.050 403.050 ;
        RECT 634.950 397.950 637.050 400.050 ;
        RECT 631.950 391.950 634.050 394.050 ;
        RECT 631.950 382.950 634.050 385.050 ;
        RECT 622.950 376.950 625.050 379.050 ;
        RECT 617.400 374.400 621.450 375.450 ;
        RECT 617.400 373.200 618.450 374.400 ;
        RECT 596.400 370.350 597.600 372.000 ;
        RECT 601.950 371.100 604.050 373.200 ;
        RECT 602.400 370.350 603.600 371.100 ;
        RECT 610.950 370.950 613.050 373.050 ;
        RECT 616.950 371.100 619.050 373.200 ;
        RECT 623.400 372.600 624.450 376.950 ;
        RECT 592.950 367.950 595.050 370.050 ;
        RECT 595.950 367.950 598.050 370.050 ;
        RECT 598.950 367.950 601.050 370.050 ;
        RECT 601.950 367.950 604.050 370.050 ;
        RECT 571.950 364.800 574.050 366.900 ;
        RECT 580.950 364.950 583.050 367.050 ;
        RECT 583.950 364.950 586.050 367.050 ;
        RECT 589.950 364.950 592.050 367.050 ;
        RECT 593.400 365.400 594.600 367.650 ;
        RECT 599.400 366.900 600.600 367.650 ;
        RECT 572.400 340.050 573.450 364.800 ;
        RECT 590.400 345.450 591.450 364.950 ;
        RECT 593.400 361.050 594.450 365.400 ;
        RECT 598.950 364.800 601.050 366.900 ;
        RECT 592.950 358.950 595.050 361.050 ;
        RECT 593.400 349.050 594.450 358.950 ;
        RECT 592.950 346.950 595.050 349.050 ;
        RECT 590.400 344.400 594.450 345.450 ;
        RECT 571.950 337.950 574.050 340.050 ;
        RECT 577.950 338.100 580.050 340.200 ;
        RECT 583.950 338.100 586.050 340.200 ;
        RECT 578.400 337.350 579.600 338.100 ;
        RECT 584.400 337.350 585.600 338.100 ;
        RECT 589.950 337.950 592.050 340.050 ;
        RECT 574.950 334.950 577.050 337.050 ;
        RECT 577.950 334.950 580.050 337.050 ;
        RECT 580.950 334.950 583.050 337.050 ;
        RECT 583.950 334.950 586.050 337.050 ;
        RECT 571.950 331.950 574.050 334.050 ;
        RECT 575.400 332.400 576.600 334.650 ;
        RECT 581.400 332.400 582.600 334.650 ;
        RECT 572.400 307.050 573.450 331.950 ;
        RECT 571.950 304.950 574.050 307.050 ;
        RECT 563.400 299.400 567.450 300.450 ;
        RECT 554.400 293.400 558.450 294.450 ;
        RECT 548.400 292.350 549.600 293.100 ;
        RECT 554.400 292.350 555.600 293.400 ;
        RECT 547.950 289.950 550.050 292.050 ;
        RECT 550.950 289.950 553.050 292.050 ;
        RECT 553.950 289.950 556.050 292.050 ;
        RECT 551.400 288.900 552.600 289.650 ;
        RECT 550.950 286.800 553.050 288.900 ;
        RECT 556.950 283.950 559.050 289.050 ;
        RECT 544.950 280.950 550.050 283.050 ;
        RECT 556.950 277.950 559.050 280.050 ;
        RECT 541.950 274.950 544.050 277.050 ;
        RECT 517.950 261.450 520.050 262.200 ;
        RECT 524.400 261.450 525.600 261.600 ;
        RECT 500.400 259.350 501.600 260.100 ;
        RECT 506.400 259.350 507.600 261.000 ;
        RECT 512.400 260.400 516.450 261.450 ;
        RECT 499.950 256.950 502.050 259.050 ;
        RECT 502.950 256.950 505.050 259.050 ;
        RECT 505.950 256.950 508.050 259.050 ;
        RECT 508.950 256.950 511.050 259.050 ;
        RECT 503.400 255.000 504.600 256.650 ;
        RECT 493.950 250.950 496.050 253.050 ;
        RECT 502.950 250.950 505.050 255.000 ;
        RECT 509.400 254.400 510.600 256.650 ;
        RECT 509.400 250.050 510.450 254.400 ;
        RECT 508.950 247.950 511.050 250.050 ;
        RECT 502.950 244.950 505.050 247.050 ;
        RECT 490.950 217.950 493.050 220.050 ;
        RECT 488.400 214.350 489.600 216.600 ;
        RECT 493.950 215.100 496.050 217.200 ;
        RECT 499.950 215.100 502.050 217.200 ;
        RECT 494.400 214.350 495.600 215.100 ;
        RECT 484.950 211.950 487.050 214.050 ;
        RECT 487.950 211.950 490.050 214.050 ;
        RECT 490.950 211.950 493.050 214.050 ;
        RECT 493.950 211.950 496.050 214.050 ;
        RECT 485.400 210.900 486.600 211.650 ;
        RECT 484.950 208.800 487.050 210.900 ;
        RECT 491.400 209.400 492.600 211.650 ;
        RECT 487.950 205.950 490.050 208.050 ;
        RECT 478.950 199.950 481.050 202.050 ;
        RECT 481.950 193.950 484.050 196.050 ;
        RECT 482.400 187.050 483.450 193.950 ;
        RECT 481.950 184.950 484.050 187.050 ;
        RECT 476.400 181.350 477.600 183.600 ;
        RECT 484.950 181.950 487.050 184.050 ;
        RECT 475.950 178.950 478.050 181.050 ;
        RECT 478.950 178.950 481.050 181.050 ;
        RECT 479.400 177.900 480.600 178.650 ;
        RECT 478.950 175.800 481.050 177.900 ;
        RECT 485.400 175.050 486.450 181.950 ;
        RECT 488.400 178.050 489.450 205.950 ;
        RECT 491.400 202.050 492.450 209.400 ;
        RECT 500.400 208.050 501.450 215.100 ;
        RECT 503.400 211.050 504.450 244.950 ;
        RECT 515.400 223.050 516.450 260.400 ;
        RECT 517.950 260.400 525.600 261.450 ;
        RECT 517.950 260.100 520.050 260.400 ;
        RECT 518.400 241.050 519.450 260.100 ;
        RECT 524.400 259.350 525.600 260.400 ;
        RECT 529.950 259.950 532.050 265.050 ;
        RECT 535.950 259.950 538.050 262.050 ;
        RECT 538.950 259.950 541.050 262.050 ;
        RECT 547.950 260.100 550.050 262.200 ;
        RECT 523.950 256.950 526.050 259.050 ;
        RECT 526.950 256.950 529.050 259.050 ;
        RECT 520.950 247.950 523.050 250.050 ;
        RECT 517.950 238.950 520.050 241.050 ;
        RECT 508.950 220.950 511.050 223.050 ;
        RECT 514.950 220.950 517.050 223.050 ;
        RECT 505.950 217.950 508.050 220.050 ;
        RECT 502.950 208.950 505.050 211.050 ;
        RECT 499.950 205.950 502.050 208.050 ;
        RECT 490.950 199.950 493.050 202.050 ;
        RECT 496.950 199.950 499.050 202.050 ;
        RECT 497.400 183.600 498.450 199.950 ;
        RECT 506.400 196.050 507.450 217.950 ;
        RECT 509.400 216.600 510.450 220.950 ;
        RECT 509.400 214.350 510.600 216.600 ;
        RECT 517.950 215.100 520.050 217.200 ;
        RECT 518.400 214.350 519.600 215.100 ;
        RECT 509.100 211.950 511.200 214.050 ;
        RECT 512.400 211.950 514.500 214.050 ;
        RECT 517.800 211.950 519.900 214.050 ;
        RECT 512.400 210.900 513.600 211.650 ;
        RECT 521.400 210.900 522.450 247.950 ;
        RECT 526.950 229.950 529.050 232.050 ;
        RECT 527.400 210.900 528.450 229.950 ;
        RECT 536.400 223.050 537.450 259.950 ;
        RECT 529.950 220.950 532.050 223.050 ;
        RECT 535.950 220.950 538.050 223.050 ;
        RECT 511.950 208.800 514.050 210.900 ;
        RECT 520.950 208.800 523.050 210.900 ;
        RECT 526.950 208.800 529.050 210.900 ;
        RECT 530.400 196.050 531.450 220.950 ;
        RECT 539.400 219.450 540.450 259.950 ;
        RECT 548.400 259.350 549.600 260.100 ;
        RECT 544.950 256.950 547.050 259.050 ;
        RECT 547.950 256.950 550.050 259.050 ;
        RECT 550.950 256.950 553.050 259.050 ;
        RECT 551.400 255.900 552.600 256.650 ;
        RECT 550.950 253.800 553.050 255.900 ;
        RECT 553.950 247.950 556.050 250.050 ;
        RECT 554.400 238.050 555.450 247.950 ;
        RECT 553.950 235.950 556.050 238.050 ;
        RECT 550.950 229.950 553.050 232.050 ;
        RECT 541.950 220.950 544.050 223.050 ;
        RECT 536.400 218.400 540.450 219.450 ;
        RECT 536.400 217.200 537.450 218.400 ;
        RECT 535.950 215.100 538.050 217.200 ;
        RECT 542.400 216.600 543.450 220.950 ;
        RECT 536.400 214.350 537.600 215.100 ;
        RECT 542.400 214.350 543.600 216.600 ;
        RECT 535.950 211.950 538.050 214.050 ;
        RECT 538.950 211.950 541.050 214.050 ;
        RECT 541.950 211.950 544.050 214.050 ;
        RECT 544.950 211.950 547.050 214.050 ;
        RECT 539.400 210.900 540.600 211.650 ;
        RECT 545.400 210.900 546.600 211.650 ;
        RECT 538.950 208.800 541.050 210.900 ;
        RECT 544.950 208.800 547.050 210.900 ;
        RECT 505.950 193.950 508.050 196.050 ;
        RECT 529.950 193.950 532.050 196.050 ;
        RECT 511.950 187.950 514.050 190.050 ;
        RECT 532.950 187.950 535.050 190.050 ;
        RECT 497.400 181.350 498.600 183.600 ;
        RECT 502.950 183.000 505.050 187.050 ;
        RECT 508.950 184.950 511.050 187.050 ;
        RECT 503.400 181.350 504.600 183.000 ;
        RECT 493.950 178.950 496.050 181.050 ;
        RECT 496.950 178.950 499.050 181.050 ;
        RECT 499.950 178.950 502.050 181.050 ;
        RECT 502.950 178.950 505.050 181.050 ;
        RECT 487.950 175.950 490.050 178.050 ;
        RECT 494.400 177.900 495.600 178.650 ;
        RECT 493.950 175.800 496.050 177.900 ;
        RECT 500.400 177.000 501.600 178.650 ;
        RECT 466.950 172.950 469.050 175.050 ;
        RECT 484.950 172.950 487.050 175.050 ;
        RECT 499.950 172.950 502.050 177.000 ;
        RECT 505.950 175.950 508.050 178.050 ;
        RECT 484.950 148.950 487.050 151.050 ;
        RECT 478.950 142.950 481.050 145.050 ;
        RECT 428.400 138.450 429.600 138.600 ;
        RECT 425.400 137.400 429.600 138.450 ;
        RECT 413.400 136.350 414.600 137.100 ;
        RECT 403.950 133.950 406.050 136.050 ;
        RECT 406.950 133.950 409.050 136.050 ;
        RECT 409.950 133.950 412.050 136.050 ;
        RECT 412.950 133.950 415.050 136.050 ;
        RECT 404.400 131.400 405.600 133.650 ;
        RECT 410.400 132.900 411.600 133.650 ;
        RECT 404.400 121.050 405.450 131.400 ;
        RECT 409.950 130.800 412.050 132.900 ;
        RECT 419.400 124.050 420.450 137.100 ;
        RECT 428.400 136.350 429.600 137.400 ;
        RECT 433.950 137.100 436.050 139.200 ;
        RECT 442.950 137.100 445.050 139.200 ;
        RECT 448.950 137.100 451.050 139.200 ;
        RECT 454.950 137.100 457.050 139.200 ;
        RECT 460.950 137.100 463.050 139.200 ;
        RECT 434.400 136.350 435.600 137.100 ;
        RECT 427.950 133.950 430.050 136.050 ;
        RECT 430.950 133.950 433.050 136.050 ;
        RECT 433.950 133.950 436.050 136.050 ;
        RECT 421.950 130.800 424.050 132.900 ;
        RECT 431.400 131.400 432.600 133.650 ;
        RECT 422.400 127.050 423.450 130.800 ;
        RECT 421.950 124.950 424.050 127.050 ;
        RECT 418.950 121.950 421.050 124.050 ;
        RECT 403.950 118.950 406.050 121.050 ;
        RECT 431.400 118.050 432.450 131.400 ;
        RECT 400.950 115.950 403.050 118.050 ;
        RECT 430.950 115.950 433.050 118.050 ;
        RECT 401.400 97.050 402.450 115.950 ;
        RECT 443.400 115.050 444.450 137.100 ;
        RECT 449.400 136.350 450.600 137.100 ;
        RECT 455.400 136.350 456.600 137.100 ;
        RECT 448.950 133.950 451.050 136.050 ;
        RECT 451.950 133.950 454.050 136.050 ;
        RECT 454.950 133.950 457.050 136.050 ;
        RECT 452.400 131.400 453.600 133.650 ;
        RECT 452.400 127.050 453.450 131.400 ;
        RECT 461.400 130.050 462.450 137.100 ;
        RECT 466.950 136.050 469.050 139.050 ;
        RECT 472.950 137.100 475.050 139.200 ;
        RECT 479.400 138.600 480.450 142.950 ;
        RECT 485.400 138.600 486.450 148.950 ;
        RECT 506.400 148.050 507.450 175.950 ;
        RECT 509.400 166.050 510.450 184.950 ;
        RECT 508.950 163.950 511.050 166.050 ;
        RECT 505.950 145.950 508.050 148.050 ;
        RECT 490.950 142.950 493.050 145.050 ;
        RECT 473.400 136.350 474.600 137.100 ;
        RECT 479.400 136.350 480.600 138.600 ;
        RECT 485.400 136.350 486.600 138.600 ;
        RECT 463.950 135.000 469.050 136.050 ;
        RECT 463.950 134.400 468.450 135.000 ;
        RECT 463.950 133.950 468.000 134.400 ;
        RECT 472.950 133.950 475.050 136.050 ;
        RECT 475.950 133.950 478.050 136.050 ;
        RECT 478.950 133.950 481.050 136.050 ;
        RECT 481.950 133.950 484.050 136.050 ;
        RECT 484.950 133.950 487.050 136.050 ;
        RECT 476.400 131.400 477.600 133.650 ;
        RECT 482.400 132.900 483.600 133.650 ;
        RECT 491.400 132.900 492.450 142.950 ;
        RECT 493.950 137.100 496.050 139.200 ;
        RECT 505.950 137.100 508.050 139.200 ;
        RECT 476.400 130.050 477.450 131.400 ;
        RECT 481.950 130.800 484.050 132.900 ;
        RECT 490.950 130.800 493.050 132.900 ;
        RECT 494.400 130.050 495.450 137.100 ;
        RECT 506.400 136.350 507.600 137.100 ;
        RECT 502.950 133.950 505.050 136.050 ;
        RECT 505.950 133.950 508.050 136.050 ;
        RECT 503.400 131.400 504.600 133.650 ;
        RECT 460.950 127.950 463.050 130.050 ;
        RECT 451.950 124.950 454.050 127.050 ;
        RECT 475.950 124.950 478.050 130.050 ;
        RECT 493.950 127.950 496.050 130.050 ;
        RECT 463.950 118.950 466.050 121.050 ;
        RECT 487.950 118.950 490.050 121.050 ;
        RECT 406.950 112.950 409.050 115.050 ;
        RECT 442.950 112.950 445.050 115.050 ;
        RECT 407.400 105.600 408.450 112.950 ;
        RECT 424.950 109.950 427.050 112.050 ;
        RECT 439.950 109.950 442.050 112.050 ;
        RECT 407.400 103.350 408.600 105.600 ;
        RECT 412.950 104.100 415.050 106.200 ;
        RECT 421.950 104.100 424.050 106.200 ;
        RECT 413.400 103.350 414.600 104.100 ;
        RECT 406.950 100.950 409.050 103.050 ;
        RECT 409.950 100.950 412.050 103.050 ;
        RECT 412.950 100.950 415.050 103.050 ;
        RECT 415.950 100.950 418.050 103.050 ;
        RECT 403.950 97.950 406.050 100.050 ;
        RECT 410.400 98.400 411.600 100.650 ;
        RECT 416.400 99.900 417.600 100.650 ;
        RECT 400.950 94.950 403.050 97.050 ;
        RECT 404.400 70.050 405.450 97.950 ;
        RECT 410.400 85.050 411.450 98.400 ;
        RECT 415.950 97.800 418.050 99.900 ;
        RECT 412.950 94.950 415.050 97.050 ;
        RECT 409.950 82.950 412.050 85.050 ;
        RECT 388.950 67.950 391.050 70.050 ;
        RECT 397.950 67.950 400.050 70.050 ;
        RECT 403.950 67.950 406.050 70.050 ;
        RECT 385.950 40.950 388.050 43.050 ;
        RECT 379.950 26.100 382.050 28.200 ;
        RECT 380.400 25.350 381.600 26.100 ;
        RECT 377.100 22.950 379.200 25.050 ;
        RECT 380.400 22.950 382.500 25.050 ;
        RECT 385.800 22.950 387.900 25.050 ;
        RECT 377.400 21.450 378.600 22.650 ;
        RECT 374.400 20.400 378.600 21.450 ;
        RECT 386.400 21.000 387.600 22.650 ;
        RECT 275.550 9.600 277.650 11.700 ;
        RECT 301.950 10.950 304.050 13.050 ;
        RECT 311.550 11.700 312.750 18.300 ;
        RECT 385.950 16.950 388.050 21.000 ;
        RECT 389.400 13.050 390.450 67.950 ;
        RECT 397.800 64.200 399.900 66.300 ;
        RECT 406.800 64.500 408.900 66.600 ;
        RECT 391.950 60.450 394.050 64.050 ;
        RECT 395.400 60.450 396.600 60.600 ;
        RECT 391.950 60.000 396.600 60.450 ;
        RECT 392.400 59.400 396.600 60.000 ;
        RECT 395.400 58.350 396.600 59.400 ;
        RECT 395.100 55.950 397.200 58.050 ;
        RECT 398.100 51.600 399.000 64.200 ;
        RECT 404.400 61.350 405.600 63.600 ;
        RECT 404.100 58.950 406.200 61.050 ;
        RECT 399.900 57.900 402.000 58.200 ;
        RECT 408.000 57.900 408.900 64.500 ;
        RECT 399.900 57.000 408.900 57.900 ;
        RECT 399.900 56.100 402.000 57.000 ;
        RECT 405.000 55.200 407.100 56.100 ;
        RECT 399.900 54.000 407.100 55.200 ;
        RECT 399.900 53.100 402.000 54.000 ;
        RECT 397.500 49.500 399.600 51.600 ;
        RECT 404.100 50.100 406.200 52.200 ;
        RECT 408.000 51.900 408.900 57.000 ;
        RECT 409.800 55.950 411.900 58.050 ;
        RECT 407.400 49.800 409.500 51.900 ;
        RECT 404.400 47.550 405.600 49.800 ;
        RECT 400.950 40.950 403.050 43.050 ;
        RECT 401.400 30.450 402.450 40.950 ;
        RECT 404.400 33.450 405.450 47.550 ;
        RECT 404.400 33.000 408.450 33.450 ;
        RECT 404.400 32.400 409.050 33.000 ;
        RECT 401.400 29.400 405.450 30.450 ;
        RECT 394.950 26.100 397.050 28.200 ;
        RECT 404.400 27.600 405.450 29.400 ;
        RECT 406.950 28.950 409.050 32.400 ;
        RECT 395.400 22.050 396.450 26.100 ;
        RECT 404.400 25.350 405.600 27.600 ;
        RECT 400.950 22.950 403.050 25.050 ;
        RECT 403.950 22.950 406.050 25.050 ;
        RECT 406.950 22.950 409.050 25.050 ;
        RECT 394.950 19.950 397.050 22.050 ;
        RECT 401.400 21.900 402.600 22.650 ;
        RECT 400.950 19.800 403.050 21.900 ;
        RECT 407.400 21.000 408.600 22.650 ;
        RECT 406.950 16.950 409.050 21.000 ;
        RECT 413.400 19.050 414.450 94.950 ;
        RECT 422.400 84.450 423.450 104.100 ;
        RECT 425.400 99.900 426.450 109.950 ;
        RECT 433.950 104.100 436.050 106.200 ;
        RECT 440.400 105.600 441.450 109.950 ;
        RECT 434.400 103.350 435.600 104.100 ;
        RECT 440.400 103.350 441.600 105.600 ;
        RECT 445.950 103.950 448.050 106.050 ;
        RECT 457.950 104.100 460.050 106.200 ;
        RECT 464.400 105.600 465.450 118.950 ;
        RECT 488.400 115.050 489.450 118.950 ;
        RECT 503.400 118.050 504.450 131.400 ;
        RECT 496.950 115.950 499.050 118.050 ;
        RECT 502.950 115.950 505.050 118.050 ;
        RECT 472.950 112.950 475.050 115.050 ;
        RECT 487.950 112.950 490.050 115.050 ;
        RECT 430.950 100.950 433.050 103.050 ;
        RECT 433.950 100.950 436.050 103.050 ;
        RECT 436.950 100.950 439.050 103.050 ;
        RECT 439.950 100.950 442.050 103.050 ;
        RECT 424.950 97.800 427.050 99.900 ;
        RECT 431.400 99.000 432.600 100.650 ;
        RECT 430.950 94.950 433.050 99.000 ;
        RECT 437.400 98.400 438.600 100.650 ;
        RECT 437.400 91.050 438.450 98.400 ;
        RECT 436.950 88.950 439.050 91.050 ;
        RECT 424.950 84.450 427.050 85.050 ;
        RECT 422.400 83.400 427.050 84.450 ;
        RECT 424.950 82.950 427.050 83.400 ;
        RECT 425.400 60.600 426.450 82.950 ;
        RECT 439.950 70.950 442.050 73.050 ;
        RECT 425.400 58.350 426.600 60.600 ;
        RECT 430.950 59.100 433.050 61.200 ;
        RECT 431.400 58.350 432.600 59.100 ;
        RECT 424.950 55.950 427.050 58.050 ;
        RECT 427.950 55.950 430.050 58.050 ;
        RECT 430.950 55.950 433.050 58.050 ;
        RECT 433.950 55.950 436.050 58.050 ;
        RECT 428.400 53.400 429.600 55.650 ;
        RECT 434.400 54.900 435.600 55.650 ;
        RECT 440.400 54.900 441.450 70.950 ;
        RECT 446.400 60.450 447.450 103.950 ;
        RECT 458.400 103.350 459.600 104.100 ;
        RECT 464.400 103.350 465.600 105.600 ;
        RECT 469.950 103.950 472.050 106.050 ;
        RECT 454.950 100.950 457.050 103.050 ;
        RECT 457.950 100.950 460.050 103.050 ;
        RECT 460.950 100.950 463.050 103.050 ;
        RECT 463.950 100.950 466.050 103.050 ;
        RECT 455.400 99.000 456.600 100.650 ;
        RECT 454.950 94.950 457.050 99.000 ;
        RECT 461.400 98.400 462.600 100.650 ;
        RECT 461.400 96.450 462.450 98.400 ;
        RECT 461.400 95.400 465.450 96.450 ;
        RECT 455.400 60.600 456.450 94.950 ;
        RECT 464.400 73.050 465.450 95.400 ;
        RECT 470.400 94.050 471.450 103.950 ;
        RECT 469.950 91.950 472.050 94.050 ;
        RECT 466.950 88.950 469.050 91.050 ;
        RECT 463.950 70.950 466.050 73.050 ;
        RECT 467.400 70.050 468.450 88.950 ;
        RECT 470.400 85.050 471.450 91.950 ;
        RECT 469.950 82.950 472.050 85.050 ;
        RECT 473.400 79.050 474.450 112.950 ;
        RECT 484.950 109.950 487.050 112.050 ;
        RECT 485.400 106.200 486.450 109.950 ;
        RECT 478.950 104.100 481.050 106.200 ;
        RECT 484.950 104.100 487.050 106.200 ;
        RECT 479.400 103.350 480.600 104.100 ;
        RECT 485.400 103.350 486.600 104.100 ;
        RECT 478.950 100.950 481.050 103.050 ;
        RECT 481.950 100.950 484.050 103.050 ;
        RECT 484.950 100.950 487.050 103.050 ;
        RECT 487.950 100.950 490.050 103.050 ;
        RECT 482.400 98.400 483.600 100.650 ;
        RECT 488.400 98.400 489.600 100.650 ;
        RECT 497.400 99.900 498.450 115.950 ;
        RECT 512.400 109.050 513.450 187.950 ;
        RECT 517.950 182.100 520.050 184.200 ;
        RECT 523.950 183.000 526.050 187.050 ;
        RECT 518.400 181.350 519.600 182.100 ;
        RECT 524.400 181.350 525.600 183.000 ;
        RECT 517.950 178.950 520.050 181.050 ;
        RECT 520.950 178.950 523.050 181.050 ;
        RECT 523.950 178.950 526.050 181.050 ;
        RECT 526.950 178.950 529.050 181.050 ;
        RECT 521.400 176.400 522.600 178.650 ;
        RECT 527.400 177.900 528.600 178.650 ;
        RECT 533.400 177.900 534.450 187.950 ;
        RECT 551.400 187.050 552.450 229.950 ;
        RECT 557.400 223.050 558.450 277.950 ;
        RECT 560.400 255.900 561.450 298.950 ;
        RECT 563.400 280.050 564.450 299.400 ;
        RECT 568.950 298.950 571.050 301.050 ;
        RECT 569.400 294.600 570.450 298.950 ;
        RECT 575.400 298.050 576.450 332.400 ;
        RECT 581.400 319.050 582.450 332.400 ;
        RECT 580.950 316.950 583.050 319.050 ;
        RECT 590.400 307.050 591.450 337.950 ;
        RECT 593.400 328.050 594.450 344.400 ;
        RECT 601.950 338.100 604.050 340.200 ;
        RECT 602.400 337.350 603.600 338.100 ;
        RECT 598.950 334.950 601.050 337.050 ;
        RECT 601.950 334.950 604.050 337.050 ;
        RECT 604.950 334.950 607.050 337.050 ;
        RECT 592.950 325.950 595.050 328.050 ;
        RECT 611.400 324.450 612.450 370.950 ;
        RECT 617.400 370.350 618.600 371.100 ;
        RECT 623.400 370.350 624.600 372.600 ;
        RECT 616.950 367.950 619.050 370.050 ;
        RECT 619.950 367.950 622.050 370.050 ;
        RECT 622.950 367.950 625.050 370.050 ;
        RECT 620.400 365.400 621.600 367.650 ;
        RECT 620.400 361.050 621.450 365.400 ;
        RECT 632.400 361.050 633.450 382.950 ;
        RECT 635.400 373.050 636.450 397.950 ;
        RECT 640.950 382.950 643.050 385.050 ;
        RECT 634.950 370.950 637.050 373.050 ;
        RECT 641.400 372.600 642.450 382.950 ;
        RECT 641.400 370.350 642.600 372.600 ;
        RECT 637.950 367.950 640.050 370.050 ;
        RECT 640.950 367.950 643.050 370.050 ;
        RECT 638.400 366.900 639.600 367.650 ;
        RECT 637.950 364.800 640.050 366.900 ;
        RECT 619.950 360.450 622.050 361.050 ;
        RECT 608.400 323.400 612.450 324.450 ;
        RECT 617.400 359.400 622.050 360.450 ;
        RECT 601.950 307.950 604.050 310.050 ;
        RECT 583.950 304.950 586.050 307.050 ;
        RECT 589.950 304.950 592.050 307.050 ;
        RECT 569.400 292.350 570.600 294.600 ;
        RECT 574.950 294.000 577.050 298.050 ;
        RECT 575.400 292.350 576.600 294.000 ;
        RECT 568.950 289.950 571.050 292.050 ;
        RECT 571.950 289.950 574.050 292.050 ;
        RECT 574.950 289.950 577.050 292.050 ;
        RECT 577.950 289.950 580.050 292.050 ;
        RECT 572.400 288.900 573.600 289.650 ;
        RECT 571.950 286.800 574.050 288.900 ;
        RECT 578.400 287.400 579.600 289.650 ;
        RECT 572.400 283.050 573.450 286.800 ;
        RECT 571.950 280.950 574.050 283.050 ;
        RECT 562.950 277.950 565.050 280.050 ;
        RECT 571.950 277.800 574.050 279.900 ;
        RECT 565.950 274.950 568.050 277.050 ;
        RECT 566.400 261.600 567.450 274.950 ;
        RECT 572.400 261.600 573.450 277.800 ;
        RECT 578.400 271.050 579.450 287.400 ;
        RECT 580.950 283.950 583.050 286.050 ;
        RECT 577.950 268.950 580.050 271.050 ;
        RECT 566.400 259.350 567.600 261.600 ;
        RECT 572.400 259.350 573.600 261.600 ;
        RECT 577.950 259.950 580.050 262.050 ;
        RECT 565.950 256.950 568.050 259.050 ;
        RECT 568.950 256.950 571.050 259.050 ;
        RECT 571.950 256.950 574.050 259.050 ;
        RECT 559.950 253.800 562.050 255.900 ;
        RECT 569.400 254.400 570.600 256.650 ;
        RECT 559.950 238.950 562.050 241.050 ;
        RECT 556.950 220.950 559.050 223.050 ;
        RECT 560.400 211.050 561.450 238.950 ;
        RECT 569.400 220.050 570.450 254.400 ;
        RECT 578.400 232.050 579.450 259.950 ;
        RECT 581.400 255.900 582.450 283.950 ;
        RECT 584.400 262.050 585.450 304.950 ;
        RECT 590.400 294.450 591.450 304.950 ;
        RECT 587.400 293.400 591.450 294.450 ;
        RECT 587.400 288.900 588.450 293.400 ;
        RECT 592.950 293.100 595.050 295.200 ;
        RECT 593.400 292.350 594.600 293.100 ;
        RECT 592.950 289.950 595.050 292.050 ;
        RECT 595.950 289.950 598.050 292.050 ;
        RECT 596.400 288.900 597.600 289.650 ;
        RECT 586.950 286.800 589.050 288.900 ;
        RECT 595.950 286.800 598.050 288.900 ;
        RECT 602.400 280.050 603.450 307.950 ;
        RECT 601.950 277.950 604.050 280.050 ;
        RECT 583.950 259.950 586.050 262.050 ;
        RECT 589.950 261.000 592.050 265.050 ;
        RECT 608.400 261.600 609.450 323.400 ;
        RECT 610.950 319.950 613.050 322.050 ;
        RECT 611.400 294.600 612.450 319.950 ;
        RECT 617.400 310.050 618.450 359.400 ;
        RECT 619.950 358.950 622.050 359.400 ;
        RECT 631.950 358.950 634.050 361.050 ;
        RECT 647.400 345.450 648.450 424.950 ;
        RECT 653.400 418.200 654.450 427.950 ;
        RECT 652.950 416.100 655.050 418.200 ;
        RECT 653.400 415.350 654.600 416.100 ;
        RECT 652.950 412.950 655.050 415.050 ;
        RECT 655.950 412.950 658.050 415.050 ;
        RECT 656.400 411.900 657.600 412.650 ;
        RECT 662.400 412.050 663.450 445.950 ;
        RECT 668.400 444.000 669.600 445.650 ;
        RECT 667.950 439.950 670.050 444.000 ;
        RECT 674.400 443.400 675.600 445.650 ;
        RECT 674.400 439.050 675.450 443.400 ;
        RECT 673.950 436.950 676.050 439.050 ;
        RECT 679.950 421.950 682.050 424.050 ;
        RECT 673.950 416.100 676.050 418.200 ;
        RECT 680.400 417.600 681.450 421.950 ;
        RECT 683.400 421.050 684.450 448.950 ;
        RECT 695.400 448.350 696.600 449.100 ;
        RECT 701.400 448.350 702.600 449.100 ;
        RECT 691.950 445.950 694.050 448.050 ;
        RECT 694.950 445.950 697.050 448.050 ;
        RECT 697.950 445.950 700.050 448.050 ;
        RECT 700.950 445.950 703.050 448.050 ;
        RECT 692.400 445.050 693.600 445.650 ;
        RECT 688.950 443.400 693.600 445.050 ;
        RECT 698.400 443.400 699.600 445.650 ;
        RECT 688.950 442.950 693.000 443.400 ;
        RECT 698.400 433.050 699.450 443.400 ;
        RECT 707.400 442.050 708.450 454.950 ;
        RECT 718.950 449.100 721.050 451.200 ;
        RECT 724.950 450.000 727.050 454.050 ;
        RECT 733.950 451.950 736.050 454.050 ;
        RECT 719.400 448.350 720.600 449.100 ;
        RECT 725.400 448.350 726.600 450.000 ;
        RECT 715.950 445.950 718.050 448.050 ;
        RECT 718.950 445.950 721.050 448.050 ;
        RECT 721.950 445.950 724.050 448.050 ;
        RECT 724.950 445.950 727.050 448.050 ;
        RECT 730.950 445.950 733.050 448.050 ;
        RECT 716.400 443.400 717.600 445.650 ;
        RECT 722.400 444.000 723.600 445.650 ;
        RECT 706.950 439.950 709.050 442.050 ;
        RECT 700.950 436.950 703.050 439.050 ;
        RECT 697.950 430.950 700.050 433.050 ;
        RECT 694.950 421.950 697.050 424.050 ;
        RECT 682.950 418.950 685.050 421.050 ;
        RECT 688.950 418.950 691.050 421.050 ;
        RECT 674.400 415.350 675.600 416.100 ;
        RECT 680.400 415.350 681.600 417.600 ;
        RECT 670.950 412.950 673.050 415.050 ;
        RECT 673.950 412.950 676.050 415.050 ;
        RECT 676.950 412.950 679.050 415.050 ;
        RECT 679.950 412.950 682.050 415.050 ;
        RECT 655.950 409.800 658.050 411.900 ;
        RECT 661.950 409.950 664.050 412.050 ;
        RECT 671.400 411.000 672.600 412.650 ;
        RECT 677.400 411.000 678.600 412.650 ;
        RECT 655.950 400.950 658.050 403.050 ;
        RECT 649.950 391.950 652.050 394.050 ;
        RECT 650.400 366.900 651.450 391.950 ;
        RECT 656.400 372.600 657.450 400.950 ;
        RECT 662.400 388.050 663.450 409.950 ;
        RECT 670.950 406.950 673.050 411.000 ;
        RECT 676.950 406.950 679.050 411.000 ;
        RECT 682.950 409.950 685.050 412.050 ;
        RECT 683.400 394.050 684.450 409.950 ;
        RECT 689.400 409.050 690.450 418.950 ;
        RECT 695.400 417.600 696.450 421.950 ;
        RECT 701.400 417.600 702.450 436.950 ;
        RECT 695.400 415.350 696.600 417.600 ;
        RECT 701.400 415.350 702.600 417.600 ;
        RECT 706.950 415.950 709.050 421.050 ;
        RECT 716.400 417.450 717.450 443.400 ;
        RECT 721.950 439.950 724.050 444.000 ;
        RECT 722.400 421.050 723.450 439.950 ;
        RECT 724.950 430.950 727.050 433.050 ;
        RECT 721.950 418.950 724.050 421.050 ;
        RECT 713.400 416.400 717.450 417.450 ;
        RECT 694.950 412.950 697.050 415.050 ;
        RECT 697.950 412.950 700.050 415.050 ;
        RECT 700.950 412.950 703.050 415.050 ;
        RECT 703.950 412.950 706.050 415.050 ;
        RECT 698.400 410.400 699.600 412.650 ;
        RECT 704.400 411.900 705.600 412.650 ;
        RECT 698.400 409.050 699.450 410.400 ;
        RECT 703.950 409.800 706.050 411.900 ;
        RECT 706.950 409.950 709.050 412.050 ;
        RECT 688.950 406.950 691.050 409.050 ;
        RECT 697.950 406.950 700.050 409.050 ;
        RECT 688.950 397.950 691.050 400.050 ;
        RECT 689.400 394.050 690.450 397.950 ;
        RECT 682.950 391.950 685.050 394.050 ;
        RECT 688.950 391.950 691.050 394.050 ;
        RECT 661.950 385.950 664.050 388.050 ;
        RECT 673.950 385.950 676.050 388.050 ;
        RECT 682.950 385.950 685.050 388.050 ;
        RECT 661.950 382.800 664.050 384.900 ;
        RECT 662.400 372.600 663.450 382.800 ;
        RECT 656.400 370.350 657.600 372.600 ;
        RECT 662.400 370.350 663.600 372.600 ;
        RECT 655.950 367.950 658.050 370.050 ;
        RECT 658.950 367.950 661.050 370.050 ;
        RECT 661.950 367.950 664.050 370.050 ;
        RECT 664.950 367.950 667.050 370.050 ;
        RECT 659.400 366.900 660.600 367.650 ;
        RECT 649.950 364.800 652.050 366.900 ;
        RECT 658.950 364.800 661.050 366.900 ;
        RECT 665.400 365.400 666.600 367.650 ;
        RECT 674.400 366.900 675.450 385.950 ;
        RECT 683.400 372.600 684.450 385.950 ;
        RECT 689.400 372.600 690.450 391.950 ;
        RECT 694.950 379.950 697.050 382.050 ;
        RECT 683.400 370.350 684.600 372.600 ;
        RECT 689.400 370.350 690.600 372.600 ;
        RECT 679.950 367.950 682.050 370.050 ;
        RECT 682.950 367.950 685.050 370.050 ;
        RECT 685.950 367.950 688.050 370.050 ;
        RECT 688.950 367.950 691.050 370.050 ;
        RECT 680.400 366.900 681.600 367.650 ;
        RECT 644.400 344.400 648.450 345.450 ;
        RECT 625.950 338.100 628.050 340.200 ;
        RECT 637.950 338.100 640.050 340.200 ;
        RECT 626.400 337.350 627.600 338.100 ;
        RECT 623.100 334.950 625.200 337.050 ;
        RECT 626.400 334.950 628.500 337.050 ;
        RECT 631.800 334.950 633.900 337.050 ;
        RECT 623.400 332.400 624.600 334.650 ;
        RECT 638.400 334.050 639.450 338.100 ;
        RECT 623.400 328.050 624.450 332.400 ;
        RECT 637.950 331.950 640.050 334.050 ;
        RECT 622.950 325.950 625.050 328.050 ;
        RECT 619.950 316.950 622.050 319.050 ;
        RECT 616.950 307.950 619.050 310.050 ;
        RECT 620.400 294.600 621.450 316.950 ;
        RECT 638.400 301.050 639.450 331.950 ;
        RECT 644.400 331.050 645.450 344.400 ;
        RECT 647.400 334.950 649.500 337.050 ;
        RECT 652.800 334.950 654.900 337.050 ;
        RECT 653.400 333.900 654.600 334.650 ;
        RECT 652.950 331.800 655.050 333.900 ;
        RECT 643.950 328.950 646.050 331.050 ;
        RECT 649.950 328.950 652.050 331.050 ;
        RECT 637.950 298.950 640.050 301.050 ;
        RECT 611.400 292.350 612.600 294.600 ;
        RECT 620.400 292.350 621.600 294.600 ;
        RECT 611.100 289.950 613.200 292.050 ;
        RECT 616.500 289.950 618.600 292.050 ;
        RECT 619.800 289.950 621.900 292.050 ;
        RECT 637.950 289.950 640.050 292.050 ;
        RECT 640.950 289.950 643.050 292.050 ;
        RECT 643.950 289.950 646.050 292.050 ;
        RECT 617.400 288.900 618.600 289.650 ;
        RECT 624.000 288.900 628.050 289.050 ;
        RECT 616.950 286.800 619.050 288.900 ;
        RECT 622.950 286.950 628.050 288.900 ;
        RECT 622.950 286.800 625.050 286.950 ;
        RECT 634.950 283.950 637.050 289.050 ;
        RECT 641.400 288.900 642.600 289.650 ;
        RECT 640.950 286.800 643.050 288.900 ;
        RECT 634.950 274.950 637.050 277.050 ;
        RECT 590.400 259.350 591.600 261.000 ;
        RECT 608.400 259.350 609.600 261.600 ;
        RECT 613.950 260.100 616.050 262.200 ;
        RECT 635.400 261.600 636.450 274.950 ;
        RECT 646.950 262.950 649.050 265.050 ;
        RECT 614.400 259.350 615.600 260.100 ;
        RECT 635.400 259.350 636.600 261.600 ;
        RECT 643.950 260.100 646.050 262.200 ;
        RECT 586.950 256.950 589.050 259.050 ;
        RECT 589.950 256.950 592.050 259.050 ;
        RECT 592.950 256.950 595.050 259.050 ;
        RECT 607.950 256.950 610.050 259.050 ;
        RECT 610.950 256.950 613.050 259.050 ;
        RECT 613.950 256.950 616.050 259.050 ;
        RECT 616.950 256.950 619.050 259.050 ;
        RECT 631.950 256.950 634.050 259.050 ;
        RECT 634.950 256.950 637.050 259.050 ;
        RECT 637.950 256.950 640.050 259.050 ;
        RECT 587.400 255.900 588.600 256.650 ;
        RECT 580.950 253.800 583.050 255.900 ;
        RECT 586.950 253.800 589.050 255.900 ;
        RECT 593.400 254.400 594.600 256.650 ;
        RECT 611.400 254.400 612.600 256.650 ;
        RECT 617.400 255.000 618.600 256.650 ;
        RECT 593.400 250.050 594.450 254.400 ;
        RECT 611.400 250.050 612.450 254.400 ;
        RECT 616.950 250.950 619.050 255.000 ;
        RECT 619.950 253.950 622.050 256.050 ;
        RECT 632.400 255.900 633.600 256.650 ;
        RECT 638.400 255.900 639.600 256.650 ;
        RECT 644.400 255.900 645.450 260.100 ;
        RECT 586.950 247.950 589.050 250.050 ;
        RECT 592.950 247.950 595.050 250.050 ;
        RECT 610.950 247.950 613.050 250.050 ;
        RECT 577.950 229.950 580.050 232.050 ;
        RECT 580.350 225.300 582.450 227.400 ;
        RECT 568.950 217.950 571.050 220.050 ;
        RECT 581.250 218.700 582.450 225.300 ;
        RECT 580.350 216.600 582.450 218.700 ;
        RECT 583.950 217.950 586.050 220.050 ;
        RECT 563.100 211.950 565.200 214.050 ;
        RECT 568.500 211.950 570.600 214.050 ;
        RECT 574.950 211.950 577.050 214.050 ;
        RECT 559.950 208.950 562.050 211.050 ;
        RECT 569.400 210.900 570.600 211.650 ;
        RECT 575.400 210.900 576.600 211.650 ;
        RECT 568.950 208.800 571.050 210.900 ;
        RECT 574.950 208.800 577.050 210.900 ;
        RECT 581.250 203.700 582.450 216.600 ;
        RECT 580.350 201.600 582.450 203.700 ;
        RECT 584.400 190.050 585.450 217.950 ;
        RECT 587.400 193.050 588.450 247.950 ;
        RECT 616.350 225.300 618.450 227.400 ;
        RECT 595.650 223.500 597.750 224.400 ;
        RECT 595.650 222.300 599.850 223.500 ;
        RECT 592.950 215.100 595.050 217.200 ;
        RECT 593.400 214.350 594.600 215.100 ;
        RECT 592.800 211.950 594.900 214.050 ;
        RECT 598.650 203.700 599.850 222.300 ;
        RECT 601.950 220.950 604.050 223.050 ;
        RECT 602.400 216.600 603.450 220.950 ;
        RECT 617.250 218.700 618.450 225.300 ;
        RECT 616.350 216.600 618.450 218.700 ;
        RECT 602.400 214.350 603.600 216.600 ;
        RECT 601.950 211.950 604.050 214.050 ;
        RECT 610.950 211.950 613.050 214.050 ;
        RECT 611.400 210.900 612.600 211.650 ;
        RECT 610.950 208.800 613.050 210.900 ;
        RECT 617.250 203.700 618.450 216.600 ;
        RECT 598.050 201.600 600.150 203.700 ;
        RECT 616.350 201.600 618.450 203.700 ;
        RECT 620.400 199.050 621.450 253.950 ;
        RECT 631.950 250.950 634.050 255.900 ;
        RECT 637.950 253.800 640.050 255.900 ;
        RECT 643.950 253.800 646.050 255.900 ;
        RECT 637.950 247.950 643.050 250.050 ;
        RECT 631.650 223.500 633.750 224.400 ;
        RECT 637.950 223.950 640.050 226.050 ;
        RECT 631.650 222.300 635.850 223.500 ;
        RECT 622.950 215.100 625.050 217.200 ;
        RECT 628.950 215.100 631.050 217.200 ;
        RECT 601.950 196.950 604.050 199.050 ;
        RECT 619.950 196.950 622.050 199.050 ;
        RECT 586.950 190.950 589.050 193.050 ;
        RECT 583.950 187.950 586.050 190.050 ;
        RECT 550.950 184.950 553.050 187.050 ;
        RECT 556.950 184.950 559.050 187.050 ;
        RECT 584.400 186.450 585.450 187.950 ;
        RECT 584.400 185.400 588.450 186.450 ;
        RECT 538.950 182.100 541.050 184.200 ;
        RECT 544.950 182.100 547.050 184.200 ;
        RECT 521.400 172.050 522.450 176.400 ;
        RECT 526.950 175.800 529.050 177.900 ;
        RECT 532.950 175.800 535.050 177.900 ;
        RECT 520.950 169.950 523.050 172.050 ;
        RECT 521.400 151.050 522.450 169.950 ;
        RECT 520.950 148.950 523.050 151.050 ;
        RECT 526.950 148.950 529.050 151.050 ;
        RECT 527.400 145.050 528.450 148.950 ;
        RECT 526.950 142.950 529.050 145.050 ;
        RECT 517.950 136.950 520.050 139.050 ;
        RECT 527.400 138.600 528.450 142.950 ;
        RECT 518.400 109.050 519.450 136.950 ;
        RECT 527.400 136.350 528.600 138.600 ;
        RECT 532.950 138.000 535.050 142.050 ;
        RECT 533.400 136.350 534.600 138.000 ;
        RECT 523.950 133.950 526.050 136.050 ;
        RECT 526.950 133.950 529.050 136.050 ;
        RECT 529.950 133.950 532.050 136.050 ;
        RECT 532.950 133.950 535.050 136.050 ;
        RECT 524.400 131.400 525.600 133.650 ;
        RECT 530.400 131.400 531.600 133.650 ;
        RECT 539.400 133.050 540.450 182.100 ;
        RECT 545.400 181.350 546.600 182.100 ;
        RECT 544.950 178.950 547.050 181.050 ;
        RECT 547.950 178.950 550.050 181.050 ;
        RECT 548.400 176.400 549.600 178.650 ;
        RECT 548.400 157.050 549.450 176.400 ;
        RECT 557.400 175.050 558.450 184.950 ;
        RECT 562.950 182.100 565.050 184.200 ;
        RECT 570.000 183.600 574.050 184.050 ;
        RECT 563.400 181.350 564.600 182.100 ;
        RECT 569.400 181.950 574.050 183.600 ;
        RECT 577.950 181.950 580.050 184.050 ;
        RECT 587.400 183.600 588.450 185.400 ;
        RECT 569.400 181.350 570.600 181.950 ;
        RECT 562.950 178.950 565.050 181.050 ;
        RECT 565.950 178.950 568.050 181.050 ;
        RECT 568.950 178.950 571.050 181.050 ;
        RECT 566.400 176.400 567.600 178.650 ;
        RECT 556.950 172.950 559.050 175.050 ;
        RECT 566.400 172.050 567.450 176.400 ;
        RECT 565.950 169.950 568.050 172.050 ;
        RECT 578.400 163.050 579.450 181.950 ;
        RECT 587.400 181.350 588.600 183.600 ;
        RECT 592.950 182.100 595.050 184.200 ;
        RECT 593.400 181.350 594.600 182.100 ;
        RECT 598.950 181.950 601.050 184.050 ;
        RECT 583.950 178.950 586.050 181.050 ;
        RECT 586.950 178.950 589.050 181.050 ;
        RECT 589.950 178.950 592.050 181.050 ;
        RECT 592.950 178.950 595.050 181.050 ;
        RECT 584.400 177.000 585.600 178.650 ;
        RECT 590.400 177.000 591.600 178.650 ;
        RECT 583.950 172.950 586.050 177.000 ;
        RECT 589.950 172.950 592.050 177.000 ;
        RECT 577.950 160.950 580.050 163.050 ;
        RECT 547.950 154.950 550.050 157.050 ;
        RECT 548.400 142.200 549.450 154.950 ;
        RECT 590.400 151.050 591.450 172.950 ;
        RECT 589.950 148.950 592.050 151.050 ;
        RECT 592.950 145.950 595.050 148.050 ;
        RECT 547.950 140.100 550.050 142.200 ;
        RECT 593.400 139.200 594.450 145.950 ;
        RECT 547.950 136.950 550.050 139.050 ;
        RECT 554.400 138.450 555.600 138.600 ;
        RECT 554.400 137.400 561.450 138.450 ;
        RECT 548.400 136.350 549.600 136.950 ;
        RECT 554.400 136.350 555.600 137.400 ;
        RECT 547.950 133.950 550.050 136.050 ;
        RECT 550.950 133.950 553.050 136.050 ;
        RECT 553.950 133.950 556.050 136.050 ;
        RECT 524.400 124.050 525.450 131.400 ;
        RECT 530.400 124.050 531.450 131.400 ;
        RECT 538.950 130.950 541.050 133.050 ;
        RECT 551.400 132.900 552.600 133.650 ;
        RECT 550.950 130.800 553.050 132.900 ;
        RECT 560.400 130.050 561.450 137.400 ;
        RECT 568.950 137.100 571.050 139.200 ;
        RECT 574.950 137.100 577.050 139.200 ;
        RECT 592.950 137.100 595.050 139.200 ;
        RECT 599.400 138.600 600.450 181.950 ;
        RECT 602.400 175.050 603.450 196.950 ;
        RECT 623.400 195.450 624.450 215.100 ;
        RECT 629.400 214.350 630.600 215.100 ;
        RECT 628.800 211.950 630.900 214.050 ;
        RECT 634.650 203.700 635.850 222.300 ;
        RECT 638.400 220.050 639.450 223.950 ;
        RECT 637.950 216.000 640.050 220.050 ;
        RECT 638.400 214.350 639.600 216.000 ;
        RECT 637.950 211.950 640.050 214.050 ;
        RECT 644.400 211.050 645.450 253.800 ;
        RECT 647.400 228.450 648.450 262.950 ;
        RECT 650.400 253.050 651.450 328.950 ;
        RECT 653.400 328.050 654.450 331.800 ;
        RECT 652.950 325.950 655.050 328.050 ;
        RECT 665.400 301.050 666.450 365.400 ;
        RECT 673.950 364.800 676.050 366.900 ;
        RECT 679.950 364.800 682.050 366.900 ;
        RECT 686.400 365.400 687.600 367.650 ;
        RECT 673.950 343.950 676.050 346.050 ;
        RECT 674.400 339.600 675.450 343.950 ;
        RECT 674.400 337.350 675.600 339.600 ;
        RECT 670.950 334.950 673.050 337.050 ;
        RECT 673.950 334.950 676.050 337.050 ;
        RECT 676.950 334.950 679.050 337.050 ;
        RECT 671.400 332.400 672.600 334.650 ;
        RECT 671.400 328.050 672.450 332.400 ;
        RECT 670.950 325.950 673.050 328.050 ;
        RECT 664.950 298.950 667.050 301.050 ;
        RECT 664.950 293.100 667.050 295.200 ;
        RECT 671.400 295.050 672.450 325.950 ;
        RECT 673.950 298.950 676.050 301.050 ;
        RECT 665.400 292.350 666.600 293.100 ;
        RECT 670.950 292.950 673.050 295.050 ;
        RECT 658.950 289.950 661.050 292.050 ;
        RECT 661.950 289.950 664.050 292.050 ;
        RECT 664.950 289.950 667.050 292.050 ;
        RECT 667.950 289.950 670.050 292.050 ;
        RECT 662.400 288.900 663.600 289.650 ;
        RECT 661.950 286.800 664.050 288.900 ;
        RECT 668.400 287.400 669.600 289.650 ;
        RECT 668.400 280.050 669.450 287.400 ;
        RECT 667.950 277.950 670.050 280.050 ;
        RECT 674.400 268.050 675.450 298.950 ;
        RECT 686.400 298.050 687.450 365.400 ;
        RECT 688.950 343.950 691.050 346.050 ;
        RECT 689.400 322.050 690.450 343.950 ;
        RECT 695.400 343.050 696.450 379.950 ;
        RECT 698.400 367.050 699.450 406.950 ;
        RECT 707.400 388.050 708.450 409.950 ;
        RECT 713.400 394.050 714.450 416.400 ;
        RECT 718.950 416.100 721.050 418.200 ;
        RECT 725.400 417.600 726.450 430.950 ;
        RECT 731.400 429.450 732.450 445.950 ;
        RECT 734.400 433.050 735.450 451.950 ;
        RECT 742.950 449.100 745.050 451.200 ;
        RECT 749.400 450.600 750.450 454.950 ;
        RECT 743.400 448.350 744.600 449.100 ;
        RECT 749.400 448.350 750.600 450.600 ;
        RECT 755.400 448.050 756.450 475.950 ;
        RECT 767.400 457.050 768.450 488.400 ;
        RECT 772.950 487.800 775.050 489.900 ;
        RECT 784.950 487.800 787.050 489.900 ;
        RECT 766.950 454.950 769.050 457.050 ;
        RECT 772.950 454.950 775.050 457.050 ;
        RECT 781.950 454.950 784.050 457.050 ;
        RECT 763.950 450.000 766.050 454.050 ;
        RECT 764.400 448.350 765.600 450.000 ;
        RECT 739.950 445.950 742.050 448.050 ;
        RECT 742.950 445.950 745.050 448.050 ;
        RECT 745.950 445.950 748.050 448.050 ;
        RECT 748.950 445.950 751.050 448.050 ;
        RECT 754.950 445.950 757.050 448.050 ;
        RECT 763.950 445.950 766.050 448.050 ;
        RECT 766.950 445.950 769.050 448.050 ;
        RECT 740.400 443.400 741.600 445.650 ;
        RECT 746.400 444.900 747.600 445.650 ;
        RECT 733.950 430.950 736.050 433.050 ;
        RECT 731.400 428.400 735.450 429.450 ;
        RECT 719.400 415.350 720.600 416.100 ;
        RECT 725.400 415.350 726.600 417.600 ;
        RECT 718.950 412.950 721.050 415.050 ;
        RECT 721.950 412.950 724.050 415.050 ;
        RECT 724.950 412.950 727.050 415.050 ;
        RECT 727.950 412.950 730.050 415.050 ;
        RECT 722.400 411.900 723.600 412.650 ;
        RECT 728.400 411.900 729.600 412.650 ;
        RECT 734.400 412.050 735.450 428.400 ;
        RECT 740.400 417.450 741.450 443.400 ;
        RECT 745.950 442.800 748.050 444.900 ;
        RECT 767.400 444.450 768.600 445.650 ;
        RECT 773.400 444.450 774.450 454.950 ;
        RECT 782.400 450.600 783.450 454.950 ;
        RECT 788.400 450.600 789.450 493.950 ;
        RECT 797.400 493.350 798.600 494.100 ;
        RECT 793.950 490.950 796.050 493.050 ;
        RECT 796.950 490.950 799.050 493.050 ;
        RECT 799.950 490.950 802.050 493.050 ;
        RECT 794.400 489.900 795.600 490.650 ;
        RECT 793.950 487.800 796.050 489.900 ;
        RECT 800.400 488.400 801.600 490.650 ;
        RECT 800.400 487.050 801.450 488.400 ;
        RECT 796.950 484.950 802.050 487.050 ;
        RECT 806.400 472.050 807.450 515.400 ;
        RECT 815.400 508.050 816.450 521.400 ;
        RECT 820.950 517.950 823.050 522.000 ;
        RECT 830.400 511.050 831.450 527.100 ;
        RECT 833.400 520.050 834.450 541.950 ;
        RECT 836.400 529.050 837.450 557.400 ;
        RECT 838.950 553.950 841.050 556.050 ;
        RECT 839.400 544.050 840.450 553.950 ;
        RECT 838.950 541.950 841.050 544.050 ;
        RECT 842.400 535.050 843.450 565.950 ;
        RECT 847.950 565.800 850.050 567.900 ;
        RECT 853.950 565.800 856.050 567.900 ;
        RECT 854.400 553.050 855.450 565.800 ;
        RECT 853.950 550.950 856.050 553.050 ;
        RECT 841.950 532.950 844.050 535.050 ;
        RECT 856.950 532.950 859.050 535.050 ;
        RECT 835.950 526.950 838.050 529.050 ;
        RECT 841.950 527.100 844.050 529.200 ;
        RECT 847.950 528.000 850.050 532.050 ;
        RECT 853.950 529.950 856.050 532.050 ;
        RECT 842.400 526.350 843.600 527.100 ;
        RECT 848.400 526.350 849.600 528.000 ;
        RECT 838.950 523.950 841.050 526.050 ;
        RECT 841.950 523.950 844.050 526.050 ;
        RECT 844.950 523.950 847.050 526.050 ;
        RECT 847.950 523.950 850.050 526.050 ;
        RECT 835.950 520.950 838.050 523.050 ;
        RECT 839.400 522.900 840.600 523.650 ;
        RECT 832.950 517.950 835.050 520.050 ;
        RECT 829.950 508.950 832.050 511.050 ;
        RECT 814.950 505.950 817.050 508.050 ;
        RECT 836.400 507.450 837.450 520.950 ;
        RECT 838.950 520.800 841.050 522.900 ;
        RECT 845.400 521.400 846.600 523.650 ;
        RECT 845.400 519.450 846.450 521.400 ;
        RECT 849.000 519.450 853.050 520.050 ;
        RECT 845.400 518.400 853.050 519.450 ;
        RECT 833.400 506.400 837.450 507.450 ;
        RECT 848.400 517.950 853.050 518.400 ;
        RECT 808.950 494.100 811.050 496.200 ;
        RECT 817.950 494.100 820.050 496.200 ;
        RECT 823.950 494.100 826.050 496.200 ;
        RECT 809.400 487.050 810.450 494.100 ;
        RECT 818.400 493.350 819.600 494.100 ;
        RECT 824.400 493.350 825.600 494.100 ;
        RECT 814.950 490.950 817.050 493.050 ;
        RECT 817.950 490.950 820.050 493.050 ;
        RECT 820.950 490.950 823.050 493.050 ;
        RECT 823.950 490.950 826.050 493.050 ;
        RECT 826.950 490.950 829.050 493.050 ;
        RECT 815.400 489.900 816.600 490.650 ;
        RECT 814.950 487.800 817.050 489.900 ;
        RECT 821.400 488.400 822.600 490.650 ;
        RECT 827.400 488.400 828.600 490.650 ;
        RECT 808.950 484.950 811.050 487.050 ;
        RECT 799.950 469.950 802.050 472.050 ;
        RECT 805.950 469.950 808.050 472.050 ;
        RECT 782.400 448.350 783.600 450.600 ;
        RECT 788.400 448.350 789.600 450.600 ;
        RECT 781.950 445.950 784.050 448.050 ;
        RECT 784.950 445.950 787.050 448.050 ;
        RECT 787.950 445.950 790.050 448.050 ;
        RECT 790.950 445.950 793.050 448.050 ;
        RECT 767.400 443.400 774.450 444.450 ;
        RECT 785.400 443.400 786.600 445.650 ;
        RECT 791.400 444.900 792.600 445.650 ;
        RECT 785.400 441.450 786.450 443.400 ;
        RECT 790.950 442.800 793.050 444.900 ;
        RECT 782.400 440.400 786.450 441.450 ;
        RECT 775.950 430.950 778.050 433.050 ;
        RECT 742.950 421.950 745.050 424.050 ;
        RECT 737.400 416.400 741.450 417.450 ;
        RECT 743.400 417.600 744.450 421.950 ;
        RECT 721.950 409.800 724.050 411.900 ;
        RECT 727.950 409.800 730.050 411.900 ;
        RECT 733.950 409.950 736.050 412.050 ;
        RECT 721.950 403.950 724.050 406.050 ;
        RECT 712.950 391.950 715.050 394.050 ;
        RECT 706.950 385.950 709.050 388.050 ;
        RECT 706.950 379.950 709.050 382.050 ;
        RECT 707.400 372.600 708.450 379.950 ;
        RECT 707.400 370.350 708.600 372.600 ;
        RECT 712.950 371.100 715.050 373.200 ;
        RECT 713.400 370.350 714.600 371.100 ;
        RECT 703.950 367.950 706.050 370.050 ;
        RECT 706.950 367.950 709.050 370.050 ;
        RECT 709.950 367.950 712.050 370.050 ;
        RECT 712.950 367.950 715.050 370.050 ;
        RECT 697.950 364.950 700.050 367.050 ;
        RECT 704.400 366.900 705.600 367.650 ;
        RECT 703.950 364.800 706.050 366.900 ;
        RECT 710.400 365.400 711.600 367.650 ;
        RECT 710.400 349.050 711.450 365.400 ;
        RECT 715.950 364.950 718.050 367.050 ;
        RECT 716.400 355.050 717.450 364.950 ;
        RECT 722.400 361.050 723.450 403.950 ;
        RECT 728.400 387.450 729.450 409.800 ;
        RECT 725.400 386.400 729.450 387.450 ;
        RECT 725.400 373.050 726.450 386.400 ;
        RECT 737.400 382.050 738.450 416.400 ;
        RECT 743.400 415.350 744.600 417.600 ;
        RECT 748.950 416.100 751.050 418.200 ;
        RECT 760.950 416.100 763.050 418.200 ;
        RECT 769.950 416.100 772.050 418.200 ;
        RECT 776.400 417.600 777.450 430.950 ;
        RECT 749.400 415.350 750.600 416.100 ;
        RECT 742.950 412.950 745.050 415.050 ;
        RECT 745.950 412.950 748.050 415.050 ;
        RECT 748.950 412.950 751.050 415.050 ;
        RECT 751.950 412.950 754.050 415.050 ;
        RECT 746.400 410.400 747.600 412.650 ;
        RECT 752.400 411.900 753.600 412.650 ;
        RECT 746.400 409.050 747.450 410.400 ;
        RECT 751.950 409.800 754.050 411.900 ;
        RECT 745.950 403.950 748.050 409.050 ;
        RECT 752.400 391.050 753.450 409.800 ;
        RECT 761.400 394.050 762.450 416.100 ;
        RECT 770.400 415.350 771.600 416.100 ;
        RECT 776.400 415.350 777.600 417.600 ;
        RECT 766.950 412.950 769.050 415.050 ;
        RECT 769.950 412.950 772.050 415.050 ;
        RECT 772.950 412.950 775.050 415.050 ;
        RECT 775.950 412.950 778.050 415.050 ;
        RECT 767.400 411.000 768.600 412.650 ;
        RECT 773.400 411.900 774.600 412.650 ;
        RECT 766.950 406.950 769.050 411.000 ;
        RECT 772.950 409.800 775.050 411.900 ;
        RECT 767.400 400.050 768.450 406.950 ;
        RECT 766.950 397.950 769.050 400.050 ;
        RECT 760.950 391.950 763.050 394.050 ;
        RECT 766.950 391.950 769.050 394.050 ;
        RECT 745.950 388.950 748.050 391.050 ;
        RECT 751.950 388.950 754.050 391.050 ;
        RECT 730.950 379.950 733.050 382.050 ;
        RECT 736.950 379.950 739.050 382.050 ;
        RECT 742.950 379.950 745.050 382.050 ;
        RECT 724.950 370.950 727.050 373.050 ;
        RECT 731.400 372.600 732.450 379.950 ;
        RECT 731.400 370.350 732.600 372.600 ;
        RECT 736.950 371.100 739.050 373.200 ;
        RECT 737.400 370.350 738.600 371.100 ;
        RECT 727.950 367.950 730.050 370.050 ;
        RECT 730.950 367.950 733.050 370.050 ;
        RECT 733.950 367.950 736.050 370.050 ;
        RECT 736.950 367.950 739.050 370.050 ;
        RECT 728.400 366.900 729.600 367.650 ;
        RECT 727.950 364.800 730.050 366.900 ;
        RECT 734.400 365.400 735.600 367.650 ;
        RECT 721.950 358.950 724.050 361.050 ;
        RECT 715.950 352.950 718.050 355.050 ;
        RECT 721.950 352.950 724.050 355.050 ;
        RECT 697.950 346.950 700.050 349.050 ;
        RECT 709.950 346.950 712.050 349.050 ;
        RECT 694.950 340.950 697.050 343.050 ;
        RECT 698.400 339.600 699.450 346.950 ;
        RECT 698.400 337.350 699.600 339.600 ;
        RECT 703.950 338.100 706.050 340.200 ;
        RECT 722.400 339.600 723.450 352.950 ;
        RECT 734.400 349.050 735.450 365.400 ;
        RECT 739.950 364.950 742.050 367.050 ;
        RECT 740.400 355.050 741.450 364.950 ;
        RECT 739.950 352.950 742.050 355.050 ;
        RECT 733.950 346.950 736.050 349.050 ;
        RECT 739.950 346.950 742.050 349.050 ;
        RECT 704.400 337.350 705.600 338.100 ;
        RECT 722.400 337.350 723.600 339.600 ;
        RECT 727.950 337.950 730.050 340.050 ;
        RECT 740.400 339.600 741.450 346.950 ;
        RECT 743.400 343.050 744.450 379.950 ;
        RECT 746.400 367.050 747.450 388.950 ;
        RECT 754.950 379.950 757.050 382.050 ;
        RECT 755.400 372.600 756.450 379.950 ;
        RECT 755.400 370.350 756.600 372.600 ;
        RECT 760.950 371.100 763.050 373.200 ;
        RECT 761.400 370.350 762.600 371.100 ;
        RECT 751.950 367.950 754.050 370.050 ;
        RECT 754.950 367.950 757.050 370.050 ;
        RECT 757.950 367.950 760.050 370.050 ;
        RECT 760.950 367.950 763.050 370.050 ;
        RECT 745.950 364.950 748.050 367.050 ;
        RECT 752.400 366.900 753.600 367.650 ;
        RECT 758.400 366.900 759.600 367.650 ;
        RECT 751.950 364.800 754.050 366.900 ;
        RECT 757.950 364.800 760.050 366.900 ;
        RECT 742.950 340.950 745.050 343.050 ;
        RECT 754.950 340.950 757.050 343.050 ;
        RECT 694.950 334.950 697.050 337.050 ;
        RECT 697.950 334.950 700.050 337.050 ;
        RECT 700.950 334.950 703.050 337.050 ;
        RECT 703.950 334.950 706.050 337.050 ;
        RECT 718.950 334.950 721.050 337.050 ;
        RECT 721.950 334.950 724.050 337.050 ;
        RECT 695.400 333.900 696.600 334.650 ;
        RECT 701.400 333.900 702.600 334.650 ;
        RECT 719.400 333.900 720.600 334.650 ;
        RECT 694.950 331.800 697.050 333.900 ;
        RECT 700.950 331.800 703.050 333.900 ;
        RECT 718.950 331.800 721.050 333.900 ;
        RECT 688.950 319.950 691.050 322.050 ;
        RECT 676.950 295.950 679.050 298.050 ;
        RECT 685.950 295.950 688.050 298.050 ;
        RECT 677.400 268.050 678.450 295.950 ;
        RECT 689.400 294.600 690.450 319.950 ;
        RECT 706.950 304.950 709.050 307.050 ;
        RECT 689.400 292.350 690.600 294.600 ;
        RECT 697.950 293.100 700.050 295.200 ;
        RECT 707.400 294.600 708.450 304.950 ;
        RECT 682.950 289.950 685.050 292.050 ;
        RECT 685.950 289.950 688.050 292.050 ;
        RECT 688.950 289.950 691.050 292.050 ;
        RECT 691.950 289.950 694.050 292.050 ;
        RECT 692.400 288.900 693.600 289.650 ;
        RECT 698.400 289.050 699.450 293.100 ;
        RECT 707.400 292.350 708.600 294.600 ;
        RECT 712.950 293.100 715.050 295.200 ;
        RECT 724.950 293.100 727.050 295.200 ;
        RECT 713.400 292.350 714.600 293.100 ;
        RECT 706.950 289.950 709.050 292.050 ;
        RECT 709.950 289.950 712.050 292.050 ;
        RECT 712.950 289.950 715.050 292.050 ;
        RECT 715.950 289.950 718.050 292.050 ;
        RECT 691.950 286.800 694.050 288.900 ;
        RECT 697.950 286.950 700.050 289.050 ;
        RECT 710.400 287.400 711.600 289.650 ;
        RECT 716.400 287.400 717.600 289.650 ;
        RECT 710.400 280.050 711.450 287.400 ;
        RECT 709.950 277.950 712.050 280.050 ;
        RECT 716.400 277.050 717.450 287.400 ;
        RECT 718.950 277.950 721.050 280.050 ;
        RECT 715.950 274.950 718.050 277.050 ;
        RECT 719.400 273.450 720.450 277.950 ;
        RECT 725.400 276.450 726.450 293.100 ;
        RECT 728.400 280.050 729.450 337.950 ;
        RECT 740.400 337.350 741.600 339.600 ;
        RECT 745.950 338.100 748.050 340.200 ;
        RECT 751.950 338.100 754.050 340.200 ;
        RECT 746.400 337.350 747.600 338.100 ;
        RECT 736.950 334.950 739.050 337.050 ;
        RECT 739.950 334.950 742.050 337.050 ;
        RECT 742.950 334.950 745.050 337.050 ;
        RECT 745.950 334.950 748.050 337.050 ;
        RECT 737.400 333.900 738.600 334.650 ;
        RECT 736.950 331.800 739.050 333.900 ;
        RECT 743.400 332.400 744.600 334.650 ;
        RECT 752.400 333.900 753.450 338.100 ;
        RECT 743.400 330.450 744.450 332.400 ;
        RECT 751.950 331.800 754.050 333.900 ;
        RECT 745.950 330.450 748.050 331.050 ;
        RECT 743.400 329.400 748.050 330.450 ;
        RECT 745.950 328.950 748.050 329.400 ;
        RECT 733.950 293.100 736.050 295.200 ;
        RECT 739.950 293.100 742.050 295.200 ;
        RECT 734.400 292.350 735.600 293.100 ;
        RECT 740.400 292.350 741.600 293.100 ;
        RECT 733.950 289.950 736.050 292.050 ;
        RECT 736.950 289.950 739.050 292.050 ;
        RECT 739.950 289.950 742.050 292.050 ;
        RECT 737.400 287.400 738.600 289.650 ;
        RECT 737.400 280.050 738.450 287.400 ;
        RECT 742.950 286.950 745.050 289.050 ;
        RECT 727.950 277.950 730.050 280.050 ;
        RECT 736.950 277.950 739.050 280.050 ;
        RECT 727.950 276.450 730.050 276.900 ;
        RECT 725.400 275.400 730.050 276.450 ;
        RECT 727.950 274.800 730.050 275.400 ;
        RECT 716.400 272.400 720.450 273.450 ;
        RECT 664.950 265.950 667.050 268.050 ;
        RECT 673.800 265.950 675.900 268.050 ;
        RECT 676.950 265.950 679.050 268.050 ;
        RECT 688.950 265.950 691.050 268.050 ;
        RECT 658.950 260.100 661.050 262.200 ;
        RECT 659.400 259.350 660.600 260.100 ;
        RECT 655.950 256.950 658.050 259.050 ;
        RECT 658.950 256.950 661.050 259.050 ;
        RECT 656.400 254.400 657.600 256.650 ;
        RECT 649.950 250.950 652.050 253.050 ;
        RECT 656.400 250.050 657.450 254.400 ;
        RECT 652.950 248.400 657.450 250.050 ;
        RECT 652.950 247.950 657.000 248.400 ;
        RECT 647.400 227.400 651.450 228.450 ;
        RECT 646.950 223.950 649.050 226.050 ;
        RECT 643.950 208.950 646.050 211.050 ;
        RECT 647.400 205.050 648.450 223.950 ;
        RECT 634.050 201.600 636.150 203.700 ;
        RECT 646.950 202.950 649.050 205.050 ;
        RECT 631.950 196.950 634.050 199.050 ;
        RECT 617.400 194.400 624.450 195.450 ;
        RECT 617.400 189.450 618.450 194.400 ;
        RECT 617.400 187.200 618.600 189.450 ;
        RECT 604.950 181.950 607.050 184.050 ;
        RECT 612.900 183.900 615.000 185.700 ;
        RECT 616.800 184.800 618.900 186.900 ;
        RECT 620.100 186.300 622.200 188.400 ;
        RECT 611.400 182.700 620.100 183.900 ;
        RECT 605.400 177.450 606.450 181.950 ;
        RECT 608.100 178.950 610.200 181.050 ;
        RECT 608.400 177.450 609.600 178.650 ;
        RECT 605.400 176.400 609.600 177.450 ;
        RECT 601.950 172.950 604.050 175.050 ;
        RECT 611.400 173.700 612.300 182.700 ;
        RECT 618.000 181.800 620.100 182.700 ;
        RECT 621.000 180.900 621.900 186.300 ;
        RECT 623.400 183.450 624.600 183.600 ;
        RECT 623.400 182.400 627.450 183.450 ;
        RECT 623.400 181.350 624.600 182.400 ;
        RECT 615.000 179.700 621.900 180.900 ;
        RECT 615.000 177.300 615.900 179.700 ;
        RECT 613.800 175.200 615.900 177.300 ;
        RECT 616.800 175.950 618.900 178.050 ;
        RECT 610.500 171.600 612.600 173.700 ;
        RECT 617.400 173.400 618.600 175.650 ;
        RECT 620.700 172.500 621.900 179.700 ;
        RECT 622.800 178.950 624.900 181.050 ;
        RECT 620.100 170.400 622.200 172.500 ;
        RECT 626.400 169.050 627.450 182.400 ;
        RECT 632.400 177.900 633.450 196.950 ;
        RECT 640.950 187.950 643.050 190.050 ;
        RECT 641.400 183.600 642.450 187.950 ;
        RECT 641.400 181.350 642.600 183.600 ;
        RECT 646.950 182.100 649.050 184.200 ;
        RECT 650.400 183.450 651.450 227.400 ;
        RECT 665.400 220.050 666.450 265.950 ;
        RECT 673.950 260.100 676.050 262.200 ;
        RECT 679.950 260.100 682.050 262.200 ;
        RECT 674.400 259.350 675.600 260.100 ;
        RECT 680.400 259.350 681.600 260.100 ;
        RECT 673.950 256.950 676.050 259.050 ;
        RECT 676.950 256.950 679.050 259.050 ;
        RECT 679.950 256.950 682.050 259.050 ;
        RECT 682.950 256.950 685.050 259.050 ;
        RECT 677.400 254.400 678.600 256.650 ;
        RECT 683.400 255.900 684.600 256.650 ;
        RECT 689.400 255.900 690.450 265.950 ;
        RECT 697.950 260.100 700.050 262.200 ;
        RECT 703.950 260.100 706.050 262.200 ;
        RECT 712.950 260.100 715.050 262.200 ;
        RECT 698.400 259.350 699.600 260.100 ;
        RECT 704.400 259.350 705.600 260.100 ;
        RECT 697.950 256.950 700.050 259.050 ;
        RECT 700.950 256.950 703.050 259.050 ;
        RECT 703.950 256.950 706.050 259.050 ;
        RECT 706.950 256.950 709.050 259.050 ;
        RECT 667.950 229.950 670.050 232.050 ;
        RECT 655.950 216.000 658.050 220.050 ;
        RECT 661.950 216.000 664.050 220.050 ;
        RECT 664.950 217.950 667.050 220.050 ;
        RECT 668.400 217.050 669.450 229.950 ;
        RECT 677.400 229.050 678.450 254.400 ;
        RECT 682.950 253.800 685.050 255.900 ;
        RECT 688.950 253.800 691.050 255.900 ;
        RECT 701.400 254.400 702.600 256.650 ;
        RECT 707.400 255.000 708.600 256.650 ;
        RECT 682.950 250.650 685.050 252.750 ;
        RECT 676.950 226.950 679.050 229.050 ;
        RECT 670.950 220.950 673.050 223.050 ;
        RECT 656.400 214.350 657.600 216.000 ;
        RECT 662.400 214.350 663.600 216.000 ;
        RECT 667.950 214.950 670.050 217.050 ;
        RECT 655.950 211.950 658.050 214.050 ;
        RECT 658.950 211.950 661.050 214.050 ;
        RECT 661.950 211.950 664.050 214.050 ;
        RECT 664.950 211.950 667.050 214.050 ;
        RECT 659.400 210.900 660.600 211.650 ;
        RECT 665.400 210.900 666.600 211.650 ;
        RECT 658.950 208.800 661.050 210.900 ;
        RECT 664.950 208.800 667.050 210.900 ;
        RECT 658.950 202.950 661.050 205.050 ;
        RECT 650.400 182.400 654.450 183.450 ;
        RECT 647.400 181.350 648.600 182.100 ;
        RECT 637.950 178.950 640.050 181.050 ;
        RECT 640.950 178.950 643.050 181.050 ;
        RECT 643.950 178.950 646.050 181.050 ;
        RECT 646.950 178.950 649.050 181.050 ;
        RECT 638.400 177.900 639.600 178.650 ;
        RECT 644.400 177.900 645.600 178.650 ;
        RECT 631.950 175.800 634.050 177.900 ;
        RECT 637.950 175.800 640.050 177.900 ;
        RECT 643.950 175.800 646.050 177.900 ;
        RECT 607.950 166.950 610.050 169.050 ;
        RECT 625.950 166.950 628.050 169.050 ;
        RECT 608.400 163.050 609.450 166.950 ;
        RECT 607.950 160.950 610.050 163.050 ;
        RECT 569.400 136.350 570.600 137.100 ;
        RECT 575.400 136.350 576.600 137.100 ;
        RECT 593.400 136.350 594.600 137.100 ;
        RECT 599.400 136.350 600.600 138.600 ;
        RECT 568.950 133.950 571.050 136.050 ;
        RECT 571.950 133.950 574.050 136.050 ;
        RECT 574.950 133.950 577.050 136.050 ;
        RECT 583.950 133.950 586.050 136.050 ;
        RECT 592.950 133.950 595.050 136.050 ;
        RECT 595.950 133.950 598.050 136.050 ;
        RECT 598.950 133.950 601.050 136.050 ;
        RECT 601.950 133.950 604.050 136.050 ;
        RECT 572.400 131.400 573.600 133.650 ;
        RECT 559.950 127.950 562.050 130.050 ;
        RECT 572.400 127.050 573.450 131.400 ;
        RECT 580.950 127.950 583.050 130.050 ;
        RECT 571.950 124.950 574.050 127.050 ;
        RECT 523.950 121.950 526.050 124.050 ;
        RECT 529.950 121.950 532.050 124.050 ;
        RECT 541.950 121.950 544.050 124.050 ;
        RECT 529.950 112.950 532.050 115.050 ;
        RECT 511.950 106.950 514.050 109.050 ;
        RECT 517.950 106.950 520.050 109.050 ;
        RECT 520.950 106.950 523.050 109.050 ;
        RECT 505.950 104.100 508.050 106.200 ;
        RECT 512.400 105.450 513.600 105.600 ;
        RECT 512.400 104.400 519.450 105.450 ;
        RECT 506.400 103.350 507.600 104.100 ;
        RECT 512.400 103.350 513.600 104.400 ;
        RECT 502.950 100.950 505.050 103.050 ;
        RECT 505.950 100.950 508.050 103.050 ;
        RECT 508.950 100.950 511.050 103.050 ;
        RECT 511.950 100.950 514.050 103.050 ;
        RECT 482.400 96.450 483.450 98.400 ;
        RECT 484.950 96.450 487.050 97.050 ;
        RECT 482.400 95.400 487.050 96.450 ;
        RECT 484.950 94.950 487.050 95.400 ;
        RECT 472.950 76.950 475.050 79.050 ;
        RECT 478.950 70.950 481.050 73.050 ;
        RECT 466.950 67.950 469.050 70.050 ;
        RECT 449.400 60.450 450.600 60.600 ;
        RECT 446.400 59.400 450.600 60.450 ;
        RECT 449.400 58.350 450.600 59.400 ;
        RECT 455.400 58.350 456.600 60.600 ;
        RECT 466.950 59.100 469.050 61.200 ;
        RECT 472.950 59.100 475.050 61.200 ;
        RECT 479.400 60.600 480.450 70.950 ;
        RECT 448.950 55.950 451.050 58.050 ;
        RECT 451.950 55.950 454.050 58.050 ;
        RECT 454.950 55.950 457.050 58.050 ;
        RECT 452.400 54.900 453.600 55.650 ;
        RECT 467.400 55.050 468.450 59.100 ;
        RECT 473.400 58.350 474.600 59.100 ;
        RECT 479.400 58.350 480.600 60.600 ;
        RECT 472.950 55.950 475.050 58.050 ;
        RECT 475.950 55.950 478.050 58.050 ;
        RECT 478.950 55.950 481.050 58.050 ;
        RECT 428.400 49.050 429.450 53.400 ;
        RECT 433.950 52.800 436.050 54.900 ;
        RECT 439.950 52.800 442.050 54.900 ;
        RECT 451.950 52.800 454.050 54.900 ;
        RECT 466.950 52.950 469.050 55.050 ;
        RECT 476.400 54.900 477.600 55.650 ;
        RECT 485.400 55.050 486.450 94.950 ;
        RECT 488.400 94.050 489.450 98.400 ;
        RECT 496.950 97.800 499.050 99.900 ;
        RECT 503.400 99.000 504.600 100.650 ;
        RECT 509.400 99.900 510.600 100.650 ;
        RECT 497.400 94.050 498.450 97.800 ;
        RECT 502.950 94.950 505.050 99.000 ;
        RECT 508.950 97.800 511.050 99.900 ;
        RECT 518.400 97.050 519.450 104.400 ;
        RECT 517.950 94.950 520.050 97.050 ;
        RECT 487.950 91.950 490.050 94.050 ;
        RECT 496.950 91.950 499.050 94.050 ;
        RECT 505.950 82.950 508.050 85.050 ;
        RECT 499.950 73.950 502.050 76.050 ;
        RECT 500.400 70.050 501.450 73.950 ;
        RECT 499.950 67.950 502.050 70.050 ;
        RECT 493.950 59.100 496.050 61.200 ;
        RECT 500.400 60.600 501.450 67.950 ;
        RECT 494.400 58.350 495.600 59.100 ;
        RECT 500.400 58.350 501.600 60.600 ;
        RECT 493.950 55.950 496.050 58.050 ;
        RECT 496.950 55.950 499.050 58.050 ;
        RECT 499.950 55.950 502.050 58.050 ;
        RECT 475.950 52.800 478.050 54.900 ;
        RECT 484.950 52.950 487.050 55.050 ;
        RECT 497.400 54.900 498.600 55.650 ;
        RECT 496.950 52.800 499.050 54.900 ;
        RECT 427.950 46.950 430.050 49.050 ;
        RECT 506.400 40.050 507.450 82.950 ;
        RECT 517.950 76.950 520.050 79.050 ;
        RECT 514.950 67.950 517.050 70.050 ;
        RECT 508.950 64.950 511.050 67.050 ;
        RECT 505.950 37.950 508.050 40.050 ;
        RECT 415.950 34.950 418.050 37.050 ;
        RECT 416.400 19.050 417.450 34.950 ;
        RECT 451.950 31.950 454.050 34.050 ;
        RECT 430.950 27.000 433.050 31.050 ;
        RECT 442.950 28.950 445.050 31.050 ;
        RECT 431.400 25.350 432.600 27.000 ;
        RECT 425.100 22.950 427.200 25.050 ;
        RECT 430.500 22.950 432.600 25.050 ;
        RECT 433.800 22.950 435.900 25.050 ;
        RECT 425.400 21.900 426.600 22.650 ;
        RECT 424.950 19.800 427.050 21.900 ;
        RECT 434.400 21.000 435.600 22.650 ;
        RECT 443.400 21.900 444.450 28.950 ;
        RECT 452.400 27.600 453.450 31.950 ;
        RECT 452.400 25.350 453.600 27.600 ;
        RECT 472.950 26.100 475.050 28.200 ;
        RECT 473.400 25.350 474.600 26.100 ;
        RECT 484.950 25.950 487.050 28.050 ;
        RECT 493.950 27.000 496.050 31.050 ;
        RECT 505.950 28.950 508.050 31.050 ;
        RECT 448.950 22.950 451.050 25.050 ;
        RECT 451.950 22.950 454.050 25.050 ;
        RECT 454.950 22.950 457.050 25.050 ;
        RECT 469.950 22.950 472.050 25.050 ;
        RECT 472.950 22.950 475.050 25.050 ;
        RECT 475.950 22.950 478.050 25.050 ;
        RECT 449.400 21.900 450.600 22.650 ;
        RECT 455.400 21.900 456.600 22.650 ;
        RECT 412.950 16.950 415.050 19.050 ;
        RECT 415.950 16.950 418.050 19.050 ;
        RECT 433.950 16.950 436.050 21.000 ;
        RECT 442.950 19.800 445.050 21.900 ;
        RECT 448.950 19.800 451.050 21.900 ;
        RECT 454.950 16.950 457.050 21.900 ;
        RECT 470.400 20.400 471.600 22.650 ;
        RECT 485.400 21.900 486.450 25.950 ;
        RECT 494.400 25.350 495.600 27.000 ;
        RECT 490.950 22.950 493.050 25.050 ;
        RECT 493.950 22.950 496.050 25.050 ;
        RECT 496.950 22.950 499.050 25.050 ;
        RECT 491.400 21.900 492.600 22.650 ;
        RECT 497.400 21.900 498.600 22.650 ;
        RECT 470.400 13.050 471.450 20.400 ;
        RECT 484.950 19.800 487.050 21.900 ;
        RECT 490.950 19.800 493.050 21.900 ;
        RECT 496.950 19.800 499.050 21.900 ;
        RECT 506.400 16.050 507.450 28.950 ;
        RECT 509.400 21.900 510.450 64.950 ;
        RECT 515.400 55.050 516.450 67.950 ;
        RECT 518.400 64.050 519.450 76.950 ;
        RECT 521.400 67.050 522.450 106.950 ;
        RECT 523.950 103.950 526.050 109.050 ;
        RECT 530.400 105.600 531.450 112.950 ;
        RECT 530.400 103.350 531.600 105.600 ;
        RECT 535.950 104.100 538.050 106.200 ;
        RECT 536.400 103.350 537.600 104.100 ;
        RECT 526.950 100.950 529.050 103.050 ;
        RECT 529.950 100.950 532.050 103.050 ;
        RECT 532.950 100.950 535.050 103.050 ;
        RECT 535.950 100.950 538.050 103.050 ;
        RECT 527.400 99.900 528.600 100.650 ;
        RECT 533.400 99.900 534.600 100.650 ;
        RECT 526.950 97.800 529.050 99.900 ;
        RECT 532.950 97.800 535.050 99.900 ;
        RECT 528.000 96.750 532.050 97.050 ;
        RECT 526.950 94.950 532.050 96.750 ;
        RECT 526.950 94.650 529.050 94.950 ;
        RECT 533.400 70.050 534.450 97.800 ;
        RECT 542.400 85.050 543.450 121.950 ;
        RECT 553.950 112.950 556.050 115.050 ;
        RECT 544.950 103.950 547.050 106.050 ;
        RECT 554.400 105.600 555.450 112.950 ;
        RECT 545.400 91.050 546.450 103.950 ;
        RECT 554.400 103.350 555.600 105.600 ;
        RECT 559.950 104.100 562.050 106.200 ;
        RECT 574.950 104.100 577.050 106.200 ;
        RECT 581.400 105.600 582.450 127.950 ;
        RECT 584.400 121.050 585.450 133.950 ;
        RECT 596.400 131.400 597.600 133.650 ;
        RECT 602.400 132.000 603.600 133.650 ;
        RECT 596.400 127.050 597.450 131.400 ;
        RECT 601.950 127.950 604.050 132.000 ;
        RECT 608.400 129.450 609.450 160.950 ;
        RECT 610.950 154.950 613.050 157.050 ;
        RECT 611.400 136.050 612.450 154.950 ;
        RECT 653.400 151.050 654.450 182.400 ;
        RECT 652.950 148.950 655.050 151.050 ;
        RECT 619.500 141.300 621.600 143.400 ;
        RECT 629.100 142.500 631.200 144.600 ;
        RECT 646.950 142.950 649.050 145.050 ;
        RECT 617.400 138.450 618.600 138.600 ;
        RECT 614.400 137.400 618.600 138.450 ;
        RECT 610.950 133.950 613.050 136.050 ;
        RECT 610.950 129.450 613.050 130.050 ;
        RECT 608.400 128.400 613.050 129.450 ;
        RECT 610.950 127.950 613.050 128.400 ;
        RECT 595.950 124.950 598.050 127.050 ;
        RECT 583.950 118.950 586.050 121.050 ;
        RECT 598.950 118.950 601.050 121.050 ;
        RECT 560.400 103.350 561.600 104.100 ;
        RECT 575.400 103.350 576.600 104.100 ;
        RECT 581.400 103.350 582.600 105.600 ;
        RECT 589.950 104.100 592.050 106.200 ;
        RECT 599.400 105.600 600.450 118.950 ;
        RECT 550.950 100.950 553.050 103.050 ;
        RECT 553.950 100.950 556.050 103.050 ;
        RECT 556.950 100.950 559.050 103.050 ;
        RECT 559.950 100.950 562.050 103.050 ;
        RECT 574.950 100.950 577.050 103.050 ;
        RECT 577.950 100.950 580.050 103.050 ;
        RECT 580.950 100.950 583.050 103.050 ;
        RECT 583.950 100.950 586.050 103.050 ;
        RECT 551.400 99.900 552.600 100.650 ;
        RECT 557.400 99.900 558.600 100.650 ;
        RECT 550.950 97.800 553.050 99.900 ;
        RECT 556.950 97.800 559.050 99.900 ;
        RECT 578.400 99.000 579.600 100.650 ;
        RECT 584.400 99.900 585.600 100.650 ;
        RECT 553.950 96.450 556.050 97.050 ;
        RECT 559.950 96.450 562.050 97.050 ;
        RECT 553.950 95.400 562.050 96.450 ;
        RECT 553.950 94.950 556.050 95.400 ;
        RECT 559.950 94.950 562.050 95.400 ;
        RECT 577.950 94.950 580.050 99.000 ;
        RECT 583.950 97.800 586.050 99.900 ;
        RECT 590.400 94.050 591.450 104.100 ;
        RECT 599.400 103.350 600.600 105.600 ;
        RECT 604.950 104.100 607.050 106.200 ;
        RECT 611.400 106.050 612.450 127.950 ;
        RECT 614.400 127.050 615.450 137.400 ;
        RECT 617.400 136.350 618.600 137.400 ;
        RECT 617.100 133.950 619.200 136.050 ;
        RECT 620.400 132.300 621.300 141.300 ;
        RECT 622.800 137.700 624.900 139.800 ;
        RECT 626.400 139.350 627.600 141.600 ;
        RECT 624.000 135.300 624.900 137.700 ;
        RECT 625.800 136.950 627.900 139.050 ;
        RECT 629.700 135.300 630.900 142.500 ;
        RECT 647.400 138.600 648.450 142.950 ;
        RECT 647.400 136.350 648.600 138.600 ;
        RECT 652.950 137.100 655.050 139.200 ;
        RECT 653.400 136.350 654.600 137.100 ;
        RECT 624.000 134.100 630.900 135.300 ;
        RECT 627.000 132.300 629.100 133.200 ;
        RECT 620.400 131.100 629.100 132.300 ;
        RECT 621.900 129.300 624.000 131.100 ;
        RECT 625.800 128.100 627.900 130.200 ;
        RECT 630.000 128.700 630.900 134.100 ;
        RECT 631.800 133.950 633.900 136.050 ;
        RECT 646.950 133.950 649.050 136.050 ;
        RECT 649.950 133.950 652.050 136.050 ;
        RECT 652.950 133.950 655.050 136.050 ;
        RECT 632.400 132.900 633.600 133.650 ;
        RECT 631.950 130.800 634.050 132.900 ;
        RECT 650.400 131.400 651.600 133.650 ;
        RECT 613.950 124.950 616.050 127.050 ;
        RECT 626.400 125.550 627.600 127.800 ;
        RECT 629.100 126.600 631.200 128.700 ;
        RECT 626.400 109.200 627.450 125.550 ;
        RECT 646.950 115.950 649.050 118.050 ;
        RECT 625.950 107.100 628.050 109.200 ;
        RECT 631.950 106.950 634.050 109.050 ;
        RECT 634.950 106.950 637.050 109.050 ;
        RECT 605.400 103.350 606.600 104.100 ;
        RECT 610.950 103.950 613.050 106.050 ;
        RECT 625.950 103.950 628.050 106.050 ;
        RECT 626.400 103.350 627.600 103.950 ;
        RECT 598.950 100.950 601.050 103.050 ;
        RECT 601.950 100.950 604.050 103.050 ;
        RECT 604.950 100.950 607.050 103.050 ;
        RECT 607.950 100.950 610.050 103.050 ;
        RECT 622.950 100.950 625.050 103.050 ;
        RECT 625.950 100.950 628.050 103.050 ;
        RECT 602.400 98.400 603.600 100.650 ;
        RECT 608.400 98.400 609.600 100.650 ;
        RECT 623.400 98.400 624.600 100.650 ;
        RECT 589.950 91.950 592.050 94.050 ;
        RECT 602.400 91.050 603.450 98.400 ;
        RECT 608.400 94.050 609.450 98.400 ;
        RECT 607.950 91.950 610.050 94.050 ;
        RECT 544.950 88.950 547.050 91.050 ;
        RECT 601.950 88.950 604.050 91.050 ;
        RECT 623.400 85.050 624.450 98.400 ;
        RECT 541.950 82.950 544.050 85.050 ;
        RECT 622.950 82.950 625.050 85.050 ;
        RECT 538.950 81.450 543.000 82.050 ;
        RECT 538.950 81.000 543.450 81.450 ;
        RECT 538.950 79.950 544.050 81.000 ;
        RECT 541.950 76.950 544.050 79.950 ;
        RECT 583.950 73.950 586.050 76.050 ;
        RECT 535.950 70.950 538.050 73.050 ;
        RECT 532.950 67.950 535.050 70.050 ;
        RECT 520.950 64.950 523.050 67.050 ;
        RECT 517.950 61.950 520.050 64.050 ;
        RECT 527.400 62.400 534.450 63.450 ;
        RECT 518.400 60.600 519.450 61.950 ;
        RECT 527.400 60.600 528.450 62.400 ;
        RECT 518.400 58.350 519.600 60.600 ;
        RECT 527.400 58.350 528.600 60.600 ;
        RECT 529.950 58.950 532.050 61.050 ;
        RECT 518.100 55.950 520.200 58.050 ;
        RECT 523.500 55.950 525.600 58.050 ;
        RECT 526.800 55.950 528.900 58.050 ;
        RECT 514.950 52.950 517.050 55.050 ;
        RECT 524.400 54.900 525.600 55.650 ;
        RECT 530.400 54.900 531.450 58.950 ;
        RECT 523.950 52.800 526.050 54.900 ;
        RECT 529.950 52.800 532.050 54.900 ;
        RECT 517.950 26.100 520.050 28.200 ;
        RECT 533.400 27.450 534.450 62.400 ;
        RECT 530.400 26.400 534.450 27.450 ;
        RECT 536.400 27.600 537.450 70.950 ;
        RECT 541.950 64.950 544.050 67.050 ;
        RECT 580.950 64.950 583.050 67.050 ;
        RECT 542.400 61.200 543.450 64.950 ;
        RECT 541.950 59.100 544.050 61.200 ;
        RECT 547.950 60.000 550.050 64.050 ;
        RECT 562.950 60.000 565.050 64.050 ;
        RECT 542.400 58.350 543.600 59.100 ;
        RECT 548.400 58.350 549.600 60.000 ;
        RECT 563.400 58.350 564.600 60.000 ;
        RECT 568.950 59.100 571.050 61.200 ;
        RECT 577.950 59.100 580.050 61.200 ;
        RECT 569.400 58.350 570.600 59.100 ;
        RECT 541.950 55.950 544.050 58.050 ;
        RECT 544.950 55.950 547.050 58.050 ;
        RECT 547.950 55.950 550.050 58.050 ;
        RECT 562.950 55.950 565.050 58.050 ;
        RECT 565.950 55.950 568.050 58.050 ;
        RECT 568.950 55.950 571.050 58.050 ;
        RECT 571.950 55.950 574.050 58.050 ;
        RECT 545.400 53.400 546.600 55.650 ;
        RECT 566.400 54.000 567.600 55.650 ;
        RECT 572.400 54.900 573.600 55.650 ;
        RECT 545.400 46.050 546.450 53.400 ;
        RECT 565.950 49.950 568.050 54.000 ;
        RECT 571.950 52.800 574.050 54.900 ;
        RECT 544.950 43.950 547.050 46.050 ;
        RECT 556.950 40.950 559.050 43.050 ;
        RECT 541.950 31.950 544.050 34.050 ;
        RECT 542.400 27.600 543.450 31.950 ;
        RECT 518.400 25.350 519.600 26.100 ;
        RECT 512.100 22.950 514.200 25.050 ;
        RECT 517.500 22.950 519.600 25.050 ;
        RECT 520.800 22.950 522.900 25.050 ;
        RECT 508.950 21.450 511.050 21.900 ;
        RECT 512.400 21.450 513.600 22.650 ;
        RECT 508.950 20.400 513.600 21.450 ;
        RECT 521.400 20.400 522.600 22.650 ;
        RECT 530.400 21.900 531.450 26.400 ;
        RECT 536.400 25.350 537.600 27.600 ;
        RECT 542.400 25.350 543.600 27.600 ;
        RECT 535.950 22.950 538.050 25.050 ;
        RECT 538.950 22.950 541.050 25.050 ;
        RECT 541.950 22.950 544.050 25.050 ;
        RECT 544.950 22.950 547.050 25.050 ;
        RECT 508.950 19.800 511.050 20.400 ;
        RECT 505.950 13.950 508.050 16.050 ;
        RECT 311.550 9.600 313.650 11.700 ;
        RECT 388.950 10.950 391.050 13.050 ;
        RECT 469.950 10.950 472.050 13.050 ;
        RECT 521.400 10.050 522.450 20.400 ;
        RECT 529.950 19.800 532.050 21.900 ;
        RECT 539.400 21.000 540.600 22.650 ;
        RECT 545.400 21.900 546.600 22.650 ;
        RECT 557.400 22.050 558.450 40.950 ;
        RECT 578.400 34.050 579.450 59.100 ;
        RECT 581.400 55.050 582.450 64.950 ;
        RECT 580.950 52.950 583.050 55.050 ;
        RECT 577.950 31.950 580.050 34.050 ;
        RECT 565.950 26.100 568.050 28.200 ;
        RECT 571.950 26.100 574.050 28.200 ;
        RECT 584.400 27.600 585.450 73.950 ;
        RECT 613.950 70.950 616.050 73.050 ;
        RECT 589.950 59.100 592.050 61.200 ;
        RECT 614.400 60.600 615.450 70.950 ;
        RECT 632.400 64.050 633.450 106.950 ;
        RECT 635.400 99.900 636.450 106.950 ;
        RECT 640.950 105.000 643.050 109.050 ;
        RECT 647.400 105.600 648.450 115.950 ;
        RECT 650.400 109.050 651.450 131.400 ;
        RECT 655.950 109.950 658.050 112.050 ;
        RECT 649.950 106.950 652.050 109.050 ;
        RECT 641.400 103.350 642.600 105.000 ;
        RECT 647.400 103.350 648.600 105.600 ;
        RECT 640.950 100.950 643.050 103.050 ;
        RECT 643.950 100.950 646.050 103.050 ;
        RECT 646.950 100.950 649.050 103.050 ;
        RECT 649.950 100.950 652.050 103.050 ;
        RECT 634.950 97.800 637.050 99.900 ;
        RECT 644.400 99.000 645.600 100.650 ;
        RECT 650.400 99.000 651.600 100.650 ;
        RECT 643.950 94.950 646.050 99.000 ;
        RECT 649.950 94.950 652.050 99.000 ;
        RECT 656.400 97.050 657.450 109.950 ;
        RECT 655.950 94.950 658.050 97.050 ;
        RECT 659.400 76.050 660.450 202.950 ;
        RECT 671.400 190.050 672.450 220.950 ;
        RECT 683.400 217.200 684.450 250.650 ;
        RECT 694.950 241.950 697.050 244.050 ;
        RECT 688.950 220.950 691.050 223.050 ;
        RECT 673.950 214.950 676.050 217.050 ;
        RECT 682.950 215.100 685.050 217.200 ;
        RECT 689.400 216.600 690.450 220.950 ;
        RECT 674.400 208.050 675.450 214.950 ;
        RECT 683.400 214.350 684.600 215.100 ;
        RECT 689.400 214.350 690.600 216.600 ;
        RECT 679.950 211.950 682.050 214.050 ;
        RECT 682.950 211.950 685.050 214.050 ;
        RECT 685.950 211.950 688.050 214.050 ;
        RECT 688.950 211.950 691.050 214.050 ;
        RECT 680.400 211.050 681.600 211.650 ;
        RECT 676.950 209.400 681.600 211.050 ;
        RECT 686.400 209.400 687.600 211.650 ;
        RECT 676.950 208.950 681.000 209.400 ;
        RECT 673.950 205.950 676.050 208.050 ;
        RECT 674.400 199.050 675.450 205.950 ;
        RECT 673.950 196.950 676.050 199.050 ;
        RECT 670.950 187.950 673.050 190.050 ;
        RECT 682.950 187.950 685.050 190.050 ;
        RECT 664.950 181.950 667.050 184.050 ;
        RECT 673.950 183.000 676.050 187.050 ;
        RECT 683.400 183.600 684.450 187.950 ;
        RECT 686.400 187.050 687.450 209.400 ;
        RECT 691.950 208.950 694.050 211.050 ;
        RECT 692.400 190.050 693.450 208.950 ;
        RECT 691.950 187.950 694.050 190.050 ;
        RECT 695.400 187.050 696.450 241.950 ;
        RECT 701.400 223.050 702.450 254.400 ;
        RECT 706.950 250.950 709.050 255.000 ;
        RECT 700.950 220.950 703.050 223.050 ;
        RECT 697.950 214.950 700.050 217.050 ;
        RECT 706.950 215.100 709.050 217.200 ;
        RECT 698.400 190.050 699.450 214.950 ;
        RECT 707.400 214.350 708.600 215.100 ;
        RECT 703.950 211.950 706.050 214.050 ;
        RECT 706.950 211.950 709.050 214.050 ;
        RECT 704.400 210.000 705.600 211.650 ;
        RECT 703.950 205.950 706.050 210.000 ;
        RECT 709.950 202.950 712.050 205.050 ;
        RECT 710.400 190.050 711.450 202.950 ;
        RECT 697.950 187.950 700.050 190.050 ;
        RECT 709.950 187.950 712.050 190.050 ;
        RECT 685.950 186.450 688.050 187.050 ;
        RECT 685.950 185.400 690.450 186.450 ;
        RECT 685.950 184.950 688.050 185.400 ;
        RECT 661.950 137.100 664.050 139.200 ;
        RECT 665.400 138.450 666.450 181.950 ;
        RECT 674.400 181.350 675.600 183.000 ;
        RECT 683.400 181.350 684.600 183.600 ;
        RECT 668.400 178.950 670.500 181.050 ;
        RECT 673.950 178.950 676.050 181.050 ;
        RECT 676.950 178.950 679.050 181.050 ;
        RECT 683.100 178.950 685.200 181.050 ;
        RECT 668.400 177.900 669.600 178.650 ;
        RECT 667.950 175.800 670.050 177.900 ;
        RECT 677.400 176.400 678.600 178.650 ;
        RECT 677.400 160.050 678.450 176.400 ;
        RECT 689.400 175.050 690.450 185.400 ;
        RECT 694.950 184.950 697.050 187.050 ;
        RECT 688.950 172.950 691.050 175.050 ;
        RECT 695.400 172.050 696.450 184.950 ;
        RECT 703.950 182.100 706.050 184.200 ;
        RECT 710.400 183.600 711.450 187.950 ;
        RECT 713.400 187.050 714.450 260.100 ;
        RECT 716.400 244.050 717.450 272.400 ;
        RECT 718.950 268.950 721.050 271.050 ;
        RECT 719.400 255.450 720.450 268.950 ;
        RECT 728.400 261.600 729.450 274.800 ;
        RECT 743.400 271.050 744.450 286.950 ;
        RECT 742.950 268.950 745.050 271.050 ;
        RECT 746.400 267.450 747.450 328.950 ;
        RECT 752.400 295.050 753.450 331.800 ;
        RECT 755.400 331.050 756.450 340.950 ;
        RECT 760.950 339.000 763.050 343.050 ;
        RECT 767.400 339.600 768.450 391.950 ;
        RECT 782.400 373.200 783.450 440.400 ;
        RECT 793.950 416.100 796.050 418.200 ;
        RECT 794.400 415.350 795.600 416.100 ;
        RECT 790.950 412.950 793.050 415.050 ;
        RECT 793.950 412.950 796.050 415.050 ;
        RECT 791.400 411.900 792.600 412.650 ;
        RECT 790.950 409.800 793.050 411.900 ;
        RECT 796.950 397.950 799.050 400.050 ;
        RECT 769.950 371.100 772.050 373.200 ;
        RECT 775.950 371.100 778.050 373.200 ;
        RECT 781.950 371.100 784.050 373.200 ;
        RECT 793.950 371.100 796.050 373.200 ;
        RECT 770.400 364.050 771.450 371.100 ;
        RECT 776.400 370.350 777.600 371.100 ;
        RECT 782.400 370.350 783.600 371.100 ;
        RECT 775.950 367.950 778.050 370.050 ;
        RECT 778.950 367.950 781.050 370.050 ;
        RECT 781.950 367.950 784.050 370.050 ;
        RECT 784.950 367.950 787.050 370.050 ;
        RECT 779.400 366.900 780.600 367.650 ;
        RECT 785.400 366.900 786.600 367.650 ;
        RECT 794.400 367.050 795.450 371.100 ;
        RECT 772.950 364.800 775.050 366.900 ;
        RECT 778.950 364.800 781.050 366.900 ;
        RECT 784.950 364.800 787.050 366.900 ;
        RECT 793.950 364.950 796.050 367.050 ;
        RECT 769.950 361.950 772.050 364.050 ;
        RECT 773.400 340.050 774.450 364.800 ;
        RECT 797.400 364.050 798.450 397.950 ;
        RECT 800.400 397.050 801.450 469.950 ;
        RECT 821.400 466.050 822.450 488.400 ;
        RECT 827.400 481.050 828.450 488.400 ;
        RECT 829.950 487.950 832.050 490.050 ;
        RECT 826.950 478.950 829.050 481.050 ;
        RECT 823.950 466.950 826.050 469.050 ;
        RECT 820.950 463.950 823.050 466.050 ;
        RECT 802.950 460.950 805.050 463.050 ;
        RECT 803.400 439.050 804.450 460.950 ;
        RECT 811.950 450.000 814.050 454.050 ;
        RECT 812.400 448.350 813.600 450.000 ;
        RECT 817.950 449.100 820.050 451.200 ;
        RECT 818.400 448.350 819.600 449.100 ;
        RECT 808.950 445.950 811.050 448.050 ;
        RECT 811.950 445.950 814.050 448.050 ;
        RECT 814.950 445.950 817.050 448.050 ;
        RECT 817.950 445.950 820.050 448.050 ;
        RECT 809.400 444.900 810.600 445.650 ;
        RECT 808.950 442.800 811.050 444.900 ;
        RECT 815.400 443.400 816.600 445.650 ;
        RECT 815.400 439.050 816.450 443.400 ;
        RECT 802.950 436.950 805.050 439.050 ;
        RECT 808.950 436.950 811.050 439.050 ;
        RECT 814.950 436.950 817.050 439.050 ;
        RECT 802.950 418.950 805.050 421.050 ;
        RECT 803.400 412.050 804.450 418.950 ;
        RECT 809.400 417.600 810.450 436.950 ;
        RECT 820.950 424.950 823.050 427.050 ;
        RECT 809.400 415.350 810.600 417.600 ;
        RECT 814.950 417.000 817.050 421.050 ;
        RECT 821.400 418.200 822.450 424.950 ;
        RECT 815.400 415.350 816.600 417.000 ;
        RECT 820.950 416.100 823.050 418.200 ;
        RECT 808.950 412.950 811.050 415.050 ;
        RECT 811.950 412.950 814.050 415.050 ;
        RECT 814.950 412.950 817.050 415.050 ;
        RECT 817.950 412.950 820.050 415.050 ;
        RECT 802.950 409.950 805.050 412.050 ;
        RECT 812.400 411.000 813.600 412.650 ;
        RECT 818.400 412.050 819.600 412.650 ;
        RECT 803.400 406.050 804.450 409.950 ;
        RECT 811.950 406.950 814.050 411.000 ;
        RECT 818.400 409.950 823.050 412.050 ;
        RECT 802.950 403.950 805.050 406.050 ;
        RECT 818.400 400.050 819.450 409.950 ;
        RECT 817.950 397.950 820.050 400.050 ;
        RECT 799.950 394.950 802.050 397.050 ;
        RECT 805.950 371.100 808.050 373.200 ;
        RECT 811.950 371.100 814.050 373.200 ;
        RECT 817.950 371.100 820.050 373.200 ;
        RECT 824.400 372.450 825.450 466.950 ;
        RECT 830.400 457.050 831.450 487.950 ;
        RECT 833.400 478.050 834.450 506.400 ;
        RECT 848.400 501.450 849.450 517.950 ;
        RECT 854.400 513.450 855.450 529.950 ;
        RECT 851.400 512.400 855.450 513.450 ;
        RECT 851.400 505.050 852.450 512.400 ;
        RECT 850.950 502.950 853.050 505.050 ;
        RECT 848.400 500.400 852.450 501.450 ;
        RECT 835.950 494.100 838.050 496.200 ;
        RECT 844.950 494.100 847.050 496.200 ;
        RECT 851.400 495.600 852.450 500.400 ;
        RECT 857.400 496.200 858.450 532.950 ;
        RECT 860.400 529.050 861.450 571.950 ;
        RECT 863.400 547.050 864.450 571.950 ;
        RECT 872.400 571.350 873.600 572.100 ;
        RECT 878.400 571.350 879.600 572.100 ;
        RECT 868.950 568.950 871.050 571.050 ;
        RECT 871.950 568.950 874.050 571.050 ;
        RECT 874.950 568.950 877.050 571.050 ;
        RECT 877.950 568.950 880.050 571.050 ;
        RECT 865.950 565.950 868.050 568.050 ;
        RECT 869.400 566.400 870.600 568.650 ;
        RECT 875.400 567.000 876.600 568.650 ;
        RECT 866.400 553.050 867.450 565.950 ;
        RECT 869.400 562.050 870.450 566.400 ;
        RECT 874.950 562.950 877.050 567.000 ;
        RECT 868.950 559.950 871.050 562.050 ;
        RECT 865.950 550.950 868.050 553.050 ;
        RECT 874.950 550.950 877.050 553.050 ;
        RECT 862.950 544.950 865.050 547.050 ;
        RECT 859.950 526.950 862.050 529.050 ;
        RECT 862.950 528.000 865.050 532.050 ;
        RECT 868.950 528.000 871.050 532.050 ;
        RECT 875.400 529.050 876.450 550.950 ;
        RECT 880.950 538.950 883.050 541.050 ;
        RECT 877.950 529.950 880.050 532.050 ;
        RECT 863.400 526.350 864.600 528.000 ;
        RECT 869.400 526.350 870.600 528.000 ;
        RECT 874.950 526.950 877.050 529.050 ;
        RECT 862.950 523.950 865.050 526.050 ;
        RECT 865.950 523.950 868.050 526.050 ;
        RECT 868.950 523.950 871.050 526.050 ;
        RECT 871.950 523.950 874.050 526.050 ;
        RECT 859.950 520.950 862.050 523.050 ;
        RECT 866.400 522.000 867.600 523.650 ;
        RECT 872.400 522.900 873.600 523.650 ;
        RECT 878.400 523.050 879.450 529.950 ;
        RECT 832.950 475.950 835.050 478.050 ;
        RECT 829.950 454.950 832.050 457.050 ;
        RECT 830.400 450.450 831.450 454.950 ;
        RECT 836.400 454.050 837.450 494.100 ;
        RECT 845.400 493.350 846.600 494.100 ;
        RECT 851.400 493.350 852.600 495.600 ;
        RECT 856.950 494.100 859.050 496.200 ;
        RECT 841.950 490.950 844.050 493.050 ;
        RECT 844.950 490.950 847.050 493.050 ;
        RECT 847.950 490.950 850.050 493.050 ;
        RECT 850.950 490.950 853.050 493.050 ;
        RECT 842.400 488.400 843.600 490.650 ;
        RECT 848.400 489.000 849.600 490.650 ;
        RECT 842.400 463.050 843.450 488.400 ;
        RECT 847.950 484.950 850.050 489.000 ;
        RECT 841.950 460.950 844.050 463.050 ;
        RECT 847.950 454.950 850.050 457.050 ;
        RECT 827.400 449.400 831.450 450.450 ;
        RECT 827.400 445.050 828.450 449.400 ;
        RECT 835.950 449.100 838.050 454.050 ;
        RECT 841.950 450.000 844.050 454.050 ;
        RECT 836.400 448.350 837.600 449.100 ;
        RECT 842.400 448.350 843.600 450.000 ;
        RECT 832.950 445.950 835.050 448.050 ;
        RECT 835.950 445.950 838.050 448.050 ;
        RECT 838.950 445.950 841.050 448.050 ;
        RECT 841.950 445.950 844.050 448.050 ;
        RECT 826.950 442.950 829.050 445.050 ;
        RECT 833.400 444.900 834.600 445.650 ;
        RECT 832.950 442.800 835.050 444.900 ;
        RECT 839.400 443.400 840.600 445.650 ;
        RECT 839.400 439.050 840.450 443.400 ;
        RECT 826.950 436.950 829.050 439.050 ;
        RECT 838.950 436.950 841.050 439.050 ;
        RECT 827.400 388.050 828.450 436.950 ;
        RECT 841.950 430.950 844.050 433.050 ;
        RECT 835.950 416.100 838.050 418.200 ;
        RECT 842.400 417.600 843.450 430.950 ;
        RECT 848.400 427.050 849.450 454.950 ;
        RECT 857.400 454.050 858.450 494.100 ;
        RECT 860.400 469.050 861.450 520.950 ;
        RECT 865.950 517.950 868.050 522.000 ;
        RECT 871.950 520.800 874.050 522.900 ;
        RECT 874.950 519.450 877.050 523.050 ;
        RECT 877.950 520.950 880.050 523.050 ;
        RECT 872.400 519.000 877.050 519.450 ;
        RECT 872.400 518.400 876.450 519.000 ;
        RECT 865.950 494.100 868.050 496.200 ;
        RECT 872.400 496.050 873.450 518.400 ;
        RECT 874.950 511.950 877.050 514.050 ;
        RECT 866.400 493.350 867.600 494.100 ;
        RECT 871.950 493.950 874.050 496.050 ;
        RECT 865.950 490.950 868.050 493.050 ;
        RECT 868.950 490.950 871.050 493.050 ;
        RECT 869.400 489.000 870.600 490.650 ;
        RECT 868.950 484.950 871.050 489.000 ;
        RECT 871.950 487.950 874.050 490.050 ;
        RECT 872.400 480.450 873.450 487.950 ;
        RECT 869.400 479.400 873.450 480.450 ;
        RECT 859.950 466.950 862.050 469.050 ;
        RECT 869.400 460.050 870.450 479.400 ;
        RECT 871.950 475.950 874.050 478.050 ;
        RECT 868.950 457.950 871.050 460.050 ;
        RECT 850.950 451.950 853.050 454.050 ;
        RECT 856.950 451.950 859.050 454.050 ;
        RECT 865.950 451.950 868.050 457.050 ;
        RECT 851.400 445.050 852.450 451.950 ;
        RECT 859.950 449.100 862.050 451.200 ;
        RECT 866.400 450.600 867.450 451.950 ;
        RECT 860.400 448.350 861.600 449.100 ;
        RECT 866.400 448.350 867.600 450.600 ;
        RECT 856.950 445.950 859.050 448.050 ;
        RECT 859.950 445.950 862.050 448.050 ;
        RECT 862.950 445.950 865.050 448.050 ;
        RECT 865.950 445.950 868.050 448.050 ;
        RECT 850.950 442.950 853.050 445.050 ;
        RECT 857.400 444.900 858.600 445.650 ;
        RECT 856.950 442.800 859.050 444.900 ;
        RECT 863.400 443.400 864.600 445.650 ;
        RECT 863.400 436.050 864.450 443.400 ;
        RECT 865.950 439.950 868.050 442.050 ;
        RECT 862.950 433.950 865.050 436.050 ;
        RECT 859.950 430.950 862.050 433.050 ;
        RECT 860.400 427.050 861.450 430.950 ;
        RECT 847.950 424.950 850.050 427.050 ;
        RECT 859.950 424.950 862.050 427.050 ;
        RECT 836.400 415.350 837.600 416.100 ;
        RECT 842.400 415.350 843.600 417.600 ;
        RECT 832.950 412.950 835.050 415.050 ;
        RECT 835.950 412.950 838.050 415.050 ;
        RECT 838.950 412.950 841.050 415.050 ;
        RECT 841.950 412.950 844.050 415.050 ;
        RECT 833.400 411.450 834.600 412.650 ;
        RECT 830.400 410.400 834.600 411.450 ;
        RECT 839.400 410.400 840.600 412.650 ;
        RECT 848.400 411.450 849.450 424.950 ;
        RECT 866.400 417.600 867.450 439.950 ;
        RECT 866.400 415.350 867.600 417.600 ;
        RECT 856.950 412.950 859.050 415.050 ;
        RECT 859.950 412.950 862.050 415.050 ;
        RECT 862.950 412.950 865.050 415.050 ;
        RECT 865.950 412.950 868.050 415.050 ;
        RECT 845.400 410.400 849.450 411.450 ;
        RECT 857.400 410.400 858.600 412.650 ;
        RECT 863.400 410.400 864.600 412.650 ;
        RECT 830.400 409.050 831.450 410.400 ;
        RECT 829.950 406.950 832.050 409.050 ;
        RECT 826.950 385.950 829.050 388.050 ;
        RECT 826.950 376.950 829.050 379.050 ;
        RECT 821.400 371.400 825.450 372.450 ;
        RECT 827.400 372.600 828.450 376.950 ;
        RECT 830.400 376.050 831.450 406.950 ;
        RECT 839.400 406.050 840.450 410.400 ;
        RECT 838.950 403.950 841.050 406.050 ;
        RECT 841.950 397.950 844.050 400.050 ;
        RECT 838.950 385.950 841.050 388.050 ;
        RECT 829.950 373.950 832.050 376.050 ;
        RECT 806.400 370.350 807.600 371.100 ;
        RECT 812.400 370.350 813.600 371.100 ;
        RECT 802.950 367.950 805.050 370.050 ;
        RECT 805.950 367.950 808.050 370.050 ;
        RECT 808.950 367.950 811.050 370.050 ;
        RECT 811.950 367.950 814.050 370.050 ;
        RECT 803.400 366.000 804.600 367.650 ;
        RECT 778.950 361.650 781.050 363.750 ;
        RECT 796.950 361.950 799.050 364.050 ;
        RECT 802.950 361.950 805.050 366.000 ;
        RECT 809.400 365.400 810.600 367.650 ;
        RECT 761.400 337.350 762.600 339.000 ;
        RECT 767.400 337.350 768.600 339.600 ;
        RECT 772.950 337.950 775.050 340.050 ;
        RECT 775.950 337.950 778.050 340.050 ;
        RECT 760.950 334.950 763.050 337.050 ;
        RECT 763.950 334.950 766.050 337.050 ;
        RECT 766.950 334.950 769.050 337.050 ;
        RECT 769.950 334.950 772.050 337.050 ;
        RECT 764.400 333.900 765.600 334.650 ;
        RECT 770.400 333.900 771.600 334.650 ;
        RECT 776.400 333.900 777.450 337.950 ;
        RECT 763.950 331.800 766.050 333.900 ;
        RECT 769.950 331.800 772.050 333.900 ;
        RECT 775.950 331.800 778.050 333.900 ;
        RECT 754.950 328.950 757.050 331.050 ;
        RECT 779.400 322.050 780.450 361.650 ;
        RECT 787.950 358.950 790.050 361.050 ;
        RECT 793.950 358.950 796.050 361.050 ;
        RECT 788.400 340.200 789.450 358.950 ;
        RECT 794.400 355.050 795.450 358.950 ;
        RECT 793.950 352.950 796.050 355.050 ;
        RECT 787.950 338.100 790.050 340.200 ;
        RECT 794.400 339.600 795.450 352.950 ;
        RECT 809.400 343.050 810.450 365.400 ;
        RECT 818.400 361.050 819.450 371.100 ;
        RECT 817.950 358.950 820.050 361.050 ;
        RECT 811.950 346.950 814.050 349.050 ;
        RECT 802.950 340.950 805.050 343.050 ;
        RECT 808.950 340.950 811.050 343.050 ;
        RECT 788.400 337.350 789.600 338.100 ;
        RECT 794.400 337.350 795.600 339.600 ;
        RECT 784.950 334.950 787.050 337.050 ;
        RECT 787.950 334.950 790.050 337.050 ;
        RECT 790.950 334.950 793.050 337.050 ;
        RECT 793.950 334.950 796.050 337.050 ;
        RECT 785.400 334.050 786.600 334.650 ;
        RECT 781.950 332.400 786.600 334.050 ;
        RECT 791.400 332.400 792.600 334.650 ;
        RECT 781.950 331.950 786.450 332.400 ;
        RECT 772.950 319.950 775.050 322.050 ;
        RECT 778.950 319.950 781.050 322.050 ;
        RECT 769.950 298.950 772.050 301.050 ;
        RECT 751.950 292.950 754.050 295.050 ;
        RECT 757.950 293.100 760.050 295.200 ;
        RECT 763.950 293.100 766.050 295.200 ;
        RECT 758.400 292.350 759.600 293.100 ;
        RECT 764.400 292.350 765.600 293.100 ;
        RECT 748.950 289.950 751.050 292.050 ;
        RECT 754.950 289.950 757.050 292.050 ;
        RECT 757.950 289.950 760.050 292.050 ;
        RECT 760.950 289.950 763.050 292.050 ;
        RECT 763.950 289.950 766.050 292.050 ;
        RECT 749.400 280.050 750.450 289.950 ;
        RECT 755.400 289.050 756.600 289.650 ;
        RECT 751.950 287.400 756.600 289.050 ;
        RECT 761.400 287.400 762.600 289.650 ;
        RECT 770.400 289.050 771.450 298.950 ;
        RECT 751.950 286.950 756.000 287.400 ;
        RECT 761.400 280.050 762.450 287.400 ;
        RECT 769.950 286.950 772.050 289.050 ;
        RECT 748.950 277.950 751.050 280.050 ;
        RECT 760.950 277.950 763.050 280.050 ;
        RECT 749.400 268.050 750.450 277.950 ;
        RECT 773.400 277.050 774.450 319.950 ;
        RECT 778.950 304.950 781.050 307.050 ;
        RECT 779.400 294.600 780.450 304.950 ;
        RECT 785.400 301.050 786.450 331.950 ;
        RECT 791.400 322.050 792.450 332.400 ;
        RECT 790.950 319.950 793.050 322.050 ;
        RECT 793.950 304.950 796.050 307.050 ;
        RECT 784.950 298.950 787.050 301.050 ;
        RECT 779.400 292.350 780.600 294.600 ;
        RECT 784.950 293.100 787.050 295.200 ;
        RECT 785.400 292.350 786.600 293.100 ;
        RECT 778.950 289.950 781.050 292.050 ;
        RECT 781.950 289.950 784.050 292.050 ;
        RECT 784.950 289.950 787.050 292.050 ;
        RECT 787.950 289.950 790.050 292.050 ;
        RECT 782.400 287.400 783.600 289.650 ;
        RECT 788.400 288.900 789.600 289.650 ;
        RECT 751.950 274.950 754.050 277.050 ;
        RECT 772.950 274.950 775.050 277.050 ;
        RECT 743.400 266.400 747.450 267.450 ;
        RECT 728.400 259.350 729.600 261.600 ;
        RECT 722.100 256.950 724.200 259.050 ;
        RECT 727.500 256.950 729.600 259.050 ;
        RECT 730.800 256.950 732.900 259.050 ;
        RECT 722.400 255.900 723.600 256.650 ;
        RECT 721.950 255.450 724.050 255.900 ;
        RECT 719.400 254.400 724.050 255.450 ;
        RECT 721.950 253.800 724.050 254.400 ;
        RECT 731.400 254.400 732.600 256.650 ;
        RECT 731.400 253.050 732.450 254.400 ;
        RECT 731.400 251.400 736.050 253.050 ;
        RECT 732.000 250.950 736.050 251.400 ;
        RECT 743.400 250.050 744.450 266.400 ;
        RECT 748.950 265.950 751.050 268.050 ;
        RECT 752.400 261.600 753.450 274.950 ;
        RECT 782.400 268.050 783.450 287.400 ;
        RECT 787.950 286.800 790.050 288.900 ;
        RECT 794.400 280.050 795.450 304.950 ;
        RECT 803.400 298.050 804.450 340.950 ;
        RECT 812.400 339.600 813.450 346.950 ;
        RECT 812.400 337.350 813.600 339.600 ;
        RECT 808.950 334.950 811.050 337.050 ;
        RECT 811.950 334.950 814.050 337.050 ;
        RECT 814.950 334.950 817.050 337.050 ;
        RECT 796.950 295.950 799.050 298.050 ;
        RECT 802.950 295.950 805.050 298.050 ;
        RECT 793.950 277.950 796.050 280.050 ;
        RECT 787.950 274.950 790.050 277.050 ;
        RECT 781.950 265.950 784.050 268.050 ;
        RECT 783.000 264.450 787.050 265.050 ;
        RECT 782.400 262.950 787.050 264.450 ;
        RECT 782.400 262.200 783.450 262.950 ;
        RECT 752.400 259.350 753.600 261.600 ;
        RECT 757.950 260.100 760.050 262.200 ;
        RECT 781.950 260.100 784.050 262.200 ;
        RECT 788.400 261.600 789.450 274.950 ;
        RECT 758.400 259.350 759.600 260.100 ;
        RECT 782.400 259.350 783.600 260.100 ;
        RECT 788.400 259.350 789.600 261.600 ;
        RECT 748.950 256.950 751.050 259.050 ;
        RECT 751.950 256.950 754.050 259.050 ;
        RECT 754.950 256.950 757.050 259.050 ;
        RECT 757.950 256.950 760.050 259.050 ;
        RECT 760.950 256.950 763.050 259.050 ;
        RECT 778.950 256.950 781.050 259.050 ;
        RECT 781.950 256.950 784.050 259.050 ;
        RECT 784.950 256.950 787.050 259.050 ;
        RECT 787.950 256.950 790.050 259.050 ;
        RECT 749.400 255.900 750.600 256.650 ;
        RECT 748.950 253.800 751.050 255.900 ;
        RECT 755.400 254.400 756.600 256.650 ;
        RECT 761.400 255.900 762.600 256.650 ;
        RECT 779.400 255.900 780.600 256.650 ;
        RECT 751.950 250.950 754.050 253.050 ;
        RECT 742.950 247.950 745.050 250.050 ;
        RECT 752.400 246.450 753.450 250.950 ;
        RECT 755.400 250.050 756.450 254.400 ;
        RECT 760.950 253.800 763.050 255.900 ;
        RECT 778.950 253.800 781.050 255.900 ;
        RECT 785.400 255.000 786.600 256.650 ;
        RECT 757.950 250.950 760.050 253.050 ;
        RECT 754.950 247.950 757.050 250.050 ;
        RECT 758.400 246.450 759.450 250.950 ;
        RECT 752.400 245.400 759.450 246.450 ;
        RECT 715.950 241.950 718.050 244.050 ;
        RECT 724.950 241.950 727.050 244.050 ;
        RECT 715.950 232.950 718.050 235.050 ;
        RECT 712.950 184.950 715.050 187.050 ;
        RECT 716.400 184.050 717.450 232.950 ;
        RECT 718.950 220.950 721.050 223.050 ;
        RECT 719.400 217.050 720.450 220.950 ;
        RECT 718.950 214.950 721.050 217.050 ;
        RECT 725.400 216.600 726.450 241.950 ;
        RECT 779.400 235.050 780.450 253.800 ;
        RECT 784.950 250.950 787.050 255.000 ;
        RECT 751.950 232.950 754.050 235.050 ;
        RECT 778.950 232.950 781.050 235.050 ;
        RECT 742.950 223.950 745.050 226.050 ;
        RECT 725.400 214.350 726.600 216.600 ;
        RECT 730.950 215.100 733.050 217.200 ;
        RECT 739.950 215.100 742.050 217.200 ;
        RECT 731.400 214.350 732.600 215.100 ;
        RECT 724.950 211.950 727.050 214.050 ;
        RECT 727.950 211.950 730.050 214.050 ;
        RECT 730.950 211.950 733.050 214.050 ;
        RECT 733.950 211.950 736.050 214.050 ;
        RECT 718.950 210.450 723.000 211.050 ;
        RECT 728.400 210.900 729.600 211.650 ;
        RECT 718.950 208.950 723.450 210.450 ;
        RECT 722.400 207.450 723.450 208.950 ;
        RECT 727.950 208.800 730.050 210.900 ;
        RECT 734.400 209.400 735.600 211.650 ;
        RECT 722.400 206.400 732.450 207.450 ;
        RECT 718.950 202.950 724.050 205.050 ;
        RECT 727.950 202.950 730.050 205.050 ;
        RECT 728.400 198.450 729.450 202.950 ;
        RECT 731.400 201.450 732.450 206.400 ;
        RECT 734.400 202.050 735.450 209.400 ;
        RECT 736.950 202.950 739.050 205.050 ;
        RECT 733.950 201.450 736.050 202.050 ;
        RECT 731.400 200.400 736.050 201.450 ;
        RECT 733.950 199.950 736.050 200.400 ;
        RECT 737.400 198.450 738.450 202.950 ;
        RECT 728.400 197.400 738.450 198.450 ;
        RECT 740.400 196.050 741.450 215.100 ;
        RECT 743.400 211.050 744.450 223.950 ;
        RECT 752.400 223.050 753.450 232.950 ;
        RECT 766.950 229.950 769.050 232.050 ;
        RECT 751.950 220.950 754.050 223.050 ;
        RECT 752.400 216.600 753.450 220.950 ;
        RECT 752.400 214.350 753.600 216.600 ;
        RECT 757.950 215.100 760.050 217.200 ;
        RECT 758.400 214.350 759.600 215.100 ;
        RECT 763.950 214.950 766.050 217.200 ;
        RECT 748.950 211.950 751.050 214.050 ;
        RECT 751.950 211.950 754.050 214.050 ;
        RECT 754.950 211.950 757.050 214.050 ;
        RECT 757.950 211.950 760.050 214.050 ;
        RECT 742.950 208.950 745.050 211.050 ;
        RECT 749.400 210.900 750.600 211.650 ;
        RECT 755.400 210.900 756.600 211.650 ;
        RECT 748.950 208.800 751.050 210.900 ;
        RECT 754.950 208.800 757.050 210.900 ;
        RECT 760.950 205.950 763.050 210.900 ;
        RECT 764.400 205.050 765.450 214.950 ;
        RECT 767.400 211.050 768.450 229.950 ;
        RECT 784.950 220.950 787.050 223.050 ;
        RECT 772.950 217.050 775.050 217.200 ;
        RECT 769.950 215.100 775.050 217.050 ;
        RECT 778.950 215.100 781.050 217.200 ;
        RECT 785.400 216.600 786.450 220.950 ;
        RECT 797.400 220.050 798.450 295.950 ;
        RECT 805.950 293.100 808.050 295.200 ;
        RECT 811.950 294.000 814.050 298.050 ;
        RECT 821.400 295.200 822.450 371.400 ;
        RECT 827.400 370.350 828.600 372.600 ;
        RECT 832.950 371.100 835.050 373.200 ;
        RECT 833.400 370.350 834.600 371.100 ;
        RECT 826.950 367.950 829.050 370.050 ;
        RECT 829.950 367.950 832.050 370.050 ;
        RECT 832.950 367.950 835.050 370.050 ;
        RECT 830.400 366.900 831.600 367.650 ;
        RECT 829.950 364.800 832.050 366.900 ;
        RECT 839.400 358.050 840.450 385.950 ;
        RECT 838.950 355.950 841.050 358.050 ;
        RECT 842.400 351.450 843.450 397.950 ;
        RECT 839.400 350.400 843.450 351.450 ;
        RECT 839.400 343.050 840.450 350.400 ;
        RECT 841.950 348.450 844.050 349.050 ;
        RECT 845.400 348.450 846.450 410.400 ;
        RECT 850.950 403.800 853.050 405.900 ;
        RECT 851.400 373.200 852.450 403.800 ;
        RECT 857.400 397.050 858.450 410.400 ;
        RECT 863.400 406.050 864.450 410.400 ;
        RECT 872.400 409.050 873.450 475.950 ;
        RECT 875.400 427.050 876.450 511.950 ;
        RECT 878.400 511.050 879.450 520.950 ;
        RECT 877.950 508.950 880.050 511.050 ;
        RECT 881.400 495.450 882.450 538.950 ;
        RECT 884.400 529.050 885.450 595.950 ;
        RECT 890.400 541.050 891.450 610.950 ;
        RECT 892.950 604.950 895.050 607.050 ;
        RECT 893.400 556.050 894.450 604.950 ;
        RECT 899.400 598.050 900.450 643.950 ;
        RECT 898.950 595.950 901.050 598.050 ;
        RECT 898.950 580.950 901.050 583.050 ;
        RECT 899.400 565.050 900.450 580.950 ;
        RECT 898.950 562.950 901.050 565.050 ;
        RECT 892.950 553.950 895.050 556.050 ;
        RECT 889.950 538.950 892.050 541.050 ;
        RECT 886.950 532.950 889.050 535.050 ;
        RECT 883.950 526.950 886.050 529.050 ;
        RECT 887.400 528.600 888.450 532.950 ;
        RECT 887.400 526.350 888.600 528.600 ;
        RECT 892.950 527.100 895.050 529.200 ;
        RECT 899.400 529.050 900.450 562.950 ;
        RECT 893.400 526.350 894.600 527.100 ;
        RECT 898.950 526.950 901.050 529.050 ;
        RECT 886.950 523.950 889.050 526.050 ;
        RECT 889.950 523.950 892.050 526.050 ;
        RECT 892.950 523.950 895.050 526.050 ;
        RECT 895.950 523.950 898.050 526.050 ;
        RECT 890.400 522.900 891.600 523.650 ;
        RECT 889.950 520.800 892.050 522.900 ;
        RECT 896.400 521.400 897.600 523.650 ;
        RECT 892.950 517.950 895.050 520.050 ;
        RECT 893.400 499.050 894.450 517.950 ;
        RECT 896.400 514.050 897.450 521.400 ;
        RECT 898.950 520.950 901.050 523.050 ;
        RECT 895.950 511.950 898.050 514.050 ;
        RECT 892.950 496.950 895.050 499.050 ;
        RECT 878.400 494.400 882.450 495.450 ;
        RECT 878.400 448.050 879.450 494.400 ;
        RECT 886.950 494.100 889.050 496.200 ;
        RECT 893.400 495.450 894.600 495.600 ;
        RECT 896.400 495.450 897.450 511.950 ;
        RECT 893.400 494.400 897.450 495.450 ;
        RECT 887.400 493.350 888.600 494.100 ;
        RECT 893.400 493.350 894.600 494.400 ;
        RECT 883.950 490.950 886.050 493.050 ;
        RECT 886.950 490.950 889.050 493.050 ;
        RECT 889.950 490.950 892.050 493.050 ;
        RECT 892.950 490.950 895.050 493.050 ;
        RECT 884.400 489.450 885.600 490.650 ;
        RECT 890.400 489.900 891.600 490.650 ;
        RECT 881.400 488.400 885.600 489.450 ;
        RECT 881.400 484.050 882.450 488.400 ;
        RECT 889.950 487.800 892.050 489.900 ;
        RECT 895.950 487.800 898.050 489.900 ;
        RECT 883.950 484.950 886.050 487.050 ;
        RECT 880.950 481.950 883.050 484.050 ;
        RECT 884.400 481.050 885.450 484.950 ;
        RECT 883.950 478.950 886.050 481.050 ;
        RECT 883.950 449.100 886.050 451.200 ;
        RECT 889.950 450.000 892.050 454.050 ;
        RECT 896.400 451.050 897.450 487.800 ;
        RECT 899.400 466.050 900.450 520.950 ;
        RECT 898.950 463.950 901.050 466.050 ;
        RECT 898.950 457.950 901.050 460.050 ;
        RECT 884.400 448.350 885.600 449.100 ;
        RECT 890.400 448.350 891.600 450.000 ;
        RECT 895.950 448.950 898.050 451.050 ;
        RECT 877.950 445.950 880.050 448.050 ;
        RECT 883.950 445.950 886.050 448.050 ;
        RECT 886.950 445.950 889.050 448.050 ;
        RECT 889.950 445.950 892.050 448.050 ;
        RECT 892.950 445.950 895.050 448.050 ;
        RECT 887.400 444.900 888.600 445.650 ;
        RECT 893.400 444.900 894.600 445.650 ;
        RECT 877.950 442.800 880.050 444.900 ;
        RECT 886.950 442.800 889.050 444.900 ;
        RECT 892.950 442.800 895.050 444.900 ;
        RECT 878.400 436.050 879.450 442.800 ;
        RECT 889.950 439.950 892.050 442.050 ;
        RECT 877.950 433.950 880.050 436.050 ;
        RECT 874.950 424.950 877.050 427.050 ;
        RECT 878.400 423.450 879.450 433.950 ;
        RECT 875.400 422.400 879.450 423.450 ;
        RECT 871.950 406.950 874.050 409.050 ;
        RECT 862.950 403.950 865.050 406.050 ;
        RECT 856.950 394.950 859.050 397.050 ;
        RECT 862.950 385.950 865.050 388.050 ;
        RECT 850.950 371.100 853.050 373.200 ;
        RECT 851.400 370.350 852.600 371.100 ;
        RECT 850.950 367.950 853.050 370.050 ;
        RECT 853.950 367.950 856.050 370.050 ;
        RECT 847.950 355.950 850.050 358.050 ;
        RECT 841.950 347.400 846.450 348.450 ;
        RECT 841.950 346.950 844.050 347.400 ;
        RECT 838.950 340.950 841.050 343.050 ;
        RECT 823.950 337.950 826.050 340.050 ;
        RECT 832.950 338.100 835.050 340.200 ;
        RECT 839.400 339.450 840.600 339.600 ;
        RECT 842.400 339.450 843.450 346.950 ;
        RECT 839.400 338.400 843.450 339.450 ;
        RECT 824.400 310.050 825.450 337.950 ;
        RECT 833.400 337.350 834.600 338.100 ;
        RECT 839.400 337.350 840.600 338.400 ;
        RECT 829.950 334.950 832.050 337.050 ;
        RECT 832.950 334.950 835.050 337.050 ;
        RECT 835.950 334.950 838.050 337.050 ;
        RECT 838.950 334.950 841.050 337.050 ;
        RECT 830.400 333.900 831.600 334.650 ;
        RECT 829.950 331.800 832.050 333.900 ;
        RECT 836.400 332.400 837.600 334.650 ;
        RECT 830.400 313.050 831.450 331.800 ;
        RECT 836.400 328.050 837.450 332.400 ;
        RECT 835.950 325.950 838.050 328.050 ;
        RECT 848.400 319.050 849.450 355.950 ;
        RECT 863.400 354.450 864.450 385.950 ;
        RECT 875.400 376.050 876.450 422.400 ;
        RECT 880.950 416.100 883.050 418.200 ;
        RECT 881.400 415.350 882.600 416.100 ;
        RECT 880.950 412.950 883.050 415.050 ;
        RECT 883.950 412.950 886.050 415.050 ;
        RECT 884.400 410.400 885.600 412.650 ;
        RECT 884.400 409.050 885.450 410.400 ;
        RECT 883.950 406.950 886.050 409.050 ;
        RECT 884.400 405.450 885.450 406.950 ;
        RECT 884.400 404.400 888.450 405.450 ;
        RECT 883.950 400.950 886.050 403.050 ;
        RECT 877.950 376.950 880.050 379.050 ;
        RECT 874.950 373.950 877.050 376.050 ;
        RECT 878.400 373.200 879.450 376.950 ;
        RECT 877.950 371.100 880.050 373.200 ;
        RECT 878.400 370.350 879.600 371.100 ;
        RECT 871.950 367.950 874.050 370.050 ;
        RECT 874.950 367.950 877.050 370.050 ;
        RECT 877.950 367.950 880.050 370.050 ;
        RECT 875.400 366.900 876.600 367.650 ;
        RECT 874.950 364.800 877.050 366.900 ;
        RECT 884.400 364.050 885.450 400.950 ;
        RECT 877.950 361.950 880.050 364.050 ;
        RECT 883.950 361.950 886.050 364.050 ;
        RECT 868.950 358.950 871.050 361.050 ;
        RECT 863.400 353.400 867.450 354.450 ;
        RECT 850.950 349.950 853.050 352.050 ;
        RECT 851.400 340.050 852.450 349.950 ;
        RECT 855.000 342.450 859.050 343.050 ;
        RECT 854.400 340.950 859.050 342.450 ;
        RECT 850.950 337.950 853.050 340.050 ;
        RECT 854.400 339.600 855.450 340.950 ;
        RECT 866.400 340.050 867.450 353.400 ;
        RECT 854.400 337.350 855.600 339.600 ;
        RECT 865.950 337.950 868.050 340.050 ;
        RECT 853.950 334.950 856.050 337.050 ;
        RECT 856.950 334.950 859.050 337.050 ;
        RECT 859.950 334.950 862.050 337.050 ;
        RECT 862.950 334.950 865.050 337.050 ;
        RECT 850.950 331.950 853.050 334.050 ;
        RECT 863.400 332.400 864.600 334.650 ;
        RECT 869.400 333.450 870.450 358.950 ;
        RECT 874.950 346.950 877.050 349.050 ;
        RECT 875.400 340.050 876.450 346.950 ;
        RECT 874.950 337.950 877.050 340.050 ;
        RECT 878.400 339.600 879.450 361.950 ;
        RECT 887.400 352.050 888.450 404.400 ;
        RECT 886.950 349.950 889.050 352.050 ;
        RECT 890.400 349.050 891.450 439.950 ;
        RECT 895.950 416.100 898.050 418.200 ;
        RECT 892.950 394.950 895.050 397.050 ;
        RECT 889.950 346.950 892.050 349.050 ;
        RECT 878.400 337.350 879.600 339.600 ;
        RECT 877.950 334.950 880.050 337.050 ;
        RECT 880.950 334.950 883.050 337.050 ;
        RECT 883.950 334.950 886.050 337.050 ;
        RECT 886.950 334.950 889.050 337.050 ;
        RECT 866.400 332.400 870.450 333.450 ;
        RECT 841.950 316.950 844.050 319.050 ;
        RECT 847.950 316.950 850.050 319.050 ;
        RECT 829.950 310.950 832.050 313.050 ;
        RECT 823.950 307.950 826.050 310.050 ;
        RECT 824.400 297.450 825.450 307.950 ;
        RECT 830.400 298.050 831.450 310.950 ;
        RECT 824.400 296.400 828.450 297.450 ;
        RECT 820.950 294.450 823.050 295.200 ;
        RECT 806.400 292.350 807.600 293.100 ;
        RECT 812.400 292.350 813.600 294.000 ;
        RECT 818.400 293.400 823.050 294.450 ;
        RECT 802.950 289.950 805.050 292.050 ;
        RECT 805.950 289.950 808.050 292.050 ;
        RECT 808.950 289.950 811.050 292.050 ;
        RECT 811.950 289.950 814.050 292.050 ;
        RECT 803.400 288.900 804.600 289.650 ;
        RECT 809.400 288.900 810.600 289.650 ;
        RECT 802.950 286.800 805.050 288.900 ;
        RECT 808.950 286.800 811.050 288.900 ;
        RECT 799.950 268.950 802.050 271.050 ;
        RECT 800.400 262.050 801.450 268.950 ;
        RECT 799.950 259.950 802.050 262.050 ;
        RECT 805.950 261.000 808.050 265.050 ;
        RECT 806.400 259.350 807.600 261.000 ;
        RECT 811.950 260.100 814.050 262.200 ;
        RECT 812.400 259.350 813.600 260.100 ;
        RECT 802.950 256.950 805.050 259.050 ;
        RECT 805.950 256.950 808.050 259.050 ;
        RECT 808.950 256.950 811.050 259.050 ;
        RECT 811.950 256.950 814.050 259.050 ;
        RECT 803.400 255.000 804.600 256.650 ;
        RECT 809.400 255.900 810.600 256.650 ;
        RECT 802.950 250.950 805.050 255.000 ;
        RECT 808.950 253.800 811.050 255.900 ;
        RECT 818.400 223.050 819.450 293.400 ;
        RECT 820.950 293.100 823.050 293.400 ;
        RECT 827.400 294.600 828.450 296.400 ;
        RECT 829.950 295.950 832.050 298.050 ;
        RECT 827.400 292.350 828.600 294.600 ;
        RECT 832.950 294.000 835.050 298.050 ;
        RECT 833.400 292.350 834.600 294.000 ;
        RECT 842.400 292.050 843.450 316.950 ;
        RECT 847.950 310.950 850.050 313.050 ;
        RECT 826.950 289.950 829.050 292.050 ;
        RECT 829.950 289.950 832.050 292.050 ;
        RECT 832.950 289.950 835.050 292.050 ;
        RECT 835.950 289.950 838.050 292.050 ;
        RECT 841.950 289.950 844.050 292.050 ;
        RECT 830.400 287.400 831.600 289.650 ;
        RECT 836.400 289.050 837.600 289.650 ;
        RECT 836.400 287.400 841.050 289.050 ;
        RECT 830.400 280.050 831.450 287.400 ;
        RECT 837.000 286.950 841.050 287.400 ;
        RECT 829.950 277.950 832.050 280.050 ;
        RECT 820.950 265.950 823.050 268.050 ;
        RECT 790.950 217.950 793.050 220.050 ;
        RECT 793.950 217.950 796.050 220.050 ;
        RECT 796.950 217.950 799.050 220.050 ;
        RECT 799.950 217.950 802.050 223.050 ;
        RECT 805.950 220.950 811.050 223.050 ;
        RECT 814.950 220.950 817.050 223.050 ;
        RECT 817.950 220.950 820.050 223.050 ;
        RECT 769.950 214.950 774.000 215.100 ;
        RECT 779.400 214.350 780.600 215.100 ;
        RECT 785.400 214.350 786.600 216.600 ;
        RECT 775.950 211.950 778.050 214.050 ;
        RECT 778.950 211.950 781.050 214.050 ;
        RECT 781.950 211.950 784.050 214.050 ;
        RECT 784.950 211.950 787.050 214.050 ;
        RECT 766.950 208.950 769.050 211.050 ;
        RECT 769.950 205.950 772.050 211.050 ;
        RECT 776.400 210.900 777.600 211.650 ;
        RECT 775.950 208.800 778.050 210.900 ;
        RECT 782.400 210.000 783.600 211.650 ;
        RECT 781.950 205.950 784.050 210.000 ;
        RECT 763.950 202.950 766.050 205.050 ;
        RECT 769.950 199.950 772.050 202.050 ;
        RECT 748.950 196.950 751.050 199.050 ;
        RECT 721.950 193.950 724.050 196.050 ;
        RECT 730.950 193.950 733.050 196.050 ;
        RECT 739.950 193.950 742.050 196.050 ;
        RECT 745.950 193.950 748.050 196.050 ;
        RECT 718.950 187.950 721.050 190.050 ;
        RECT 704.400 181.350 705.600 182.100 ;
        RECT 710.400 181.350 711.600 183.600 ;
        RECT 715.950 181.950 718.050 184.050 ;
        RECT 700.950 178.950 703.050 181.050 ;
        RECT 703.950 178.950 706.050 181.050 ;
        RECT 706.950 178.950 709.050 181.050 ;
        RECT 709.950 178.950 712.050 181.050 ;
        RECT 701.400 177.000 702.600 178.650 ;
        RECT 700.950 172.950 703.050 177.000 ;
        RECT 707.400 176.400 708.600 178.650 ;
        RECT 694.950 169.950 697.050 172.050 ;
        RECT 676.950 157.950 679.050 160.050 ;
        RECT 707.400 154.050 708.450 176.400 ;
        RECT 712.950 175.950 715.050 178.050 ;
        RECT 706.950 151.950 709.050 154.050 ;
        RECT 694.950 148.950 697.050 151.050 ;
        RECT 682.950 142.950 685.050 145.050 ;
        RECT 668.400 138.450 669.600 138.600 ;
        RECT 665.400 137.400 669.600 138.450 ;
        RECT 662.400 133.050 663.450 137.100 ;
        RECT 668.400 136.350 669.600 137.400 ;
        RECT 673.950 137.100 676.050 139.200 ;
        RECT 674.400 136.350 675.600 137.100 ;
        RECT 667.950 133.950 670.050 136.050 ;
        RECT 670.950 133.950 673.050 136.050 ;
        RECT 673.950 133.950 676.050 136.050 ;
        RECT 676.950 133.950 679.050 136.050 ;
        RECT 661.950 130.950 664.050 133.050 ;
        RECT 671.400 132.900 672.600 133.650 ;
        RECT 670.950 130.800 673.050 132.900 ;
        RECT 677.400 131.400 678.600 133.650 ;
        RECT 677.400 124.050 678.450 131.400 ;
        RECT 683.400 127.050 684.450 142.950 ;
        RECT 695.400 141.450 696.450 148.950 ;
        RECT 713.400 148.050 714.450 175.950 ;
        RECT 719.400 160.050 720.450 187.950 ;
        RECT 718.950 157.950 721.050 160.050 ;
        RECT 722.400 157.050 723.450 193.950 ;
        RECT 731.400 190.050 732.450 193.950 ;
        RECT 742.950 190.950 745.050 193.050 ;
        RECT 730.950 187.950 733.050 190.050 ;
        RECT 736.950 186.450 739.050 190.050 ;
        RECT 734.400 186.000 739.050 186.450 ;
        RECT 734.400 185.400 738.450 186.000 ;
        RECT 724.950 183.600 729.000 184.050 ;
        RECT 734.400 183.600 735.450 185.400 ;
        RECT 724.950 181.950 729.600 183.600 ;
        RECT 728.400 181.350 729.600 181.950 ;
        RECT 734.400 181.350 735.600 183.600 ;
        RECT 727.950 178.950 730.050 181.050 ;
        RECT 730.950 178.950 733.050 181.050 ;
        RECT 733.950 178.950 736.050 181.050 ;
        RECT 736.950 178.950 739.050 181.050 ;
        RECT 731.400 177.900 732.600 178.650 ;
        RECT 737.400 177.900 738.600 178.650 ;
        RECT 724.950 175.800 727.050 177.900 ;
        RECT 730.950 175.800 733.050 177.900 ;
        RECT 736.950 175.800 739.050 177.900 ;
        RECT 725.400 172.050 726.450 175.800 ;
        RECT 724.950 169.950 727.050 172.050 ;
        RECT 730.950 169.950 733.050 172.050 ;
        RECT 731.400 166.050 732.450 169.950 ;
        RECT 737.400 166.050 738.450 175.800 ;
        RECT 730.950 163.950 733.050 166.050 ;
        RECT 736.950 163.950 739.050 166.050 ;
        RECT 721.950 154.950 724.050 157.050 ;
        RECT 739.950 154.950 742.050 157.050 ;
        RECT 712.950 145.950 715.050 148.050 ;
        RECT 721.950 145.950 724.050 148.050 ;
        RECT 697.950 141.450 700.050 142.050 ;
        RECT 695.400 140.400 700.050 141.450 ;
        RECT 697.950 139.950 700.050 140.400 ;
        RECT 712.950 139.950 715.050 142.050 ;
        RECT 685.950 137.100 688.050 139.200 ;
        RECT 698.400 138.600 699.450 139.950 ;
        RECT 686.400 133.050 687.450 137.100 ;
        RECT 698.400 136.350 699.600 138.600 ;
        RECT 703.950 137.100 706.050 139.200 ;
        RECT 709.950 137.100 712.050 139.200 ;
        RECT 704.400 136.350 705.600 137.100 ;
        RECT 694.950 133.950 697.050 136.050 ;
        RECT 697.950 133.950 700.050 136.050 ;
        RECT 700.950 133.950 703.050 136.050 ;
        RECT 703.950 133.950 706.050 136.050 ;
        RECT 685.950 130.950 688.050 133.050 ;
        RECT 695.400 132.900 696.600 133.650 ;
        RECT 694.950 130.800 697.050 132.900 ;
        RECT 701.400 131.400 702.600 133.650 ;
        RECT 710.400 132.450 711.450 137.100 ;
        RECT 707.400 131.400 711.450 132.450 ;
        RECT 682.950 124.950 685.050 127.050 ;
        RECT 676.950 121.950 679.050 124.050 ;
        RECT 701.400 115.050 702.450 131.400 ;
        RECT 707.400 118.050 708.450 131.400 ;
        RECT 709.950 124.950 712.050 127.050 ;
        RECT 710.400 121.050 711.450 124.950 ;
        RECT 709.950 118.950 712.050 121.050 ;
        RECT 706.950 115.950 709.050 118.050 ;
        RECT 667.950 112.950 670.050 115.050 ;
        RECT 700.950 112.950 703.050 115.050 ;
        RECT 668.400 105.600 669.450 112.950 ;
        RECT 701.400 108.450 702.450 112.950 ;
        RECT 701.400 107.400 705.450 108.450 ;
        RECT 668.400 103.350 669.600 105.600 ;
        RECT 673.950 103.950 676.050 106.050 ;
        RECT 688.950 104.100 691.050 106.200 ;
        RECT 694.950 104.100 697.050 106.200 ;
        RECT 700.950 104.100 703.050 106.200 ;
        RECT 664.950 100.950 667.050 103.050 ;
        RECT 667.950 100.950 670.050 103.050 ;
        RECT 665.400 98.400 666.600 100.650 ;
        RECT 665.400 97.050 666.450 98.400 ;
        RECT 661.950 95.400 666.450 97.050 ;
        RECT 661.950 94.950 666.000 95.400 ;
        RECT 674.400 94.050 675.450 103.950 ;
        RECT 689.400 103.350 690.600 104.100 ;
        RECT 695.400 103.350 696.600 104.100 ;
        RECT 685.950 100.950 688.050 103.050 ;
        RECT 688.950 100.950 691.050 103.050 ;
        RECT 691.950 100.950 694.050 103.050 ;
        RECT 694.950 100.950 697.050 103.050 ;
        RECT 686.400 98.400 687.600 100.650 ;
        RECT 692.400 98.400 693.600 100.650 ;
        RECT 673.950 91.950 676.050 94.050 ;
        RECT 686.400 91.050 687.450 98.400 ;
        RECT 685.950 88.950 688.050 91.050 ;
        RECT 643.950 73.950 646.050 76.050 ;
        RECT 658.950 73.950 661.050 76.050 ;
        RECT 625.950 61.950 628.050 64.050 ;
        RECT 631.950 61.950 634.050 64.050 ;
        RECT 596.400 60.450 597.600 60.600 ;
        RECT 596.400 59.400 603.450 60.450 ;
        RECT 590.400 58.350 591.600 59.100 ;
        RECT 596.400 58.350 597.600 59.400 ;
        RECT 589.950 55.950 592.050 58.050 ;
        RECT 592.950 55.950 595.050 58.050 ;
        RECT 595.950 55.950 598.050 58.050 ;
        RECT 586.950 52.950 589.050 55.050 ;
        RECT 593.400 54.000 594.600 55.650 ;
        RECT 587.400 31.050 588.450 52.950 ;
        RECT 592.950 49.950 595.050 54.000 ;
        RECT 602.400 46.050 603.450 59.400 ;
        RECT 614.400 58.350 615.600 60.600 ;
        RECT 604.950 55.950 607.050 58.050 ;
        RECT 610.950 55.950 613.050 58.050 ;
        RECT 613.950 55.950 616.050 58.050 ;
        RECT 616.950 55.950 619.050 58.050 ;
        RECT 605.400 52.050 606.450 55.950 ;
        RECT 611.400 53.400 612.600 55.650 ;
        RECT 617.400 54.900 618.600 55.650 ;
        RECT 626.400 55.050 627.450 61.950 ;
        RECT 634.950 59.100 637.050 61.200 ;
        RECT 635.400 58.350 636.600 59.100 ;
        RECT 631.950 55.950 634.050 58.050 ;
        RECT 634.950 55.950 637.050 58.050 ;
        RECT 637.950 55.950 640.050 58.050 ;
        RECT 604.950 49.950 607.050 52.050 ;
        RECT 611.400 46.050 612.450 53.400 ;
        RECT 616.950 52.800 619.050 54.900 ;
        RECT 625.950 52.950 628.050 55.050 ;
        RECT 632.400 54.450 633.600 55.650 ;
        RECT 629.400 53.400 633.600 54.450 ;
        RECT 638.400 53.400 639.600 55.650 ;
        RECT 617.400 49.050 618.450 52.800 ;
        RECT 616.950 46.950 619.050 49.050 ;
        RECT 589.950 43.950 592.050 46.050 ;
        RECT 601.950 43.950 604.050 46.050 ;
        RECT 610.950 43.950 613.050 46.050 ;
        RECT 586.950 28.950 589.050 31.050 ;
        RECT 590.400 27.600 591.450 43.950 ;
        RECT 629.400 43.050 630.450 53.400 ;
        RECT 631.950 46.950 634.050 49.050 ;
        RECT 628.950 40.950 631.050 43.050 ;
        RECT 632.400 33.450 633.450 46.950 ;
        RECT 638.400 37.050 639.450 53.400 ;
        RECT 640.950 52.950 643.050 55.050 ;
        RECT 637.950 34.950 640.050 37.050 ;
        RECT 641.400 34.050 642.450 52.950 ;
        RECT 644.400 40.050 645.450 73.950 ;
        RECT 652.950 64.950 655.050 67.050 ;
        RECT 658.950 64.950 664.050 67.050 ;
        RECT 670.950 64.950 673.050 67.050 ;
        RECT 682.950 64.950 685.050 67.050 ;
        RECT 646.950 58.950 649.050 61.050 ;
        RECT 653.400 60.600 654.450 64.950 ;
        RECT 647.400 46.050 648.450 58.950 ;
        RECT 653.400 58.350 654.600 60.600 ;
        RECT 658.950 60.000 661.050 63.900 ;
        RECT 659.400 58.350 660.600 60.000 ;
        RECT 667.950 59.100 670.050 61.200 ;
        RECT 652.950 55.950 655.050 58.050 ;
        RECT 655.950 55.950 658.050 58.050 ;
        RECT 658.950 55.950 661.050 58.050 ;
        RECT 661.950 55.950 664.050 58.050 ;
        RECT 656.400 54.900 657.600 55.650 ;
        RECT 662.400 54.900 663.600 55.650 ;
        RECT 655.950 52.800 658.050 54.900 ;
        RECT 661.950 52.800 664.050 54.900 ;
        RECT 656.400 49.050 657.450 52.800 ;
        RECT 668.400 49.050 669.450 59.100 ;
        RECT 671.400 52.050 672.450 64.950 ;
        RECT 676.950 59.100 679.050 61.200 ;
        RECT 683.400 60.600 684.450 64.950 ;
        RECT 686.400 64.050 687.450 88.950 ;
        RECT 685.950 61.950 688.050 64.050 ;
        RECT 677.400 58.350 678.600 59.100 ;
        RECT 683.400 58.350 684.600 60.600 ;
        RECT 676.950 55.950 679.050 58.050 ;
        RECT 679.950 55.950 682.050 58.050 ;
        RECT 682.950 55.950 685.050 58.050 ;
        RECT 685.950 55.950 688.050 58.050 ;
        RECT 680.400 54.900 681.600 55.650 ;
        RECT 670.950 49.950 673.050 52.050 ;
        RECT 679.950 49.950 682.050 54.900 ;
        RECT 686.400 54.000 687.600 55.650 ;
        RECT 685.950 49.950 688.050 54.000 ;
        RECT 692.400 52.050 693.450 98.400 ;
        RECT 701.400 97.050 702.450 104.100 ;
        RECT 700.950 94.950 703.050 97.050 ;
        RECT 704.400 91.050 705.450 107.400 ;
        RECT 707.400 100.050 708.450 115.950 ;
        RECT 713.400 112.050 714.450 139.950 ;
        RECT 722.400 138.600 723.450 145.950 ;
        RECT 740.400 145.050 741.450 154.950 ;
        RECT 739.950 142.950 742.050 145.050 ;
        RECT 722.400 136.350 723.600 138.600 ;
        RECT 727.950 137.100 730.050 139.200 ;
        RECT 728.400 136.350 729.600 137.100 ;
        RECT 718.950 133.950 721.050 136.050 ;
        RECT 721.950 133.950 724.050 136.050 ;
        RECT 724.950 133.950 727.050 136.050 ;
        RECT 727.950 133.950 730.050 136.050 ;
        RECT 719.400 132.000 720.600 133.650 ;
        RECT 718.950 127.950 721.050 132.000 ;
        RECT 725.400 131.400 726.600 133.650 ;
        RECT 721.950 124.950 724.050 127.050 ;
        RECT 712.950 109.950 715.050 112.050 ;
        RECT 713.400 108.450 714.450 109.950 ;
        RECT 713.400 107.400 717.450 108.450 ;
        RECT 716.400 106.200 717.450 107.400 ;
        RECT 715.950 104.100 718.050 106.200 ;
        RECT 722.400 105.600 723.450 124.950 ;
        RECT 725.400 118.050 726.450 131.400 ;
        RECT 730.950 130.950 733.050 133.050 ;
        RECT 740.400 132.900 741.450 142.950 ;
        RECT 743.400 139.200 744.450 190.950 ;
        RECT 746.400 172.050 747.450 193.950 ;
        RECT 749.400 184.050 750.450 196.950 ;
        RECT 766.950 187.950 769.050 190.050 ;
        RECT 748.950 181.950 751.050 184.050 ;
        RECT 751.950 182.100 754.050 184.200 ;
        RECT 757.950 182.100 760.050 184.200 ;
        RECT 752.400 181.350 753.600 182.100 ;
        RECT 758.400 181.350 759.600 182.100 ;
        RECT 751.950 178.950 754.050 181.050 ;
        RECT 754.950 178.950 757.050 181.050 ;
        RECT 757.950 178.950 760.050 181.050 ;
        RECT 760.950 178.950 763.050 181.050 ;
        RECT 748.950 175.950 751.050 178.050 ;
        RECT 755.400 176.400 756.600 178.650 ;
        RECT 761.400 177.000 762.600 178.650 ;
        RECT 745.950 169.950 748.050 172.050 ;
        RECT 749.400 154.050 750.450 175.950 ;
        RECT 755.400 174.450 756.450 176.400 ;
        RECT 757.950 174.450 760.050 175.050 ;
        RECT 755.400 173.400 760.050 174.450 ;
        RECT 757.950 172.950 760.050 173.400 ;
        RECT 760.950 172.950 763.050 177.000 ;
        RECT 767.400 175.050 768.450 187.950 ;
        RECT 770.400 178.050 771.450 199.950 ;
        RECT 775.950 196.950 778.050 199.050 ;
        RECT 776.400 183.600 777.450 196.950 ;
        RECT 776.400 181.350 777.600 183.600 ;
        RECT 781.950 182.100 784.050 184.200 ;
        RECT 782.400 181.350 783.600 182.100 ;
        RECT 775.950 178.950 778.050 181.050 ;
        RECT 778.950 178.950 781.050 181.050 ;
        RECT 781.950 178.950 784.050 181.050 ;
        RECT 784.950 178.950 787.050 181.050 ;
        RECT 769.950 175.950 772.050 178.050 ;
        RECT 779.400 177.000 780.600 178.650 ;
        RECT 766.950 172.950 769.050 175.050 ;
        RECT 778.950 172.950 781.050 177.000 ;
        RECT 785.400 176.400 786.600 178.650 ;
        RECT 758.400 157.050 759.450 172.950 ;
        RECT 778.950 163.950 781.050 166.050 ;
        RECT 757.950 154.950 760.050 157.050 ;
        RECT 748.950 151.950 751.050 154.050 ;
        RECT 742.950 137.100 745.050 139.200 ;
        RECT 752.400 138.450 753.600 138.600 ;
        RECT 752.400 137.400 756.450 138.450 ;
        RECT 743.400 136.350 744.600 137.100 ;
        RECT 752.400 136.350 753.600 137.400 ;
        RECT 743.100 133.950 745.200 136.050 ;
        RECT 748.500 133.950 750.600 136.050 ;
        RECT 751.800 133.950 753.900 136.050 ;
        RECT 749.400 132.900 750.600 133.650 ;
        RECT 731.400 127.050 732.450 130.950 ;
        RECT 739.950 130.800 742.050 132.900 ;
        RECT 748.950 127.950 751.050 132.900 ;
        RECT 730.950 124.950 733.050 127.050 ;
        RECT 724.950 115.950 727.050 118.050 ;
        RECT 751.950 115.950 754.050 118.050 ;
        RECT 752.400 108.450 753.450 115.950 ;
        RECT 755.400 112.050 756.450 137.400 ;
        RECT 758.400 127.050 759.450 154.950 ;
        RECT 772.950 142.950 775.050 145.050 ;
        RECT 766.950 137.100 769.050 139.200 ;
        RECT 773.400 138.600 774.450 142.950 ;
        RECT 767.400 136.350 768.600 137.100 ;
        RECT 773.400 136.350 774.600 138.600 ;
        RECT 766.950 133.950 769.050 136.050 ;
        RECT 769.950 133.950 772.050 136.050 ;
        RECT 772.950 133.950 775.050 136.050 ;
        RECT 770.400 132.900 771.600 133.650 ;
        RECT 769.950 130.800 772.050 132.900 ;
        RECT 779.400 127.050 780.450 163.950 ;
        RECT 785.400 157.050 786.450 176.400 ;
        RECT 787.950 175.950 790.050 178.050 ;
        RECT 784.950 154.950 787.050 157.050 ;
        RECT 788.400 151.050 789.450 175.950 ;
        RECT 791.400 175.050 792.450 217.950 ;
        RECT 794.400 208.050 795.450 217.950 ;
        RECT 802.950 215.100 805.050 217.200 ;
        RECT 808.950 216.000 811.050 219.900 ;
        RECT 803.400 214.350 804.600 215.100 ;
        RECT 809.400 214.350 810.600 216.000 ;
        RECT 799.950 211.950 802.050 214.050 ;
        RECT 802.950 211.950 805.050 214.050 ;
        RECT 805.950 211.950 808.050 214.050 ;
        RECT 808.950 211.950 811.050 214.050 ;
        RECT 796.950 208.950 799.050 211.050 ;
        RECT 800.400 209.400 801.600 211.650 ;
        RECT 806.400 210.900 807.600 211.650 ;
        RECT 815.400 211.050 816.450 220.950 ;
        RECT 817.950 217.800 820.050 219.900 ;
        RECT 793.950 205.950 796.050 208.050 ;
        RECT 797.400 202.050 798.450 208.950 ;
        RECT 796.950 199.950 799.050 202.050 ;
        RECT 800.400 196.050 801.450 209.400 ;
        RECT 805.950 208.800 808.050 210.900 ;
        RECT 814.950 208.950 817.050 211.050 ;
        RECT 793.950 193.950 796.050 196.050 ;
        RECT 799.950 193.950 802.050 196.050 ;
        RECT 790.950 172.950 793.050 175.050 ;
        RECT 794.400 160.050 795.450 193.950 ;
        RECT 805.950 190.950 808.050 193.050 ;
        RECT 806.400 184.200 807.450 190.950 ;
        RECT 818.400 186.450 819.450 217.800 ;
        RECT 821.400 217.050 822.450 265.950 ;
        RECT 842.400 262.200 843.450 289.950 ;
        RECT 826.950 260.100 829.050 262.200 ;
        RECT 832.950 260.100 835.050 262.200 ;
        RECT 841.950 260.100 844.050 262.200 ;
        RECT 848.400 261.450 849.450 310.950 ;
        RECT 851.400 295.050 852.450 331.950 ;
        RECT 856.950 325.950 859.050 330.750 ;
        RECT 863.400 325.050 864.450 332.400 ;
        RECT 862.950 322.950 865.050 325.050 ;
        RECT 856.800 300.000 858.900 301.050 ;
        RECT 856.800 298.950 859.050 300.000 ;
        RECT 856.950 295.950 859.050 298.950 ;
        RECT 866.400 295.050 867.450 332.400 ;
        RECT 874.950 331.950 877.050 334.050 ;
        RECT 887.400 332.400 888.600 334.650 ;
        RECT 868.950 328.950 871.050 331.050 ;
        RECT 850.950 292.950 853.050 295.050 ;
        RECT 865.950 292.950 868.050 295.050 ;
        RECT 853.950 289.950 856.050 292.050 ;
        RECT 856.950 289.950 859.050 292.050 ;
        RECT 859.950 289.950 862.050 292.050 ;
        RECT 862.950 289.950 865.050 292.050 ;
        RECT 863.400 288.900 864.600 289.650 ;
        RECT 862.950 286.800 865.050 288.900 ;
        RECT 853.950 283.950 856.050 286.050 ;
        RECT 854.400 277.050 855.450 283.950 ;
        RECT 853.950 274.950 856.050 277.050 ;
        RECT 850.950 268.950 853.050 271.050 ;
        RECT 845.400 260.400 849.450 261.450 ;
        RECT 851.400 261.600 852.450 268.950 ;
        RECT 827.400 259.350 828.600 260.100 ;
        RECT 833.400 259.350 834.600 260.100 ;
        RECT 826.950 256.950 829.050 259.050 ;
        RECT 829.950 256.950 832.050 259.050 ;
        RECT 832.950 256.950 835.050 259.050 ;
        RECT 835.950 256.950 838.050 259.050 ;
        RECT 830.400 254.400 831.600 256.650 ;
        RECT 836.400 256.050 837.600 256.650 ;
        RECT 845.400 256.050 846.450 260.400 ;
        RECT 851.400 259.350 852.600 261.600 ;
        RECT 856.950 261.000 859.050 265.050 ;
        RECT 857.400 259.350 858.600 261.000 ;
        RECT 865.950 259.950 868.050 262.050 ;
        RECT 850.950 256.950 853.050 259.050 ;
        RECT 853.950 256.950 856.050 259.050 ;
        RECT 856.950 256.950 859.050 259.050 ;
        RECT 859.950 256.950 862.050 259.050 ;
        RECT 836.400 254.400 841.050 256.050 ;
        RECT 830.400 250.050 831.450 254.400 ;
        RECT 837.000 253.950 841.050 254.400 ;
        RECT 844.950 253.950 847.050 256.050 ;
        RECT 854.400 255.900 855.600 256.650 ;
        RECT 829.950 247.950 832.050 250.050 ;
        RECT 839.400 241.050 840.450 253.950 ;
        RECT 853.950 253.800 856.050 255.900 ;
        RECT 860.400 254.400 861.600 256.650 ;
        RECT 844.950 250.800 847.050 252.900 ;
        RECT 823.950 238.950 826.050 241.050 ;
        RECT 838.950 238.950 841.050 241.050 ;
        RECT 824.400 220.050 825.450 238.950 ;
        RECT 841.950 232.950 844.050 235.050 ;
        RECT 823.950 217.950 826.050 220.050 ;
        RECT 820.950 214.950 823.050 217.050 ;
        RECT 826.950 216.000 829.050 220.050 ;
        RECT 832.950 217.950 838.050 220.050 ;
        RECT 842.400 217.050 843.450 232.950 ;
        RECT 845.400 217.050 846.450 250.800 ;
        RECT 854.400 250.050 855.450 253.800 ;
        RECT 853.950 247.950 856.050 250.050 ;
        RECT 860.400 241.050 861.450 254.400 ;
        RECT 859.950 238.950 862.050 241.050 ;
        RECT 859.950 220.950 862.050 223.050 ;
        RECT 847.950 219.450 852.000 220.050 ;
        RECT 847.950 217.950 852.450 219.450 ;
        RECT 834.000 216.900 837.000 217.050 ;
        RECT 834.000 216.600 838.050 216.900 ;
        RECT 827.400 214.350 828.600 216.000 ;
        RECT 833.400 214.950 838.050 216.600 ;
        RECT 841.950 214.950 844.050 217.050 ;
        RECT 844.950 214.950 847.050 217.050 ;
        RECT 851.400 216.600 852.450 217.950 ;
        RECT 833.400 214.350 834.600 214.950 ;
        RECT 835.950 214.800 838.050 214.950 ;
        RECT 823.950 211.950 826.050 214.050 ;
        RECT 826.950 211.950 829.050 214.050 ;
        RECT 829.950 211.950 832.050 214.050 ;
        RECT 832.950 211.950 835.050 214.050 ;
        RECT 838.950 211.950 841.050 214.050 ;
        RECT 824.400 210.900 825.600 211.650 ;
        RECT 823.950 208.800 826.050 210.900 ;
        RECT 830.400 209.400 831.600 211.650 ;
        RECT 820.950 187.950 823.050 190.050 ;
        RECT 815.400 185.400 819.450 186.450 ;
        RECT 799.950 182.100 802.050 184.200 ;
        RECT 805.950 182.100 808.050 184.200 ;
        RECT 800.400 181.350 801.600 182.100 ;
        RECT 806.400 181.350 807.600 182.100 ;
        RECT 799.950 178.950 802.050 181.050 ;
        RECT 802.950 178.950 805.050 181.050 ;
        RECT 805.950 178.950 808.050 181.050 ;
        RECT 808.950 178.950 811.050 181.050 ;
        RECT 803.400 177.000 804.600 178.650 ;
        RECT 802.950 172.950 805.050 177.000 ;
        RECT 809.400 176.400 810.600 178.650 ;
        RECT 809.400 166.050 810.450 176.400 ;
        RECT 815.400 175.050 816.450 185.400 ;
        RECT 821.400 184.050 822.450 187.950 ;
        RECT 830.400 187.050 831.450 209.400 ;
        RECT 839.400 189.450 840.450 211.950 ;
        RECT 842.400 205.050 843.450 214.950 ;
        RECT 851.400 214.350 852.600 216.600 ;
        RECT 847.950 211.950 850.050 214.050 ;
        RECT 850.950 211.950 853.050 214.050 ;
        RECT 853.950 211.950 856.050 214.050 ;
        RECT 848.400 210.000 849.600 211.650 ;
        RECT 854.400 210.000 855.600 211.650 ;
        RECT 847.950 205.950 850.050 210.000 ;
        RECT 853.950 205.950 856.050 210.000 ;
        RECT 860.400 208.050 861.450 220.950 ;
        RECT 866.400 220.050 867.450 259.950 ;
        RECT 869.400 255.900 870.450 328.950 ;
        RECT 871.950 307.950 874.050 310.050 ;
        RECT 872.400 262.050 873.450 307.950 ;
        RECT 875.400 298.050 876.450 331.950 ;
        RECT 887.400 325.050 888.450 332.400 ;
        RECT 893.400 325.050 894.450 394.950 ;
        RECT 896.400 361.050 897.450 416.100 ;
        RECT 899.400 388.050 900.450 457.950 ;
        RECT 898.950 385.950 901.050 388.050 ;
        RECT 898.950 371.100 901.050 373.200 ;
        RECT 895.950 358.950 898.050 361.050 ;
        RECT 886.950 322.950 889.050 325.050 ;
        RECT 892.950 322.950 895.050 325.050 ;
        RECT 887.400 298.200 888.450 322.950 ;
        RECT 874.950 295.950 877.050 298.050 ;
        RECT 886.950 296.100 889.050 298.200 ;
        RECT 892.950 295.800 895.050 297.900 ;
        RECT 899.400 297.450 900.450 371.100 ;
        RECT 896.400 296.400 900.450 297.450 ;
        RECT 877.950 289.950 880.050 292.050 ;
        RECT 880.950 289.950 883.050 292.050 ;
        RECT 883.950 289.950 886.050 292.050 ;
        RECT 886.950 289.950 889.050 292.050 ;
        RECT 878.400 288.900 879.600 289.650 ;
        RECT 877.950 286.800 880.050 288.900 ;
        RECT 878.400 268.050 879.450 286.800 ;
        RECT 877.950 265.950 880.050 268.050 ;
        RECT 889.950 265.950 892.050 268.050 ;
        RECT 871.950 259.950 874.050 262.050 ;
        RECT 877.950 260.100 880.050 262.200 ;
        RECT 878.400 259.350 879.600 260.100 ;
        RECT 874.950 256.950 877.050 259.050 ;
        RECT 877.950 256.950 880.050 259.050 ;
        RECT 880.950 256.950 883.050 259.050 ;
        RECT 875.400 255.900 876.600 256.650 ;
        RECT 868.950 253.800 871.050 255.900 ;
        RECT 874.950 253.800 877.050 255.900 ;
        RECT 881.400 255.000 882.600 256.650 ;
        RECT 880.950 252.450 883.050 255.000 ;
        RECT 890.400 253.050 891.450 265.950 ;
        RECT 880.950 251.400 885.450 252.450 ;
        RECT 880.950 250.950 883.050 251.400 ;
        RECT 877.950 220.950 880.050 223.050 ;
        RECT 865.950 217.950 868.050 220.050 ;
        RECT 866.400 208.050 867.450 217.950 ;
        RECT 871.950 216.000 874.050 220.050 ;
        RECT 878.400 216.600 879.450 220.950 ;
        RECT 872.400 214.350 873.600 216.000 ;
        RECT 878.400 214.350 879.600 216.600 ;
        RECT 871.950 211.950 874.050 214.050 ;
        RECT 874.950 211.950 877.050 214.050 ;
        RECT 877.950 211.950 880.050 214.050 ;
        RECT 875.400 209.400 876.600 211.650 ;
        RECT 859.950 205.950 862.050 208.050 ;
        RECT 865.950 205.950 868.050 208.050 ;
        RECT 875.400 205.050 876.450 209.400 ;
        RECT 841.950 202.950 844.050 205.050 ;
        RECT 874.950 202.950 877.050 205.050 ;
        RECT 836.400 188.400 840.450 189.450 ;
        RECT 829.950 184.950 832.050 187.050 ;
        RECT 817.950 181.950 820.050 184.050 ;
        RECT 820.950 181.950 823.050 184.050 ;
        RECT 826.950 182.100 829.050 184.200 ;
        RECT 818.400 177.900 819.450 181.950 ;
        RECT 827.400 181.350 828.600 182.100 ;
        RECT 832.950 181.950 835.050 187.050 ;
        RECT 823.950 178.950 826.050 181.050 ;
        RECT 826.950 178.950 829.050 181.050 ;
        RECT 829.950 178.950 832.050 181.050 ;
        RECT 817.950 175.800 820.050 177.900 ;
        RECT 820.950 175.950 823.050 178.050 ;
        RECT 824.400 177.000 825.600 178.650 ;
        RECT 830.400 177.900 831.600 178.650 ;
        RECT 814.950 172.950 817.050 175.050 ;
        RECT 808.950 163.950 811.050 166.050 ;
        RECT 793.950 157.950 796.050 160.050 ;
        RECT 787.950 148.950 790.050 151.050 ;
        RECT 781.950 139.950 784.050 142.050 ;
        RECT 790.950 139.950 793.050 145.050 ;
        RECT 782.400 133.050 783.450 139.950 ;
        RECT 787.950 137.100 790.050 139.200 ;
        RECT 794.400 138.600 795.450 157.950 ;
        RECT 808.950 148.950 811.050 151.050 ;
        RECT 788.400 136.350 789.600 137.100 ;
        RECT 794.400 136.350 795.600 138.600 ;
        RECT 800.400 138.450 801.600 138.600 ;
        RECT 800.400 137.400 807.450 138.450 ;
        RECT 800.400 136.350 801.600 137.400 ;
        RECT 787.950 133.950 790.050 136.050 ;
        RECT 790.950 133.950 793.050 136.050 ;
        RECT 793.950 133.950 796.050 136.050 ;
        RECT 796.950 133.950 799.050 136.050 ;
        RECT 799.950 133.950 802.050 136.050 ;
        RECT 781.950 130.950 784.050 133.050 ;
        RECT 791.400 132.000 792.600 133.650 ;
        RECT 797.400 132.000 798.600 133.650 ;
        RECT 757.950 124.950 760.050 127.050 ;
        RECT 769.950 124.950 772.050 127.050 ;
        RECT 778.950 124.950 781.050 127.050 ;
        RECT 754.950 109.950 757.050 112.050 ;
        RECT 752.400 107.400 756.450 108.450 ;
        RECT 716.400 103.350 717.600 104.100 ;
        RECT 722.400 103.350 723.600 105.600 ;
        RECT 736.950 104.100 739.050 106.200 ;
        RECT 748.950 104.100 751.050 106.200 ;
        RECT 755.400 105.600 756.450 107.400 ;
        RECT 737.400 103.350 738.600 104.100 ;
        RECT 712.950 100.950 715.050 103.050 ;
        RECT 715.950 100.950 718.050 103.050 ;
        RECT 718.950 100.950 721.050 103.050 ;
        RECT 721.950 100.950 724.050 103.050 ;
        RECT 736.950 100.950 739.050 103.050 ;
        RECT 739.950 100.950 742.050 103.050 ;
        RECT 706.950 97.950 709.050 100.050 ;
        RECT 713.400 98.400 714.600 100.650 ;
        RECT 719.400 99.900 720.600 100.650 ;
        RECT 713.400 91.050 714.450 98.400 ;
        RECT 718.950 97.800 721.050 99.900 ;
        RECT 740.400 99.000 741.600 100.650 ;
        RECT 719.400 96.450 720.450 97.800 ;
        RECT 719.400 95.400 723.450 96.450 ;
        RECT 703.950 88.950 706.050 91.050 ;
        RECT 712.950 88.950 715.050 91.050 ;
        RECT 715.950 85.950 718.050 88.050 ;
        RECT 706.950 76.950 709.050 79.050 ;
        RECT 694.950 59.100 697.050 61.200 ;
        RECT 700.950 59.100 703.050 61.200 ;
        RECT 707.400 60.600 708.450 76.950 ;
        RECT 695.400 55.050 696.450 59.100 ;
        RECT 701.400 58.350 702.600 59.100 ;
        RECT 707.400 58.350 708.600 60.600 ;
        RECT 700.950 55.950 703.050 58.050 ;
        RECT 703.950 55.950 706.050 58.050 ;
        RECT 706.950 55.950 709.050 58.050 ;
        RECT 709.950 55.950 712.050 58.050 ;
        RECT 694.950 52.950 697.050 55.050 ;
        RECT 704.400 53.400 705.600 55.650 ;
        RECT 710.400 54.900 711.600 55.650 ;
        RECT 716.400 55.050 717.450 85.950 ;
        RECT 718.950 61.950 721.050 64.050 ;
        RECT 691.950 49.950 694.050 52.050 ;
        RECT 700.950 49.950 703.050 52.050 ;
        RECT 655.950 46.950 658.050 49.050 ;
        RECT 667.950 46.950 670.050 49.050 ;
        RECT 701.400 46.050 702.450 49.950 ;
        RECT 704.400 49.050 705.450 53.400 ;
        RECT 709.950 52.800 712.050 54.900 ;
        RECT 715.950 52.950 718.050 55.050 ;
        RECT 719.400 52.050 720.450 61.950 ;
        RECT 722.400 61.050 723.450 95.400 ;
        RECT 739.950 94.950 742.050 99.000 ;
        RECT 749.400 88.050 750.450 104.100 ;
        RECT 755.400 103.350 756.600 105.600 ;
        RECT 760.950 104.100 763.050 106.200 ;
        RECT 761.400 103.350 762.600 104.100 ;
        RECT 754.950 100.950 757.050 103.050 ;
        RECT 757.950 100.950 760.050 103.050 ;
        RECT 760.950 100.950 763.050 103.050 ;
        RECT 763.950 100.950 766.050 103.050 ;
        RECT 758.400 98.400 759.600 100.650 ;
        RECT 764.400 99.000 765.600 100.650 ;
        RECT 758.400 91.050 759.450 98.400 ;
        RECT 763.950 94.950 766.050 99.000 ;
        RECT 757.950 88.950 760.050 91.050 ;
        RECT 748.950 85.950 751.050 88.050 ;
        RECT 724.950 76.950 727.050 79.050 ;
        RECT 721.950 58.950 724.050 61.050 ;
        RECT 725.400 60.600 726.450 76.950 ;
        RECT 758.400 76.050 759.450 88.950 ;
        RECT 757.950 73.950 760.050 76.050 ;
        RECT 763.950 73.950 766.050 76.050 ;
        RECT 739.950 70.950 742.050 73.050 ;
        RECT 725.400 58.350 726.600 60.600 ;
        RECT 730.950 60.000 733.050 64.050 ;
        RECT 731.400 58.350 732.600 60.000 ;
        RECT 724.950 55.950 727.050 58.050 ;
        RECT 727.950 55.950 730.050 58.050 ;
        RECT 730.950 55.950 733.050 58.050 ;
        RECT 733.950 55.950 736.050 58.050 ;
        RECT 728.400 54.000 729.600 55.650 ;
        RECT 734.400 54.900 735.600 55.650 ;
        RECT 740.400 54.900 741.450 70.950 ;
        RECT 757.950 64.950 760.050 67.050 ;
        RECT 751.950 60.000 754.050 64.050 ;
        RECT 758.400 61.200 759.450 64.950 ;
        RECT 752.400 58.350 753.600 60.000 ;
        RECT 757.950 59.100 760.050 61.200 ;
        RECT 758.400 58.350 759.600 59.100 ;
        RECT 748.950 55.950 751.050 58.050 ;
        RECT 751.950 55.950 754.050 58.050 ;
        RECT 754.950 55.950 757.050 58.050 ;
        RECT 757.950 55.950 760.050 58.050 ;
        RECT 749.400 54.900 750.600 55.650 ;
        RECT 755.400 54.900 756.600 55.650 ;
        RECT 764.400 55.050 765.450 73.950 ;
        RECT 770.400 66.450 771.450 124.950 ;
        RECT 778.950 118.950 781.050 121.050 ;
        RECT 779.400 105.600 780.450 118.950 ;
        RECT 782.400 109.050 783.450 130.950 ;
        RECT 790.950 127.950 793.050 132.000 ;
        RECT 796.950 127.950 799.050 132.000 ;
        RECT 806.400 129.450 807.450 137.400 ;
        RECT 809.400 133.050 810.450 148.950 ;
        RECT 817.950 142.950 820.050 145.050 ;
        RECT 818.400 138.600 819.450 142.950 ;
        RECT 821.400 142.050 822.450 175.950 ;
        RECT 823.950 172.950 826.050 177.000 ;
        RECT 829.950 175.800 832.050 177.900 ;
        RECT 829.950 148.950 832.050 151.050 ;
        RECT 820.950 139.950 823.050 142.050 ;
        RECT 818.400 136.350 819.600 138.600 ;
        RECT 823.950 137.100 826.050 139.200 ;
        RECT 824.400 136.350 825.600 137.100 ;
        RECT 814.950 133.950 817.050 136.050 ;
        RECT 817.950 133.950 820.050 136.050 ;
        RECT 820.950 133.950 823.050 136.050 ;
        RECT 823.950 133.950 826.050 136.050 ;
        RECT 808.950 130.950 811.050 133.050 ;
        RECT 815.400 132.900 816.600 133.650 ;
        RECT 821.400 132.900 822.600 133.650 ;
        RECT 814.950 130.800 817.050 132.900 ;
        RECT 820.950 130.800 823.050 132.900 ;
        RECT 826.950 130.800 829.050 132.900 ;
        RECT 806.400 128.400 810.450 129.450 ;
        RECT 802.950 124.950 805.050 127.050 ;
        RECT 803.400 112.050 804.450 124.950 ;
        RECT 809.400 121.050 810.450 128.400 ;
        RECT 817.950 127.950 820.050 130.050 ;
        RECT 808.950 118.950 811.050 121.050 ;
        RECT 784.950 109.050 787.050 112.050 ;
        RECT 802.950 109.950 805.050 112.050 ;
        RECT 781.950 106.950 784.050 109.050 ;
        RECT 784.950 108.000 790.050 109.050 ;
        RECT 785.400 107.400 790.050 108.000 ;
        RECT 786.000 106.950 790.050 107.400 ;
        RECT 793.950 106.950 796.050 109.050 ;
        RECT 779.400 103.350 780.600 105.600 ;
        RECT 784.950 104.100 787.050 106.200 ;
        RECT 785.400 103.350 786.600 104.100 ;
        RECT 778.950 100.950 781.050 103.050 ;
        RECT 781.950 100.950 784.050 103.050 ;
        RECT 784.950 100.950 787.050 103.050 ;
        RECT 787.950 100.950 790.050 103.050 ;
        RECT 782.400 99.000 783.600 100.650 ;
        RECT 781.950 94.950 784.050 99.000 ;
        RECT 788.400 98.400 789.600 100.650 ;
        RECT 788.400 91.050 789.450 98.400 ;
        RECT 787.950 88.950 790.050 91.050 ;
        RECT 772.950 73.950 775.050 76.050 ;
        RECT 767.400 65.400 771.450 66.450 ;
        RECT 718.950 49.950 721.050 52.050 ;
        RECT 727.950 49.950 730.050 54.000 ;
        RECT 733.950 52.800 736.050 54.900 ;
        RECT 739.950 52.800 742.050 54.900 ;
        RECT 748.950 52.800 751.050 54.900 ;
        RECT 754.950 52.800 757.050 54.900 ;
        RECT 763.950 52.950 766.050 55.050 ;
        RECT 767.400 52.050 768.450 65.400 ;
        RECT 773.400 60.600 774.450 73.950 ;
        RECT 794.400 61.200 795.450 106.950 ;
        RECT 796.950 103.950 799.050 106.050 ;
        RECT 802.950 104.100 805.050 106.200 ;
        RECT 809.400 105.600 810.450 118.950 ;
        RECT 797.400 79.050 798.450 103.950 ;
        RECT 803.400 103.350 804.600 104.100 ;
        RECT 809.400 103.350 810.600 105.600 ;
        RECT 802.950 100.950 805.050 103.050 ;
        RECT 805.950 100.950 808.050 103.050 ;
        RECT 808.950 100.950 811.050 103.050 ;
        RECT 811.950 100.950 814.050 103.050 ;
        RECT 806.400 98.400 807.600 100.650 ;
        RECT 812.400 100.050 813.600 100.650 ;
        RECT 812.400 98.400 817.050 100.050 ;
        RECT 796.950 76.950 799.050 79.050 ;
        RECT 806.400 64.050 807.450 98.400 ;
        RECT 813.000 97.950 817.050 98.400 ;
        RECT 818.400 76.050 819.450 127.950 ;
        RECT 820.950 127.650 823.050 129.750 ;
        RECT 817.950 73.950 820.050 76.050 ;
        RECT 773.400 58.350 774.600 60.600 ;
        RECT 778.950 59.100 781.050 61.200 ;
        RECT 793.950 60.450 796.050 61.200 ;
        RECT 797.400 60.450 798.600 60.600 ;
        RECT 793.950 59.400 798.600 60.450 ;
        RECT 802.950 60.000 805.050 64.050 ;
        RECT 805.950 61.950 808.050 64.050 ;
        RECT 811.950 61.950 814.050 64.050 ;
        RECT 793.950 59.100 796.050 59.400 ;
        RECT 779.400 58.350 780.600 59.100 ;
        RECT 797.400 58.350 798.600 59.400 ;
        RECT 803.400 58.350 804.600 60.000 ;
        RECT 772.950 55.950 775.050 58.050 ;
        RECT 775.950 55.950 778.050 58.050 ;
        RECT 778.950 55.950 781.050 58.050 ;
        RECT 781.950 55.950 784.050 58.050 ;
        RECT 796.950 55.950 799.050 58.050 ;
        RECT 799.950 55.950 802.050 58.050 ;
        RECT 802.950 55.950 805.050 58.050 ;
        RECT 805.950 55.950 808.050 58.050 ;
        RECT 776.400 54.900 777.600 55.650 ;
        RECT 782.400 54.900 783.600 55.650 ;
        RECT 775.950 52.800 778.050 54.900 ;
        RECT 781.950 52.800 784.050 54.900 ;
        RECT 800.400 54.000 801.600 55.650 ;
        RECT 806.400 54.900 807.600 55.650 ;
        RECT 766.950 49.950 769.050 52.050 ;
        RECT 799.950 49.950 802.050 54.000 ;
        RECT 805.950 52.800 808.050 54.900 ;
        RECT 703.950 46.950 706.050 49.050 ;
        RECT 646.950 43.950 649.050 46.050 ;
        RECT 652.950 45.450 655.050 46.050 ;
        RECT 658.950 45.450 661.050 46.050 ;
        RECT 652.950 44.400 661.050 45.450 ;
        RECT 652.950 43.950 655.050 44.400 ;
        RECT 658.950 43.950 661.050 44.400 ;
        RECT 700.950 43.950 703.050 46.050 ;
        RECT 812.400 43.050 813.450 61.950 ;
        RECT 821.400 61.050 822.450 127.650 ;
        RECT 827.400 127.050 828.450 130.800 ;
        RECT 826.950 124.950 829.050 127.050 ;
        RECT 830.400 115.050 831.450 148.950 ;
        RECT 832.950 142.950 835.050 145.050 ;
        RECT 829.950 112.950 832.050 115.050 ;
        RECT 833.400 112.050 834.450 142.950 ;
        RECT 836.400 139.200 837.450 188.400 ;
        RECT 847.950 187.950 850.050 190.050 ;
        RECT 856.950 187.950 859.050 190.050 ;
        RECT 871.950 187.950 874.050 190.050 ;
        RECT 838.950 184.950 841.050 187.050 ;
        RECT 839.400 151.050 840.450 184.950 ;
        RECT 848.400 183.600 849.450 187.950 ;
        RECT 857.400 184.050 858.450 187.950 ;
        RECT 872.400 187.200 873.600 187.950 ;
        RECT 868.500 185.100 870.600 187.200 ;
        RECT 848.400 181.350 849.600 183.600 ;
        RECT 856.950 181.950 859.050 184.050 ;
        RECT 859.950 181.950 862.050 184.050 ;
        RECT 844.950 178.950 847.050 181.050 ;
        RECT 847.950 178.950 850.050 181.050 ;
        RECT 850.950 178.950 853.050 181.050 ;
        RECT 856.950 178.800 859.050 180.900 ;
        RECT 841.950 175.950 844.050 178.050 ;
        RECT 845.400 176.400 846.600 178.650 ;
        RECT 842.400 151.050 843.450 175.950 ;
        RECT 845.400 169.050 846.450 176.400 ;
        RECT 853.950 175.950 856.050 178.050 ;
        RECT 844.950 166.950 847.050 169.050 ;
        RECT 854.400 166.050 855.450 175.950 ;
        RECT 853.950 163.950 856.050 166.050 ;
        RECT 838.800 148.950 840.900 151.050 ;
        RECT 841.950 148.950 844.050 151.050 ;
        RECT 857.400 142.050 858.450 178.800 ;
        RECT 860.400 169.050 861.450 181.950 ;
        RECT 866.100 178.950 868.200 181.050 ;
        RECT 869.100 180.000 870.000 185.100 ;
        RECT 871.800 184.800 873.900 186.900 ;
        RECT 878.400 185.400 880.500 187.500 ;
        RECT 876.000 183.000 878.100 183.900 ;
        RECT 870.900 181.800 878.100 183.000 ;
        RECT 870.900 180.900 873.000 181.800 ;
        RECT 876.000 180.000 878.100 180.900 ;
        RECT 869.100 179.100 878.100 180.000 ;
        RECT 869.100 172.500 870.000 179.100 ;
        RECT 876.000 178.800 878.100 179.100 ;
        RECT 871.800 175.950 873.900 178.050 ;
        RECT 872.400 173.400 873.600 175.650 ;
        RECT 879.000 172.800 879.900 185.400 ;
        RECT 880.800 178.950 882.900 181.050 ;
        RECT 881.400 177.450 882.600 178.650 ;
        RECT 884.400 177.450 885.450 251.400 ;
        RECT 889.950 250.950 892.050 253.050 ;
        RECT 881.400 176.400 885.450 177.450 ;
        RECT 869.100 170.400 871.200 172.500 ;
        RECT 878.100 170.700 880.200 172.800 ;
        RECT 859.950 166.950 862.050 169.050 ;
        RECT 893.400 166.050 894.450 295.800 ;
        RECT 874.950 163.950 877.050 166.050 ;
        RECT 892.950 163.950 895.050 166.050 ;
        RECT 862.950 148.950 865.050 151.050 ;
        RECT 835.950 137.100 838.050 139.200 ;
        RECT 841.950 137.100 844.050 142.050 ;
        RECT 847.950 138.000 850.050 142.050 ;
        RECT 853.950 139.950 856.050 142.050 ;
        RECT 856.950 139.950 859.050 142.050 ;
        RECT 842.400 136.350 843.600 137.100 ;
        RECT 848.400 136.350 849.600 138.000 ;
        RECT 838.950 133.950 841.050 136.050 ;
        RECT 841.950 133.950 844.050 136.050 ;
        RECT 844.950 133.950 847.050 136.050 ;
        RECT 847.950 133.950 850.050 136.050 ;
        RECT 839.400 131.400 840.600 133.650 ;
        RECT 845.400 131.400 846.600 133.650 ;
        RECT 839.400 127.050 840.450 131.400 ;
        RECT 838.950 124.950 841.050 127.050 ;
        RECT 845.400 124.050 846.450 131.400 ;
        RECT 850.950 130.950 853.050 133.050 ;
        RECT 844.950 121.950 847.050 124.050 ;
        RECT 838.950 118.950 841.050 121.050 ;
        RECT 826.950 109.950 829.050 112.050 ;
        RECT 832.950 109.950 835.050 112.050 ;
        RECT 827.400 105.600 828.450 109.950 ;
        RECT 827.400 103.350 828.600 105.600 ;
        RECT 832.950 104.100 835.050 106.200 ;
        RECT 839.400 106.050 840.450 118.950 ;
        RECT 844.950 112.950 847.050 115.050 ;
        RECT 841.950 109.950 844.050 112.050 ;
        RECT 833.400 103.350 834.600 104.100 ;
        RECT 838.950 103.950 841.050 106.050 ;
        RECT 826.950 100.950 829.050 103.050 ;
        RECT 829.950 100.950 832.050 103.050 ;
        RECT 832.950 100.950 835.050 103.050 ;
        RECT 835.950 100.950 838.050 103.050 ;
        RECT 830.400 99.900 831.600 100.650 ;
        RECT 829.950 97.800 832.050 99.900 ;
        RECT 836.400 99.450 837.600 100.650 ;
        RECT 836.400 98.400 840.450 99.450 ;
        RECT 839.400 76.050 840.450 98.400 ;
        RECT 838.950 73.950 841.050 76.050 ;
        RECT 826.950 67.950 829.050 70.050 ;
        RECT 814.950 58.950 817.050 61.050 ;
        RECT 820.950 58.950 823.050 61.050 ;
        RECT 827.400 60.600 828.450 67.950 ;
        RECT 811.950 40.950 814.050 43.050 ;
        RECT 643.950 37.950 646.050 40.050 ;
        RECT 673.950 37.950 676.050 40.050 ;
        RECT 628.800 30.300 630.900 32.400 ;
        RECT 632.400 31.200 633.600 33.450 ;
        RECT 640.950 31.950 643.050 34.050 ;
        RECT 566.400 25.350 567.600 26.100 ;
        RECT 562.950 22.950 565.050 25.050 ;
        RECT 565.950 22.950 568.050 25.050 ;
        RECT 538.950 16.950 541.050 21.000 ;
        RECT 544.950 19.800 547.050 21.900 ;
        RECT 556.950 19.950 559.050 22.050 ;
        RECT 563.400 21.000 564.600 22.650 ;
        RECT 562.950 16.950 565.050 21.000 ;
        RECT 520.950 7.950 523.050 10.050 ;
        RECT 572.400 7.050 573.450 26.100 ;
        RECT 584.400 25.350 585.600 27.600 ;
        RECT 590.400 25.350 591.600 27.600 ;
        RECT 598.950 25.950 601.050 28.050 ;
        RECT 607.950 26.100 610.050 28.200 ;
        RECT 626.400 27.450 627.600 27.600 ;
        RECT 623.400 27.000 627.600 27.450 ;
        RECT 622.950 26.400 627.600 27.000 ;
        RECT 580.950 22.950 583.050 25.050 ;
        RECT 583.950 22.950 586.050 25.050 ;
        RECT 586.950 22.950 589.050 25.050 ;
        RECT 589.950 22.950 592.050 25.050 ;
        RECT 595.950 22.950 598.050 25.050 ;
        RECT 581.400 20.400 582.600 22.650 ;
        RECT 587.400 21.900 588.600 22.650 ;
        RECT 581.400 7.050 582.450 20.400 ;
        RECT 586.950 19.800 589.050 21.900 ;
        RECT 592.950 16.950 595.050 19.050 ;
        RECT 593.400 10.050 594.450 16.950 ;
        RECT 596.400 16.050 597.450 22.950 ;
        RECT 595.950 13.950 598.050 16.050 ;
        RECT 592.950 7.950 595.050 10.050 ;
        RECT 599.400 7.050 600.450 25.950 ;
        RECT 608.400 25.350 609.600 26.100 ;
        RECT 604.950 22.950 607.050 25.050 ;
        RECT 607.950 22.950 610.050 25.050 ;
        RECT 610.950 22.950 613.050 25.050 ;
        RECT 622.950 22.950 625.050 26.400 ;
        RECT 626.400 25.350 627.600 26.400 ;
        RECT 626.100 22.950 628.200 25.050 ;
        RECT 629.100 24.900 630.000 30.300 ;
        RECT 632.100 28.800 634.200 30.900 ;
        RECT 636.000 27.900 638.100 29.700 ;
        RECT 630.900 26.700 639.600 27.900 ;
        RECT 630.900 25.800 633.000 26.700 ;
        RECT 629.100 23.700 636.000 24.900 ;
        RECT 605.400 21.000 606.600 22.650 ;
        RECT 611.400 21.000 612.600 22.650 ;
        RECT 604.950 16.950 607.050 21.000 ;
        RECT 610.950 16.950 613.050 21.000 ;
        RECT 605.400 10.050 606.450 16.950 ;
        RECT 629.100 16.500 630.300 23.700 ;
        RECT 632.100 19.950 634.200 22.050 ;
        RECT 635.100 21.300 636.000 23.700 ;
        RECT 632.400 17.400 633.600 19.650 ;
        RECT 635.100 19.200 637.200 21.300 ;
        RECT 638.700 17.700 639.600 26.700 ;
        RECT 658.950 26.100 661.050 28.200 ;
        RECT 659.400 25.350 660.600 26.100 ;
        RECT 670.950 25.950 673.050 28.050 ;
        RECT 640.800 22.950 642.900 25.050 ;
        RECT 655.950 22.950 658.050 25.050 ;
        RECT 658.950 22.950 661.050 25.050 ;
        RECT 661.950 22.950 664.050 25.050 ;
        RECT 641.400 21.450 642.600 22.650 ;
        RECT 656.400 21.900 657.600 22.650 ;
        RECT 641.400 21.000 645.450 21.450 ;
        RECT 641.400 20.400 646.050 21.000 ;
        RECT 628.800 14.400 630.900 16.500 ;
        RECT 638.400 15.600 640.500 17.700 ;
        RECT 643.950 16.950 646.050 20.400 ;
        RECT 655.950 19.800 658.050 21.900 ;
        RECT 662.400 20.400 663.600 22.650 ;
        RECT 671.400 21.900 672.450 25.950 ;
        RECT 662.400 19.050 663.450 20.400 ;
        RECT 670.950 19.800 673.050 21.900 ;
        RECT 661.950 16.950 664.050 19.050 ;
        RECT 662.400 13.050 663.450 16.950 ;
        RECT 674.400 16.050 675.450 37.950 ;
        RECT 682.950 34.950 685.050 37.050 ;
        RECT 676.950 31.950 679.050 34.050 ;
        RECT 677.400 28.050 678.450 31.950 ;
        RECT 676.950 25.950 679.050 28.050 ;
        RECT 683.400 27.600 684.450 34.950 ;
        RECT 695.850 33.300 697.950 35.400 ;
        RECT 713.550 33.300 715.650 35.400 ;
        RECT 731.850 33.300 733.950 35.400 ;
        RECT 749.550 33.300 751.650 35.400 ;
        RECT 683.400 25.350 684.600 27.600 ;
        RECT 679.950 22.950 682.050 25.050 ;
        RECT 682.950 22.950 685.050 25.050 ;
        RECT 685.950 22.950 688.050 25.050 ;
        RECT 691.950 22.950 694.050 25.050 ;
        RECT 680.400 21.900 681.600 22.650 ;
        RECT 679.950 19.800 682.050 21.900 ;
        RECT 686.400 20.400 687.600 22.650 ;
        RECT 692.400 20.400 693.600 22.650 ;
        RECT 673.950 13.950 676.050 16.050 ;
        RECT 661.950 10.950 664.050 13.050 ;
        RECT 604.950 7.950 607.050 10.050 ;
        RECT 658.950 9.450 661.050 10.050 ;
        RECT 664.950 9.450 667.050 10.050 ;
        RECT 658.950 8.400 667.050 9.450 ;
        RECT 658.950 7.950 661.050 8.400 ;
        RECT 664.950 7.950 667.050 8.400 ;
        RECT 686.400 7.050 687.450 20.400 ;
        RECT 692.400 16.050 693.450 20.400 ;
        RECT 691.950 13.950 694.050 16.050 ;
        RECT 696.150 14.700 697.350 33.300 ;
        RECT 706.950 25.950 709.050 28.050 ;
        RECT 701.100 22.950 703.200 25.050 ;
        RECT 701.400 21.900 702.600 22.650 ;
        RECT 707.400 21.900 708.450 25.950 ;
        RECT 700.950 19.800 703.050 21.900 ;
        RECT 706.950 19.800 709.050 21.900 ;
        RECT 713.550 20.400 714.750 33.300 ;
        RECT 718.950 26.100 721.050 28.200 ;
        RECT 719.400 25.350 720.600 26.100 ;
        RECT 718.950 22.950 721.050 25.050 ;
        RECT 727.950 22.950 730.050 25.050 ;
        RECT 728.400 20.400 729.600 22.650 ;
        RECT 713.550 18.300 715.650 20.400 ;
        RECT 696.150 13.500 700.350 14.700 ;
        RECT 698.250 12.600 700.350 13.500 ;
        RECT 713.550 11.700 714.750 18.300 ;
        RECT 728.400 16.050 729.450 20.400 ;
        RECT 727.950 13.950 730.050 16.050 ;
        RECT 732.150 14.700 733.350 33.300 ;
        RECT 737.100 22.950 739.200 25.050 ;
        RECT 737.400 21.900 738.600 22.650 ;
        RECT 736.950 19.800 739.050 21.900 ;
        RECT 749.550 20.400 750.750 33.300 ;
        RECT 799.950 31.950 802.050 34.050 ;
        RECT 754.950 26.100 757.050 28.200 ;
        RECT 772.950 26.100 775.050 28.200 ;
        RECT 755.400 25.350 756.600 26.100 ;
        RECT 773.400 25.350 774.600 26.100 ;
        RECT 781.950 25.950 784.050 28.050 ;
        RECT 793.950 26.100 796.050 28.200 ;
        RECT 800.400 27.600 801.450 31.950 ;
        RECT 754.950 22.950 757.050 25.050 ;
        RECT 773.400 22.950 775.500 25.050 ;
        RECT 778.800 22.950 780.900 25.050 ;
        RECT 749.550 18.300 751.650 20.400 ;
        RECT 732.150 13.500 736.350 14.700 ;
        RECT 734.250 12.600 736.350 13.500 ;
        RECT 749.550 11.700 750.750 18.300 ;
        RECT 713.550 9.600 715.650 11.700 ;
        RECT 749.550 9.600 751.650 11.700 ;
        RECT 782.400 7.050 783.450 25.950 ;
        RECT 794.400 25.350 795.600 26.100 ;
        RECT 800.400 25.350 801.600 27.600 ;
        RECT 808.950 25.950 811.050 28.050 ;
        RECT 815.400 27.450 816.450 58.950 ;
        RECT 827.400 58.350 828.600 60.600 ;
        RECT 832.950 59.100 835.050 61.200 ;
        RECT 833.400 58.350 834.600 59.100 ;
        RECT 823.950 55.950 826.050 58.050 ;
        RECT 826.950 55.950 829.050 58.050 ;
        RECT 829.950 55.950 832.050 58.050 ;
        RECT 832.950 55.950 835.050 58.050 ;
        RECT 824.400 54.900 825.600 55.650 ;
        RECT 830.400 54.900 831.600 55.650 ;
        RECT 823.950 52.800 826.050 54.900 ;
        RECT 829.950 52.800 832.050 54.900 ;
        RECT 839.400 52.050 840.450 73.950 ;
        RECT 842.400 61.200 843.450 109.950 ;
        RECT 845.400 99.900 846.450 112.950 ;
        RECT 851.400 111.450 852.450 130.950 ;
        RECT 854.400 115.050 855.450 139.950 ;
        RECT 863.400 138.600 864.450 148.950 ;
        RECT 863.400 136.350 864.600 138.600 ;
        RECT 868.950 137.100 871.050 139.200 ;
        RECT 869.400 136.350 870.600 137.100 ;
        RECT 862.950 133.950 865.050 136.050 ;
        RECT 865.950 133.950 868.050 136.050 ;
        RECT 868.950 133.950 871.050 136.050 ;
        RECT 866.400 131.400 867.600 133.650 ;
        RECT 875.400 132.900 876.450 163.950 ;
        RECT 889.950 137.100 892.050 139.200 ;
        RECT 890.400 136.350 891.600 137.100 ;
        RECT 886.950 133.950 889.050 136.050 ;
        RECT 889.950 133.950 892.050 136.050 ;
        RECT 887.400 132.900 888.600 133.650 ;
        RECT 866.400 124.050 867.450 131.400 ;
        RECT 874.950 130.800 877.050 132.900 ;
        RECT 886.950 130.800 889.050 132.900 ;
        RECT 865.950 123.450 868.050 124.050 ;
        RECT 863.400 122.400 868.050 123.450 ;
        RECT 853.950 112.950 856.050 115.050 ;
        RECT 851.400 110.400 855.450 111.450 ;
        RECT 854.400 105.600 855.450 110.400 ;
        RECT 854.400 103.350 855.600 105.600 ;
        RECT 863.400 103.050 864.450 122.400 ;
        RECT 865.950 121.950 868.050 122.400 ;
        RECT 865.950 112.950 868.050 115.050 ;
        RECT 850.950 100.950 853.050 103.050 ;
        RECT 853.950 100.950 856.050 103.050 ;
        RECT 856.950 100.950 859.050 103.050 ;
        RECT 862.950 100.950 865.050 103.050 ;
        RECT 851.400 99.900 852.600 100.650 ;
        RECT 844.950 97.800 847.050 99.900 ;
        RECT 850.950 97.800 853.050 99.900 ;
        RECT 857.400 98.400 858.600 100.650 ;
        RECT 851.400 70.050 852.450 97.800 ;
        RECT 857.400 82.050 858.450 98.400 ;
        RECT 859.950 97.950 862.050 100.050 ;
        RECT 866.400 99.900 867.450 112.950 ;
        RECT 874.950 104.100 877.050 106.200 ;
        RECT 875.400 103.350 876.600 104.100 ;
        RECT 871.950 100.950 874.050 103.050 ;
        RECT 874.950 100.950 877.050 103.050 ;
        RECT 877.950 100.950 880.050 103.050 ;
        RECT 872.400 99.900 873.600 100.650 ;
        RECT 865.950 99.450 868.050 99.900 ;
        RECT 863.400 98.400 868.050 99.450 ;
        RECT 856.950 79.950 859.050 82.050 ;
        RECT 850.950 67.950 853.050 70.050 ;
        RECT 856.950 67.950 859.050 70.050 ;
        RECT 841.950 59.100 844.050 61.200 ;
        RECT 851.400 60.600 852.450 67.950 ;
        RECT 857.400 64.050 858.450 67.950 ;
        RECT 838.950 49.950 841.050 52.050 ;
        RECT 842.400 34.050 843.450 59.100 ;
        RECT 851.400 58.350 852.600 60.600 ;
        RECT 856.950 60.000 859.050 64.050 ;
        RECT 860.400 61.200 861.450 97.950 ;
        RECT 857.400 58.350 858.600 60.000 ;
        RECT 859.950 59.100 862.050 61.200 ;
        RECT 847.950 55.950 850.050 58.050 ;
        RECT 850.950 55.950 853.050 58.050 ;
        RECT 853.950 55.950 856.050 58.050 ;
        RECT 856.950 55.950 859.050 58.050 ;
        RECT 848.400 54.000 849.600 55.650 ;
        RECT 854.400 54.900 855.600 55.650 ;
        RECT 847.950 49.950 850.050 54.000 ;
        RECT 853.950 52.800 856.050 54.900 ;
        RECT 844.950 43.950 847.050 46.050 ;
        RECT 829.950 31.950 832.050 34.050 ;
        RECT 841.950 31.950 844.050 34.050 ;
        RECT 812.400 26.400 816.450 27.450 ;
        RECT 793.950 22.950 796.050 25.050 ;
        RECT 796.950 22.950 799.050 25.050 ;
        RECT 799.950 22.950 802.050 25.050 ;
        RECT 802.950 22.950 805.050 25.050 ;
        RECT 797.400 20.400 798.600 22.650 ;
        RECT 803.400 21.900 804.600 22.650 ;
        RECT 797.400 10.050 798.450 20.400 ;
        RECT 802.950 19.800 805.050 21.900 ;
        RECT 809.400 13.050 810.450 25.950 ;
        RECT 812.400 21.900 813.450 26.400 ;
        RECT 820.950 26.100 823.050 28.200 ;
        RECT 821.400 25.350 822.600 26.100 ;
        RECT 817.950 22.950 820.050 25.050 ;
        RECT 820.950 22.950 823.050 25.050 ;
        RECT 823.950 22.950 826.050 25.050 ;
        RECT 811.950 19.800 814.050 21.900 ;
        RECT 818.400 21.000 819.600 22.650 ;
        RECT 812.400 16.050 813.450 19.800 ;
        RECT 817.950 16.950 820.050 21.000 ;
        RECT 824.400 20.400 825.600 22.650 ;
        RECT 824.400 18.450 825.450 20.400 ;
        RECT 830.400 19.050 831.450 31.950 ;
        RECT 845.400 30.450 846.450 43.950 ;
        RECT 850.950 40.950 853.050 43.050 ;
        RECT 842.400 29.400 846.450 30.450 ;
        RECT 842.400 27.600 843.450 29.400 ;
        RECT 842.400 25.350 843.600 27.600 ;
        RECT 838.950 22.950 841.050 25.050 ;
        RECT 841.950 22.950 844.050 25.050 ;
        RECT 844.950 22.950 847.050 25.050 ;
        RECT 845.400 21.000 846.600 22.650 ;
        RECT 851.400 22.050 852.450 40.950 ;
        RECT 863.400 30.450 864.450 98.400 ;
        RECT 865.950 97.800 868.050 98.400 ;
        RECT 871.950 97.800 874.050 99.900 ;
        RECT 878.400 98.400 879.600 100.650 ;
        RECT 878.400 82.050 879.450 98.400 ;
        RECT 865.950 79.950 868.050 82.050 ;
        RECT 877.950 79.950 880.050 82.050 ;
        RECT 866.400 37.050 867.450 79.950 ;
        RECT 880.950 67.950 883.050 70.050 ;
        RECT 874.950 59.100 877.050 61.200 ;
        RECT 881.400 60.600 882.450 67.950 ;
        RECT 875.400 58.350 876.600 59.100 ;
        RECT 881.400 58.350 882.600 60.600 ;
        RECT 874.950 55.950 877.050 58.050 ;
        RECT 877.950 55.950 880.050 58.050 ;
        RECT 880.950 55.950 883.050 58.050 ;
        RECT 878.400 53.400 879.600 55.650 ;
        RECT 878.400 37.050 879.450 53.400 ;
        RECT 896.400 46.050 897.450 296.400 ;
        RECT 898.950 274.950 901.050 277.050 ;
        RECT 899.400 184.050 900.450 274.950 ;
        RECT 898.950 181.950 901.050 184.050 ;
        RECT 898.950 163.950 901.050 166.050 ;
        RECT 895.950 43.950 898.050 46.050 ;
        RECT 865.950 34.950 868.050 37.050 ;
        RECT 877.950 34.950 880.050 37.050 ;
        RECT 860.400 29.400 864.450 30.450 ;
        RECT 860.400 27.600 861.450 29.400 ;
        RECT 866.400 27.600 867.450 34.950 ;
        RECT 860.400 25.350 861.600 27.600 ;
        RECT 866.400 25.350 867.600 27.600 ;
        RECT 859.950 22.950 862.050 25.050 ;
        RECT 862.950 22.950 865.050 25.050 ;
        RECT 865.950 22.950 868.050 25.050 ;
        RECT 881.100 22.950 883.200 25.050 ;
        RECT 886.500 22.950 888.600 25.050 ;
        RECT 821.400 17.400 825.450 18.450 ;
        RECT 821.400 16.050 822.450 17.400 ;
        RECT 829.950 16.950 832.050 19.050 ;
        RECT 844.950 16.950 847.050 21.000 ;
        RECT 850.950 19.950 853.050 22.050 ;
        RECT 863.400 21.900 864.600 22.650 ;
        RECT 862.950 19.800 865.050 21.900 ;
        RECT 881.400 21.000 882.600 22.650 ;
        RECT 880.950 16.950 883.050 21.000 ;
        RECT 899.400 19.050 900.450 163.950 ;
        RECT 898.950 16.950 901.050 19.050 ;
        RECT 811.950 13.950 814.050 16.050 ;
        RECT 819.000 15.900 822.450 16.050 ;
        RECT 817.950 14.400 822.450 15.900 ;
        RECT 817.950 13.950 822.000 14.400 ;
        RECT 817.950 13.800 820.050 13.950 ;
        RECT 808.950 10.950 811.050 13.050 ;
        RECT 796.950 7.950 799.050 10.050 ;
        RECT 571.950 4.950 574.050 7.050 ;
        RECT 580.950 4.950 583.050 7.050 ;
        RECT 598.950 4.950 601.050 7.050 ;
        RECT 685.950 4.950 688.050 7.050 ;
        RECT 781.950 4.950 784.050 7.050 ;
      LAYER via2 ;
        RECT 19.950 730.950 22.050 733.050 ;
        RECT 94.950 808.950 97.050 811.050 ;
        RECT 25.950 730.950 28.050 733.050 ;
        RECT 211.950 763.950 214.050 766.050 ;
        RECT 277.950 811.950 280.050 814.050 ;
        RECT 223.950 685.950 226.050 688.050 ;
        RECT 307.950 763.950 310.050 766.050 ;
        RECT 265.950 730.950 268.050 733.050 ;
        RECT 253.950 685.950 256.050 688.050 ;
        RECT 346.950 761.100 349.050 763.200 ;
        RECT 70.950 574.950 73.050 577.050 ;
        RECT 76.950 574.950 79.050 577.050 ;
        RECT 136.950 610.950 139.050 613.050 ;
        RECT 79.950 529.950 82.050 532.050 ;
        RECT 154.950 610.950 157.050 613.050 ;
        RECT 178.950 529.950 181.050 532.050 ;
        RECT 61.950 418.950 64.050 421.050 ;
        RECT 103.950 418.950 106.050 421.050 ;
        RECT 319.950 730.950 322.050 733.050 ;
        RECT 343.950 721.800 346.050 723.900 ;
        RECT 313.950 652.950 316.050 655.050 ;
        RECT 355.950 652.950 358.050 655.050 ;
        RECT 304.950 607.950 307.050 610.050 ;
        RECT 331.950 607.950 334.050 610.050 ;
        RECT 481.950 841.950 484.050 844.050 ;
        RECT 517.950 841.950 520.050 844.050 ;
        RECT 568.950 841.950 571.050 844.050 ;
        RECT 586.950 841.950 589.050 844.050 ;
        RECT 514.950 799.800 517.050 801.900 ;
        RECT 499.950 763.950 502.050 766.050 ;
        RECT 520.950 763.950 523.050 766.050 ;
        RECT 493.950 730.950 496.050 733.050 ;
        RECT 385.950 652.950 388.050 655.050 ;
        RECT 505.950 652.950 508.050 655.050 ;
        RECT 364.950 574.950 367.050 577.050 ;
        RECT 568.950 808.950 571.050 811.050 ;
        RECT 598.950 808.950 601.050 811.050 ;
        RECT 595.950 763.950 598.050 766.050 ;
        RECT 619.950 763.950 622.050 766.050 ;
        RECT 664.950 841.950 667.050 844.050 ;
        RECT 679.950 841.950 682.050 844.050 ;
        RECT 655.950 799.800 658.050 801.900 ;
        RECT 580.950 685.950 583.050 688.050 ;
        RECT 649.950 733.950 652.050 736.050 ;
        RECT 673.950 730.950 676.050 733.050 ;
        RECT 637.950 685.950 640.050 688.050 ;
        RECT 706.950 685.950 709.050 688.050 ;
        RECT 364.950 529.950 367.050 532.050 ;
        RECT 394.950 529.950 397.050 532.050 ;
        RECT 322.950 496.950 325.050 499.050 ;
        RECT 262.950 418.950 265.050 421.050 ;
        RECT 22.950 340.950 25.050 343.050 ;
        RECT 103.950 340.950 106.050 343.050 ;
        RECT 40.950 262.950 43.050 265.050 ;
        RECT 286.950 418.950 289.050 421.050 ;
        RECT 70.950 253.950 73.050 256.050 ;
        RECT 37.950 184.950 40.050 187.050 ;
        RECT 22.950 106.950 25.050 109.050 ;
        RECT 43.950 106.950 46.050 109.050 ;
        RECT 124.950 184.950 127.050 187.050 ;
        RECT 82.950 61.950 85.050 64.050 ;
        RECT 130.950 109.950 133.050 112.050 ;
        RECT 340.950 496.950 343.050 499.050 ;
        RECT 421.950 499.950 424.050 502.050 ;
        RECT 385.950 451.950 388.050 454.050 ;
        RECT 262.950 295.950 265.050 298.050 ;
        RECT 178.950 184.950 181.050 187.050 ;
        RECT 409.950 454.950 412.050 457.050 ;
        RECT 403.950 451.950 406.050 454.050 ;
        RECT 409.950 418.950 412.050 421.050 ;
        RECT 406.950 409.800 409.050 411.900 ;
        RECT 550.950 610.950 553.050 613.050 ;
        RECT 541.950 607.800 544.050 609.900 ;
        RECT 577.950 607.950 580.050 610.050 ;
        RECT 556.950 574.950 559.050 577.050 ;
        RECT 562.950 574.950 565.050 577.050 ;
        RECT 604.950 607.950 607.050 610.050 ;
        RECT 610.950 607.950 613.050 610.050 ;
        RECT 745.950 721.800 748.050 723.900 ;
        RECT 808.950 799.800 811.050 801.900 ;
        RECT 853.950 808.950 856.050 811.050 ;
        RECT 847.950 763.950 850.050 766.050 ;
        RECT 817.950 730.950 820.050 733.050 ;
        RECT 820.950 721.800 823.050 723.900 ;
        RECT 766.950 676.950 769.050 679.050 ;
        RECT 568.950 523.950 571.050 526.050 ;
        RECT 541.950 496.950 544.050 499.050 ;
        RECT 451.950 418.950 454.050 421.050 ;
        RECT 448.950 373.950 451.050 376.050 ;
        RECT 397.950 343.950 400.050 346.050 ;
        RECT 331.950 295.950 334.050 298.050 ;
        RECT 286.950 262.800 289.050 264.900 ;
        RECT 355.950 295.950 358.050 298.050 ;
        RECT 373.950 295.950 376.050 298.050 ;
        RECT 250.950 217.950 253.050 220.050 ;
        RECT 298.950 217.950 301.050 220.050 ;
        RECT 319.950 217.950 322.050 220.050 ;
        RECT 268.950 184.950 271.050 187.050 ;
        RECT 286.950 142.950 289.050 145.050 ;
        RECT 289.950 139.950 292.050 142.050 ;
        RECT 313.950 139.950 316.050 142.050 ;
        RECT 343.950 142.950 346.050 145.050 ;
        RECT 499.950 340.950 502.050 343.050 ;
        RECT 526.950 373.950 529.050 376.050 ;
        RECT 469.950 295.800 472.050 297.900 ;
        RECT 448.950 262.950 451.050 265.050 ;
        RECT 412.950 232.950 415.050 235.050 ;
        RECT 415.950 184.950 418.050 187.050 ;
        RECT 346.950 106.950 349.050 109.050 ;
        RECT 370.950 103.950 373.050 106.050 ;
        RECT 328.950 61.950 331.050 64.050 ;
        RECT 391.950 106.950 394.050 109.050 ;
        RECT 289.950 19.800 292.050 21.900 ;
        RECT 361.950 28.950 364.050 31.050 ;
        RECT 505.950 262.950 508.050 265.050 ;
        RECT 556.950 340.950 559.050 343.050 ;
        RECT 826.950 685.950 829.050 688.050 ;
        RECT 772.950 577.950 775.050 580.050 ;
        RECT 667.950 529.950 670.050 532.050 ;
        RECT 625.950 451.950 628.050 454.050 ;
        RECT 697.950 529.950 700.050 532.050 ;
        RECT 655.950 496.950 658.050 499.050 ;
        RECT 646.950 451.950 649.050 454.050 ;
        RECT 667.950 451.950 670.050 454.050 ;
        RECT 670.950 451.950 673.050 454.050 ;
        RECT 745.950 529.950 748.050 532.050 ;
        RECT 865.950 685.950 868.050 688.050 ;
        RECT 889.950 685.950 892.050 688.050 ;
        RECT 778.950 520.950 781.050 523.050 ;
        RECT 769.950 496.950 772.050 499.050 ;
        RECT 862.950 604.950 865.050 607.050 ;
        RECT 637.950 409.800 640.050 411.900 ;
        RECT 556.950 286.950 559.050 289.050 ;
        RECT 547.950 280.950 550.050 283.050 ;
        RECT 529.950 262.950 532.050 265.050 ;
        RECT 502.950 184.950 505.050 187.050 ;
        RECT 466.950 136.950 469.050 139.050 ;
        RECT 391.950 61.950 394.050 64.050 ;
        RECT 523.950 184.950 526.050 187.050 ;
        RECT 589.950 262.950 592.050 265.050 ;
        RECT 634.950 286.950 637.050 289.050 ;
        RECT 631.950 253.800 634.050 255.900 ;
        RECT 637.950 217.950 640.050 220.050 ;
        RECT 763.950 451.950 766.050 454.050 ;
        RECT 760.950 340.950 763.050 343.050 ;
        RECT 655.950 217.950 658.050 220.050 ;
        RECT 430.950 28.950 433.050 31.050 ;
        RECT 493.950 28.950 496.050 31.050 ;
        RECT 454.950 19.800 457.050 21.900 ;
        RECT 529.950 94.950 532.050 97.050 ;
        RECT 640.950 106.950 643.050 109.050 ;
        RECT 547.950 61.950 550.050 64.050 ;
        RECT 562.950 61.950 565.050 64.050 ;
        RECT 811.950 451.950 814.050 454.050 ;
        RECT 814.950 418.950 817.050 421.050 ;
        RECT 820.950 409.950 823.050 412.050 ;
        RECT 862.950 529.950 865.050 532.050 ;
        RECT 841.950 451.950 844.050 454.050 ;
        RECT 865.950 454.950 868.050 457.050 ;
        RECT 811.950 295.950 814.050 298.050 ;
        RECT 784.950 262.950 787.050 265.050 ;
        RECT 721.950 202.950 724.050 205.050 ;
        RECT 763.950 215.100 766.050 217.200 ;
        RECT 760.950 208.800 763.050 210.900 ;
        RECT 772.950 215.100 775.050 217.200 ;
        RECT 805.950 262.950 808.050 265.050 ;
        RECT 799.950 220.950 802.050 223.050 ;
        RECT 736.950 187.950 739.050 190.050 ;
        RECT 661.950 64.950 664.050 67.050 ;
        RECT 658.950 61.800 661.050 63.900 ;
        RECT 679.950 52.800 682.050 54.900 ;
        RECT 748.950 130.800 751.050 132.900 ;
        RECT 808.950 217.800 811.050 219.900 ;
        RECT 856.950 262.950 859.050 265.050 ;
        RECT 826.950 217.950 829.050 220.050 ;
        RECT 832.950 184.950 835.050 187.050 ;
        RECT 790.950 142.950 793.050 145.050 ;
        RECT 730.950 61.950 733.050 64.050 ;
        RECT 751.950 61.950 754.050 64.050 ;
        RECT 784.950 109.950 787.050 112.050 ;
        RECT 787.950 106.950 790.050 109.050 ;
        RECT 814.950 97.950 817.050 100.050 ;
        RECT 802.950 61.950 805.050 64.050 ;
        RECT 847.950 139.950 850.050 142.050 ;
        RECT 856.950 61.950 859.050 64.050 ;
      LAYER metal3 ;
        RECT 709.950 891.600 712.050 892.050 ;
        RECT 760.950 891.600 763.050 892.050 ;
        RECT 709.950 890.400 763.050 891.600 ;
        RECT 709.950 889.950 712.050 890.400 ;
        RECT 760.950 889.950 763.050 890.400 ;
        RECT 40.950 885.600 43.050 886.200 ;
        RECT 52.950 885.600 55.050 886.050 ;
        RECT 40.950 884.400 55.050 885.600 ;
        RECT 40.950 884.100 43.050 884.400 ;
        RECT 52.950 883.950 55.050 884.400 ;
        RECT 64.950 885.600 67.050 886.200 ;
        RECT 70.950 885.600 73.050 886.200 ;
        RECT 64.950 884.400 73.050 885.600 ;
        RECT 64.950 884.100 67.050 884.400 ;
        RECT 70.950 884.100 73.050 884.400 ;
        RECT 160.950 885.600 163.050 886.200 ;
        RECT 166.950 885.600 169.050 886.200 ;
        RECT 160.950 884.400 169.050 885.600 ;
        RECT 160.950 884.100 163.050 884.400 ;
        RECT 166.950 884.100 169.050 884.400 ;
        RECT 229.950 885.600 232.050 886.200 ;
        RECT 247.950 885.600 250.050 886.200 ;
        RECT 229.950 884.400 250.050 885.600 ;
        RECT 229.950 884.100 232.050 884.400 ;
        RECT 247.950 884.100 250.050 884.400 ;
        RECT 280.950 885.750 283.050 886.200 ;
        RECT 286.950 885.750 289.050 886.200 ;
        RECT 280.950 884.550 289.050 885.750 ;
        RECT 280.950 884.100 283.050 884.550 ;
        RECT 286.950 884.100 289.050 884.550 ;
        RECT 322.950 885.600 325.050 886.200 ;
        RECT 343.950 885.600 346.050 886.200 ;
        RECT 322.950 884.400 346.050 885.600 ;
        RECT 322.950 884.100 325.050 884.400 ;
        RECT 343.950 884.100 346.050 884.400 ;
        RECT 361.950 885.600 364.050 886.050 ;
        RECT 367.950 885.600 370.050 886.200 ;
        RECT 361.950 884.400 370.050 885.600 ;
        RECT 361.950 883.950 364.050 884.400 ;
        RECT 367.950 884.100 370.050 884.400 ;
        RECT 382.950 885.600 385.050 886.050 ;
        RECT 391.950 885.600 394.050 886.200 ;
        RECT 382.950 884.400 394.050 885.600 ;
        RECT 382.950 883.950 385.050 884.400 ;
        RECT 391.950 884.100 394.050 884.400 ;
        RECT 421.950 885.600 424.050 886.200 ;
        RECT 427.950 885.600 430.050 886.200 ;
        RECT 421.950 884.400 430.050 885.600 ;
        RECT 421.950 884.100 424.050 884.400 ;
        RECT 427.950 884.100 430.050 884.400 ;
        RECT 502.950 885.600 505.050 886.200 ;
        RECT 508.950 885.600 511.050 886.200 ;
        RECT 502.950 884.400 511.050 885.600 ;
        RECT 502.950 884.100 505.050 884.400 ;
        RECT 508.950 884.100 511.050 884.400 ;
        RECT 571.950 885.600 574.050 886.200 ;
        RECT 592.950 885.600 595.050 886.200 ;
        RECT 571.950 884.400 595.050 885.600 ;
        RECT 571.950 884.100 574.050 884.400 ;
        RECT 592.950 884.100 595.050 884.400 ;
        RECT 655.950 885.750 658.050 886.200 ;
        RECT 664.950 885.750 667.050 886.200 ;
        RECT 655.950 884.550 667.050 885.750 ;
        RECT 655.950 884.100 658.050 884.550 ;
        RECT 664.950 884.100 667.050 884.550 ;
        RECT 670.950 885.600 673.050 886.200 ;
        RECT 682.950 885.600 685.050 886.050 ;
        RECT 670.950 884.400 685.050 885.600 ;
        RECT 670.950 884.100 673.050 884.400 ;
        RECT 682.950 883.950 685.050 884.400 ;
        RECT 730.950 885.600 733.050 886.200 ;
        RECT 739.800 885.600 741.900 886.050 ;
        RECT 730.950 884.400 741.900 885.600 ;
        RECT 730.950 884.100 733.050 884.400 ;
        RECT 739.800 883.950 741.900 884.400 ;
        RECT 742.950 885.600 745.050 886.050 ;
        RECT 751.950 885.600 754.050 886.200 ;
        RECT 742.950 884.400 754.050 885.600 ;
        RECT 742.950 883.950 745.050 884.400 ;
        RECT 751.950 884.100 754.050 884.400 ;
        RECT 793.950 885.600 796.050 886.200 ;
        RECT 802.950 885.600 805.050 886.050 ;
        RECT 793.950 884.400 805.050 885.600 ;
        RECT 793.950 884.100 796.050 884.400 ;
        RECT 802.950 883.950 805.050 884.400 ;
        RECT 808.950 885.600 811.050 886.050 ;
        RECT 817.950 885.600 820.050 886.200 ;
        RECT 808.950 884.400 820.050 885.600 ;
        RECT 808.950 883.950 811.050 884.400 ;
        RECT 817.950 884.100 820.050 884.400 ;
        RECT 829.950 885.750 832.050 886.200 ;
        RECT 835.950 885.750 838.050 886.200 ;
        RECT 829.950 884.550 838.050 885.750 ;
        RECT 829.950 884.100 832.050 884.550 ;
        RECT 835.950 884.100 838.050 884.550 ;
        RECT 841.950 885.750 844.050 886.200 ;
        RECT 847.950 885.750 850.050 886.200 ;
        RECT 841.950 884.550 850.050 885.750 ;
        RECT 841.950 884.100 844.050 884.550 ;
        RECT 847.950 884.100 850.050 884.550 ;
        RECT 862.950 885.750 865.050 886.200 ;
        RECT 868.950 885.750 871.050 886.200 ;
        RECT 862.950 884.550 871.050 885.750 ;
        RECT 862.950 884.100 865.050 884.550 ;
        RECT 868.950 884.100 871.050 884.550 ;
        RECT 16.950 879.600 19.050 879.900 ;
        RECT 25.950 879.600 28.050 880.050 ;
        RECT 37.950 879.600 40.050 879.900 ;
        RECT 16.950 878.400 40.050 879.600 ;
        RECT 16.950 877.800 19.050 878.400 ;
        RECT 25.950 877.950 28.050 878.400 ;
        RECT 37.950 877.800 40.050 878.400 ;
        RECT 97.950 879.600 100.050 879.900 ;
        RECT 118.950 879.600 121.050 879.900 ;
        RECT 97.950 878.400 121.050 879.600 ;
        RECT 97.950 877.800 100.050 878.400 ;
        RECT 118.950 877.800 121.050 878.400 ;
        RECT 193.950 879.600 196.050 879.900 ;
        RECT 202.950 879.600 205.050 879.900 ;
        RECT 193.950 878.400 205.050 879.600 ;
        RECT 193.950 877.800 196.050 878.400 ;
        RECT 202.950 877.800 205.050 878.400 ;
        RECT 535.950 879.600 538.050 879.900 ;
        RECT 544.950 879.600 547.050 879.900 ;
        RECT 535.950 878.400 547.050 879.600 ;
        RECT 535.950 877.800 538.050 878.400 ;
        RECT 544.950 877.800 547.050 878.400 ;
        RECT 712.950 879.600 715.050 879.900 ;
        RECT 727.950 879.600 730.050 879.900 ;
        RECT 712.950 879.450 730.050 879.600 ;
        RECT 742.950 879.450 745.050 879.900 ;
        RECT 712.950 878.400 745.050 879.450 ;
        RECT 712.950 877.800 715.050 878.400 ;
        RECT 727.950 878.250 745.050 878.400 ;
        RECT 727.950 877.800 730.050 878.250 ;
        RECT 742.950 877.800 745.050 878.250 ;
        RECT 754.950 879.600 757.050 879.900 ;
        RECT 775.950 879.600 778.050 879.900 ;
        RECT 754.950 878.400 778.050 879.600 ;
        RECT 754.950 877.800 757.050 878.400 ;
        RECT 775.950 877.800 778.050 878.400 ;
        RECT 802.950 879.450 805.050 879.900 ;
        RECT 814.950 879.450 817.050 879.900 ;
        RECT 802.950 878.250 817.050 879.450 ;
        RECT 802.950 877.800 805.050 878.250 ;
        RECT 814.950 877.800 817.050 878.250 ;
        RECT 88.950 876.600 91.050 877.050 ;
        RECT 211.950 876.600 214.050 877.050 ;
        RECT 247.950 876.600 250.050 877.050 ;
        RECT 88.950 875.400 96.600 876.600 ;
        RECT 88.950 874.950 91.050 875.400 ;
        RECT 95.400 873.600 96.600 875.400 ;
        RECT 211.950 875.400 250.050 876.600 ;
        RECT 211.950 874.950 214.050 875.400 ;
        RECT 247.950 874.950 250.050 875.400 ;
        RECT 289.950 876.600 292.050 877.050 ;
        RECT 310.950 876.600 313.050 877.050 ;
        RECT 289.950 875.400 313.050 876.600 ;
        RECT 289.950 874.950 292.050 875.400 ;
        RECT 310.950 874.950 313.050 875.400 ;
        RECT 349.950 876.600 352.050 877.050 ;
        RECT 376.950 876.600 379.050 877.050 ;
        RECT 400.950 876.600 403.050 877.050 ;
        RECT 472.950 876.600 475.050 877.050 ;
        RECT 349.950 875.400 475.050 876.600 ;
        RECT 349.950 874.950 352.050 875.400 ;
        RECT 376.950 874.950 379.050 875.400 ;
        RECT 400.950 874.950 403.050 875.400 ;
        RECT 472.950 874.950 475.050 875.400 ;
        RECT 553.950 876.600 556.050 877.050 ;
        RECT 613.950 876.600 616.050 877.050 ;
        RECT 655.950 876.600 658.050 877.050 ;
        RECT 553.950 875.400 658.050 876.600 ;
        RECT 553.950 874.950 556.050 875.400 ;
        RECT 613.950 874.950 616.050 875.400 ;
        RECT 655.950 874.950 658.050 875.400 ;
        RECT 688.950 876.600 691.050 877.050 ;
        RECT 706.950 876.600 709.050 877.050 ;
        RECT 688.950 875.400 709.050 876.600 ;
        RECT 688.950 874.950 691.050 875.400 ;
        RECT 706.950 874.950 709.050 875.400 ;
        RECT 847.950 876.600 850.050 877.050 ;
        RECT 862.950 876.600 865.050 877.050 ;
        RECT 871.950 876.600 874.050 877.050 ;
        RECT 847.950 875.400 874.050 876.600 ;
        RECT 847.950 874.950 850.050 875.400 ;
        RECT 862.950 874.950 865.050 875.400 ;
        RECT 871.950 874.950 874.050 875.400 ;
        RECT 142.950 873.600 145.050 874.050 ;
        RECT 95.400 872.400 145.050 873.600 ;
        RECT 142.950 871.950 145.050 872.400 ;
        RECT 202.950 873.600 205.050 874.050 ;
        RECT 295.950 873.600 298.050 874.050 ;
        RECT 346.950 873.600 349.050 874.050 ;
        RECT 202.950 872.400 349.050 873.600 ;
        RECT 202.950 871.950 205.050 872.400 ;
        RECT 295.950 871.950 298.050 872.400 ;
        RECT 346.950 871.950 349.050 872.400 ;
        RECT 667.950 873.600 670.050 874.050 ;
        RECT 689.400 873.600 690.600 874.950 ;
        RECT 667.950 872.400 690.600 873.600 ;
        RECT 775.950 873.600 778.050 874.050 ;
        RECT 784.950 873.600 787.050 874.050 ;
        RECT 796.950 873.600 799.050 874.050 ;
        RECT 775.950 872.400 799.050 873.600 ;
        RECT 667.950 871.950 670.050 872.400 ;
        RECT 775.950 871.950 778.050 872.400 ;
        RECT 784.950 871.950 787.050 872.400 ;
        RECT 796.950 871.950 799.050 872.400 ;
        RECT 829.950 873.600 832.050 874.050 ;
        RECT 838.950 873.600 841.050 874.050 ;
        RECT 829.950 872.400 841.050 873.600 ;
        RECT 829.950 871.950 832.050 872.400 ;
        RECT 838.950 871.950 841.050 872.400 ;
        RECT 454.950 870.600 457.050 871.050 ;
        RECT 481.950 870.600 484.050 871.050 ;
        RECT 454.950 869.400 484.050 870.600 ;
        RECT 454.950 868.950 457.050 869.400 ;
        RECT 481.950 868.950 484.050 869.400 ;
        RECT 280.950 867.600 283.050 868.050 ;
        RECT 289.950 867.600 292.050 868.050 ;
        RECT 361.950 867.600 364.050 868.050 ;
        RECT 412.950 867.600 415.050 868.050 ;
        RECT 280.950 866.400 415.050 867.600 ;
        RECT 280.950 865.950 283.050 866.400 ;
        RECT 289.950 865.950 292.050 866.400 ;
        RECT 361.950 865.950 364.050 866.400 ;
        RECT 412.950 865.950 415.050 866.400 ;
        RECT 472.950 867.600 475.050 868.050 ;
        RECT 661.950 867.600 664.050 868.050 ;
        RECT 472.950 866.400 664.050 867.600 ;
        RECT 472.950 865.950 475.050 866.400 ;
        RECT 661.950 865.950 664.050 866.400 ;
        RECT 748.950 864.600 751.050 865.050 ;
        RECT 769.950 864.600 772.050 865.050 ;
        RECT 689.400 863.400 772.050 864.600 ;
        RECT 643.950 861.600 646.050 862.050 ;
        RECT 689.400 861.600 690.600 863.400 ;
        RECT 748.950 862.950 751.050 863.400 ;
        RECT 769.950 862.950 772.050 863.400 ;
        RECT 643.950 860.400 690.600 861.600 ;
        RECT 643.950 859.950 646.050 860.400 ;
        RECT 814.950 858.600 817.050 859.050 ;
        RECT 871.950 858.600 874.050 859.050 ;
        RECT 814.950 857.400 874.050 858.600 ;
        RECT 814.950 856.950 817.050 857.400 ;
        RECT 871.950 856.950 874.050 857.400 ;
        RECT 277.950 855.600 280.050 856.050 ;
        RECT 298.950 855.600 301.050 856.050 ;
        RECT 382.950 855.600 385.050 856.050 ;
        RECT 277.950 854.400 385.050 855.600 ;
        RECT 277.950 853.950 280.050 854.400 ;
        RECT 298.950 853.950 301.050 854.400 ;
        RECT 382.950 853.950 385.050 854.400 ;
        RECT 715.950 855.600 718.050 856.050 ;
        RECT 739.950 855.600 742.050 856.050 ;
        RECT 715.950 854.400 742.050 855.600 ;
        RECT 715.950 853.950 718.050 854.400 ;
        RECT 739.950 853.950 742.050 854.400 ;
        RECT 118.950 852.600 121.050 853.050 ;
        RECT 187.950 852.600 190.050 853.050 ;
        RECT 202.950 852.600 205.050 853.050 ;
        RECT 118.950 851.400 205.050 852.600 ;
        RECT 118.950 850.950 121.050 851.400 ;
        RECT 187.950 850.950 190.050 851.400 ;
        RECT 202.950 850.950 205.050 851.400 ;
        RECT 307.950 852.600 310.050 853.050 ;
        RECT 364.950 852.600 367.050 853.050 ;
        RECT 307.950 851.400 367.050 852.600 ;
        RECT 307.950 850.950 310.050 851.400 ;
        RECT 364.950 850.950 367.050 851.400 ;
        RECT 625.950 852.600 628.050 853.050 ;
        RECT 667.950 852.600 670.050 853.050 ;
        RECT 625.950 851.400 670.050 852.600 ;
        RECT 625.950 850.950 628.050 851.400 ;
        RECT 667.950 850.950 670.050 851.400 ;
        RECT 790.950 852.600 793.050 853.050 ;
        RECT 835.950 852.600 838.050 853.050 ;
        RECT 790.950 851.400 838.050 852.600 ;
        RECT 790.950 850.950 793.050 851.400 ;
        RECT 835.950 850.950 838.050 851.400 ;
        RECT 43.950 849.600 46.050 850.050 ;
        RECT 76.950 849.600 79.050 850.050 ;
        RECT 100.950 849.600 103.050 850.050 ;
        RECT 349.950 849.600 352.050 850.050 ;
        RECT 43.950 848.400 352.050 849.600 ;
        RECT 43.950 847.950 46.050 848.400 ;
        RECT 76.950 847.950 79.050 848.400 ;
        RECT 100.950 847.950 103.050 848.400 ;
        RECT 349.950 847.950 352.050 848.400 ;
        RECT 382.950 849.600 385.050 850.050 ;
        RECT 406.950 849.600 409.050 850.050 ;
        RECT 382.950 848.400 409.050 849.600 ;
        RECT 382.950 847.950 385.050 848.400 ;
        RECT 406.950 847.950 409.050 848.400 ;
        RECT 442.950 849.600 445.050 850.050 ;
        RECT 475.950 849.600 478.050 850.050 ;
        RECT 442.950 848.400 478.050 849.600 ;
        RECT 442.950 847.950 445.050 848.400 ;
        RECT 475.950 847.950 478.050 848.400 ;
        RECT 682.950 849.600 685.050 850.050 ;
        RECT 709.950 849.600 712.050 850.050 ;
        RECT 727.950 849.600 730.050 850.050 ;
        RECT 682.950 848.400 730.050 849.600 ;
        RECT 682.950 847.950 685.050 848.400 ;
        RECT 709.950 847.950 712.050 848.400 ;
        RECT 727.950 847.950 730.050 848.400 ;
        RECT 856.950 849.600 859.050 850.050 ;
        RECT 877.950 849.600 880.050 850.050 ;
        RECT 856.950 848.400 880.050 849.600 ;
        RECT 856.950 847.950 859.050 848.400 ;
        RECT 877.950 847.950 880.050 848.400 ;
        RECT 145.950 846.600 148.050 847.050 ;
        RECT 208.950 846.600 211.050 847.050 ;
        RECT 235.950 846.600 238.050 847.050 ;
        RECT 145.950 845.400 238.050 846.600 ;
        RECT 145.950 844.950 148.050 845.400 ;
        RECT 208.950 844.950 211.050 845.400 ;
        RECT 235.950 844.950 238.050 845.400 ;
        RECT 262.950 846.600 265.050 847.050 ;
        RECT 289.950 846.600 292.050 847.050 ;
        RECT 262.950 845.400 292.050 846.600 ;
        RECT 262.950 844.950 265.050 845.400 ;
        RECT 289.950 844.950 292.050 845.400 ;
        RECT 346.950 846.600 349.050 847.050 ;
        RECT 382.950 846.600 385.050 846.900 ;
        RECT 346.950 845.400 385.050 846.600 ;
        RECT 346.950 844.950 349.050 845.400 ;
        RECT 382.950 844.800 385.050 845.400 ;
        RECT 616.950 846.600 619.050 847.050 ;
        RECT 637.950 846.600 640.050 847.050 ;
        RECT 649.950 846.600 652.050 847.050 ;
        RECT 616.950 845.400 652.050 846.600 ;
        RECT 616.950 844.950 619.050 845.400 ;
        RECT 637.950 844.950 640.050 845.400 ;
        RECT 649.950 844.950 652.050 845.400 ;
        RECT 667.950 846.600 670.050 847.050 ;
        RECT 745.950 846.600 748.050 847.050 ;
        RECT 667.950 845.400 748.050 846.600 ;
        RECT 667.950 844.950 670.050 845.400 ;
        RECT 745.950 844.950 748.050 845.400 ;
        RECT 472.950 843.600 475.050 844.050 ;
        RECT 481.950 843.600 484.050 844.050 ;
        RECT 517.950 843.600 520.050 844.050 ;
        RECT 535.950 843.600 538.050 844.050 ;
        RECT 472.950 842.400 538.050 843.600 ;
        RECT 472.950 841.950 475.050 842.400 ;
        RECT 481.950 841.950 484.050 842.400 ;
        RECT 517.950 841.950 520.050 842.400 ;
        RECT 535.950 841.950 538.050 842.400 ;
        RECT 568.950 843.600 571.050 844.050 ;
        RECT 586.950 843.600 589.050 844.050 ;
        RECT 568.950 842.400 589.050 843.600 ;
        RECT 568.950 841.950 571.050 842.400 ;
        RECT 586.950 841.950 589.050 842.400 ;
        RECT 664.950 843.600 667.050 844.050 ;
        RECT 679.950 843.600 682.050 844.050 ;
        RECT 664.950 842.400 682.050 843.600 ;
        RECT 664.950 841.950 667.050 842.400 ;
        RECT 679.950 841.950 682.050 842.400 ;
        RECT 16.950 840.600 19.050 841.200 ;
        RECT 28.950 840.600 31.050 841.050 ;
        RECT 34.950 840.600 37.050 841.200 ;
        RECT 16.950 839.400 37.050 840.600 ;
        RECT 16.950 839.100 19.050 839.400 ;
        RECT 28.950 838.950 31.050 839.400 ;
        RECT 34.950 839.100 37.050 839.400 ;
        RECT 40.950 840.750 43.050 841.200 ;
        RECT 52.950 840.750 55.050 841.200 ;
        RECT 40.950 839.550 55.050 840.750 ;
        RECT 40.950 839.100 43.050 839.550 ;
        RECT 52.950 839.100 55.050 839.550 ;
        RECT 118.950 840.750 121.050 841.200 ;
        RECT 127.950 840.750 130.050 841.200 ;
        RECT 118.950 839.550 130.050 840.750 ;
        RECT 118.950 839.100 121.050 839.550 ;
        RECT 127.950 839.100 130.050 839.550 ;
        RECT 133.950 840.600 136.050 841.200 ;
        RECT 151.950 840.600 154.050 841.200 ;
        RECT 133.950 839.400 154.050 840.600 ;
        RECT 133.950 839.100 136.050 839.400 ;
        RECT 151.950 839.100 154.050 839.400 ;
        RECT 178.950 839.100 181.050 841.200 ;
        RECT 214.950 839.100 217.050 841.200 ;
        RECT 223.950 840.750 226.050 841.200 ;
        RECT 229.950 840.750 232.050 841.200 ;
        RECT 223.950 839.550 232.050 840.750 ;
        RECT 223.950 839.100 226.050 839.550 ;
        RECT 229.950 839.100 232.050 839.550 ;
        RECT 256.950 840.750 259.050 841.200 ;
        RECT 268.950 840.750 271.050 841.200 ;
        RECT 256.950 840.600 271.050 840.750 ;
        RECT 283.950 840.600 286.050 841.200 ;
        RECT 256.950 839.550 286.050 840.600 ;
        RECT 256.950 839.100 259.050 839.550 ;
        RECT 268.950 839.400 286.050 839.550 ;
        RECT 268.950 839.100 271.050 839.400 ;
        RECT 283.950 839.100 286.050 839.400 ;
        RECT 295.950 840.750 298.050 841.200 ;
        RECT 304.950 840.750 307.050 841.200 ;
        RECT 295.950 839.550 307.050 840.750 ;
        RECT 295.950 839.100 298.050 839.550 ;
        RECT 304.950 839.100 307.050 839.550 ;
        RECT 310.950 840.600 313.050 841.200 ;
        RECT 328.800 840.600 330.900 841.050 ;
        RECT 310.950 839.400 330.900 840.600 ;
        RECT 310.950 839.100 313.050 839.400 ;
        RECT 79.950 834.600 82.050 834.900 ;
        RECT 103.950 834.600 106.050 834.900 ;
        RECT 79.950 833.400 106.050 834.600 ;
        RECT 79.950 832.800 82.050 833.400 ;
        RECT 103.950 832.800 106.050 833.400 ;
        RECT 136.950 834.600 139.050 834.900 ;
        RECT 145.950 834.600 148.050 835.050 ;
        RECT 136.950 833.400 148.050 834.600 ;
        RECT 136.950 832.800 139.050 833.400 ;
        RECT 145.950 832.950 148.050 833.400 ;
        RECT 179.400 832.050 180.600 839.100 ;
        RECT 215.400 834.600 216.600 839.100 ;
        RECT 328.800 838.950 330.900 839.400 ;
        RECT 331.950 840.750 334.050 841.200 ;
        RECT 337.950 840.750 340.050 841.200 ;
        RECT 331.950 839.550 340.050 840.750 ;
        RECT 331.950 839.100 334.050 839.550 ;
        RECT 337.950 839.100 340.050 839.550 ;
        RECT 373.950 840.600 376.050 841.200 ;
        RECT 427.950 840.600 430.050 841.050 ;
        RECT 373.950 839.400 430.050 840.600 ;
        RECT 373.950 839.100 376.050 839.400 ;
        RECT 427.950 838.950 430.050 839.400 ;
        RECT 508.950 840.600 511.050 841.200 ;
        RECT 538.950 840.600 541.050 841.200 ;
        RECT 508.950 839.400 541.050 840.600 ;
        RECT 508.950 839.100 511.050 839.400 ;
        RECT 538.950 839.100 541.050 839.400 ;
        RECT 547.950 840.750 550.050 841.200 ;
        RECT 562.950 840.750 565.050 841.200 ;
        RECT 547.950 839.550 565.050 840.750 ;
        RECT 547.950 839.100 550.050 839.550 ;
        RECT 562.950 839.100 565.050 839.550 ;
        RECT 574.950 840.750 577.050 841.200 ;
        RECT 592.950 840.750 595.050 841.200 ;
        RECT 574.950 839.550 595.050 840.750 ;
        RECT 574.950 839.100 577.050 839.550 ;
        RECT 592.950 839.100 595.050 839.550 ;
        RECT 604.950 840.750 607.050 841.200 ;
        RECT 610.950 840.750 613.050 841.200 ;
        RECT 604.950 839.550 613.050 840.750 ;
        RECT 604.950 839.100 607.050 839.550 ;
        RECT 610.950 839.100 613.050 839.550 ;
        RECT 643.950 840.600 646.050 841.200 ;
        RECT 661.950 840.600 664.050 841.200 ;
        RECT 643.950 839.400 664.050 840.600 ;
        RECT 643.950 839.100 646.050 839.400 ;
        RECT 661.950 839.100 664.050 839.400 ;
        RECT 685.950 840.750 688.050 841.200 ;
        RECT 691.800 840.750 693.900 841.200 ;
        RECT 685.950 839.550 693.900 840.750 ;
        RECT 685.950 839.100 688.050 839.550 ;
        RECT 691.800 839.100 693.900 839.550 ;
        RECT 694.950 840.750 697.050 841.200 ;
        RECT 703.950 840.750 706.050 841.200 ;
        RECT 694.950 840.600 706.050 840.750 ;
        RECT 733.950 840.600 736.050 841.200 ;
        RECT 694.950 839.550 736.050 840.600 ;
        RECT 694.950 839.100 697.050 839.550 ;
        RECT 703.950 839.400 736.050 839.550 ;
        RECT 703.950 839.100 706.050 839.400 ;
        RECT 733.950 839.100 736.050 839.400 ;
        RECT 754.950 839.100 757.050 841.200 ;
        RECT 760.950 840.600 763.050 841.200 ;
        RECT 766.950 840.600 769.050 840.900 ;
        RECT 760.950 839.400 769.050 840.600 ;
        RECT 760.950 839.100 763.050 839.400 ;
        RECT 247.950 837.600 250.050 838.050 ;
        RECT 247.950 836.400 321.600 837.600 ;
        RECT 247.950 835.950 250.050 836.400 ;
        RECT 320.400 834.900 321.600 836.400 ;
        RECT 232.950 834.600 235.050 834.900 ;
        RECT 253.950 834.600 256.050 834.900 ;
        RECT 215.400 833.400 256.050 834.600 ;
        RECT 232.950 832.800 235.050 833.400 ;
        RECT 253.950 832.800 256.050 833.400 ;
        RECT 298.950 834.450 301.050 834.900 ;
        RECT 313.950 834.450 316.050 834.900 ;
        RECT 298.950 833.250 316.050 834.450 ;
        RECT 298.950 832.800 301.050 833.250 ;
        RECT 313.950 832.800 316.050 833.250 ;
        RECT 319.950 832.800 322.050 834.900 ;
        RECT 355.950 834.450 358.050 834.900 ;
        RECT 364.950 834.450 367.050 834.900 ;
        RECT 355.950 833.250 367.050 834.450 ;
        RECT 355.950 832.800 358.050 833.250 ;
        RECT 364.950 832.800 367.050 833.250 ;
        RECT 391.950 834.450 394.050 834.900 ;
        RECT 403.950 834.450 406.050 834.900 ;
        RECT 430.950 834.600 433.050 834.900 ;
        RECT 391.950 833.250 406.050 834.450 ;
        RECT 391.950 832.800 394.050 833.250 ;
        RECT 403.950 832.800 406.050 833.250 ;
        RECT 428.400 833.400 433.050 834.600 ;
        RECT 178.950 829.950 181.050 832.050 ;
        RECT 331.950 831.600 334.050 832.050 ;
        RECT 346.950 831.600 349.050 832.050 ;
        RECT 331.950 830.400 349.050 831.600 ;
        RECT 331.950 829.950 334.050 830.400 ;
        RECT 346.950 829.950 349.050 830.400 ;
        RECT 406.950 831.600 409.050 832.050 ;
        RECT 428.400 831.600 429.600 833.400 ;
        RECT 430.950 832.800 433.050 833.400 ;
        RECT 475.950 834.450 478.050 834.900 ;
        RECT 490.950 834.450 493.050 834.900 ;
        RECT 475.950 833.250 493.050 834.450 ;
        RECT 475.950 832.800 478.050 833.250 ;
        RECT 490.950 832.800 493.050 833.250 ;
        RECT 619.950 834.450 622.050 834.900 ;
        RECT 625.950 834.600 628.050 834.900 ;
        RECT 634.950 834.600 637.050 834.900 ;
        RECT 625.950 834.450 637.050 834.600 ;
        RECT 619.950 833.400 637.050 834.450 ;
        RECT 619.950 833.250 628.050 833.400 ;
        RECT 619.950 832.800 622.050 833.250 ;
        RECT 625.950 832.800 628.050 833.250 ;
        RECT 634.950 832.800 637.050 833.400 ;
        RECT 649.950 834.600 652.050 835.050 ;
        RECT 700.950 834.600 703.050 834.900 ;
        RECT 649.950 833.400 703.050 834.600 ;
        RECT 649.950 832.950 652.050 833.400 ;
        RECT 700.950 832.800 703.050 833.400 ;
        RECT 712.950 834.600 715.050 835.050 ;
        RECT 724.950 834.600 727.050 834.900 ;
        RECT 712.950 833.400 727.050 834.600 ;
        RECT 712.950 832.950 715.050 833.400 ;
        RECT 724.950 832.800 727.050 833.400 ;
        RECT 730.950 834.450 733.050 834.900 ;
        RECT 739.950 834.450 742.050 834.900 ;
        RECT 730.950 833.250 742.050 834.450 ;
        RECT 730.950 832.800 733.050 833.250 ;
        RECT 739.950 832.800 742.050 833.250 ;
        RECT 745.950 834.600 748.050 835.050 ;
        RECT 751.950 834.600 754.050 834.900 ;
        RECT 745.950 833.400 754.050 834.600 ;
        RECT 745.950 832.950 748.050 833.400 ;
        RECT 751.950 832.800 754.050 833.400 ;
        RECT 755.400 832.050 756.600 839.100 ;
        RECT 766.950 838.800 769.050 839.400 ;
        RECT 784.950 840.600 787.050 841.200 ;
        RECT 808.950 840.600 811.050 841.050 ;
        RECT 832.950 840.600 835.050 841.200 ;
        RECT 847.950 840.600 850.050 841.200 ;
        RECT 784.950 839.400 850.050 840.600 ;
        RECT 784.950 839.100 787.050 839.400 ;
        RECT 808.950 838.950 811.050 839.400 ;
        RECT 832.950 839.100 835.050 839.400 ;
        RECT 847.950 839.100 850.050 839.400 ;
        RECT 877.950 840.600 880.050 841.200 ;
        RECT 892.950 840.600 895.050 841.200 ;
        RECT 877.950 839.400 895.050 840.600 ;
        RECT 877.950 839.100 880.050 839.400 ;
        RECT 892.950 839.100 895.050 839.400 ;
        RECT 769.950 834.450 772.050 834.900 ;
        RECT 781.950 834.450 784.050 834.900 ;
        RECT 769.950 833.250 784.050 834.450 ;
        RECT 769.950 832.800 772.050 833.250 ;
        RECT 781.950 832.800 784.050 833.250 ;
        RECT 406.950 830.400 429.600 831.600 ;
        RECT 406.950 829.950 409.050 830.400 ;
        RECT 754.950 829.950 757.050 832.050 ;
        RECT 25.950 828.600 28.050 829.050 ;
        RECT 79.950 828.600 82.050 829.050 ;
        RECT 25.950 827.400 82.050 828.600 ;
        RECT 25.950 826.950 28.050 827.400 ;
        RECT 79.950 826.950 82.050 827.400 ;
        RECT 109.950 828.600 112.050 829.050 ;
        RECT 127.950 828.600 130.050 829.050 ;
        RECT 109.950 827.400 130.050 828.600 ;
        RECT 109.950 826.950 112.050 827.400 ;
        RECT 127.950 826.950 130.050 827.400 ;
        RECT 142.950 828.600 145.050 829.050 ;
        RECT 160.950 828.600 163.050 829.050 ;
        RECT 142.950 827.400 163.050 828.600 ;
        RECT 142.950 826.950 145.050 827.400 ;
        RECT 160.950 826.950 163.050 827.400 ;
        RECT 427.950 828.600 430.050 829.050 ;
        RECT 436.950 828.600 439.050 829.050 ;
        RECT 427.950 827.400 439.050 828.600 ;
        RECT 427.950 826.950 430.050 827.400 ;
        RECT 436.950 826.950 439.050 827.400 ;
        RECT 523.950 828.600 526.050 829.050 ;
        RECT 556.950 828.600 559.050 829.050 ;
        RECT 523.950 827.400 559.050 828.600 ;
        RECT 523.950 826.950 526.050 827.400 ;
        RECT 556.950 826.950 559.050 827.400 ;
        RECT 598.950 828.600 601.050 829.050 ;
        RECT 613.950 828.600 616.050 829.050 ;
        RECT 598.950 827.400 616.050 828.600 ;
        RECT 598.950 826.950 601.050 827.400 ;
        RECT 613.950 826.950 616.050 827.400 ;
        RECT 625.950 828.600 628.050 829.050 ;
        RECT 658.950 828.600 661.050 829.050 ;
        RECT 625.950 827.400 661.050 828.600 ;
        RECT 625.950 826.950 628.050 827.400 ;
        RECT 658.950 826.950 661.050 827.400 ;
        RECT 781.950 828.600 784.050 829.050 ;
        RECT 805.950 828.600 808.050 829.050 ;
        RECT 781.950 827.400 808.050 828.600 ;
        RECT 781.950 826.950 784.050 827.400 ;
        RECT 805.950 826.950 808.050 827.400 ;
        RECT 862.950 828.600 865.050 829.050 ;
        RECT 898.950 828.600 901.050 829.050 ;
        RECT 862.950 827.400 901.050 828.600 ;
        RECT 862.950 826.950 865.050 827.400 ;
        RECT 898.950 826.950 901.050 827.400 ;
        RECT 103.950 825.600 106.050 826.050 ;
        RECT 130.950 825.600 133.050 826.050 ;
        RECT 103.950 824.400 133.050 825.600 ;
        RECT 103.950 823.950 106.050 824.400 ;
        RECT 130.950 823.950 133.050 824.400 ;
        RECT 310.950 825.600 313.050 826.050 ;
        RECT 328.950 825.600 331.050 826.050 ;
        RECT 310.950 824.400 331.050 825.600 ;
        RECT 310.950 823.950 313.050 824.400 ;
        RECT 328.950 823.950 331.050 824.400 ;
        RECT 490.950 825.600 493.050 826.050 ;
        RECT 535.950 825.600 538.050 826.050 ;
        RECT 490.950 824.400 538.050 825.600 ;
        RECT 490.950 823.950 493.050 824.400 ;
        RECT 535.950 823.950 538.050 824.400 ;
        RECT 565.950 825.600 568.050 826.050 ;
        RECT 589.950 825.600 592.050 826.050 ;
        RECT 676.950 825.600 679.050 826.050 ;
        RECT 565.950 824.400 679.050 825.600 ;
        RECT 565.950 823.950 568.050 824.400 ;
        RECT 589.950 823.950 592.050 824.400 ;
        RECT 676.950 823.950 679.050 824.400 ;
        RECT 751.950 825.600 754.050 826.050 ;
        RECT 775.950 825.600 778.050 826.050 ;
        RECT 751.950 824.400 778.050 825.600 ;
        RECT 751.950 823.950 754.050 824.400 ;
        RECT 775.950 823.950 778.050 824.400 ;
        RECT 808.950 825.600 811.050 826.050 ;
        RECT 823.950 825.600 826.050 826.050 ;
        RECT 808.950 824.400 826.050 825.600 ;
        RECT 808.950 823.950 811.050 824.400 ;
        RECT 823.950 823.950 826.050 824.400 ;
        RECT 118.950 822.600 121.050 823.050 ;
        RECT 145.950 822.600 148.050 823.050 ;
        RECT 118.950 821.400 148.050 822.600 ;
        RECT 118.950 820.950 121.050 821.400 ;
        RECT 145.950 820.950 148.050 821.400 ;
        RECT 172.950 822.600 175.050 823.050 ;
        RECT 181.950 822.600 184.050 823.050 ;
        RECT 172.950 821.400 184.050 822.600 ;
        RECT 172.950 820.950 175.050 821.400 ;
        RECT 181.950 820.950 184.050 821.400 ;
        RECT 211.950 822.600 214.050 823.050 ;
        RECT 223.950 822.600 226.050 823.050 ;
        RECT 307.950 822.600 310.050 823.050 ;
        RECT 211.950 821.400 310.050 822.600 ;
        RECT 211.950 820.950 214.050 821.400 ;
        RECT 223.950 820.950 226.050 821.400 ;
        RECT 307.950 820.950 310.050 821.400 ;
        RECT 436.950 822.600 439.050 823.050 ;
        RECT 448.950 822.600 451.050 823.050 ;
        RECT 436.950 821.400 451.050 822.600 ;
        RECT 436.950 820.950 439.050 821.400 ;
        RECT 448.950 820.950 451.050 821.400 ;
        RECT 514.950 822.600 517.050 823.050 ;
        RECT 559.950 822.600 562.050 823.050 ;
        RECT 514.950 821.400 562.050 822.600 ;
        RECT 514.950 820.950 517.050 821.400 ;
        RECT 559.950 820.950 562.050 821.400 ;
        RECT 655.950 822.600 658.050 823.050 ;
        RECT 682.950 822.600 685.050 823.050 ;
        RECT 712.950 822.600 715.050 823.050 ;
        RECT 655.950 821.400 715.050 822.600 ;
        RECT 655.950 820.950 658.050 821.400 ;
        RECT 682.950 820.950 685.050 821.400 ;
        RECT 712.950 820.950 715.050 821.400 ;
        RECT 37.950 819.600 40.050 820.050 ;
        RECT 91.950 819.600 94.050 820.050 ;
        RECT 37.950 818.400 94.050 819.600 ;
        RECT 37.950 817.950 40.050 818.400 ;
        RECT 91.950 817.950 94.050 818.400 ;
        RECT 259.950 819.600 262.050 820.050 ;
        RECT 286.950 819.600 289.050 820.050 ;
        RECT 319.950 819.600 322.050 820.050 ;
        RECT 259.950 818.400 322.050 819.600 ;
        RECT 259.950 817.950 262.050 818.400 ;
        RECT 286.950 817.950 289.050 818.400 ;
        RECT 319.950 817.950 322.050 818.400 ;
        RECT 523.950 819.600 526.050 820.050 ;
        RECT 604.950 819.600 607.050 820.050 ;
        RECT 625.950 819.600 628.050 820.050 ;
        RECT 523.950 818.400 628.050 819.600 ;
        RECT 523.950 817.950 526.050 818.400 ;
        RECT 604.950 817.950 607.050 818.400 ;
        RECT 625.950 817.950 628.050 818.400 ;
        RECT 688.950 819.600 691.050 820.050 ;
        RECT 694.950 819.600 697.050 820.050 ;
        RECT 733.950 819.600 736.050 820.050 ;
        RECT 748.950 819.600 751.050 820.050 ;
        RECT 688.950 818.400 751.050 819.600 ;
        RECT 688.950 817.950 691.050 818.400 ;
        RECT 694.950 817.950 697.050 818.400 ;
        RECT 733.950 817.950 736.050 818.400 ;
        RECT 748.950 817.950 751.050 818.400 ;
        RECT 757.950 819.600 760.050 820.050 ;
        RECT 763.950 819.600 766.050 820.050 ;
        RECT 799.950 819.600 802.050 820.050 ;
        RECT 757.950 818.400 802.050 819.600 ;
        RECT 757.950 817.950 760.050 818.400 ;
        RECT 763.950 817.950 766.050 818.400 ;
        RECT 799.950 817.950 802.050 818.400 ;
        RECT 805.950 819.600 808.050 820.050 ;
        RECT 817.950 819.600 820.050 820.050 ;
        RECT 805.950 818.400 820.050 819.600 ;
        RECT 805.950 817.950 808.050 818.400 ;
        RECT 817.950 817.950 820.050 818.400 ;
        RECT 868.950 819.600 871.050 820.050 ;
        RECT 880.950 819.600 883.050 820.050 ;
        RECT 868.950 818.400 883.050 819.600 ;
        RECT 868.950 817.950 871.050 818.400 ;
        RECT 880.950 817.950 883.050 818.400 ;
        RECT 94.950 816.600 97.050 817.050 ;
        RECT 124.950 816.600 127.050 817.050 ;
        RECT 154.950 816.600 157.050 817.050 ;
        RECT 169.950 816.600 172.050 817.050 ;
        RECT 94.950 815.400 172.050 816.600 ;
        RECT 94.950 814.950 97.050 815.400 ;
        RECT 124.950 814.950 127.050 815.400 ;
        RECT 154.950 814.950 157.050 815.400 ;
        RECT 169.950 814.950 172.050 815.400 ;
        RECT 175.950 816.600 178.050 817.050 ;
        RECT 259.950 816.600 262.050 816.900 ;
        RECT 265.950 816.600 268.050 817.050 ;
        RECT 175.950 815.400 268.050 816.600 ;
        RECT 175.950 814.950 178.050 815.400 ;
        RECT 259.950 814.800 262.050 815.400 ;
        RECT 265.950 814.950 268.050 815.400 ;
        RECT 289.950 816.600 292.050 817.050 ;
        RECT 295.950 816.600 298.050 817.050 ;
        RECT 313.950 816.600 316.050 817.050 ;
        RECT 289.950 815.400 316.050 816.600 ;
        RECT 289.950 814.950 292.050 815.400 ;
        RECT 295.950 814.950 298.050 815.400 ;
        RECT 313.950 814.950 316.050 815.400 ;
        RECT 547.950 816.600 550.050 817.050 ;
        RECT 574.950 816.600 577.050 817.050 ;
        RECT 592.950 816.600 595.050 817.050 ;
        RECT 547.950 815.400 595.050 816.600 ;
        RECT 547.950 814.950 550.050 815.400 ;
        RECT 574.950 814.950 577.050 815.400 ;
        RECT 592.950 814.950 595.050 815.400 ;
        RECT 643.950 816.600 646.050 817.050 ;
        RECT 664.950 816.600 667.050 817.050 ;
        RECT 691.950 816.600 694.050 817.050 ;
        RECT 706.950 816.600 709.050 817.050 ;
        RECT 643.950 815.400 709.050 816.600 ;
        RECT 643.950 814.950 646.050 815.400 ;
        RECT 664.950 814.950 667.050 815.400 ;
        RECT 691.950 814.950 694.050 815.400 ;
        RECT 706.950 814.950 709.050 815.400 ;
        RECT 724.950 816.600 727.050 817.050 ;
        RECT 754.950 816.600 757.050 817.050 ;
        RECT 724.950 815.400 757.050 816.600 ;
        RECT 724.950 814.950 727.050 815.400 ;
        RECT 754.950 814.950 757.050 815.400 ;
        RECT 19.950 813.600 22.050 814.050 ;
        RECT 25.950 813.600 28.050 814.050 ;
        RECT 19.950 812.400 28.050 813.600 ;
        RECT 19.950 811.950 22.050 812.400 ;
        RECT 25.950 811.950 28.050 812.400 ;
        RECT 52.950 813.600 55.050 814.050 ;
        RECT 76.950 813.600 79.050 814.050 ;
        RECT 52.950 812.400 79.050 813.600 ;
        RECT 52.950 811.950 55.050 812.400 ;
        RECT 76.950 811.950 79.050 812.400 ;
        RECT 127.950 813.600 130.050 814.050 ;
        RECT 148.950 813.600 151.050 814.050 ;
        RECT 127.950 812.400 151.050 813.600 ;
        RECT 127.950 811.950 130.050 812.400 ;
        RECT 148.950 811.950 151.050 812.400 ;
        RECT 190.950 813.600 193.050 814.050 ;
        RECT 205.950 813.600 208.050 814.050 ;
        RECT 190.950 812.400 208.050 813.600 ;
        RECT 190.950 811.950 193.050 812.400 ;
        RECT 205.950 811.950 208.050 812.400 ;
        RECT 250.950 813.600 253.050 814.050 ;
        RECT 277.950 813.600 280.050 814.050 ;
        RECT 250.950 812.400 280.050 813.600 ;
        RECT 250.950 811.950 253.050 812.400 ;
        RECT 277.950 811.950 280.050 812.400 ;
        RECT 298.950 813.600 301.050 814.050 ;
        RECT 304.950 813.600 307.050 814.050 ;
        RECT 298.950 812.400 307.050 813.600 ;
        RECT 298.950 811.950 301.050 812.400 ;
        RECT 304.950 811.950 307.050 812.400 ;
        RECT 370.950 813.600 373.050 814.050 ;
        RECT 406.950 813.600 409.050 814.050 ;
        RECT 370.950 812.400 409.050 813.600 ;
        RECT 370.950 811.950 373.050 812.400 ;
        RECT 406.950 811.950 409.050 812.400 ;
        RECT 541.950 813.600 544.050 814.050 ;
        RECT 559.950 813.600 562.050 814.050 ;
        RECT 541.950 812.400 562.050 813.600 ;
        RECT 541.950 811.950 544.050 812.400 ;
        RECT 559.950 811.950 562.050 812.400 ;
        RECT 631.950 813.600 634.050 814.050 ;
        RECT 640.950 813.600 643.050 814.050 ;
        RECT 631.950 812.400 643.050 813.600 ;
        RECT 631.950 811.950 634.050 812.400 ;
        RECT 640.950 811.950 643.050 812.400 ;
        RECT 721.950 813.600 724.050 814.050 ;
        RECT 757.950 813.600 760.050 814.050 ;
        RECT 721.950 812.400 760.050 813.600 ;
        RECT 721.950 811.950 724.050 812.400 ;
        RECT 757.950 811.950 760.050 812.400 ;
        RECT 775.950 813.600 778.050 814.050 ;
        RECT 814.950 813.600 817.050 814.050 ;
        RECT 868.950 813.600 871.050 814.050 ;
        RECT 775.950 812.400 871.050 813.600 ;
        RECT 775.950 811.950 778.050 812.400 ;
        RECT 814.950 811.950 817.050 812.400 ;
        RECT 868.950 811.950 871.050 812.400 ;
        RECT 874.950 813.600 877.050 814.050 ;
        RECT 883.950 813.600 886.050 814.050 ;
        RECT 874.950 812.400 886.050 813.600 ;
        RECT 874.950 811.950 877.050 812.400 ;
        RECT 883.950 811.950 886.050 812.400 ;
        RECT 85.950 810.600 88.050 811.050 ;
        RECT 94.950 810.600 97.050 811.050 ;
        RECT 85.950 809.400 97.050 810.600 ;
        RECT 85.950 808.950 88.050 809.400 ;
        RECT 94.950 808.950 97.050 809.400 ;
        RECT 178.950 808.950 181.050 811.050 ;
        RECT 409.950 810.600 412.050 811.050 ;
        RECT 523.950 810.600 526.050 811.050 ;
        RECT 409.950 809.400 526.050 810.600 ;
        RECT 409.950 808.950 412.050 809.400 ;
        RECT 523.950 808.950 526.050 809.400 ;
        RECT 538.950 810.600 541.050 811.050 ;
        RECT 568.950 810.600 571.050 811.050 ;
        RECT 538.950 809.400 571.050 810.600 ;
        RECT 538.950 808.950 541.050 809.400 ;
        RECT 568.950 808.950 571.050 809.400 ;
        RECT 598.950 810.600 601.050 811.050 ;
        RECT 607.950 810.600 610.050 811.050 ;
        RECT 598.950 809.400 610.050 810.600 ;
        RECT 598.950 808.950 601.050 809.400 ;
        RECT 607.950 808.950 610.050 809.400 ;
        RECT 751.950 808.950 754.050 811.050 ;
        RECT 835.950 810.600 838.050 811.050 ;
        RECT 853.950 810.600 856.050 811.050 ;
        RECT 835.950 809.400 856.050 810.600 ;
        RECT 835.950 808.950 838.050 809.400 ;
        RECT 853.950 808.950 856.050 809.400 ;
        RECT 13.950 807.600 16.050 808.200 ;
        RECT 31.950 807.600 34.050 808.050 ;
        RECT 37.950 807.600 40.050 808.200 ;
        RECT 13.950 806.400 34.050 807.600 ;
        RECT 13.950 806.100 16.050 806.400 ;
        RECT 31.950 805.950 34.050 806.400 ;
        RECT 35.400 806.400 40.050 807.600 ;
        RECT 35.400 802.050 36.600 806.400 ;
        RECT 37.950 806.100 40.050 806.400 ;
        RECT 43.950 807.600 46.050 808.200 ;
        RECT 58.950 807.750 61.050 808.200 ;
        RECT 67.950 807.750 70.050 808.200 ;
        RECT 58.950 807.600 70.050 807.750 ;
        RECT 43.950 806.550 70.050 807.600 ;
        RECT 43.950 806.400 61.050 806.550 ;
        RECT 43.950 806.100 46.050 806.400 ;
        RECT 58.950 806.100 61.050 806.400 ;
        RECT 67.950 806.100 70.050 806.550 ;
        RECT 73.950 807.600 76.050 808.200 ;
        RECT 82.950 807.600 85.050 808.050 ;
        RECT 73.950 806.400 85.050 807.600 ;
        RECT 73.950 806.100 76.050 806.400 ;
        RECT 82.950 805.950 85.050 806.400 ;
        RECT 106.950 807.600 109.050 808.050 ;
        RECT 112.950 807.600 115.050 808.200 ;
        RECT 118.950 807.600 121.050 808.200 ;
        RECT 106.950 806.400 115.050 807.600 ;
        RECT 106.950 805.950 109.050 806.400 ;
        RECT 112.950 806.100 115.050 806.400 ;
        RECT 116.400 806.400 121.050 807.600 ;
        RECT 116.400 804.600 117.600 806.400 ;
        RECT 118.950 806.100 121.050 806.400 ;
        RECT 130.950 807.750 133.050 808.200 ;
        RECT 136.950 807.750 139.050 808.200 ;
        RECT 130.950 807.600 139.050 807.750 ;
        RECT 154.950 807.600 157.050 808.200 ;
        RECT 130.950 806.550 157.050 807.600 ;
        RECT 130.950 806.100 133.050 806.550 ;
        RECT 136.950 806.400 157.050 806.550 ;
        RECT 136.950 806.100 139.050 806.400 ;
        RECT 154.950 806.100 157.050 806.400 ;
        RECT 160.950 807.600 163.050 808.200 ;
        RECT 175.950 807.600 178.050 808.050 ;
        RECT 160.950 806.400 178.050 807.600 ;
        RECT 160.950 806.100 163.050 806.400 ;
        RECT 175.950 805.950 178.050 806.400 ;
        RECT 92.400 803.400 117.600 804.600 ;
        RECT 16.950 801.450 19.050 801.900 ;
        RECT 28.950 801.450 31.050 801.900 ;
        RECT 16.950 800.250 31.050 801.450 ;
        RECT 16.950 799.800 19.050 800.250 ;
        RECT 28.950 799.800 31.050 800.250 ;
        RECT 34.950 799.950 37.050 802.050 ;
        RECT 92.400 801.900 93.600 803.400 ;
        RECT 91.950 799.800 94.050 801.900 ;
        RECT 97.950 801.450 100.050 801.900 ;
        RECT 103.950 801.600 106.050 801.900 ;
        RECT 115.950 801.600 118.050 801.900 ;
        RECT 103.950 801.450 118.050 801.600 ;
        RECT 97.950 800.400 118.050 801.450 ;
        RECT 97.950 800.250 106.050 800.400 ;
        RECT 97.950 799.800 100.050 800.250 ;
        RECT 103.950 799.800 106.050 800.250 ;
        RECT 115.950 799.800 118.050 800.400 ;
        RECT 121.950 801.450 124.050 801.900 ;
        RECT 127.950 801.450 130.050 801.900 ;
        RECT 121.950 800.250 130.050 801.450 ;
        RECT 121.950 799.800 124.050 800.250 ;
        RECT 127.950 799.800 130.050 800.250 ;
        RECT 139.950 801.600 142.050 801.900 ;
        RECT 145.800 801.600 147.900 802.050 ;
        RECT 179.400 801.900 180.600 808.950 ;
        RECT 202.950 807.600 205.050 808.200 ;
        RECT 200.400 806.400 205.050 807.600 ;
        RECT 200.400 802.050 201.600 806.400 ;
        RECT 202.950 806.100 205.050 806.400 ;
        RECT 208.950 807.600 211.050 808.200 ;
        RECT 217.950 807.600 220.050 808.050 ;
        RECT 208.950 806.400 220.050 807.600 ;
        RECT 208.950 806.100 211.050 806.400 ;
        RECT 217.950 805.950 220.050 806.400 ;
        RECT 229.950 806.100 232.050 808.200 ;
        RECT 235.950 807.600 238.050 808.050 ;
        RECT 244.950 807.600 247.050 808.200 ;
        RECT 235.950 806.400 247.050 807.600 ;
        RECT 230.400 802.050 231.600 806.100 ;
        RECT 235.950 805.950 238.050 806.400 ;
        RECT 244.950 806.100 247.050 806.400 ;
        RECT 262.950 807.600 265.050 808.050 ;
        RECT 271.950 807.600 274.050 808.200 ;
        RECT 262.950 806.400 274.050 807.600 ;
        RECT 262.950 805.950 265.050 806.400 ;
        RECT 271.950 806.100 274.050 806.400 ;
        RECT 289.950 807.600 292.050 808.050 ;
        RECT 298.950 807.600 301.050 808.200 ;
        RECT 289.950 806.400 301.050 807.600 ;
        RECT 289.950 805.950 292.050 806.400 ;
        RECT 298.950 806.100 301.050 806.400 ;
        RECT 319.950 807.600 322.050 808.200 ;
        RECT 391.950 807.600 394.050 808.200 ;
        RECT 319.950 806.400 394.050 807.600 ;
        RECT 319.950 806.100 322.050 806.400 ;
        RECT 391.950 806.100 394.050 806.400 ;
        RECT 415.950 807.750 418.050 808.200 ;
        RECT 427.950 807.750 430.050 808.200 ;
        RECT 415.950 806.550 430.050 807.750 ;
        RECT 415.950 806.100 418.050 806.550 ;
        RECT 427.950 806.100 430.050 806.550 ;
        RECT 445.950 807.750 448.050 808.200 ;
        RECT 454.950 807.750 457.050 808.200 ;
        RECT 445.950 806.550 457.050 807.750 ;
        RECT 445.950 806.100 448.050 806.550 ;
        RECT 454.950 806.100 457.050 806.550 ;
        RECT 463.950 807.600 466.050 808.050 ;
        RECT 499.950 807.600 502.050 808.200 ;
        RECT 463.950 806.400 502.050 807.600 ;
        RECT 463.950 805.950 466.050 806.400 ;
        RECT 499.950 806.100 502.050 806.400 ;
        RECT 505.950 807.750 508.050 808.200 ;
        RECT 511.950 807.750 514.050 808.200 ;
        RECT 505.950 807.600 514.050 807.750 ;
        RECT 520.950 807.600 523.050 808.200 ;
        RECT 505.950 806.550 523.050 807.600 ;
        RECT 505.950 806.100 508.050 806.550 ;
        RECT 511.950 806.400 523.050 806.550 ;
        RECT 511.950 806.100 514.050 806.400 ;
        RECT 520.950 806.100 523.050 806.400 ;
        RECT 526.950 807.750 529.050 808.200 ;
        RECT 535.950 807.750 538.050 808.200 ;
        RECT 526.950 806.550 538.050 807.750 ;
        RECT 526.950 806.100 529.050 806.550 ;
        RECT 535.950 806.100 538.050 806.550 ;
        RECT 574.950 806.100 577.050 808.200 ;
        RECT 613.950 807.750 616.050 808.200 ;
        RECT 619.950 807.750 622.050 808.200 ;
        RECT 613.950 806.550 622.050 807.750 ;
        RECT 637.950 807.600 640.050 808.200 ;
        RECT 613.950 806.100 616.050 806.550 ;
        RECT 619.950 806.100 622.050 806.550 ;
        RECT 623.400 806.400 640.050 807.600 ;
        RECT 139.950 800.400 147.900 801.600 ;
        RECT 139.950 799.800 142.050 800.400 ;
        RECT 145.800 799.950 147.900 800.400 ;
        RECT 148.950 801.450 151.050 801.900 ;
        RECT 157.950 801.450 160.050 801.900 ;
        RECT 148.950 800.250 160.050 801.450 ;
        RECT 148.950 799.800 151.050 800.250 ;
        RECT 157.950 799.800 160.050 800.250 ;
        RECT 178.950 799.800 181.050 801.900 ;
        RECT 199.950 799.950 202.050 802.050 ;
        RECT 211.950 801.600 214.050 801.900 ;
        RECT 226.950 801.600 229.050 801.900 ;
        RECT 211.950 800.400 229.050 801.600 ;
        RECT 230.400 800.400 235.050 802.050 ;
        RECT 211.950 799.800 214.050 800.400 ;
        RECT 226.950 799.800 229.050 800.400 ;
        RECT 231.000 799.950 235.050 800.400 ;
        RECT 253.950 801.450 256.050 801.900 ;
        RECT 259.950 801.450 262.050 801.900 ;
        RECT 253.950 800.250 262.050 801.450 ;
        RECT 253.950 799.800 256.050 800.250 ;
        RECT 259.950 799.800 262.050 800.250 ;
        RECT 265.950 801.450 268.050 801.900 ;
        RECT 274.950 801.450 277.050 801.900 ;
        RECT 265.950 800.250 277.050 801.450 ;
        RECT 265.950 799.800 268.050 800.250 ;
        RECT 274.950 799.800 277.050 800.250 ;
        RECT 280.950 801.450 283.050 801.900 ;
        RECT 289.950 801.450 292.050 801.900 ;
        RECT 280.950 800.250 292.050 801.450 ;
        RECT 280.950 799.800 283.050 800.250 ;
        RECT 289.950 799.800 292.050 800.250 ;
        RECT 301.950 801.450 304.050 801.900 ;
        RECT 310.800 801.450 312.900 801.900 ;
        RECT 301.950 800.250 312.900 801.450 ;
        RECT 301.950 799.800 304.050 800.250 ;
        RECT 310.800 799.800 312.900 800.250 ;
        RECT 313.950 801.600 316.050 802.050 ;
        RECT 322.950 801.600 325.050 801.900 ;
        RECT 313.950 800.400 325.050 801.600 ;
        RECT 313.950 799.950 316.050 800.400 ;
        RECT 322.950 799.800 325.050 800.400 ;
        RECT 355.950 801.450 358.050 801.900 ;
        RECT 367.950 801.450 370.050 801.900 ;
        RECT 355.950 800.250 370.050 801.450 ;
        RECT 355.950 799.800 358.050 800.250 ;
        RECT 367.950 799.800 370.050 800.250 ;
        RECT 514.950 801.450 517.050 801.900 ;
        RECT 523.950 801.450 526.050 801.900 ;
        RECT 514.950 800.250 526.050 801.450 ;
        RECT 514.950 799.800 517.050 800.250 ;
        RECT 523.950 799.800 526.050 800.250 ;
        RECT 538.950 801.450 541.050 801.900 ;
        RECT 544.950 801.450 547.050 801.900 ;
        RECT 538.950 800.250 547.050 801.450 ;
        RECT 575.400 801.600 576.600 806.100 ;
        RECT 623.400 804.600 624.600 806.400 ;
        RECT 637.950 806.100 640.050 806.400 ;
        RECT 658.950 807.600 663.000 808.050 ;
        RECT 658.950 805.950 663.600 807.600 ;
        RECT 670.950 806.100 673.050 808.200 ;
        RECT 712.950 807.750 715.050 808.200 ;
        RECT 724.950 807.750 727.050 808.200 ;
        RECT 712.950 806.550 727.050 807.750 ;
        RECT 712.950 806.100 715.050 806.550 ;
        RECT 724.950 806.100 727.050 806.550 ;
        RECT 662.400 804.600 663.600 805.950 ;
        RECT 617.400 803.400 624.600 804.600 ;
        RECT 641.400 803.400 663.600 804.600 ;
        RECT 580.950 801.600 583.050 802.050 ;
        RECT 575.400 800.400 583.050 801.600 ;
        RECT 538.950 799.800 541.050 800.250 ;
        RECT 544.950 799.800 547.050 800.250 ;
        RECT 580.950 799.950 583.050 800.400 ;
        RECT 595.950 801.600 598.050 801.900 ;
        RECT 617.400 801.600 618.600 803.400 ;
        RECT 641.400 801.900 642.600 803.400 ;
        RECT 662.400 801.900 663.600 803.400 ;
        RECT 671.400 802.050 672.600 806.100 ;
        RECT 595.950 800.400 618.600 801.600 ;
        RECT 595.950 799.800 598.050 800.400 ;
        RECT 640.950 799.800 643.050 801.900 ;
        RECT 646.950 801.450 649.050 801.900 ;
        RECT 655.950 801.450 658.050 801.900 ;
        RECT 646.950 800.250 658.050 801.450 ;
        RECT 646.950 799.800 649.050 800.250 ;
        RECT 655.950 799.800 658.050 800.250 ;
        RECT 661.950 799.800 664.050 801.900 ;
        RECT 671.400 800.400 676.050 802.050 ;
        RECT 672.000 799.950 676.050 800.400 ;
        RECT 715.950 801.450 718.050 801.900 ;
        RECT 721.800 801.450 723.900 801.900 ;
        RECT 715.950 800.250 723.900 801.450 ;
        RECT 715.950 799.800 718.050 800.250 ;
        RECT 721.800 799.800 723.900 800.250 ;
        RECT 724.950 801.600 727.050 802.050 ;
        RECT 752.400 801.900 753.600 808.950 ;
        RECT 754.950 806.100 757.050 808.200 ;
        RECT 775.950 807.600 778.050 808.200 ;
        RECT 799.950 807.750 802.050 808.200 ;
        RECT 805.950 807.750 808.050 808.200 ;
        RECT 775.950 806.400 798.600 807.600 ;
        RECT 775.950 806.100 778.050 806.400 ;
        RECT 755.400 804.600 756.600 806.100 ;
        RECT 755.400 803.400 777.600 804.600 ;
        RECT 730.950 801.600 733.050 801.900 ;
        RECT 724.950 800.400 733.050 801.600 ;
        RECT 724.950 799.950 727.050 800.400 ;
        RECT 730.950 799.800 733.050 800.400 ;
        RECT 751.950 799.800 754.050 801.900 ;
        RECT 757.950 801.450 760.050 801.900 ;
        RECT 763.950 801.450 766.050 801.900 ;
        RECT 757.950 800.250 766.050 801.450 ;
        RECT 776.400 801.600 777.600 803.400 ;
        RECT 790.950 801.600 793.050 802.050 ;
        RECT 797.400 801.900 798.600 806.400 ;
        RECT 799.950 806.550 808.050 807.750 ;
        RECT 799.950 806.100 802.050 806.550 ;
        RECT 805.950 806.100 808.050 806.550 ;
        RECT 814.950 807.600 819.000 808.050 ;
        RECT 826.950 807.750 829.050 808.200 ;
        RECT 832.950 807.750 835.050 808.200 ;
        RECT 814.950 805.950 819.600 807.600 ;
        RECT 826.950 806.550 835.050 807.750 ;
        RECT 826.950 806.100 829.050 806.550 ;
        RECT 832.950 806.100 835.050 806.550 ;
        RECT 862.950 807.600 865.050 808.050 ;
        RECT 874.950 807.600 877.050 808.200 ;
        RECT 862.950 806.400 877.050 807.600 ;
        RECT 862.950 805.950 865.050 806.400 ;
        RECT 874.950 806.100 877.050 806.400 ;
        RECT 880.950 805.950 883.050 808.050 ;
        RECT 818.400 801.900 819.600 805.950 ;
        RECT 881.400 802.050 882.600 805.950 ;
        RECT 776.400 800.400 793.050 801.600 ;
        RECT 757.950 799.800 760.050 800.250 ;
        RECT 763.950 799.800 766.050 800.250 ;
        RECT 790.950 799.950 793.050 800.400 ;
        RECT 796.950 799.800 799.050 801.900 ;
        RECT 802.950 801.450 805.050 801.900 ;
        RECT 808.950 801.450 811.050 801.900 ;
        RECT 802.950 800.250 811.050 801.450 ;
        RECT 802.950 799.800 805.050 800.250 ;
        RECT 808.950 799.800 811.050 800.250 ;
        RECT 817.950 799.800 820.050 801.900 ;
        RECT 880.950 799.950 883.050 802.050 ;
        RECT 40.950 798.600 43.050 799.050 ;
        RECT 64.950 798.600 67.050 799.050 ;
        RECT 79.950 798.600 82.050 799.050 ;
        RECT 130.950 798.600 133.050 799.050 ;
        RECT 40.950 797.400 133.050 798.600 ;
        RECT 40.950 796.950 43.050 797.400 ;
        RECT 64.950 796.950 67.050 797.400 ;
        RECT 79.950 796.950 82.050 797.400 ;
        RECT 130.950 796.950 133.050 797.400 ;
        RECT 241.950 798.600 244.050 799.050 ;
        RECT 262.950 798.600 265.050 799.050 ;
        RECT 241.950 797.400 265.050 798.600 ;
        RECT 241.950 796.950 244.050 797.400 ;
        RECT 262.950 796.950 265.050 797.400 ;
        RECT 388.950 798.600 391.050 799.050 ;
        RECT 394.950 798.600 397.050 799.050 ;
        RECT 388.950 797.400 397.050 798.600 ;
        RECT 388.950 796.950 391.050 797.400 ;
        RECT 394.950 796.950 397.050 797.400 ;
        RECT 511.950 798.600 514.050 799.050 ;
        RECT 571.950 798.600 574.050 799.050 ;
        RECT 511.950 797.400 574.050 798.600 ;
        RECT 511.950 796.950 514.050 797.400 ;
        RECT 571.950 796.950 574.050 797.400 ;
        RECT 709.950 798.600 712.050 799.050 ;
        RECT 766.950 798.600 769.050 799.050 ;
        RECT 709.950 797.400 769.050 798.600 ;
        RECT 709.950 796.950 712.050 797.400 ;
        RECT 766.950 796.950 769.050 797.400 ;
        RECT 844.950 798.600 847.050 799.050 ;
        RECT 859.950 798.600 862.050 799.050 ;
        RECT 844.950 797.400 862.050 798.600 ;
        RECT 844.950 796.950 847.050 797.400 ;
        RECT 859.950 796.950 862.050 797.400 ;
        RECT 865.950 798.600 868.050 799.050 ;
        RECT 877.950 798.600 880.050 799.050 ;
        RECT 865.950 797.400 880.050 798.600 ;
        RECT 865.950 796.950 868.050 797.400 ;
        RECT 877.950 796.950 880.050 797.400 ;
        RECT 31.950 795.600 34.050 796.050 ;
        RECT 37.950 795.600 40.050 796.050 ;
        RECT 31.950 794.400 40.050 795.600 ;
        RECT 31.950 793.950 34.050 794.400 ;
        RECT 37.950 793.950 40.050 794.400 ;
        RECT 85.950 795.600 88.050 796.050 ;
        RECT 172.950 795.600 175.050 796.050 ;
        RECT 85.950 794.400 175.050 795.600 ;
        RECT 85.950 793.950 88.050 794.400 ;
        RECT 172.950 793.950 175.050 794.400 ;
        RECT 187.950 795.600 190.050 796.050 ;
        RECT 211.950 795.600 214.050 796.050 ;
        RECT 187.950 794.400 214.050 795.600 ;
        RECT 187.950 793.950 190.050 794.400 ;
        RECT 211.950 793.950 214.050 794.400 ;
        RECT 232.950 795.600 235.050 796.050 ;
        RECT 373.950 795.600 376.050 796.050 ;
        RECT 232.950 794.400 376.050 795.600 ;
        RECT 232.950 793.950 235.050 794.400 ;
        RECT 373.950 793.950 376.050 794.400 ;
        RECT 427.950 795.600 430.050 796.050 ;
        RECT 499.950 795.600 502.050 796.050 ;
        RECT 427.950 794.400 502.050 795.600 ;
        RECT 427.950 793.950 430.050 794.400 ;
        RECT 499.950 793.950 502.050 794.400 ;
        RECT 544.950 795.600 547.050 796.050 ;
        RECT 550.950 795.600 553.050 796.050 ;
        RECT 565.950 795.600 568.050 796.050 ;
        RECT 544.950 794.400 568.050 795.600 ;
        RECT 544.950 793.950 547.050 794.400 ;
        RECT 550.950 793.950 553.050 794.400 ;
        RECT 565.950 793.950 568.050 794.400 ;
        RECT 577.950 795.600 580.050 796.050 ;
        RECT 601.950 795.600 604.050 796.050 ;
        RECT 613.950 795.600 616.050 796.050 ;
        RECT 673.950 795.600 676.050 796.050 ;
        RECT 577.950 794.400 676.050 795.600 ;
        RECT 577.950 793.950 580.050 794.400 ;
        RECT 601.950 793.950 604.050 794.400 ;
        RECT 613.950 793.950 616.050 794.400 ;
        RECT 673.950 793.950 676.050 794.400 ;
        RECT 790.950 795.600 793.050 796.050 ;
        RECT 820.950 795.600 823.050 796.050 ;
        RECT 790.950 794.400 823.050 795.600 ;
        RECT 790.950 793.950 793.050 794.400 ;
        RECT 820.950 793.950 823.050 794.400 ;
        RECT 247.950 792.600 250.050 793.050 ;
        RECT 280.950 792.600 283.050 793.050 ;
        RECT 247.950 791.400 283.050 792.600 ;
        RECT 247.950 790.950 250.050 791.400 ;
        RECT 280.950 790.950 283.050 791.400 ;
        RECT 427.950 792.600 430.050 792.900 ;
        RECT 529.950 792.600 532.050 793.050 ;
        RECT 427.950 791.400 532.050 792.600 ;
        RECT 427.950 790.800 430.050 791.400 ;
        RECT 529.950 790.950 532.050 791.400 ;
        RECT 574.950 792.600 577.050 793.050 ;
        RECT 631.950 792.600 634.050 793.050 ;
        RECT 574.950 791.400 634.050 792.600 ;
        RECT 574.950 790.950 577.050 791.400 ;
        RECT 631.950 790.950 634.050 791.400 ;
        RECT 76.950 789.600 79.050 790.050 ;
        RECT 232.950 789.600 235.050 790.050 ;
        RECT 76.950 788.400 235.050 789.600 ;
        RECT 76.950 787.950 79.050 788.400 ;
        RECT 232.950 787.950 235.050 788.400 ;
        RECT 367.950 789.600 370.050 790.050 ;
        RECT 418.950 789.600 421.050 790.050 ;
        RECT 433.950 789.600 436.050 790.050 ;
        RECT 367.950 788.400 436.050 789.600 ;
        RECT 367.950 787.950 370.050 788.400 ;
        RECT 418.950 787.950 421.050 788.400 ;
        RECT 433.950 787.950 436.050 788.400 ;
        RECT 874.950 789.600 877.050 790.050 ;
        RECT 883.950 789.600 886.050 790.050 ;
        RECT 874.950 788.400 886.050 789.600 ;
        RECT 874.950 787.950 877.050 788.400 ;
        RECT 883.950 787.950 886.050 788.400 ;
        RECT 256.950 786.600 259.050 787.050 ;
        RECT 322.950 786.600 325.050 787.050 ;
        RECT 355.950 786.600 358.050 787.050 ;
        RECT 256.950 785.400 358.050 786.600 ;
        RECT 256.950 784.950 259.050 785.400 ;
        RECT 322.950 784.950 325.050 785.400 ;
        RECT 355.950 784.950 358.050 785.400 ;
        RECT 376.950 786.600 379.050 787.050 ;
        RECT 406.950 786.600 409.050 787.050 ;
        RECT 463.950 786.600 466.050 787.050 ;
        RECT 376.950 785.400 466.050 786.600 ;
        RECT 376.950 784.950 379.050 785.400 ;
        RECT 406.950 784.950 409.050 785.400 ;
        RECT 463.950 784.950 466.050 785.400 ;
        RECT 835.950 786.600 838.050 787.050 ;
        RECT 871.950 786.600 874.050 787.050 ;
        RECT 835.950 785.400 874.050 786.600 ;
        RECT 835.950 784.950 838.050 785.400 ;
        RECT 871.950 784.950 874.050 785.400 ;
        RECT 217.950 783.600 220.050 784.050 ;
        RECT 334.950 783.600 337.050 784.050 ;
        RECT 217.950 782.400 337.050 783.600 ;
        RECT 217.950 781.950 220.050 782.400 ;
        RECT 334.950 781.950 337.050 782.400 ;
        RECT 607.950 783.600 610.050 784.050 ;
        RECT 769.950 783.600 772.050 784.050 ;
        RECT 607.950 782.400 772.050 783.600 ;
        RECT 607.950 781.950 610.050 782.400 ;
        RECT 769.950 781.950 772.050 782.400 ;
        RECT 232.950 780.600 235.050 781.050 ;
        RECT 241.950 780.600 244.050 781.050 ;
        RECT 232.950 779.400 244.050 780.600 ;
        RECT 232.950 778.950 235.050 779.400 ;
        RECT 241.950 778.950 244.050 779.400 ;
        RECT 250.950 780.600 253.050 781.050 ;
        RECT 331.950 780.600 334.050 781.050 ;
        RECT 250.950 779.400 334.050 780.600 ;
        RECT 250.950 778.950 253.050 779.400 ;
        RECT 331.950 778.950 334.050 779.400 ;
        RECT 448.950 780.600 451.050 781.050 ;
        RECT 466.950 780.600 469.050 781.050 ;
        RECT 583.950 780.600 586.050 781.050 ;
        RECT 448.950 779.400 586.050 780.600 ;
        RECT 448.950 778.950 451.050 779.400 ;
        RECT 466.950 778.950 469.050 779.400 ;
        RECT 583.950 778.950 586.050 779.400 ;
        RECT 862.950 780.600 865.050 781.050 ;
        RECT 883.950 780.600 886.050 781.050 ;
        RECT 862.950 779.400 886.050 780.600 ;
        RECT 862.950 778.950 865.050 779.400 ;
        RECT 883.950 778.950 886.050 779.400 ;
        RECT 223.950 777.600 226.050 778.050 ;
        RECT 427.950 777.600 430.050 778.050 ;
        RECT 223.950 776.400 430.050 777.600 ;
        RECT 223.950 775.950 226.050 776.400 ;
        RECT 427.950 775.950 430.050 776.400 ;
        RECT 820.950 777.600 823.050 778.050 ;
        RECT 895.950 777.600 898.050 778.050 ;
        RECT 820.950 776.400 898.050 777.600 ;
        RECT 820.950 775.950 823.050 776.400 ;
        RECT 895.950 775.950 898.050 776.400 ;
        RECT 130.950 774.600 133.050 775.050 ;
        RECT 139.950 774.600 142.050 775.050 ;
        RECT 199.950 774.600 202.050 775.050 ;
        RECT 130.950 773.400 202.050 774.600 ;
        RECT 130.950 772.950 133.050 773.400 ;
        RECT 139.950 772.950 142.050 773.400 ;
        RECT 199.950 772.950 202.050 773.400 ;
        RECT 331.950 774.600 334.050 775.050 ;
        RECT 409.950 774.600 412.050 775.050 ;
        RECT 331.950 773.400 412.050 774.600 ;
        RECT 331.950 772.950 334.050 773.400 ;
        RECT 409.950 772.950 412.050 773.400 ;
        RECT 472.950 774.600 475.050 775.050 ;
        RECT 487.950 774.600 490.050 775.050 ;
        RECT 472.950 773.400 490.050 774.600 ;
        RECT 472.950 772.950 475.050 773.400 ;
        RECT 487.950 772.950 490.050 773.400 ;
        RECT 841.950 774.600 844.050 775.050 ;
        RECT 862.950 774.600 865.050 775.050 ;
        RECT 841.950 773.400 865.050 774.600 ;
        RECT 841.950 772.950 844.050 773.400 ;
        RECT 862.950 772.950 865.050 773.400 ;
        RECT 328.950 771.600 331.050 772.050 ;
        RECT 412.950 771.600 415.050 772.050 ;
        RECT 445.950 771.600 448.050 772.050 ;
        RECT 328.950 770.400 448.050 771.600 ;
        RECT 328.950 769.950 331.050 770.400 ;
        RECT 412.950 769.950 415.050 770.400 ;
        RECT 445.950 769.950 448.050 770.400 ;
        RECT 505.950 771.600 508.050 772.050 ;
        RECT 526.950 771.600 529.050 772.050 ;
        RECT 556.950 771.600 559.050 771.900 ;
        RECT 505.950 770.400 559.050 771.600 ;
        RECT 505.950 769.950 508.050 770.400 ;
        RECT 526.950 769.950 529.050 770.400 ;
        RECT 556.950 769.800 559.050 770.400 ;
        RECT 34.950 768.600 37.050 769.050 ;
        RECT 40.950 768.600 43.050 769.050 ;
        RECT 34.950 767.400 43.050 768.600 ;
        RECT 34.950 766.950 37.050 767.400 ;
        RECT 40.950 766.950 43.050 767.400 ;
        RECT 166.950 768.600 169.050 769.050 ;
        RECT 181.950 768.600 184.050 769.050 ;
        RECT 235.950 768.600 238.050 769.050 ;
        RECT 241.950 768.600 244.050 768.900 ;
        RECT 358.950 768.600 361.050 769.050 ;
        RECT 166.950 767.400 244.050 768.600 ;
        RECT 166.950 766.950 169.050 767.400 ;
        RECT 181.950 766.950 184.050 767.400 ;
        RECT 235.950 766.950 238.050 767.400 ;
        RECT 241.950 766.800 244.050 767.400 ;
        RECT 350.400 767.400 361.050 768.600 ;
        RECT 211.950 765.600 214.050 766.050 ;
        RECT 238.950 765.600 241.050 766.050 ;
        RECT 211.950 764.400 241.050 765.600 ;
        RECT 211.950 763.950 214.050 764.400 ;
        RECT 238.950 763.950 241.050 764.400 ;
        RECT 307.950 765.600 310.050 766.050 ;
        RECT 350.400 765.600 351.600 767.400 ;
        RECT 358.950 766.950 361.050 767.400 ;
        RECT 409.950 768.600 412.050 769.050 ;
        RECT 454.950 768.600 457.050 769.050 ;
        RECT 478.950 768.600 481.050 769.050 ;
        RECT 496.950 768.600 499.050 769.050 ;
        RECT 409.950 767.400 499.050 768.600 ;
        RECT 409.950 766.950 412.050 767.400 ;
        RECT 454.950 766.950 457.050 767.400 ;
        RECT 478.950 766.950 481.050 767.400 ;
        RECT 496.950 766.950 499.050 767.400 ;
        RECT 604.950 768.600 607.050 769.050 ;
        RECT 613.950 768.600 616.050 769.050 ;
        RECT 604.950 767.400 616.050 768.600 ;
        RECT 604.950 766.950 607.050 767.400 ;
        RECT 613.950 766.950 616.050 767.400 ;
        RECT 769.950 768.600 772.050 769.050 ;
        RECT 805.950 768.600 808.050 769.050 ;
        RECT 769.950 767.400 808.050 768.600 ;
        RECT 769.950 766.950 772.050 767.400 ;
        RECT 805.950 766.950 808.050 767.400 ;
        RECT 811.950 768.600 814.050 769.050 ;
        RECT 826.950 768.600 829.050 769.050 ;
        RECT 811.950 767.400 829.050 768.600 ;
        RECT 811.950 766.950 814.050 767.400 ;
        RECT 826.950 766.950 829.050 767.400 ;
        RECT 868.950 768.600 871.050 769.050 ;
        RECT 877.950 768.600 880.050 769.050 ;
        RECT 868.950 767.400 880.050 768.600 ;
        RECT 868.950 766.950 871.050 767.400 ;
        RECT 877.950 766.950 880.050 767.400 ;
        RECT 307.950 764.400 351.600 765.600 ;
        RECT 499.950 765.600 502.050 766.050 ;
        RECT 520.950 765.600 523.050 766.050 ;
        RECT 499.950 764.400 523.050 765.600 ;
        RECT 307.950 763.950 310.050 764.400 ;
        RECT 499.950 763.950 502.050 764.400 ;
        RECT 520.950 763.950 523.050 764.400 ;
        RECT 595.950 765.600 598.050 766.050 ;
        RECT 619.950 765.600 622.050 766.050 ;
        RECT 595.950 764.400 622.050 765.600 ;
        RECT 595.950 763.950 598.050 764.400 ;
        RECT 619.950 763.950 622.050 764.400 ;
        RECT 847.950 765.600 850.050 766.050 ;
        RECT 880.950 765.600 883.050 766.050 ;
        RECT 847.950 764.400 883.050 765.600 ;
        RECT 847.950 763.950 850.050 764.400 ;
        RECT 13.950 762.600 16.050 763.200 ;
        RECT 34.950 762.600 37.050 763.200 ;
        RECT 13.950 761.400 37.050 762.600 ;
        RECT 13.950 761.100 16.050 761.400 ;
        RECT 34.950 761.100 37.050 761.400 ;
        RECT 67.950 762.750 70.050 763.200 ;
        RECT 88.950 762.750 91.050 763.200 ;
        RECT 67.950 761.550 91.050 762.750 ;
        RECT 67.950 761.100 70.050 761.550 ;
        RECT 88.950 761.100 91.050 761.550 ;
        RECT 97.950 761.100 100.050 763.200 ;
        RECT 103.950 762.750 106.050 763.200 ;
        RECT 109.950 762.750 112.050 763.200 ;
        RECT 103.950 761.550 112.050 762.750 ;
        RECT 121.950 762.600 124.050 763.200 ;
        RECT 148.950 762.600 151.050 763.050 ;
        RECT 103.950 761.100 106.050 761.550 ;
        RECT 109.950 761.100 112.050 761.550 ;
        RECT 113.400 761.400 151.050 762.600 ;
        RECT 98.400 759.600 99.600 761.100 ;
        RECT 113.400 759.600 114.600 761.400 ;
        RECT 121.950 761.100 124.050 761.400 ;
        RECT 148.950 760.950 151.050 761.400 ;
        RECT 160.950 762.600 163.050 763.200 ;
        RECT 187.950 762.600 190.050 763.200 ;
        RECT 205.950 762.600 208.050 763.050 ;
        RECT 160.950 761.400 208.050 762.600 ;
        RECT 160.950 761.100 163.050 761.400 ;
        RECT 187.950 761.100 190.050 761.400 ;
        RECT 205.950 760.950 208.050 761.400 ;
        RECT 274.950 762.750 277.050 763.200 ;
        RECT 280.950 762.750 283.050 763.200 ;
        RECT 274.950 761.550 283.050 762.750 ;
        RECT 274.950 761.100 277.050 761.550 ;
        RECT 280.950 761.100 283.050 761.550 ;
        RECT 286.950 762.750 289.050 763.200 ;
        RECT 295.950 762.750 298.050 763.200 ;
        RECT 286.950 761.550 298.050 762.750 ;
        RECT 286.950 761.100 289.050 761.550 ;
        RECT 295.950 761.100 298.050 761.550 ;
        RECT 346.950 762.750 349.050 763.200 ;
        RECT 352.950 762.750 355.050 763.200 ;
        RECT 346.950 761.550 355.050 762.750 ;
        RECT 346.950 761.100 349.050 761.550 ;
        RECT 352.950 761.100 355.050 761.550 ;
        RECT 382.950 762.600 385.050 763.200 ;
        RECT 400.950 762.750 403.050 763.200 ;
        RECT 418.950 762.750 421.050 763.200 ;
        RECT 400.950 762.600 421.050 762.750 ;
        RECT 382.950 761.550 421.050 762.600 ;
        RECT 382.950 761.400 403.050 761.550 ;
        RECT 382.950 761.100 385.050 761.400 ;
        RECT 400.950 761.100 403.050 761.400 ;
        RECT 418.950 761.100 421.050 761.550 ;
        RECT 433.950 762.600 436.050 763.200 ;
        RECT 448.950 762.600 451.050 763.200 ;
        RECT 472.950 762.600 475.050 763.200 ;
        RECT 553.950 762.600 556.050 763.200 ;
        RECT 571.950 762.600 574.050 763.200 ;
        RECT 634.950 762.600 637.050 763.200 ;
        RECT 433.950 761.400 451.050 762.600 ;
        RECT 433.950 761.100 436.050 761.400 ;
        RECT 448.950 761.100 451.050 761.400 ;
        RECT 452.400 761.400 501.600 762.600 ;
        RECT 71.400 758.400 114.600 759.600 ;
        RECT 71.400 756.900 72.600 758.400 ;
        RECT 43.950 756.450 46.050 756.900 ;
        RECT 52.950 756.450 55.050 756.900 ;
        RECT 43.950 755.250 55.050 756.450 ;
        RECT 43.950 754.800 46.050 755.250 ;
        RECT 52.950 754.800 55.050 755.250 ;
        RECT 70.950 754.800 73.050 756.900 ;
        RECT 85.950 756.600 88.050 757.050 ;
        RECT 100.950 756.600 103.050 756.900 ;
        RECT 85.950 755.400 103.050 756.600 ;
        RECT 85.950 754.950 88.050 755.400 ;
        RECT 100.950 754.800 103.050 755.400 ;
        RECT 118.950 756.450 121.050 756.900 ;
        RECT 130.950 756.450 133.050 756.900 ;
        RECT 118.950 755.250 133.050 756.450 ;
        RECT 118.950 754.800 121.050 755.250 ;
        RECT 130.950 754.800 133.050 755.250 ;
        RECT 163.950 756.600 166.050 756.900 ;
        RECT 208.950 756.600 211.050 756.900 ;
        RECT 163.950 755.400 211.050 756.600 ;
        RECT 163.950 754.800 166.050 755.400 ;
        RECT 208.950 754.800 211.050 755.400 ;
        RECT 214.950 756.600 217.050 756.900 ;
        RECT 223.950 756.600 226.050 757.050 ;
        RECT 214.950 755.400 226.050 756.600 ;
        RECT 214.950 754.800 217.050 755.400 ;
        RECT 223.950 754.950 226.050 755.400 ;
        RECT 235.950 756.600 238.050 756.900 ;
        RECT 250.950 756.600 253.050 757.050 ;
        RECT 235.950 755.400 253.050 756.600 ;
        RECT 235.950 754.800 238.050 755.400 ;
        RECT 250.950 754.950 253.050 755.400 ;
        RECT 289.950 756.600 292.050 756.900 ;
        RECT 304.950 756.600 307.050 756.900 ;
        RECT 289.950 755.400 307.050 756.600 ;
        RECT 289.950 754.800 292.050 755.400 ;
        RECT 304.950 754.800 307.050 755.400 ;
        RECT 331.950 756.600 334.050 756.900 ;
        RECT 355.950 756.600 358.050 756.900 ;
        RECT 331.950 755.400 358.050 756.600 ;
        RECT 331.950 754.800 334.050 755.400 ;
        RECT 355.950 754.800 358.050 755.400 ;
        RECT 361.950 756.600 364.050 756.900 ;
        RECT 367.950 756.600 370.050 757.050 ;
        RECT 452.400 756.900 453.600 761.400 ;
        RECT 472.950 761.100 475.050 761.400 ;
        RECT 500.400 759.600 501.600 761.400 ;
        RECT 553.950 761.400 637.050 762.600 ;
        RECT 553.950 761.100 556.050 761.400 ;
        RECT 571.950 761.100 574.050 761.400 ;
        RECT 634.950 761.100 637.050 761.400 ;
        RECT 655.950 762.750 658.050 763.200 ;
        RECT 664.950 762.750 667.050 763.200 ;
        RECT 655.950 761.550 667.050 762.750 ;
        RECT 655.950 761.100 658.050 761.550 ;
        RECT 664.950 761.100 667.050 761.550 ;
        RECT 676.950 762.750 679.050 763.200 ;
        RECT 685.950 762.750 688.050 763.200 ;
        RECT 676.950 761.550 688.050 762.750 ;
        RECT 676.950 761.100 679.050 761.550 ;
        RECT 685.950 761.100 688.050 761.550 ;
        RECT 691.950 762.600 694.050 763.200 ;
        RECT 712.950 762.600 715.050 763.200 ;
        RECT 691.950 761.400 715.050 762.600 ;
        RECT 691.950 761.100 694.050 761.400 ;
        RECT 712.950 761.100 715.050 761.400 ;
        RECT 724.950 762.600 727.050 763.050 ;
        RECT 733.950 762.600 736.050 763.200 ;
        RECT 724.950 761.400 736.050 762.600 ;
        RECT 724.950 760.950 727.050 761.400 ;
        RECT 733.950 761.100 736.050 761.400 ;
        RECT 739.950 762.600 742.050 763.200 ;
        RECT 748.950 762.600 751.050 763.050 ;
        RECT 739.950 761.400 751.050 762.600 ;
        RECT 739.950 761.100 742.050 761.400 ;
        RECT 748.950 760.950 751.050 761.400 ;
        RECT 760.950 762.600 763.050 763.200 ;
        RECT 778.950 762.600 781.050 763.200 ;
        RECT 760.950 761.400 781.050 762.600 ;
        RECT 760.950 761.100 763.050 761.400 ;
        RECT 778.950 761.100 781.050 761.400 ;
        RECT 799.950 762.750 802.050 763.200 ;
        RECT 811.950 762.750 814.050 763.200 ;
        RECT 799.950 761.550 814.050 762.750 ;
        RECT 868.950 762.600 871.050 763.200 ;
        RECT 799.950 761.100 802.050 761.550 ;
        RECT 811.950 761.100 814.050 761.550 ;
        RECT 851.400 761.400 871.050 762.600 ;
        RECT 500.400 758.400 528.600 759.600 ;
        RECT 361.950 755.400 370.050 756.600 ;
        RECT 361.950 754.800 364.050 755.400 ;
        RECT 367.950 754.950 370.050 755.400 ;
        RECT 403.950 756.600 406.050 756.900 ;
        RECT 424.950 756.600 427.050 756.900 ;
        RECT 403.950 755.400 427.050 756.600 ;
        RECT 403.950 754.800 406.050 755.400 ;
        RECT 424.950 754.800 427.050 755.400 ;
        RECT 430.950 756.600 433.050 756.900 ;
        RECT 451.950 756.600 454.050 756.900 ;
        RECT 430.950 755.400 454.050 756.600 ;
        RECT 430.950 754.800 433.050 755.400 ;
        RECT 451.950 754.800 454.050 755.400 ;
        RECT 466.950 756.450 469.050 756.900 ;
        RECT 475.950 756.450 478.050 756.900 ;
        RECT 466.950 755.250 478.050 756.450 ;
        RECT 466.950 754.800 469.050 755.250 ;
        RECT 475.950 754.800 478.050 755.250 ;
        RECT 490.950 756.600 493.050 757.050 ;
        RECT 496.950 756.600 499.050 756.900 ;
        RECT 490.950 755.400 499.050 756.600 ;
        RECT 527.400 756.600 528.600 758.400 ;
        RECT 568.950 756.600 571.050 756.900 ;
        RECT 527.400 755.400 571.050 756.600 ;
        RECT 490.950 754.950 493.050 755.400 ;
        RECT 496.950 754.800 499.050 755.400 ;
        RECT 568.950 754.800 571.050 755.400 ;
        RECT 574.950 756.600 577.050 756.900 ;
        RECT 628.950 756.600 631.050 756.900 ;
        RECT 574.950 756.450 631.050 756.600 ;
        RECT 637.950 756.450 640.050 756.900 ;
        RECT 574.950 755.400 640.050 756.450 ;
        RECT 574.950 754.800 577.050 755.400 ;
        RECT 628.950 755.250 640.050 755.400 ;
        RECT 628.950 754.800 631.050 755.250 ;
        RECT 637.950 754.800 640.050 755.250 ;
        RECT 643.950 756.600 646.050 756.900 ;
        RECT 682.950 756.600 685.050 757.050 ;
        RECT 643.950 755.400 685.050 756.600 ;
        RECT 643.950 754.800 646.050 755.400 ;
        RECT 682.950 754.950 685.050 755.400 ;
        RECT 748.950 756.450 751.050 756.900 ;
        RECT 757.950 756.450 760.050 756.900 ;
        RECT 748.950 755.250 760.050 756.450 ;
        RECT 748.950 754.800 751.050 755.250 ;
        RECT 757.950 754.800 760.050 755.250 ;
        RECT 832.950 756.600 835.050 757.050 ;
        RECT 838.950 756.600 841.050 757.050 ;
        RECT 851.400 756.900 852.600 761.400 ;
        RECT 868.950 761.100 871.050 761.400 ;
        RECT 872.400 756.900 873.600 764.400 ;
        RECT 880.950 763.950 883.050 764.400 ;
        RECT 832.950 755.400 841.050 756.600 ;
        RECT 832.950 754.950 835.050 755.400 ;
        RECT 838.950 754.950 841.050 755.400 ;
        RECT 850.950 754.800 853.050 756.900 ;
        RECT 871.950 754.800 874.050 756.900 ;
        RECT 79.950 753.600 82.050 754.050 ;
        RECT 124.950 753.600 127.050 754.050 ;
        RECT 79.950 752.400 127.050 753.600 ;
        RECT 79.950 751.950 82.050 752.400 ;
        RECT 124.950 751.950 127.050 752.400 ;
        RECT 259.950 753.600 262.050 754.050 ;
        RECT 274.950 753.600 277.050 754.050 ;
        RECT 280.800 753.600 282.900 754.050 ;
        RECT 259.950 752.400 282.900 753.600 ;
        RECT 259.950 751.950 262.050 752.400 ;
        RECT 274.950 751.950 277.050 752.400 ;
        RECT 280.800 751.950 282.900 752.400 ;
        RECT 283.950 753.600 286.050 754.050 ;
        RECT 325.950 753.600 328.050 754.050 ;
        RECT 283.950 752.400 328.050 753.600 ;
        RECT 283.950 751.950 286.050 752.400 ;
        RECT 325.950 751.950 328.050 752.400 ;
        RECT 385.950 753.600 388.050 754.050 ;
        RECT 397.950 753.600 400.050 754.050 ;
        RECT 486.000 753.600 490.050 754.050 ;
        RECT 385.950 752.400 400.050 753.600 ;
        RECT 385.950 751.950 388.050 752.400 ;
        RECT 397.950 751.950 400.050 752.400 ;
        RECT 485.400 751.950 490.050 753.600 ;
        RECT 502.950 753.600 505.050 754.050 ;
        RECT 523.950 753.600 526.050 754.050 ;
        RECT 502.950 752.400 526.050 753.600 ;
        RECT 502.950 751.950 505.050 752.400 ;
        RECT 523.950 751.950 526.050 752.400 ;
        RECT 721.950 753.600 724.050 754.050 ;
        RECT 736.950 753.600 739.050 754.050 ;
        RECT 781.950 753.600 784.050 754.050 ;
        RECT 796.950 753.600 799.050 754.050 ;
        RECT 721.950 752.400 799.050 753.600 ;
        RECT 721.950 751.950 724.050 752.400 ;
        RECT 736.950 751.950 739.050 752.400 ;
        RECT 781.950 751.950 784.050 752.400 ;
        RECT 796.950 751.950 799.050 752.400 ;
        RECT 136.950 750.600 139.050 751.050 ;
        RECT 145.950 750.600 148.050 751.050 ;
        RECT 119.400 749.400 148.050 750.600 ;
        RECT 37.950 747.600 40.050 748.050 ;
        RECT 119.400 747.600 120.600 749.400 ;
        RECT 136.950 748.950 139.050 749.400 ;
        RECT 145.950 748.950 148.050 749.400 ;
        RECT 184.950 750.600 187.050 751.050 ;
        RECT 229.950 750.600 232.050 751.050 ;
        RECT 184.950 749.400 232.050 750.600 ;
        RECT 184.950 748.950 187.050 749.400 ;
        RECT 229.950 748.950 232.050 749.400 ;
        RECT 346.950 750.600 349.050 751.050 ;
        RECT 415.950 750.600 418.050 751.050 ;
        RECT 346.950 749.400 418.050 750.600 ;
        RECT 346.950 748.950 349.050 749.400 ;
        RECT 415.950 748.950 418.050 749.400 ;
        RECT 478.950 750.600 481.050 751.050 ;
        RECT 485.400 750.600 486.600 751.950 ;
        RECT 478.950 749.400 486.600 750.600 ;
        RECT 526.950 750.600 529.050 751.050 ;
        RECT 541.950 750.600 544.050 751.050 ;
        RECT 526.950 749.400 544.050 750.600 ;
        RECT 478.950 748.950 481.050 749.400 ;
        RECT 526.950 748.950 529.050 749.400 ;
        RECT 541.950 748.950 544.050 749.400 ;
        RECT 550.950 750.600 553.050 751.050 ;
        RECT 565.950 750.600 568.050 751.050 ;
        RECT 592.950 750.600 595.050 751.050 ;
        RECT 550.950 749.400 595.050 750.600 ;
        RECT 550.950 748.950 553.050 749.400 ;
        RECT 565.950 748.950 568.050 749.400 ;
        RECT 592.950 748.950 595.050 749.400 ;
        RECT 616.950 750.600 619.050 751.050 ;
        RECT 661.950 750.600 664.050 751.050 ;
        RECT 616.950 749.400 664.050 750.600 ;
        RECT 616.950 748.950 619.050 749.400 ;
        RECT 661.950 748.950 664.050 749.400 ;
        RECT 685.950 750.600 688.050 751.050 ;
        RECT 700.950 750.600 703.050 751.050 ;
        RECT 715.950 750.600 718.050 751.050 ;
        RECT 685.950 749.400 718.050 750.600 ;
        RECT 685.950 748.950 688.050 749.400 ;
        RECT 700.950 748.950 703.050 749.400 ;
        RECT 715.950 748.950 718.050 749.400 ;
        RECT 724.950 750.600 727.050 751.050 ;
        RECT 730.950 750.600 733.050 751.050 ;
        RECT 724.950 749.400 733.050 750.600 ;
        RECT 724.950 748.950 727.050 749.400 ;
        RECT 730.950 748.950 733.050 749.400 ;
        RECT 763.950 750.600 766.050 751.050 ;
        RECT 769.950 750.600 772.050 751.050 ;
        RECT 763.950 749.400 772.050 750.600 ;
        RECT 763.950 748.950 766.050 749.400 ;
        RECT 769.950 748.950 772.050 749.400 ;
        RECT 829.950 750.600 832.050 751.050 ;
        RECT 844.950 750.600 847.050 751.050 ;
        RECT 829.950 749.400 847.050 750.600 ;
        RECT 829.950 748.950 832.050 749.400 ;
        RECT 844.950 748.950 847.050 749.400 ;
        RECT 37.950 746.400 120.600 747.600 ;
        RECT 148.950 747.600 151.050 748.050 ;
        RECT 283.950 747.600 286.050 748.050 ;
        RECT 148.950 746.400 286.050 747.600 ;
        RECT 37.950 745.950 40.050 746.400 ;
        RECT 148.950 745.950 151.050 746.400 ;
        RECT 283.950 745.950 286.050 746.400 ;
        RECT 355.950 747.600 358.050 748.050 ;
        RECT 391.950 747.600 394.050 748.050 ;
        RECT 355.950 746.400 394.050 747.600 ;
        RECT 355.950 745.950 358.050 746.400 ;
        RECT 391.950 745.950 394.050 746.400 ;
        RECT 418.950 747.600 421.050 748.050 ;
        RECT 487.950 747.600 490.050 748.050 ;
        RECT 418.950 746.400 490.050 747.600 ;
        RECT 418.950 745.950 421.050 746.400 ;
        RECT 487.950 745.950 490.050 746.400 ;
        RECT 634.950 747.600 637.050 748.050 ;
        RECT 649.950 747.600 652.050 748.050 ;
        RECT 634.950 746.400 652.050 747.600 ;
        RECT 634.950 745.950 637.050 746.400 ;
        RECT 649.950 745.950 652.050 746.400 ;
        RECT 682.950 747.600 685.050 748.050 ;
        RECT 736.950 747.600 739.050 748.050 ;
        RECT 682.950 746.400 739.050 747.600 ;
        RECT 682.950 745.950 685.050 746.400 ;
        RECT 736.950 745.950 739.050 746.400 ;
        RECT 127.950 744.600 130.050 745.050 ;
        RECT 199.950 744.600 202.050 745.050 ;
        RECT 127.950 743.400 202.050 744.600 ;
        RECT 127.950 742.950 130.050 743.400 ;
        RECT 199.950 742.950 202.050 743.400 ;
        RECT 223.950 744.600 226.050 745.050 ;
        RECT 277.950 744.600 280.050 745.050 ;
        RECT 223.950 743.400 280.050 744.600 ;
        RECT 223.950 742.950 226.050 743.400 ;
        RECT 277.950 742.950 280.050 743.400 ;
        RECT 415.950 744.600 418.050 745.050 ;
        RECT 550.950 744.600 553.050 745.050 ;
        RECT 415.950 743.400 553.050 744.600 ;
        RECT 415.950 742.950 418.050 743.400 ;
        RECT 550.950 742.950 553.050 743.400 ;
        RECT 562.950 744.600 565.050 745.050 ;
        RECT 568.950 744.600 571.050 745.050 ;
        RECT 562.950 743.400 571.050 744.600 ;
        RECT 562.950 742.950 565.050 743.400 ;
        RECT 568.950 742.950 571.050 743.400 ;
        RECT 637.950 744.600 640.050 745.050 ;
        RECT 646.950 744.600 649.050 745.050 ;
        RECT 637.950 743.400 649.050 744.600 ;
        RECT 637.950 742.950 640.050 743.400 ;
        RECT 646.950 742.950 649.050 743.400 ;
        RECT 658.950 744.600 661.050 745.050 ;
        RECT 688.950 744.600 691.050 745.050 ;
        RECT 658.950 743.400 691.050 744.600 ;
        RECT 658.950 742.950 661.050 743.400 ;
        RECT 688.950 742.950 691.050 743.400 ;
        RECT 703.950 744.600 706.050 745.050 ;
        RECT 709.950 744.600 712.050 745.050 ;
        RECT 703.950 743.400 712.050 744.600 ;
        RECT 703.950 742.950 706.050 743.400 ;
        RECT 709.950 742.950 712.050 743.400 ;
        RECT 16.950 741.600 19.050 742.050 ;
        RECT 58.950 741.600 61.050 742.050 ;
        RECT 16.950 740.400 61.050 741.600 ;
        RECT 16.950 739.950 19.050 740.400 ;
        RECT 58.950 739.950 61.050 740.400 ;
        RECT 142.950 741.600 145.050 742.050 ;
        RECT 160.950 741.600 163.050 742.050 ;
        RECT 142.950 740.400 163.050 741.600 ;
        RECT 142.950 739.950 145.050 740.400 ;
        RECT 160.950 739.950 163.050 740.400 ;
        RECT 280.950 741.600 283.050 742.050 ;
        RECT 340.950 741.600 343.050 742.050 ;
        RECT 280.950 740.400 343.050 741.600 ;
        RECT 280.950 739.950 283.050 740.400 ;
        RECT 340.950 739.950 343.050 740.400 ;
        RECT 379.950 741.600 382.050 742.050 ;
        RECT 403.950 741.600 406.050 742.050 ;
        RECT 379.950 740.400 406.050 741.600 ;
        RECT 379.950 739.950 382.050 740.400 ;
        RECT 403.950 739.950 406.050 740.400 ;
        RECT 481.950 741.600 484.050 742.050 ;
        RECT 499.950 741.600 502.050 742.050 ;
        RECT 481.950 740.400 502.050 741.600 ;
        RECT 481.950 739.950 484.050 740.400 ;
        RECT 499.950 739.950 502.050 740.400 ;
        RECT 505.950 741.600 508.050 742.050 ;
        RECT 538.950 741.600 541.050 742.050 ;
        RECT 547.950 741.600 550.050 742.050 ;
        RECT 643.950 741.600 646.050 742.050 ;
        RECT 505.950 740.400 550.050 741.600 ;
        RECT 505.950 739.950 508.050 740.400 ;
        RECT 538.950 739.950 541.050 740.400 ;
        RECT 547.950 739.950 550.050 740.400 ;
        RECT 566.400 740.400 646.050 741.600 ;
        RECT 566.400 739.050 567.600 740.400 ;
        RECT 643.950 739.950 646.050 740.400 ;
        RECT 88.950 738.600 91.050 739.050 ;
        RECT 94.950 738.600 97.050 739.050 ;
        RECT 169.950 738.600 172.050 739.050 ;
        RECT 88.950 737.400 172.050 738.600 ;
        RECT 88.950 736.950 91.050 737.400 ;
        RECT 94.950 736.950 97.050 737.400 ;
        RECT 169.950 736.950 172.050 737.400 ;
        RECT 235.950 738.600 238.050 739.050 ;
        RECT 271.950 738.600 274.050 739.050 ;
        RECT 235.950 737.400 274.050 738.600 ;
        RECT 235.950 736.950 238.050 737.400 ;
        RECT 271.950 736.950 274.050 737.400 ;
        RECT 310.950 738.600 313.050 739.050 ;
        RECT 346.950 738.600 349.050 739.050 ;
        RECT 310.950 737.400 349.050 738.600 ;
        RECT 310.950 736.950 313.050 737.400 ;
        RECT 346.950 736.950 349.050 737.400 ;
        RECT 379.950 738.600 382.050 738.900 ;
        RECT 394.950 738.600 397.050 739.050 ;
        RECT 379.950 737.400 397.050 738.600 ;
        RECT 379.950 736.800 382.050 737.400 ;
        RECT 394.950 736.950 397.050 737.400 ;
        RECT 406.950 738.600 409.050 739.050 ;
        RECT 418.950 738.600 421.050 739.050 ;
        RECT 406.950 737.400 421.050 738.600 ;
        RECT 406.950 736.950 409.050 737.400 ;
        RECT 418.950 736.950 421.050 737.400 ;
        RECT 454.950 738.600 457.050 739.050 ;
        RECT 463.950 738.600 466.050 739.050 ;
        RECT 454.950 737.400 466.050 738.600 ;
        RECT 454.950 736.950 457.050 737.400 ;
        RECT 463.950 736.950 466.050 737.400 ;
        RECT 469.950 738.600 472.050 739.050 ;
        RECT 502.950 738.600 505.050 739.050 ;
        RECT 514.950 738.600 517.050 739.050 ;
        RECT 469.950 737.400 517.050 738.600 ;
        RECT 469.950 736.950 472.050 737.400 ;
        RECT 502.950 736.950 505.050 737.400 ;
        RECT 514.950 736.950 517.050 737.400 ;
        RECT 562.950 737.400 567.600 739.050 ;
        RECT 604.950 738.600 607.050 739.050 ;
        RECT 613.950 738.600 616.050 739.050 ;
        RECT 604.950 737.400 616.050 738.600 ;
        RECT 562.950 736.950 567.000 737.400 ;
        RECT 604.950 736.950 607.050 737.400 ;
        RECT 613.950 736.950 616.050 737.400 ;
        RECT 640.950 738.600 643.050 739.050 ;
        RECT 673.950 738.600 676.050 739.050 ;
        RECT 640.950 737.400 676.050 738.600 ;
        RECT 640.950 736.950 643.050 737.400 ;
        RECT 673.950 736.950 676.050 737.400 ;
        RECT 724.950 738.600 727.050 739.050 ;
        RECT 757.950 738.600 760.050 739.050 ;
        RECT 772.950 738.600 775.050 739.050 ;
        RECT 724.950 737.400 775.050 738.600 ;
        RECT 724.950 736.950 727.050 737.400 ;
        RECT 757.950 736.950 760.050 737.400 ;
        RECT 772.950 736.950 775.050 737.400 ;
        RECT 811.950 738.600 814.050 739.050 ;
        RECT 823.950 738.600 826.050 739.050 ;
        RECT 811.950 737.400 826.050 738.600 ;
        RECT 811.950 736.950 814.050 737.400 ;
        RECT 823.950 736.950 826.050 737.400 ;
        RECT 838.950 738.600 841.050 739.050 ;
        RECT 865.950 738.600 868.050 739.050 ;
        RECT 838.950 737.400 868.050 738.600 ;
        RECT 838.950 736.950 841.050 737.400 ;
        RECT 865.950 736.950 868.050 737.400 ;
        RECT 73.950 735.600 76.050 736.050 ;
        RECT 97.950 735.600 100.050 736.050 ;
        RECT 112.950 735.600 115.050 736.050 ;
        RECT 73.950 734.400 115.050 735.600 ;
        RECT 73.950 733.950 76.050 734.400 ;
        RECT 97.950 733.950 100.050 734.400 ;
        RECT 112.950 733.950 115.050 734.400 ;
        RECT 190.950 735.600 193.050 736.050 ;
        RECT 223.950 735.600 226.050 736.050 ;
        RECT 190.950 734.400 226.050 735.600 ;
        RECT 190.950 733.950 193.050 734.400 ;
        RECT 223.950 733.950 226.050 734.400 ;
        RECT 280.950 735.600 283.050 736.050 ;
        RECT 289.950 735.600 292.050 736.050 ;
        RECT 280.950 734.400 292.050 735.600 ;
        RECT 280.950 733.950 283.050 734.400 ;
        RECT 289.950 733.950 292.050 734.400 ;
        RECT 529.950 735.600 532.050 736.050 ;
        RECT 541.950 735.600 544.050 736.050 ;
        RECT 529.950 734.400 544.050 735.600 ;
        RECT 529.950 733.950 532.050 734.400 ;
        RECT 541.950 733.950 544.050 734.400 ;
        RECT 547.950 735.600 550.050 736.050 ;
        RECT 559.950 735.600 562.050 736.050 ;
        RECT 547.950 734.400 562.050 735.600 ;
        RECT 547.950 733.950 550.050 734.400 ;
        RECT 559.950 733.950 562.050 734.400 ;
        RECT 649.950 735.600 652.050 736.050 ;
        RECT 667.950 735.600 670.050 736.050 ;
        RECT 649.950 734.400 670.050 735.600 ;
        RECT 649.950 733.950 652.050 734.400 ;
        RECT 667.950 733.950 670.050 734.400 ;
        RECT 676.950 735.600 679.050 736.050 ;
        RECT 682.950 735.600 685.050 736.050 ;
        RECT 676.950 734.400 685.050 735.600 ;
        RECT 676.950 733.950 679.050 734.400 ;
        RECT 682.950 733.950 685.050 734.400 ;
        RECT 688.950 735.600 691.050 736.050 ;
        RECT 694.950 735.600 697.050 736.050 ;
        RECT 688.950 734.400 697.050 735.600 ;
        RECT 688.950 733.950 691.050 734.400 ;
        RECT 694.950 733.950 697.050 734.400 ;
        RECT 766.950 735.600 769.050 736.050 ;
        RECT 787.950 735.600 790.050 736.050 ;
        RECT 766.950 734.400 790.050 735.600 ;
        RECT 766.950 733.950 769.050 734.400 ;
        RECT 787.950 733.950 790.050 734.400 ;
        RECT 19.950 732.600 22.050 733.050 ;
        RECT 25.950 732.600 28.050 733.050 ;
        RECT 19.950 731.400 28.050 732.600 ;
        RECT 19.950 730.950 22.050 731.400 ;
        RECT 25.950 730.950 28.050 731.400 ;
        RECT 82.950 732.600 85.050 733.050 ;
        RECT 88.950 732.600 91.050 733.050 ;
        RECT 82.950 731.400 91.050 732.600 ;
        RECT 82.950 730.950 85.050 731.400 ;
        RECT 88.950 730.950 91.050 731.400 ;
        RECT 244.950 732.600 247.050 733.050 ;
        RECT 265.950 732.600 268.050 733.050 ;
        RECT 244.950 731.400 268.050 732.600 ;
        RECT 244.950 730.950 247.050 731.400 ;
        RECT 265.950 730.950 268.050 731.400 ;
        RECT 277.950 732.600 280.050 733.050 ;
        RECT 319.950 732.600 322.050 733.050 ;
        RECT 277.950 731.400 322.050 732.600 ;
        RECT 277.950 730.950 280.050 731.400 ;
        RECT 319.950 730.950 322.050 731.400 ;
        RECT 430.950 732.600 433.050 733.050 ;
        RECT 442.950 732.600 445.050 733.050 ;
        RECT 430.950 731.400 445.050 732.600 ;
        RECT 430.950 730.950 433.050 731.400 ;
        RECT 442.950 730.950 445.050 731.400 ;
        RECT 457.950 732.600 460.050 733.050 ;
        RECT 493.950 732.600 496.050 733.050 ;
        RECT 520.950 732.600 523.050 733.050 ;
        RECT 457.950 731.400 471.600 732.600 ;
        RECT 457.950 730.950 460.050 731.400 ;
        RECT 470.400 730.200 471.600 731.400 ;
        RECT 493.950 731.400 523.050 732.600 ;
        RECT 493.950 730.950 496.050 731.400 ;
        RECT 520.950 730.950 523.050 731.400 ;
        RECT 610.950 732.600 613.050 733.050 ;
        RECT 616.950 732.600 619.050 733.050 ;
        RECT 610.950 731.400 619.050 732.600 ;
        RECT 610.950 730.950 613.050 731.400 ;
        RECT 616.950 730.950 619.050 731.400 ;
        RECT 673.950 732.600 676.050 733.050 ;
        RECT 703.950 732.600 706.050 733.050 ;
        RECT 723.000 732.600 727.050 733.050 ;
        RECT 802.950 732.600 805.050 733.050 ;
        RECT 817.950 732.600 820.050 733.050 ;
        RECT 673.950 731.400 706.050 732.600 ;
        RECT 673.950 730.950 676.050 731.400 ;
        RECT 703.950 730.950 706.050 731.400 ;
        RECT 722.400 730.950 727.050 732.600 ;
        RECT 758.400 731.400 820.050 732.600 ;
        RECT 22.950 727.950 25.050 730.050 ;
        RECT 103.950 729.600 106.050 730.200 ;
        RECT 112.950 729.600 115.050 730.050 ;
        RECT 103.950 728.400 115.050 729.600 ;
        RECT 103.950 728.100 106.050 728.400 ;
        RECT 112.950 727.950 115.050 728.400 ;
        RECT 151.950 729.600 154.050 730.200 ;
        RECT 175.950 729.600 178.050 730.200 ;
        RECT 205.950 729.600 208.050 730.050 ;
        RECT 217.950 729.600 220.050 730.200 ;
        RECT 247.950 729.600 250.050 730.200 ;
        RECT 151.950 728.400 220.050 729.600 ;
        RECT 151.950 728.100 154.050 728.400 ;
        RECT 175.950 728.100 178.050 728.400 ;
        RECT 205.950 727.950 208.050 728.400 ;
        RECT 217.950 728.100 220.050 728.400 ;
        RECT 230.400 728.400 250.050 729.600 ;
        RECT 23.400 724.050 24.600 727.950 ;
        RECT 230.400 724.050 231.600 728.400 ;
        RECT 247.950 728.100 250.050 728.400 ;
        RECT 271.950 729.600 274.050 730.200 ;
        RECT 307.950 729.600 310.050 730.050 ;
        RECT 271.950 728.400 310.050 729.600 ;
        RECT 271.950 728.100 274.050 728.400 ;
        RECT 307.950 727.950 310.050 728.400 ;
        RECT 325.950 729.600 328.050 730.200 ;
        RECT 334.950 729.600 337.050 730.050 ;
        RECT 325.950 728.400 337.050 729.600 ;
        RECT 325.950 728.100 328.050 728.400 ;
        RECT 334.950 727.950 337.050 728.400 ;
        RECT 355.950 729.750 358.050 730.200 ;
        RECT 367.950 729.750 370.050 730.200 ;
        RECT 355.950 728.550 370.050 729.750 ;
        RECT 355.950 728.100 358.050 728.550 ;
        RECT 367.950 728.100 370.050 728.550 ;
        RECT 373.950 729.600 376.050 730.200 ;
        RECT 382.950 729.600 385.050 730.050 ;
        RECT 373.950 728.400 385.050 729.600 ;
        RECT 373.950 728.100 376.050 728.400 ;
        RECT 382.950 727.950 385.050 728.400 ;
        RECT 409.950 729.750 412.050 730.200 ;
        RECT 421.950 729.750 424.050 730.200 ;
        RECT 409.950 728.550 424.050 729.750 ;
        RECT 409.950 728.100 412.050 728.550 ;
        RECT 421.950 728.100 424.050 728.550 ;
        RECT 433.950 729.600 436.050 730.050 ;
        RECT 439.950 729.600 442.050 730.200 ;
        RECT 433.950 728.400 442.050 729.600 ;
        RECT 433.950 727.950 436.050 728.400 ;
        RECT 439.950 728.100 442.050 728.400 ;
        RECT 445.950 729.600 448.050 730.050 ;
        RECT 469.950 729.600 472.050 730.200 ;
        RECT 445.950 728.400 472.050 729.600 ;
        RECT 445.950 727.950 448.050 728.400 ;
        RECT 469.950 728.100 472.050 728.400 ;
        RECT 484.950 729.600 487.050 730.050 ;
        RECT 499.950 729.600 502.050 730.050 ;
        RECT 532.950 729.600 535.050 730.200 ;
        RECT 484.950 728.400 492.600 729.600 ;
        RECT 484.950 727.950 487.050 728.400 ;
        RECT 22.950 721.950 25.050 724.050 ;
        RECT 58.950 723.450 61.050 723.900 ;
        RECT 70.950 723.450 73.050 723.900 ;
        RECT 58.950 722.250 73.050 723.450 ;
        RECT 58.950 721.800 61.050 722.250 ;
        RECT 70.950 721.800 73.050 722.250 ;
        RECT 76.950 723.600 79.050 723.900 ;
        RECT 88.950 723.600 91.050 723.900 ;
        RECT 76.950 723.450 91.050 723.600 ;
        RECT 94.950 723.450 97.050 723.900 ;
        RECT 76.950 722.400 97.050 723.450 ;
        RECT 76.950 721.800 79.050 722.400 ;
        RECT 88.950 722.250 97.050 722.400 ;
        RECT 88.950 721.800 91.050 722.250 ;
        RECT 94.950 721.800 97.050 722.250 ;
        RECT 160.950 723.600 163.050 724.050 ;
        RECT 166.950 723.600 169.050 723.900 ;
        RECT 160.950 723.450 169.050 723.600 ;
        RECT 172.950 723.450 175.050 723.900 ;
        RECT 160.950 722.400 175.050 723.450 ;
        RECT 160.950 721.950 163.050 722.400 ;
        RECT 166.950 722.250 175.050 722.400 ;
        RECT 166.950 721.800 169.050 722.250 ;
        RECT 172.950 721.800 175.050 722.250 ;
        RECT 178.950 723.450 181.050 723.900 ;
        RECT 190.950 723.450 193.050 723.900 ;
        RECT 178.950 722.250 193.050 723.450 ;
        RECT 178.950 721.800 181.050 722.250 ;
        RECT 190.950 721.800 193.050 722.250 ;
        RECT 199.950 723.450 202.050 723.900 ;
        RECT 205.950 723.450 208.050 723.900 ;
        RECT 199.950 722.250 208.050 723.450 ;
        RECT 199.950 721.800 202.050 722.250 ;
        RECT 205.950 721.800 208.050 722.250 ;
        RECT 229.950 721.950 232.050 724.050 ;
        RECT 491.400 723.900 492.600 728.400 ;
        RECT 499.950 728.400 535.050 729.600 ;
        RECT 499.950 727.950 502.050 728.400 ;
        RECT 532.950 728.100 535.050 728.400 ;
        RECT 538.950 729.600 541.050 730.200 ;
        RECT 538.950 728.400 543.600 729.600 ;
        RECT 538.950 728.100 541.050 728.400 ;
        RECT 542.400 724.050 543.600 728.400 ;
        RECT 565.950 727.950 568.050 730.050 ;
        RECT 571.950 729.600 574.050 730.050 ;
        RECT 577.950 729.600 580.050 730.200 ;
        RECT 571.950 728.400 580.050 729.600 ;
        RECT 571.950 727.950 574.050 728.400 ;
        RECT 577.950 728.100 580.050 728.400 ;
        RECT 595.950 729.750 598.050 730.200 ;
        RECT 604.950 729.750 607.050 730.200 ;
        RECT 595.950 728.550 607.050 729.750 ;
        RECT 595.950 728.100 598.050 728.550 ;
        RECT 604.950 728.100 607.050 728.550 ;
        RECT 619.950 729.750 622.050 730.200 ;
        RECT 625.950 729.750 628.050 730.200 ;
        RECT 619.950 728.550 628.050 729.750 ;
        RECT 619.950 728.100 622.050 728.550 ;
        RECT 625.950 728.100 628.050 728.550 ;
        RECT 640.950 727.950 643.050 730.050 ;
        RECT 658.950 729.600 661.050 730.050 ;
        RECT 670.950 729.600 673.050 730.200 ;
        RECT 694.950 729.600 697.050 730.200 ;
        RECT 715.950 729.600 718.050 730.200 ;
        RECT 722.400 729.600 723.600 730.950 ;
        RECT 758.400 730.200 759.600 731.400 ;
        RECT 802.950 730.950 805.050 731.400 ;
        RECT 817.950 730.950 820.050 731.400 ;
        RECT 898.950 732.600 903.000 733.050 ;
        RECT 898.950 730.950 903.600 732.600 ;
        RECT 658.950 728.400 673.050 729.600 ;
        RECT 658.950 727.950 661.050 728.400 ;
        RECT 670.950 728.100 673.050 728.400 ;
        RECT 680.400 728.400 697.050 729.600 ;
        RECT 244.950 723.600 247.050 723.900 ;
        RECT 256.950 723.600 259.050 723.900 ;
        RECT 244.950 723.450 259.050 723.600 ;
        RECT 268.950 723.450 271.050 723.900 ;
        RECT 244.950 722.400 271.050 723.450 ;
        RECT 244.950 721.800 247.050 722.400 ;
        RECT 256.950 722.250 271.050 722.400 ;
        RECT 256.950 721.800 259.050 722.250 ;
        RECT 268.950 721.800 271.050 722.250 ;
        RECT 307.950 723.450 310.050 723.900 ;
        RECT 316.950 723.450 319.050 723.900 ;
        RECT 307.950 722.250 319.050 723.450 ;
        RECT 307.950 721.800 310.050 722.250 ;
        RECT 316.950 721.800 319.050 722.250 ;
        RECT 334.950 723.450 337.050 723.900 ;
        RECT 343.950 723.450 346.050 723.900 ;
        RECT 334.950 722.250 346.050 723.450 ;
        RECT 334.950 721.800 337.050 722.250 ;
        RECT 343.950 721.800 346.050 722.250 ;
        RECT 382.950 723.450 385.050 723.900 ;
        RECT 388.950 723.450 391.050 723.900 ;
        RECT 382.950 722.250 391.050 723.450 ;
        RECT 382.950 721.800 385.050 722.250 ;
        RECT 388.950 721.800 391.050 722.250 ;
        RECT 424.950 723.450 427.050 723.900 ;
        RECT 430.950 723.450 433.050 723.900 ;
        RECT 424.950 722.250 433.050 723.450 ;
        RECT 424.950 721.800 427.050 722.250 ;
        RECT 430.950 721.800 433.050 722.250 ;
        RECT 448.950 723.600 451.050 723.900 ;
        RECT 466.950 723.600 469.050 723.900 ;
        RECT 448.950 723.450 469.050 723.600 ;
        RECT 481.950 723.450 484.050 723.900 ;
        RECT 448.950 722.400 484.050 723.450 ;
        RECT 448.950 721.800 451.050 722.400 ;
        RECT 466.950 722.250 484.050 722.400 ;
        RECT 466.950 721.800 469.050 722.250 ;
        RECT 481.950 721.800 484.050 722.250 ;
        RECT 490.950 721.800 493.050 723.900 ;
        RECT 496.950 723.450 499.050 723.900 ;
        RECT 502.950 723.450 505.050 723.900 ;
        RECT 496.950 722.250 505.050 723.450 ;
        RECT 496.950 721.800 499.050 722.250 ;
        RECT 502.950 721.800 505.050 722.250 ;
        RECT 511.950 723.600 514.050 723.900 ;
        RECT 535.950 723.600 538.050 723.900 ;
        RECT 511.950 722.400 538.050 723.600 ;
        RECT 511.950 721.800 514.050 722.400 ;
        RECT 535.950 721.800 538.050 722.400 ;
        RECT 541.950 721.950 544.050 724.050 ;
        RECT 553.950 723.600 556.050 723.900 ;
        RECT 566.400 723.600 567.600 727.950 ;
        RECT 553.950 722.400 567.600 723.600 ;
        RECT 580.950 723.600 583.050 723.900 ;
        RECT 601.950 723.600 604.050 723.900 ;
        RECT 619.950 723.600 622.050 724.050 ;
        RECT 580.950 722.400 622.050 723.600 ;
        RECT 553.950 721.800 556.050 722.400 ;
        RECT 580.950 721.800 583.050 722.400 ;
        RECT 601.950 721.800 604.050 722.400 ;
        RECT 619.950 721.950 622.050 722.400 ;
        RECT 628.950 723.600 631.050 723.900 ;
        RECT 641.400 723.600 642.600 727.950 ;
        RECT 680.400 724.050 681.600 728.400 ;
        RECT 694.950 728.100 697.050 728.400 ;
        RECT 713.400 728.400 718.050 729.600 ;
        RECT 713.400 724.050 714.600 728.400 ;
        RECT 715.950 728.100 718.050 728.400 ;
        RECT 719.400 728.400 723.600 729.600 ;
        RECT 748.950 729.750 751.050 730.200 ;
        RECT 757.950 729.750 760.050 730.200 ;
        RECT 748.950 728.550 760.050 729.750 ;
        RECT 646.950 723.600 649.050 723.900 ;
        RECT 628.950 722.400 649.050 723.600 ;
        RECT 628.950 721.800 631.050 722.400 ;
        RECT 646.950 721.800 649.050 722.400 ;
        RECT 652.950 723.450 655.050 723.900 ;
        RECT 658.950 723.450 661.050 723.900 ;
        RECT 652.950 722.250 661.050 723.450 ;
        RECT 652.950 721.800 655.050 722.250 ;
        RECT 658.950 721.800 661.050 722.250 ;
        RECT 679.950 721.950 682.050 724.050 ;
        RECT 712.950 721.950 715.050 724.050 ;
        RECT 719.400 723.900 720.600 728.400 ;
        RECT 748.950 728.100 751.050 728.550 ;
        RECT 757.950 728.100 760.050 728.550 ;
        RECT 778.950 729.600 781.050 730.200 ;
        RECT 793.950 729.600 796.050 730.200 ;
        RECT 778.950 728.400 796.050 729.600 ;
        RECT 778.950 728.100 781.050 728.400 ;
        RECT 793.950 728.100 796.050 728.400 ;
        RECT 814.950 729.600 817.050 730.050 ;
        RECT 835.950 729.750 838.050 730.200 ;
        RECT 847.950 729.750 850.050 730.200 ;
        RECT 814.950 728.400 831.600 729.600 ;
        RECT 814.950 727.950 817.050 728.400 ;
        RECT 830.400 726.600 831.600 728.400 ;
        RECT 835.950 728.550 850.050 729.750 ;
        RECT 835.950 728.100 838.050 728.550 ;
        RECT 847.950 728.100 850.050 728.550 ;
        RECT 856.950 729.750 859.050 730.200 ;
        RECT 862.950 729.750 865.050 730.050 ;
        RECT 871.950 729.750 874.050 730.200 ;
        RECT 856.950 728.550 874.050 729.750 ;
        RECT 856.950 728.100 859.050 728.550 ;
        RECT 862.950 727.950 865.050 728.550 ;
        RECT 871.950 728.100 874.050 728.550 ;
        RECT 877.950 727.950 880.050 730.050 ;
        RECT 895.950 728.100 898.050 730.200 ;
        RECT 830.400 725.400 846.600 726.600 ;
        RECT 718.950 721.800 721.050 723.900 ;
        RECT 724.950 723.450 727.050 723.900 ;
        RECT 730.950 723.450 733.050 723.900 ;
        RECT 724.950 722.250 733.050 723.450 ;
        RECT 724.950 721.800 727.050 722.250 ;
        RECT 730.950 721.800 733.050 722.250 ;
        RECT 736.950 723.450 739.050 723.900 ;
        RECT 745.950 723.450 748.050 723.900 ;
        RECT 736.950 722.250 748.050 723.450 ;
        RECT 736.950 721.800 739.050 722.250 ;
        RECT 745.950 721.800 748.050 722.250 ;
        RECT 757.950 723.600 760.050 724.050 ;
        RECT 790.950 723.600 793.050 724.050 ;
        RECT 845.400 723.900 846.600 725.400 ;
        RECT 757.950 722.400 793.050 723.600 ;
        RECT 757.950 721.950 760.050 722.400 ;
        RECT 790.950 721.950 793.050 722.400 ;
        RECT 802.950 723.450 805.050 723.900 ;
        RECT 811.800 723.450 813.900 723.900 ;
        RECT 820.950 723.600 823.050 723.900 ;
        RECT 802.950 722.250 813.900 723.450 ;
        RECT 815.400 723.000 823.050 723.600 ;
        RECT 802.950 721.800 805.050 722.250 ;
        RECT 811.800 721.800 813.900 722.250 ;
        RECT 814.950 722.400 823.050 723.000 ;
        RECT 283.950 720.600 286.050 721.050 ;
        RECT 298.950 720.600 301.050 721.050 ;
        RECT 283.950 719.400 301.050 720.600 ;
        RECT 283.950 718.950 286.050 719.400 ;
        RECT 298.950 718.950 301.050 719.400 ;
        RECT 325.950 720.600 328.050 721.050 ;
        RECT 349.950 720.600 352.050 721.050 ;
        RECT 355.950 720.600 358.050 721.050 ;
        RECT 325.950 719.400 358.050 720.600 ;
        RECT 325.950 718.950 328.050 719.400 ;
        RECT 349.950 718.950 352.050 719.400 ;
        RECT 355.950 718.950 358.050 719.400 ;
        RECT 682.950 720.600 685.050 721.050 ;
        RECT 697.950 720.600 700.050 721.050 ;
        RECT 682.950 719.400 700.050 720.600 ;
        RECT 682.950 718.950 685.050 719.400 ;
        RECT 697.950 718.950 700.050 719.400 ;
        RECT 814.950 718.950 817.050 722.400 ;
        RECT 820.950 721.800 823.050 722.400 ;
        RECT 844.950 721.800 847.050 723.900 ;
        RECT 874.950 723.600 877.050 723.900 ;
        RECT 878.400 723.600 879.600 727.950 ;
        RECT 874.950 722.400 879.600 723.600 ;
        RECT 889.950 723.600 892.050 724.050 ;
        RECT 896.400 723.600 897.600 728.100 ;
        RECT 902.400 724.050 903.600 730.950 ;
        RECT 889.950 722.400 897.600 723.600 ;
        RECT 898.950 722.400 903.600 724.050 ;
        RECT 874.950 721.800 877.050 722.400 ;
        RECT 889.950 721.950 892.050 722.400 ;
        RECT 898.950 721.950 903.000 722.400 ;
        RECT 847.950 720.600 850.050 721.050 ;
        RECT 859.950 720.600 862.050 721.050 ;
        RECT 892.950 720.600 895.050 721.050 ;
        RECT 847.950 719.400 862.050 720.600 ;
        RECT 878.400 720.000 895.050 720.600 ;
        RECT 847.950 718.950 850.050 719.400 ;
        RECT 859.950 718.950 862.050 719.400 ;
        RECT 877.950 719.400 895.050 720.000 ;
        RECT 61.950 717.600 64.050 718.050 ;
        RECT 94.950 717.600 97.050 718.050 ;
        RECT 109.950 717.600 112.050 718.050 ;
        RECT 61.950 716.400 112.050 717.600 ;
        RECT 61.950 715.950 64.050 716.400 ;
        RECT 94.950 715.950 97.050 716.400 ;
        RECT 109.950 715.950 112.050 716.400 ;
        RECT 232.950 717.600 235.050 718.050 ;
        RECT 250.950 717.600 253.050 718.050 ;
        RECT 232.950 716.400 253.050 717.600 ;
        RECT 232.950 715.950 235.050 716.400 ;
        RECT 250.950 715.950 253.050 716.400 ;
        RECT 331.950 717.600 334.050 718.050 ;
        RECT 370.950 717.600 373.050 718.050 ;
        RECT 331.950 716.400 373.050 717.600 ;
        RECT 331.950 715.950 334.050 716.400 ;
        RECT 370.950 715.950 373.050 716.400 ;
        RECT 394.950 717.600 397.050 718.050 ;
        RECT 433.950 717.600 436.050 718.050 ;
        RECT 394.950 716.400 436.050 717.600 ;
        RECT 394.950 715.950 397.050 716.400 ;
        RECT 433.950 715.950 436.050 716.400 ;
        RECT 460.950 717.600 463.050 718.050 ;
        RECT 580.950 717.600 583.050 718.050 ;
        RECT 460.950 716.400 583.050 717.600 ;
        RECT 460.950 715.950 463.050 716.400 ;
        RECT 580.950 715.950 583.050 716.400 ;
        RECT 595.950 717.600 598.050 718.050 ;
        RECT 679.950 717.600 682.050 718.050 ;
        RECT 595.950 716.400 682.050 717.600 ;
        RECT 595.950 715.950 598.050 716.400 ;
        RECT 679.950 715.950 682.050 716.400 ;
        RECT 832.950 717.600 835.050 718.050 ;
        RECT 871.950 717.600 874.050 718.050 ;
        RECT 832.950 716.400 874.050 717.600 ;
        RECT 832.950 715.950 835.050 716.400 ;
        RECT 871.950 715.950 874.050 716.400 ;
        RECT 877.950 715.950 880.050 719.400 ;
        RECT 892.950 718.950 895.050 719.400 ;
        RECT 70.950 714.600 73.050 715.050 ;
        RECT 82.800 714.600 84.900 715.050 ;
        RECT 70.950 713.400 84.900 714.600 ;
        RECT 70.950 712.950 73.050 713.400 ;
        RECT 82.800 712.950 84.900 713.400 ;
        RECT 85.950 714.600 88.050 715.050 ;
        RECT 100.950 714.600 103.050 715.050 ;
        RECT 142.950 714.600 145.050 715.050 ;
        RECT 85.950 713.400 145.050 714.600 ;
        RECT 85.950 712.950 88.050 713.400 ;
        RECT 100.950 712.950 103.050 713.400 ;
        RECT 142.950 712.950 145.050 713.400 ;
        RECT 157.950 714.600 160.050 715.050 ;
        RECT 217.950 714.600 220.050 715.050 ;
        RECT 157.950 713.400 220.050 714.600 ;
        RECT 157.950 712.950 160.050 713.400 ;
        RECT 217.950 712.950 220.050 713.400 ;
        RECT 487.950 714.600 490.050 715.050 ;
        RECT 505.950 714.600 508.050 715.050 ;
        RECT 487.950 713.400 508.050 714.600 ;
        RECT 487.950 712.950 490.050 713.400 ;
        RECT 505.950 712.950 508.050 713.400 ;
        RECT 547.950 714.600 550.050 715.050 ;
        RECT 562.950 714.600 565.050 715.050 ;
        RECT 547.950 713.400 565.050 714.600 ;
        RECT 547.950 712.950 550.050 713.400 ;
        RECT 562.950 712.950 565.050 713.400 ;
        RECT 796.950 714.600 799.050 715.050 ;
        RECT 820.950 714.600 823.050 715.050 ;
        RECT 796.950 713.400 823.050 714.600 ;
        RECT 796.950 712.950 799.050 713.400 ;
        RECT 820.950 712.950 823.050 713.400 ;
        RECT 850.950 714.600 853.050 715.050 ;
        RECT 868.950 714.600 871.050 715.050 ;
        RECT 850.950 713.400 871.050 714.600 ;
        RECT 850.950 712.950 853.050 713.400 ;
        RECT 868.950 712.950 871.050 713.400 ;
        RECT 208.950 711.600 211.050 712.050 ;
        RECT 274.950 711.600 277.050 712.050 ;
        RECT 208.950 710.400 277.050 711.600 ;
        RECT 208.950 709.950 211.050 710.400 ;
        RECT 274.950 709.950 277.050 710.400 ;
        RECT 763.950 711.600 766.050 712.050 ;
        RECT 778.950 711.600 781.050 712.050 ;
        RECT 763.950 710.400 781.050 711.600 ;
        RECT 763.950 709.950 766.050 710.400 ;
        RECT 778.950 709.950 781.050 710.400 ;
        RECT 220.950 708.600 223.050 709.050 ;
        RECT 247.950 708.600 250.050 709.050 ;
        RECT 220.950 707.400 250.050 708.600 ;
        RECT 220.950 706.950 223.050 707.400 ;
        RECT 247.950 706.950 250.050 707.400 ;
        RECT 262.950 708.600 265.050 709.050 ;
        RECT 322.950 708.600 325.050 709.050 ;
        RECT 262.950 707.400 325.050 708.600 ;
        RECT 262.950 706.950 265.050 707.400 ;
        RECT 322.950 706.950 325.050 707.400 ;
        RECT 355.950 708.600 358.050 709.050 ;
        RECT 418.950 708.600 421.050 709.050 ;
        RECT 355.950 707.400 421.050 708.600 ;
        RECT 355.950 706.950 358.050 707.400 ;
        RECT 418.950 706.950 421.050 707.400 ;
        RECT 586.950 708.600 589.050 709.050 ;
        RECT 607.950 708.600 610.050 709.050 ;
        RECT 643.950 708.600 646.050 709.050 ;
        RECT 586.950 707.400 646.050 708.600 ;
        RECT 586.950 706.950 589.050 707.400 ;
        RECT 607.950 706.950 610.050 707.400 ;
        RECT 643.950 706.950 646.050 707.400 ;
        RECT 751.950 708.600 754.050 709.050 ;
        RECT 811.950 708.600 814.050 709.050 ;
        RECT 751.950 707.400 814.050 708.600 ;
        RECT 751.950 706.950 754.050 707.400 ;
        RECT 811.950 706.950 814.050 707.400 ;
        RECT 145.950 705.600 148.050 706.050 ;
        RECT 178.950 705.600 181.050 706.050 ;
        RECT 145.950 704.400 181.050 705.600 ;
        RECT 145.950 703.950 148.050 704.400 ;
        RECT 178.950 703.950 181.050 704.400 ;
        RECT 250.950 705.600 253.050 706.050 ;
        RECT 334.950 705.600 337.050 706.050 ;
        RECT 250.950 704.400 337.050 705.600 ;
        RECT 250.950 703.950 253.050 704.400 ;
        RECT 334.950 703.950 337.050 704.400 ;
        RECT 433.950 705.600 436.050 706.050 ;
        RECT 442.950 705.600 445.050 706.050 ;
        RECT 472.950 705.600 475.050 706.050 ;
        RECT 529.950 705.600 532.050 706.050 ;
        RECT 433.950 704.400 532.050 705.600 ;
        RECT 433.950 703.950 436.050 704.400 ;
        RECT 442.950 703.950 445.050 704.400 ;
        RECT 472.950 703.950 475.050 704.400 ;
        RECT 529.950 703.950 532.050 704.400 ;
        RECT 142.950 702.600 145.050 703.050 ;
        RECT 181.950 702.600 184.050 703.050 ;
        RECT 214.950 702.600 217.050 703.050 ;
        RECT 142.950 701.400 217.050 702.600 ;
        RECT 142.950 700.950 145.050 701.400 ;
        RECT 181.950 700.950 184.050 701.400 ;
        RECT 214.950 700.950 217.050 701.400 ;
        RECT 253.950 702.600 256.050 703.050 ;
        RECT 280.950 702.600 283.050 703.050 ;
        RECT 331.950 702.600 334.050 703.050 ;
        RECT 253.950 701.400 334.050 702.600 ;
        RECT 253.950 700.950 256.050 701.400 ;
        RECT 280.950 700.950 283.050 701.400 ;
        RECT 331.950 700.950 334.050 701.400 ;
        RECT 850.950 702.600 853.050 703.050 ;
        RECT 883.950 702.600 886.050 703.050 ;
        RECT 850.950 701.400 886.050 702.600 ;
        RECT 850.950 700.950 853.050 701.400 ;
        RECT 883.950 700.950 886.050 701.400 ;
        RECT 13.950 699.600 16.050 700.050 ;
        RECT 22.950 699.600 25.050 700.050 ;
        RECT 13.950 698.400 25.050 699.600 ;
        RECT 13.950 697.950 16.050 698.400 ;
        RECT 22.950 697.950 25.050 698.400 ;
        RECT 112.950 699.600 115.050 700.050 ;
        RECT 142.950 699.600 145.050 699.900 ;
        RECT 169.950 699.600 172.050 700.050 ;
        RECT 112.950 698.400 172.050 699.600 ;
        RECT 112.950 697.950 115.050 698.400 ;
        RECT 142.950 697.800 145.050 698.400 ;
        RECT 169.950 697.950 172.050 698.400 ;
        RECT 178.950 699.600 181.050 700.050 ;
        RECT 262.950 699.600 265.050 700.050 ;
        RECT 178.950 698.400 265.050 699.600 ;
        RECT 178.950 697.950 181.050 698.400 ;
        RECT 262.950 697.950 265.050 698.400 ;
        RECT 268.950 699.600 271.050 700.050 ;
        RECT 292.950 699.600 295.050 700.050 ;
        RECT 301.950 699.600 304.050 700.050 ;
        RECT 268.950 698.400 304.050 699.600 ;
        RECT 268.950 697.950 271.050 698.400 ;
        RECT 292.950 697.950 295.050 698.400 ;
        RECT 301.950 697.950 304.050 698.400 ;
        RECT 520.950 699.600 523.050 700.050 ;
        RECT 541.950 699.600 544.050 700.050 ;
        RECT 655.950 699.600 658.050 700.050 ;
        RECT 667.950 699.600 670.050 700.050 ;
        RECT 520.950 698.400 528.600 699.600 ;
        RECT 520.950 697.950 523.050 698.400 ;
        RECT 274.950 696.600 277.050 697.050 ;
        RECT 289.950 696.600 292.050 697.050 ;
        RECT 274.950 695.400 292.050 696.600 ;
        RECT 274.950 694.950 277.050 695.400 ;
        RECT 289.950 694.950 292.050 695.400 ;
        RECT 352.950 696.600 355.050 697.050 ;
        RECT 454.950 696.600 457.050 697.050 ;
        RECT 352.950 695.400 457.050 696.600 ;
        RECT 352.950 694.950 355.050 695.400 ;
        RECT 454.950 694.950 457.050 695.400 ;
        RECT 478.950 696.600 481.050 697.050 ;
        RECT 505.950 696.600 508.050 697.050 ;
        RECT 511.950 696.600 514.050 697.050 ;
        RECT 478.950 695.400 514.050 696.600 ;
        RECT 527.400 696.600 528.600 698.400 ;
        RECT 541.950 698.400 670.050 699.600 ;
        RECT 541.950 697.950 544.050 698.400 ;
        RECT 655.950 697.950 658.050 698.400 ;
        RECT 667.950 697.950 670.050 698.400 ;
        RECT 778.950 699.600 781.050 700.050 ;
        RECT 805.950 699.600 808.050 700.050 ;
        RECT 778.950 698.400 808.050 699.600 ;
        RECT 778.950 697.950 781.050 698.400 ;
        RECT 805.950 697.950 808.050 698.400 ;
        RECT 679.950 696.600 682.050 697.050 ;
        RECT 527.400 695.400 682.050 696.600 ;
        RECT 478.950 694.950 481.050 695.400 ;
        RECT 505.950 694.950 508.050 695.400 ;
        RECT 511.950 694.950 514.050 695.400 ;
        RECT 679.950 694.950 682.050 695.400 ;
        RECT 697.950 696.600 700.050 697.050 ;
        RECT 721.950 696.600 724.050 697.050 ;
        RECT 697.950 695.400 724.050 696.600 ;
        RECT 697.950 694.950 700.050 695.400 ;
        RECT 721.950 694.950 724.050 695.400 ;
        RECT 775.950 696.600 778.050 697.050 ;
        RECT 832.950 696.600 835.050 697.050 ;
        RECT 775.950 695.400 835.050 696.600 ;
        RECT 775.950 694.950 778.050 695.400 ;
        RECT 832.950 694.950 835.050 695.400 ;
        RECT 523.950 693.600 526.050 694.050 ;
        RECT 586.950 693.600 589.050 694.050 ;
        RECT 523.950 692.400 589.050 693.600 ;
        RECT 523.950 691.950 526.050 692.400 ;
        RECT 586.950 691.950 589.050 692.400 ;
        RECT 619.950 693.600 622.050 694.050 ;
        RECT 634.950 693.600 637.050 694.050 ;
        RECT 619.950 692.400 637.050 693.600 ;
        RECT 619.950 691.950 622.050 692.400 ;
        RECT 634.950 691.950 637.050 692.400 ;
        RECT 661.950 693.600 664.050 694.050 ;
        RECT 784.950 693.600 787.050 694.050 ;
        RECT 796.950 693.600 799.050 694.050 ;
        RECT 661.950 692.400 672.600 693.600 ;
        RECT 661.950 691.950 664.050 692.400 ;
        RECT 133.950 690.600 136.050 691.050 ;
        RECT 148.950 690.600 151.050 691.050 ;
        RECT 196.950 690.600 199.050 691.050 ;
        RECT 133.950 689.400 199.050 690.600 ;
        RECT 133.950 688.950 136.050 689.400 ;
        RECT 148.950 688.950 151.050 689.400 ;
        RECT 196.950 688.950 199.050 689.400 ;
        RECT 277.950 690.600 280.050 691.050 ;
        RECT 316.950 690.600 319.050 691.050 ;
        RECT 277.950 689.400 319.050 690.600 ;
        RECT 277.950 688.950 280.050 689.400 ;
        RECT 316.950 688.950 319.050 689.400 ;
        RECT 358.950 690.600 361.050 691.050 ;
        RECT 409.950 690.600 412.050 691.050 ;
        RECT 451.950 690.600 454.050 691.050 ;
        RECT 358.950 689.400 454.050 690.600 ;
        RECT 358.950 688.950 361.050 689.400 ;
        RECT 409.950 688.950 412.050 689.400 ;
        RECT 451.950 688.950 454.050 689.400 ;
        RECT 511.950 690.600 514.050 691.050 ;
        RECT 541.950 690.600 544.050 691.050 ;
        RECT 511.950 689.400 544.050 690.600 ;
        RECT 671.400 690.600 672.600 692.400 ;
        RECT 784.950 692.400 799.050 693.600 ;
        RECT 784.950 691.950 787.050 692.400 ;
        RECT 796.950 691.950 799.050 692.400 ;
        RECT 685.950 690.600 688.050 691.050 ;
        RECT 712.950 690.600 715.050 691.050 ;
        RECT 671.400 689.400 715.050 690.600 ;
        RECT 511.950 688.950 514.050 689.400 ;
        RECT 541.950 688.950 544.050 689.400 ;
        RECT 685.950 688.950 688.050 689.400 ;
        RECT 712.950 688.950 715.050 689.400 ;
        RECT 733.950 690.600 736.050 691.050 ;
        RECT 742.950 690.600 745.050 691.050 ;
        RECT 733.950 689.400 745.050 690.600 ;
        RECT 733.950 688.950 736.050 689.400 ;
        RECT 742.950 688.950 745.050 689.400 ;
        RECT 193.950 687.600 196.050 688.050 ;
        RECT 223.950 687.600 226.050 688.050 ;
        RECT 253.950 687.600 256.050 688.050 ;
        RECT 193.950 686.400 256.050 687.600 ;
        RECT 193.950 685.950 196.050 686.400 ;
        RECT 223.950 685.950 226.050 686.400 ;
        RECT 253.950 685.950 256.050 686.400 ;
        RECT 544.950 687.600 547.050 688.050 ;
        RECT 571.950 687.600 574.050 688.050 ;
        RECT 580.950 687.600 583.050 688.050 ;
        RECT 544.950 686.400 583.050 687.600 ;
        RECT 544.950 685.950 547.050 686.400 ;
        RECT 571.950 685.950 574.050 686.400 ;
        RECT 580.950 685.950 583.050 686.400 ;
        RECT 637.950 687.600 640.050 688.050 ;
        RECT 667.950 687.600 670.050 688.050 ;
        RECT 637.950 686.400 670.050 687.600 ;
        RECT 637.950 685.950 640.050 686.400 ;
        RECT 667.950 685.950 670.050 686.400 ;
        RECT 691.950 687.600 694.050 688.050 ;
        RECT 706.950 687.600 709.050 688.050 ;
        RECT 691.950 686.400 709.050 687.600 ;
        RECT 691.950 685.950 694.050 686.400 ;
        RECT 706.950 685.950 709.050 686.400 ;
        RECT 787.950 687.600 790.050 688.050 ;
        RECT 793.950 687.600 796.050 688.050 ;
        RECT 787.950 686.400 796.050 687.600 ;
        RECT 787.950 685.950 790.050 686.400 ;
        RECT 793.950 685.950 796.050 686.400 ;
        RECT 817.950 687.600 820.050 688.050 ;
        RECT 826.950 687.600 829.050 688.050 ;
        RECT 817.950 686.400 829.050 687.600 ;
        RECT 817.950 685.950 820.050 686.400 ;
        RECT 826.950 685.950 829.050 686.400 ;
        RECT 865.950 687.600 868.050 688.050 ;
        RECT 889.950 687.600 892.050 688.050 ;
        RECT 865.950 686.400 892.050 687.600 ;
        RECT 865.950 685.950 868.050 686.400 ;
        RECT 889.950 685.950 892.050 686.400 ;
        RECT 13.950 683.100 16.050 685.200 ;
        RECT 37.950 683.100 40.050 685.200 ;
        RECT 43.950 683.100 46.050 685.200 ;
        RECT 88.950 684.600 91.050 685.200 ;
        RECT 97.950 684.600 100.050 685.050 ;
        RECT 88.950 683.400 100.050 684.600 ;
        RECT 88.950 683.100 91.050 683.400 ;
        RECT 14.400 681.600 15.600 683.100 ;
        RECT 14.400 680.400 21.600 681.600 ;
        RECT 20.400 678.600 21.600 680.400 ;
        RECT 38.400 679.050 39.600 683.100 ;
        RECT 44.400 681.600 45.600 683.100 ;
        RECT 97.950 682.950 100.050 683.400 ;
        RECT 109.950 684.600 112.050 685.200 ;
        RECT 127.950 684.600 130.050 685.200 ;
        RECT 136.950 684.600 139.050 685.050 ;
        RECT 109.950 683.400 130.050 684.600 ;
        RECT 109.950 683.100 112.050 683.400 ;
        RECT 127.950 683.100 130.050 683.400 ;
        RECT 131.400 683.400 139.050 684.600 ;
        RECT 55.950 681.600 58.050 682.050 ;
        RECT 44.400 680.400 58.050 681.600 ;
        RECT 55.950 679.950 58.050 680.400 ;
        RECT 25.950 678.600 28.050 679.050 ;
        RECT 20.400 677.400 28.050 678.600 ;
        RECT 25.950 676.950 28.050 677.400 ;
        RECT 34.950 677.400 39.600 679.050 ;
        RECT 131.400 678.900 132.600 683.400 ;
        RECT 136.950 682.950 139.050 683.400 ;
        RECT 157.950 683.100 160.050 685.200 ;
        RECT 158.400 679.050 159.600 683.100 ;
        RECT 169.950 681.600 172.050 685.050 ;
        RECT 175.950 683.100 178.050 685.200 ;
        RECT 205.950 683.100 208.050 685.200 ;
        RECT 229.950 684.600 232.050 685.200 ;
        RECT 247.950 684.600 250.050 685.200 ;
        RECT 229.950 683.400 250.050 684.600 ;
        RECT 229.950 683.100 232.050 683.400 ;
        RECT 247.950 683.100 250.050 683.400 ;
        RECT 286.950 684.750 289.050 685.200 ;
        RECT 295.950 684.750 298.050 685.200 ;
        RECT 286.950 684.600 298.050 684.750 ;
        RECT 310.950 684.600 313.050 685.050 ;
        RECT 286.950 683.550 313.050 684.600 ;
        RECT 286.950 683.100 289.050 683.550 ;
        RECT 295.950 683.400 313.050 683.550 ;
        RECT 295.950 683.100 298.050 683.400 ;
        RECT 169.950 681.000 174.600 681.600 ;
        RECT 170.400 680.400 174.600 681.000 ;
        RECT 46.950 678.600 49.050 678.900 ;
        RECT 67.950 678.600 70.050 678.900 ;
        RECT 85.950 678.600 88.050 678.900 ;
        RECT 46.950 677.400 88.050 678.600 ;
        RECT 34.950 676.950 39.000 677.400 ;
        RECT 46.950 676.800 49.050 677.400 ;
        RECT 67.950 676.800 70.050 677.400 ;
        RECT 85.950 676.800 88.050 677.400 ;
        RECT 100.950 678.450 103.050 678.900 ;
        RECT 106.950 678.450 109.050 678.900 ;
        RECT 100.950 677.250 109.050 678.450 ;
        RECT 100.950 676.800 103.050 677.250 ;
        RECT 106.950 676.800 109.050 677.250 ;
        RECT 130.950 676.800 133.050 678.900 ;
        RECT 142.950 678.450 145.050 678.900 ;
        RECT 148.950 678.450 151.050 678.900 ;
        RECT 142.950 677.250 151.050 678.450 ;
        RECT 158.400 677.400 163.050 679.050 ;
        RECT 173.400 678.900 174.600 680.400 ;
        RECT 142.950 676.800 145.050 677.250 ;
        RECT 148.950 676.800 151.050 677.250 ;
        RECT 159.000 676.950 163.050 677.400 ;
        RECT 172.950 676.800 175.050 678.900 ;
        RECT 176.400 678.600 177.600 683.100 ;
        RECT 206.400 681.600 207.600 683.100 ;
        RECT 310.950 682.950 313.050 683.400 ;
        RECT 367.950 684.600 370.050 685.200 ;
        RECT 376.950 684.600 379.050 685.050 ;
        RECT 367.950 683.400 379.050 684.600 ;
        RECT 367.950 683.100 370.050 683.400 ;
        RECT 376.950 682.950 379.050 683.400 ;
        RECT 400.950 684.750 403.050 685.200 ;
        RECT 415.950 684.750 418.050 685.200 ;
        RECT 400.950 683.550 418.050 684.750 ;
        RECT 400.950 683.100 403.050 683.550 ;
        RECT 415.950 683.100 418.050 683.550 ;
        RECT 436.950 684.750 439.050 685.200 ;
        RECT 445.950 684.750 448.050 685.200 ;
        RECT 436.950 683.550 448.050 684.750 ;
        RECT 436.950 683.100 439.050 683.550 ;
        RECT 445.950 683.100 448.050 683.550 ;
        RECT 490.950 684.600 493.050 685.050 ;
        RECT 496.950 684.600 499.050 685.200 ;
        RECT 490.950 683.400 499.050 684.600 ;
        RECT 490.950 682.950 493.050 683.400 ;
        RECT 496.950 683.100 499.050 683.400 ;
        RECT 532.950 684.750 535.050 685.200 ;
        RECT 550.950 684.750 553.050 685.200 ;
        RECT 532.950 683.550 553.050 684.750 ;
        RECT 532.950 683.100 535.050 683.550 ;
        RECT 550.950 683.100 553.050 683.550 ;
        RECT 586.950 684.750 589.050 685.200 ;
        RECT 595.950 684.750 598.050 685.050 ;
        RECT 616.950 684.750 619.050 685.200 ;
        RECT 586.950 683.550 619.050 684.750 ;
        RECT 586.950 683.100 589.050 683.550 ;
        RECT 595.950 682.950 598.050 683.550 ;
        RECT 616.950 683.100 619.050 683.550 ;
        RECT 631.950 683.100 634.050 685.200 ;
        RECT 724.950 684.600 727.050 685.050 ;
        RECT 716.400 683.400 727.050 684.600 ;
        RECT 283.950 681.600 286.050 682.050 ;
        RECT 206.400 680.400 286.050 681.600 ;
        RECT 632.400 681.600 633.600 683.100 ;
        RECT 667.950 681.600 670.050 682.050 ;
        RECT 632.400 680.400 657.600 681.600 ;
        RECT 283.950 679.950 286.050 680.400 ;
        RECT 193.950 678.600 196.050 678.900 ;
        RECT 176.400 677.400 196.050 678.600 ;
        RECT 193.950 676.800 196.050 677.400 ;
        RECT 217.950 678.450 220.050 678.900 ;
        RECT 226.950 678.600 229.050 678.900 ;
        RECT 250.950 678.600 253.050 678.900 ;
        RECT 226.950 678.450 253.050 678.600 ;
        RECT 217.950 677.400 253.050 678.450 ;
        RECT 217.950 677.250 229.050 677.400 ;
        RECT 217.950 676.800 220.050 677.250 ;
        RECT 226.950 676.800 229.050 677.250 ;
        RECT 250.950 676.800 253.050 677.400 ;
        RECT 256.950 678.600 259.050 678.900 ;
        RECT 268.950 678.600 271.050 679.050 ;
        RECT 256.950 677.400 271.050 678.600 ;
        RECT 256.950 676.800 259.050 677.400 ;
        RECT 268.950 676.950 271.050 677.400 ;
        RECT 358.950 678.600 361.050 679.050 ;
        RECT 364.950 678.600 367.050 678.900 ;
        RECT 358.950 678.450 367.050 678.600 ;
        RECT 370.950 678.450 373.050 678.900 ;
        RECT 358.950 677.400 373.050 678.450 ;
        RECT 358.950 676.950 361.050 677.400 ;
        RECT 364.950 677.250 373.050 677.400 ;
        RECT 364.950 676.800 367.050 677.250 ;
        RECT 370.950 676.800 373.050 677.250 ;
        RECT 376.950 678.450 379.050 678.900 ;
        RECT 382.950 678.450 385.050 678.900 ;
        RECT 376.950 677.250 385.050 678.450 ;
        RECT 376.950 676.800 379.050 677.250 ;
        RECT 382.950 676.800 385.050 677.250 ;
        RECT 409.950 678.450 412.050 678.900 ;
        RECT 430.950 678.450 433.050 678.900 ;
        RECT 409.950 677.250 433.050 678.450 ;
        RECT 409.950 676.800 412.050 677.250 ;
        RECT 430.950 676.800 433.050 677.250 ;
        RECT 448.950 678.450 451.050 678.900 ;
        RECT 460.950 678.450 463.050 678.900 ;
        RECT 448.950 677.250 463.050 678.450 ;
        RECT 448.950 676.800 451.050 677.250 ;
        RECT 460.950 676.800 463.050 677.250 ;
        RECT 565.950 678.450 568.050 678.900 ;
        RECT 571.950 678.450 574.050 678.900 ;
        RECT 565.950 677.250 574.050 678.450 ;
        RECT 565.950 676.800 568.050 677.250 ;
        RECT 571.950 676.800 574.050 677.250 ;
        RECT 595.950 678.450 598.050 678.900 ;
        RECT 604.950 678.450 607.050 678.900 ;
        RECT 595.950 677.250 607.050 678.450 ;
        RECT 595.950 676.800 598.050 677.250 ;
        RECT 604.950 676.800 607.050 677.250 ;
        RECT 643.950 678.600 646.050 679.050 ;
        RECT 652.950 678.600 655.050 678.900 ;
        RECT 643.950 677.400 655.050 678.600 ;
        RECT 656.400 678.600 657.600 680.400 ;
        RECT 667.950 680.400 684.600 681.600 ;
        RECT 667.950 679.950 670.050 680.400 ;
        RECT 676.950 678.600 679.050 678.900 ;
        RECT 656.400 677.400 679.050 678.600 ;
        RECT 683.400 678.600 684.600 680.400 ;
        RECT 716.400 679.050 717.600 683.400 ;
        RECT 724.950 682.950 727.050 683.400 ;
        RECT 736.950 684.600 739.050 685.200 ;
        RECT 757.950 684.600 760.050 685.200 ;
        RECT 736.950 683.400 760.050 684.600 ;
        RECT 736.950 683.100 739.050 683.400 ;
        RECT 757.950 683.100 760.050 683.400 ;
        RECT 763.950 684.600 766.050 685.200 ;
        RECT 769.950 684.600 772.050 685.050 ;
        RECT 763.950 683.400 772.050 684.600 ;
        RECT 763.950 683.100 766.050 683.400 ;
        RECT 769.950 682.950 772.050 683.400 ;
        RECT 775.950 684.600 778.050 685.050 ;
        RECT 775.950 683.400 789.600 684.600 ;
        RECT 775.950 682.950 778.050 683.400 ;
        RECT 703.950 678.600 706.050 678.900 ;
        RECT 683.400 677.400 706.050 678.600 ;
        RECT 643.950 676.950 646.050 677.400 ;
        RECT 652.950 676.800 655.050 677.400 ;
        RECT 676.950 676.800 679.050 677.400 ;
        RECT 703.950 676.800 706.050 677.400 ;
        RECT 715.950 676.950 718.050 679.050 ;
        RECT 733.950 678.600 736.050 678.900 ;
        RECT 760.950 678.600 763.050 678.900 ;
        RECT 766.950 678.600 769.050 679.050 ;
        RECT 788.400 678.900 789.600 683.400 ;
        RECT 790.950 682.950 793.050 685.050 ;
        RECT 811.950 684.600 814.050 685.200 ;
        RECT 838.950 684.750 841.050 685.200 ;
        RECT 844.950 684.750 847.050 685.200 ;
        RECT 811.950 683.400 819.600 684.600 ;
        RECT 811.950 683.100 814.050 683.400 ;
        RECT 733.950 677.400 769.050 678.600 ;
        RECT 733.950 676.800 736.050 677.400 ;
        RECT 760.950 676.800 763.050 677.400 ;
        RECT 766.950 676.950 769.050 677.400 ;
        RECT 772.950 678.450 775.050 678.900 ;
        RECT 781.950 678.450 784.050 678.900 ;
        RECT 772.950 677.250 784.050 678.450 ;
        RECT 772.950 676.800 775.050 677.250 ;
        RECT 781.950 676.800 784.050 677.250 ;
        RECT 787.950 676.800 790.050 678.900 ;
        RECT 791.400 678.600 792.600 682.950 ;
        RECT 808.950 678.600 811.050 678.900 ;
        RECT 791.400 677.400 811.050 678.600 ;
        RECT 808.950 676.800 811.050 677.400 ;
        RECT 818.400 676.050 819.600 683.400 ;
        RECT 838.950 683.550 847.050 684.750 ;
        RECT 838.950 683.100 841.050 683.550 ;
        RECT 844.950 683.100 847.050 683.550 ;
        RECT 859.950 684.600 862.050 685.200 ;
        RECT 883.950 684.600 886.050 685.200 ;
        RECT 859.950 683.400 886.050 684.600 ;
        RECT 859.950 683.100 862.050 683.400 ;
        RECT 883.950 683.100 886.050 683.400 ;
        RECT 835.950 678.600 838.050 678.900 ;
        RECT 856.950 678.600 859.050 678.900 ;
        RECT 835.950 677.400 859.050 678.600 ;
        RECT 835.950 676.800 838.050 677.400 ;
        RECT 856.950 676.800 859.050 677.400 ;
        RECT 874.950 678.600 877.050 679.050 ;
        RECT 886.950 678.600 889.050 678.900 ;
        RECT 874.950 677.400 889.050 678.600 ;
        RECT 874.950 676.950 877.050 677.400 ;
        RECT 886.950 676.800 889.050 677.400 ;
        RECT 166.950 675.600 169.050 676.050 ;
        RECT 181.950 675.600 184.050 676.050 ;
        RECT 166.950 674.400 184.050 675.600 ;
        RECT 166.950 673.950 169.050 674.400 ;
        RECT 181.950 673.950 184.050 674.400 ;
        RECT 283.950 675.600 286.050 676.050 ;
        RECT 304.950 675.600 307.050 676.050 ;
        RECT 322.950 675.600 325.050 676.050 ;
        RECT 283.950 674.400 325.050 675.600 ;
        RECT 283.950 673.950 286.050 674.400 ;
        RECT 304.950 673.950 307.050 674.400 ;
        RECT 322.950 673.950 325.050 674.400 ;
        RECT 472.950 675.600 475.050 676.050 ;
        RECT 478.950 675.600 481.050 676.050 ;
        RECT 472.950 674.400 481.050 675.600 ;
        RECT 472.950 673.950 475.050 674.400 ;
        RECT 478.950 673.950 481.050 674.400 ;
        RECT 490.950 675.600 493.050 676.050 ;
        RECT 514.950 675.600 517.050 676.050 ;
        RECT 490.950 674.400 517.050 675.600 ;
        RECT 490.950 673.950 493.050 674.400 ;
        RECT 514.950 673.950 517.050 674.400 ;
        RECT 817.950 673.950 820.050 676.050 ;
        RECT 865.950 675.600 868.050 676.050 ;
        RECT 871.950 675.600 874.050 676.050 ;
        RECT 865.950 674.400 874.050 675.600 ;
        RECT 865.950 673.950 868.050 674.400 ;
        RECT 871.950 673.950 874.050 674.400 ;
        RECT 40.950 672.600 43.050 673.050 ;
        RECT 58.950 672.600 61.050 673.050 ;
        RECT 40.950 671.400 61.050 672.600 ;
        RECT 40.950 670.950 43.050 671.400 ;
        RECT 58.950 670.950 61.050 671.400 ;
        RECT 124.950 672.600 127.050 673.050 ;
        RECT 139.950 672.600 142.050 673.050 ;
        RECT 124.950 671.400 142.050 672.600 ;
        RECT 124.950 670.950 127.050 671.400 ;
        RECT 139.950 670.950 142.050 671.400 ;
        RECT 178.950 672.600 181.050 673.050 ;
        RECT 184.950 672.600 187.050 673.050 ;
        RECT 178.950 671.400 187.050 672.600 ;
        RECT 178.950 670.950 181.050 671.400 ;
        RECT 184.950 670.950 187.050 671.400 ;
        RECT 193.950 672.600 196.050 673.050 ;
        RECT 268.950 672.600 271.050 673.050 ;
        RECT 193.950 671.400 271.050 672.600 ;
        RECT 193.950 670.950 196.050 671.400 ;
        RECT 268.950 670.950 271.050 671.400 ;
        RECT 424.950 672.600 427.050 673.050 ;
        RECT 433.950 672.600 436.050 673.050 ;
        RECT 424.950 671.400 436.050 672.600 ;
        RECT 424.950 670.950 427.050 671.400 ;
        RECT 433.950 670.950 436.050 671.400 ;
        RECT 514.950 672.600 517.050 672.900 ;
        RECT 526.950 672.600 529.050 673.050 ;
        RECT 514.950 671.400 529.050 672.600 ;
        RECT 160.950 669.600 163.050 670.050 ;
        RECT 194.400 669.600 195.600 670.950 ;
        RECT 514.950 670.800 517.050 671.400 ;
        RECT 526.950 670.950 529.050 671.400 ;
        RECT 712.950 672.600 715.050 673.050 ;
        RECT 754.950 672.600 757.050 673.050 ;
        RECT 712.950 671.400 757.050 672.600 ;
        RECT 712.950 670.950 715.050 671.400 ;
        RECT 754.950 670.950 757.050 671.400 ;
        RECT 862.950 672.600 865.050 673.050 ;
        RECT 874.950 672.600 877.050 673.050 ;
        RECT 862.950 671.400 877.050 672.600 ;
        RECT 862.950 670.950 865.050 671.400 ;
        RECT 874.950 670.950 877.050 671.400 ;
        RECT 160.950 668.400 195.600 669.600 ;
        RECT 199.950 669.600 202.050 670.050 ;
        RECT 280.950 669.600 283.050 670.050 ;
        RECT 361.950 669.600 364.050 670.050 ;
        RECT 199.950 668.400 364.050 669.600 ;
        RECT 160.950 667.950 163.050 668.400 ;
        RECT 199.950 667.950 202.050 668.400 ;
        RECT 280.950 667.950 283.050 668.400 ;
        RECT 361.950 667.950 364.050 668.400 ;
        RECT 400.950 669.600 403.050 670.050 ;
        RECT 436.950 669.600 439.050 670.050 ;
        RECT 400.950 668.400 439.050 669.600 ;
        RECT 400.950 667.950 403.050 668.400 ;
        RECT 436.950 667.950 439.050 668.400 ;
        RECT 562.950 669.600 565.050 670.050 ;
        RECT 583.950 669.600 586.050 670.050 ;
        RECT 562.950 668.400 586.050 669.600 ;
        RECT 562.950 667.950 565.050 668.400 ;
        RECT 583.950 667.950 586.050 668.400 ;
        RECT 658.950 669.600 661.050 670.050 ;
        RECT 682.950 669.600 685.050 670.050 ;
        RECT 709.950 669.600 712.050 670.050 ;
        RECT 658.950 668.400 712.050 669.600 ;
        RECT 658.950 667.950 661.050 668.400 ;
        RECT 682.950 667.950 685.050 668.400 ;
        RECT 709.950 667.950 712.050 668.400 ;
        RECT 784.950 669.600 787.050 670.050 ;
        RECT 802.950 669.600 805.050 670.050 ;
        RECT 784.950 668.400 805.050 669.600 ;
        RECT 784.950 667.950 787.050 668.400 ;
        RECT 802.950 667.950 805.050 668.400 ;
        RECT 832.950 669.600 835.050 670.050 ;
        RECT 847.950 669.600 850.050 670.050 ;
        RECT 832.950 668.400 850.050 669.600 ;
        RECT 832.950 667.950 835.050 668.400 ;
        RECT 847.950 667.950 850.050 668.400 ;
        RECT 232.950 666.600 235.050 667.050 ;
        RECT 298.950 666.600 301.050 667.050 ;
        RECT 355.950 666.600 358.050 667.050 ;
        RECT 232.950 665.400 279.600 666.600 ;
        RECT 232.950 664.950 235.050 665.400 ;
        RECT 22.950 663.600 25.050 664.050 ;
        RECT 55.950 663.600 58.050 664.050 ;
        RECT 79.950 663.600 82.050 664.050 ;
        RECT 22.950 662.400 82.050 663.600 ;
        RECT 22.950 661.950 25.050 662.400 ;
        RECT 55.950 661.950 58.050 662.400 ;
        RECT 79.950 661.950 82.050 662.400 ;
        RECT 154.950 663.600 157.050 664.050 ;
        RECT 190.950 663.600 193.050 664.050 ;
        RECT 154.950 662.400 193.050 663.600 ;
        RECT 278.400 663.600 279.600 665.400 ;
        RECT 298.950 665.400 358.050 666.600 ;
        RECT 298.950 664.950 301.050 665.400 ;
        RECT 355.950 664.950 358.050 665.400 ;
        RECT 388.950 666.600 391.050 667.050 ;
        RECT 412.950 666.600 415.050 667.050 ;
        RECT 388.950 665.400 415.050 666.600 ;
        RECT 388.950 664.950 391.050 665.400 ;
        RECT 412.950 664.950 415.050 665.400 ;
        RECT 439.950 666.600 442.050 667.050 ;
        RECT 487.950 666.600 490.050 667.050 ;
        RECT 439.950 665.400 490.050 666.600 ;
        RECT 439.950 664.950 442.050 665.400 ;
        RECT 487.950 664.950 490.050 665.400 ;
        RECT 286.950 663.600 289.050 664.050 ;
        RECT 278.400 662.400 289.050 663.600 ;
        RECT 154.950 661.950 157.050 662.400 ;
        RECT 190.950 661.950 193.050 662.400 ;
        RECT 286.950 661.950 289.050 662.400 ;
        RECT 574.950 663.600 577.050 664.050 ;
        RECT 625.950 663.600 628.050 664.050 ;
        RECT 574.950 662.400 628.050 663.600 ;
        RECT 574.950 661.950 577.050 662.400 ;
        RECT 625.950 661.950 628.050 662.400 ;
        RECT 676.950 663.600 679.050 664.050 ;
        RECT 691.950 663.600 694.050 664.050 ;
        RECT 676.950 662.400 694.050 663.600 ;
        RECT 676.950 661.950 679.050 662.400 ;
        RECT 691.950 661.950 694.050 662.400 ;
        RECT 799.950 663.600 802.050 664.050 ;
        RECT 820.950 663.600 823.050 664.050 ;
        RECT 862.950 663.600 865.050 664.050 ;
        RECT 799.950 662.400 865.050 663.600 ;
        RECT 799.950 661.950 802.050 662.400 ;
        RECT 820.950 661.950 823.050 662.400 ;
        RECT 862.950 661.950 865.050 662.400 ;
        RECT 655.950 660.600 658.050 661.050 ;
        RECT 703.950 660.600 706.050 661.050 ;
        RECT 655.950 659.400 706.050 660.600 ;
        RECT 655.950 658.950 658.050 659.400 ;
        RECT 703.950 658.950 706.050 659.400 ;
        RECT 742.950 660.600 745.050 661.050 ;
        RECT 763.950 660.600 766.050 661.050 ;
        RECT 742.950 659.400 766.050 660.600 ;
        RECT 742.950 658.950 745.050 659.400 ;
        RECT 763.950 658.950 766.050 659.400 ;
        RECT 37.950 657.600 40.050 658.050 ;
        RECT 103.950 657.600 106.050 658.050 ;
        RECT 37.950 656.400 106.050 657.600 ;
        RECT 37.950 655.950 40.050 656.400 ;
        RECT 103.950 655.950 106.050 656.400 ;
        RECT 109.950 657.600 112.050 658.050 ;
        RECT 130.950 657.600 133.050 658.050 ;
        RECT 151.950 657.600 154.050 658.050 ;
        RECT 109.950 656.400 154.050 657.600 ;
        RECT 109.950 655.950 112.050 656.400 ;
        RECT 130.950 655.950 133.050 656.400 ;
        RECT 151.950 655.950 154.050 656.400 ;
        RECT 166.950 657.600 169.050 658.050 ;
        RECT 229.950 657.600 232.050 658.050 ;
        RECT 166.950 656.400 232.050 657.600 ;
        RECT 166.950 655.950 169.050 656.400 ;
        RECT 229.950 655.950 232.050 656.400 ;
        RECT 316.950 657.600 319.050 658.050 ;
        RECT 379.950 657.600 382.050 658.050 ;
        RECT 409.950 657.600 412.050 658.050 ;
        RECT 424.950 657.600 427.050 658.050 ;
        RECT 316.950 656.400 427.050 657.600 ;
        RECT 316.950 655.950 319.050 656.400 ;
        RECT 379.950 655.950 382.050 656.400 ;
        RECT 409.950 655.950 412.050 656.400 ;
        RECT 424.950 655.950 427.050 656.400 ;
        RECT 535.950 657.600 538.050 658.050 ;
        RECT 580.950 657.600 583.050 658.050 ;
        RECT 535.950 656.400 583.050 657.600 ;
        RECT 535.950 655.950 538.050 656.400 ;
        RECT 580.950 655.950 583.050 656.400 ;
        RECT 607.950 657.600 610.050 658.050 ;
        RECT 637.950 657.600 640.050 658.050 ;
        RECT 685.950 657.600 688.050 658.050 ;
        RECT 607.950 656.400 688.050 657.600 ;
        RECT 607.950 655.950 610.050 656.400 ;
        RECT 637.950 655.950 640.050 656.400 ;
        RECT 685.950 655.950 688.050 656.400 ;
        RECT 748.950 657.600 753.000 658.050 ;
        RECT 850.950 657.600 853.050 658.050 ;
        RECT 859.950 657.600 862.050 658.050 ;
        RECT 748.950 655.950 753.600 657.600 ;
        RECT 850.950 656.400 862.050 657.600 ;
        RECT 850.950 655.950 853.050 656.400 ;
        RECT 859.950 655.950 862.050 656.400 ;
        RECT 313.950 654.600 316.050 655.050 ;
        RECT 302.400 653.400 316.050 654.600 ;
        RECT 22.950 651.600 25.050 652.200 ;
        RECT 37.950 651.600 40.050 652.200 ;
        RECT 22.950 650.400 40.050 651.600 ;
        RECT 22.950 650.100 25.050 650.400 ;
        RECT 37.950 650.100 40.050 650.400 ;
        RECT 61.950 651.600 64.050 652.200 ;
        RECT 118.950 651.600 121.050 652.050 ;
        RECT 124.950 651.600 127.050 652.200 ;
        RECT 61.950 650.400 121.050 651.600 ;
        RECT 61.950 650.100 64.050 650.400 ;
        RECT 118.950 649.950 121.050 650.400 ;
        RECT 122.400 650.400 127.050 651.600 ;
        RECT 122.400 646.050 123.600 650.400 ;
        RECT 124.950 650.100 127.050 650.400 ;
        RECT 157.950 651.600 160.050 652.200 ;
        RECT 166.800 651.600 168.900 652.050 ;
        RECT 157.950 650.400 168.900 651.600 ;
        RECT 157.950 650.100 160.050 650.400 ;
        RECT 166.800 649.950 168.900 650.400 ;
        RECT 169.950 651.750 172.050 652.200 ;
        RECT 175.950 651.750 178.050 652.200 ;
        RECT 169.950 650.550 178.050 651.750 ;
        RECT 169.950 650.100 172.050 650.550 ;
        RECT 175.950 650.100 178.050 650.550 ;
        RECT 211.950 651.600 214.050 652.050 ;
        RECT 223.950 651.600 226.050 652.200 ;
        RECT 211.950 650.400 226.050 651.600 ;
        RECT 211.950 649.950 214.050 650.400 ;
        RECT 223.950 650.100 226.050 650.400 ;
        RECT 229.950 651.600 232.050 652.200 ;
        RECT 247.950 651.600 250.050 652.200 ;
        RECT 229.950 650.400 250.050 651.600 ;
        RECT 229.950 650.100 232.050 650.400 ;
        RECT 247.950 650.100 250.050 650.400 ;
        RECT 256.950 651.600 259.050 652.050 ;
        RECT 274.950 651.600 277.050 652.200 ;
        RECT 302.400 651.600 303.600 653.400 ;
        RECT 313.950 652.950 316.050 653.400 ;
        RECT 322.950 654.600 325.050 655.050 ;
        RECT 355.950 654.600 358.050 655.050 ;
        RECT 322.950 653.400 358.050 654.600 ;
        RECT 322.950 652.950 325.050 653.400 ;
        RECT 355.950 652.950 358.050 653.400 ;
        RECT 385.950 654.600 388.050 655.050 ;
        RECT 400.950 654.600 403.050 655.050 ;
        RECT 385.950 653.400 403.050 654.600 ;
        RECT 385.950 652.950 388.050 653.400 ;
        RECT 400.950 652.950 403.050 653.400 ;
        RECT 493.950 654.600 496.050 655.050 ;
        RECT 505.950 654.600 508.050 655.050 ;
        RECT 493.950 653.400 508.050 654.600 ;
        RECT 752.400 654.600 753.600 655.950 ;
        RECT 769.950 654.600 772.050 655.050 ;
        RECT 752.400 653.400 772.050 654.600 ;
        RECT 493.950 652.950 496.050 653.400 ;
        RECT 505.950 652.950 508.050 653.400 ;
        RECT 769.950 652.950 772.050 653.400 ;
        RECT 796.950 654.600 799.050 655.050 ;
        RECT 808.950 654.600 811.050 655.050 ;
        RECT 796.950 653.400 811.050 654.600 ;
        RECT 796.950 652.950 799.050 653.400 ;
        RECT 808.950 652.950 811.050 653.400 ;
        RECT 256.950 650.400 303.600 651.600 ;
        RECT 343.950 651.750 346.050 652.200 ;
        RECT 379.950 651.750 382.050 652.200 ;
        RECT 343.950 650.550 382.050 651.750 ;
        RECT 256.950 649.950 259.050 650.400 ;
        RECT 274.950 650.100 277.050 650.400 ;
        RECT 343.950 650.100 346.050 650.550 ;
        RECT 379.950 650.100 382.050 650.550 ;
        RECT 415.950 651.600 418.050 652.200 ;
        RECT 433.950 651.600 436.050 652.200 ;
        RECT 415.950 650.400 436.050 651.600 ;
        RECT 415.950 650.100 418.050 650.400 ;
        RECT 433.950 650.100 436.050 650.400 ;
        RECT 445.950 651.600 448.050 652.050 ;
        RECT 454.950 651.600 457.050 652.200 ;
        RECT 445.950 650.400 457.050 651.600 ;
        RECT 445.950 649.950 448.050 650.400 ;
        RECT 454.950 650.100 457.050 650.400 ;
        RECT 481.950 651.600 484.050 652.200 ;
        RECT 490.950 651.600 493.050 652.050 ;
        RECT 481.950 650.400 493.050 651.600 ;
        RECT 481.950 650.100 484.050 650.400 ;
        RECT 490.950 649.950 493.050 650.400 ;
        RECT 499.950 650.100 502.050 652.200 ;
        RECT 526.950 651.750 529.050 652.200 ;
        RECT 538.950 651.750 541.050 652.200 ;
        RECT 526.950 650.550 541.050 651.750 ;
        RECT 526.950 650.100 529.050 650.550 ;
        RECT 538.950 650.100 541.050 650.550 ;
        RECT 544.950 651.600 547.050 652.200 ;
        RECT 574.950 651.600 577.050 652.200 ;
        RECT 544.950 650.400 577.050 651.600 ;
        RECT 544.950 650.100 547.050 650.400 ;
        RECT 574.950 650.100 577.050 650.400 ;
        RECT 586.950 650.100 589.050 652.200 ;
        RECT 646.950 651.600 649.050 652.200 ;
        RECT 658.950 651.600 661.050 652.050 ;
        RECT 664.950 651.600 667.050 652.200 ;
        RECT 646.950 650.400 667.050 651.600 ;
        RECT 646.950 650.100 649.050 650.400 ;
        RECT 500.400 648.600 501.600 650.100 ;
        RECT 431.400 647.400 501.600 648.600 ;
        RECT 40.950 645.600 43.050 645.900 ;
        RECT 58.950 645.600 61.050 645.900 ;
        RECT 40.950 644.400 61.050 645.600 ;
        RECT 40.950 643.800 43.050 644.400 ;
        RECT 58.950 643.800 61.050 644.400 ;
        RECT 64.950 645.450 67.050 645.900 ;
        RECT 70.950 645.450 73.050 645.900 ;
        RECT 64.950 644.250 73.050 645.450 ;
        RECT 64.950 643.800 67.050 644.250 ;
        RECT 70.950 643.800 73.050 644.250 ;
        RECT 91.950 645.450 94.050 645.900 ;
        RECT 100.950 645.450 103.050 645.900 ;
        RECT 91.950 644.250 103.050 645.450 ;
        RECT 91.950 643.800 94.050 644.250 ;
        RECT 100.950 643.800 103.050 644.250 ;
        RECT 121.950 643.950 124.050 646.050 ;
        RECT 133.950 645.600 136.050 645.900 ;
        RECT 154.950 645.600 157.050 645.900 ;
        RECT 133.950 644.400 157.050 645.600 ;
        RECT 133.950 643.800 136.050 644.400 ;
        RECT 154.950 643.800 157.050 644.400 ;
        RECT 166.950 645.450 169.050 645.900 ;
        RECT 178.950 645.450 181.050 645.900 ;
        RECT 166.950 644.250 181.050 645.450 ;
        RECT 166.950 643.800 169.050 644.250 ;
        RECT 178.950 643.800 181.050 644.250 ;
        RECT 265.950 645.450 268.050 645.900 ;
        RECT 280.950 645.450 283.050 646.050 ;
        RECT 265.950 644.250 283.050 645.450 ;
        RECT 265.950 643.800 268.050 644.250 ;
        RECT 280.950 643.950 283.050 644.250 ;
        RECT 343.950 645.450 346.050 645.900 ;
        RECT 364.950 645.450 367.050 645.900 ;
        RECT 343.950 644.250 367.050 645.450 ;
        RECT 343.950 643.800 346.050 644.250 ;
        RECT 364.950 643.800 367.050 644.250 ;
        RECT 412.950 645.600 415.050 645.900 ;
        RECT 431.400 645.600 432.600 647.400 ;
        RECT 412.950 644.400 432.600 645.600 ;
        RECT 436.950 645.450 439.050 645.900 ;
        RECT 445.950 645.450 448.050 645.900 ;
        RECT 412.950 643.800 415.050 644.400 ;
        RECT 436.950 644.250 448.050 645.450 ;
        RECT 436.950 643.800 439.050 644.250 ;
        RECT 445.950 643.800 448.050 644.250 ;
        RECT 457.950 645.600 460.050 645.900 ;
        RECT 490.950 645.600 493.050 645.900 ;
        RECT 457.950 645.450 493.050 645.600 ;
        RECT 502.950 645.450 505.050 645.900 ;
        RECT 457.950 644.400 505.050 645.450 ;
        RECT 457.950 643.800 460.050 644.400 ;
        RECT 490.950 644.250 505.050 644.400 ;
        RECT 490.950 643.800 493.050 644.250 ;
        RECT 502.950 643.800 505.050 644.250 ;
        RECT 508.950 645.600 511.050 645.900 ;
        RECT 514.950 645.600 517.050 646.050 ;
        RECT 508.950 644.400 517.050 645.600 ;
        RECT 508.950 643.800 511.050 644.400 ;
        RECT 514.950 643.950 517.050 644.400 ;
        RECT 565.950 645.450 568.050 645.900 ;
        RECT 577.950 645.450 580.050 645.900 ;
        RECT 565.950 644.250 580.050 645.450 ;
        RECT 587.400 645.600 588.600 650.100 ;
        RECT 658.950 649.950 661.050 650.400 ;
        RECT 664.950 650.100 667.050 650.400 ;
        RECT 691.950 651.750 694.050 652.200 ;
        RECT 697.950 651.750 700.050 652.200 ;
        RECT 691.950 650.550 700.050 651.750 ;
        RECT 691.950 650.100 694.050 650.550 ;
        RECT 697.950 650.100 700.050 650.550 ;
        RECT 775.950 651.600 778.050 652.200 ;
        RECT 787.950 651.600 790.050 652.050 ;
        RECT 775.950 650.400 790.050 651.600 ;
        RECT 775.950 650.100 778.050 650.400 ;
        RECT 787.950 649.950 790.050 650.400 ;
        RECT 814.950 649.950 817.050 652.050 ;
        RECT 823.950 651.600 826.050 652.200 ;
        RECT 844.950 651.600 847.050 652.200 ;
        RECT 823.950 650.400 847.050 651.600 ;
        RECT 823.950 650.100 826.050 650.400 ;
        RECT 844.950 650.100 847.050 650.400 ;
        RECT 850.950 650.100 853.050 652.200 ;
        RECT 856.950 651.600 859.050 652.050 ;
        RECT 868.950 651.600 871.050 652.200 ;
        RECT 856.950 650.400 871.050 651.600 ;
        RECT 784.950 648.600 787.050 649.050 ;
        RECT 773.400 647.400 787.050 648.600 ;
        RECT 604.950 645.600 607.050 645.900 ;
        RECT 587.400 644.400 607.050 645.600 ;
        RECT 565.950 643.800 568.050 644.250 ;
        RECT 577.950 643.800 580.050 644.250 ;
        RECT 604.950 643.800 607.050 644.400 ;
        RECT 613.950 645.600 616.050 646.050 ;
        RECT 622.950 645.600 625.050 645.900 ;
        RECT 613.950 644.400 625.050 645.600 ;
        RECT 613.950 643.950 616.050 644.400 ;
        RECT 622.950 643.800 625.050 644.400 ;
        RECT 628.950 645.450 631.050 645.900 ;
        RECT 637.950 645.450 640.050 645.900 ;
        RECT 628.950 644.250 640.050 645.450 ;
        RECT 628.950 643.800 631.050 644.250 ;
        RECT 637.950 643.800 640.050 644.250 ;
        RECT 649.950 645.600 652.050 645.900 ;
        RECT 655.950 645.600 658.050 646.050 ;
        RECT 773.400 645.900 774.600 647.400 ;
        RECT 784.950 646.950 787.050 647.400 ;
        RECT 649.950 644.400 658.050 645.600 ;
        RECT 649.950 643.800 652.050 644.400 ;
        RECT 655.950 643.950 658.050 644.400 ;
        RECT 706.950 645.600 709.050 645.900 ;
        RECT 739.950 645.600 742.050 645.900 ;
        RECT 706.950 644.400 742.050 645.600 ;
        RECT 706.950 643.800 709.050 644.400 ;
        RECT 739.950 643.800 742.050 644.400 ;
        RECT 772.950 643.800 775.050 645.900 ;
        RECT 796.950 645.600 799.050 645.900 ;
        RECT 815.400 645.600 816.600 649.950 ;
        RECT 851.400 648.600 852.600 650.100 ;
        RECT 856.950 649.950 859.050 650.400 ;
        RECT 868.950 650.100 871.050 650.400 ;
        RECT 880.950 651.600 883.050 652.050 ;
        RECT 889.950 651.600 892.050 652.200 ;
        RECT 880.950 650.400 892.050 651.600 ;
        RECT 851.400 648.000 855.600 648.600 ;
        RECT 851.400 647.400 856.050 648.000 ;
        RECT 796.950 644.400 816.600 645.600 ;
        RECT 796.950 643.800 799.050 644.400 ;
        RECT 853.950 643.950 856.050 647.400 ;
        RECT 869.400 645.600 870.600 650.100 ;
        RECT 880.950 649.950 883.050 650.400 ;
        RECT 889.950 650.100 892.050 650.400 ;
        RECT 898.950 649.950 901.050 652.050 ;
        RECT 899.400 646.050 900.600 649.950 ;
        RECT 886.950 645.600 889.050 645.900 ;
        RECT 869.400 644.400 889.050 645.600 ;
        RECT 886.950 643.800 889.050 644.400 ;
        RECT 898.950 643.950 901.050 646.050 ;
        RECT 118.950 642.600 121.050 643.050 ;
        RECT 127.950 642.600 130.050 643.050 ;
        RECT 118.950 641.400 130.050 642.600 ;
        RECT 118.950 640.950 121.050 641.400 ;
        RECT 127.950 640.950 130.050 641.400 ;
        RECT 202.950 642.600 205.050 643.050 ;
        RECT 226.950 642.600 229.050 643.050 ;
        RECT 202.950 641.400 229.050 642.600 ;
        RECT 202.950 640.950 205.050 641.400 ;
        RECT 226.950 640.950 229.050 641.400 ;
        RECT 280.950 642.600 283.050 642.900 ;
        RECT 295.950 642.600 298.050 643.050 ;
        RECT 280.950 641.400 298.050 642.600 ;
        RECT 280.950 640.800 283.050 641.400 ;
        RECT 295.950 640.950 298.050 641.400 ;
        RECT 424.950 642.600 427.050 643.050 ;
        RECT 478.950 642.600 481.050 643.050 ;
        RECT 523.950 642.600 526.050 643.050 ;
        RECT 424.950 641.400 526.050 642.600 ;
        RECT 424.950 640.950 427.050 641.400 ;
        RECT 478.950 640.950 481.050 641.400 ;
        RECT 523.950 640.950 526.050 641.400 ;
        RECT 583.950 642.600 586.050 643.050 ;
        RECT 598.950 642.600 601.050 643.050 ;
        RECT 583.950 641.400 601.050 642.600 ;
        RECT 583.950 640.950 586.050 641.400 ;
        RECT 598.950 640.950 601.050 641.400 ;
        RECT 676.950 642.600 679.050 643.050 ;
        RECT 682.950 642.600 685.050 643.050 ;
        RECT 676.950 641.400 685.050 642.600 ;
        RECT 676.950 640.950 679.050 641.400 ;
        RECT 682.950 640.950 685.050 641.400 ;
        RECT 763.950 642.600 766.050 643.050 ;
        RECT 778.950 642.600 781.050 643.050 ;
        RECT 763.950 641.400 781.050 642.600 ;
        RECT 763.950 640.950 766.050 641.400 ;
        RECT 778.950 640.950 781.050 641.400 ;
        RECT 331.950 639.600 334.050 640.050 ;
        RECT 388.950 639.600 391.050 640.050 ;
        RECT 331.950 638.400 391.050 639.600 ;
        RECT 331.950 637.950 334.050 638.400 ;
        RECT 388.950 637.950 391.050 638.400 ;
        RECT 820.950 639.600 823.050 639.900 ;
        RECT 832.950 639.600 835.050 640.050 ;
        RECT 820.950 638.400 835.050 639.600 ;
        RECT 820.950 637.800 823.050 638.400 ;
        RECT 832.950 637.950 835.050 638.400 ;
        RECT 862.950 639.600 865.050 640.050 ;
        RECT 892.950 639.600 895.050 640.050 ;
        RECT 862.950 638.400 895.050 639.600 ;
        RECT 862.950 637.950 865.050 638.400 ;
        RECT 892.950 637.950 895.050 638.400 ;
        RECT 121.950 636.600 124.050 637.050 ;
        RECT 175.950 636.600 178.050 637.050 ;
        RECT 184.950 636.600 187.050 637.050 ;
        RECT 190.950 636.600 193.050 637.050 ;
        RECT 121.950 635.400 193.050 636.600 ;
        RECT 121.950 634.950 124.050 635.400 ;
        RECT 175.950 634.950 178.050 635.400 ;
        RECT 184.950 634.950 187.050 635.400 ;
        RECT 190.950 634.950 193.050 635.400 ;
        RECT 205.950 636.600 208.050 637.050 ;
        RECT 220.950 636.600 223.050 637.050 ;
        RECT 271.950 636.600 274.050 637.050 ;
        RECT 205.950 635.400 274.050 636.600 ;
        RECT 205.950 634.950 208.050 635.400 ;
        RECT 220.950 634.950 223.050 635.400 ;
        RECT 271.950 634.950 274.050 635.400 ;
        RECT 382.950 636.600 385.050 637.050 ;
        RECT 412.950 636.600 415.050 637.050 ;
        RECT 382.950 635.400 415.050 636.600 ;
        RECT 382.950 634.950 385.050 635.400 ;
        RECT 412.950 634.950 415.050 635.400 ;
        RECT 493.950 636.600 496.050 637.050 ;
        RECT 649.950 636.600 652.050 637.050 ;
        RECT 493.950 635.400 652.050 636.600 ;
        RECT 493.950 634.950 496.050 635.400 ;
        RECT 649.950 634.950 652.050 635.400 ;
        RECT 847.950 636.600 850.050 637.050 ;
        RECT 871.950 636.600 874.050 637.050 ;
        RECT 847.950 635.400 874.050 636.600 ;
        RECT 847.950 634.950 850.050 635.400 ;
        RECT 871.950 634.950 874.050 635.400 ;
        RECT 13.950 633.600 16.050 634.050 ;
        RECT 34.950 633.600 37.050 634.050 ;
        RECT 199.950 633.600 202.050 634.050 ;
        RECT 349.950 633.600 352.050 634.050 ;
        RECT 13.950 632.400 352.050 633.600 ;
        RECT 13.950 631.950 16.050 632.400 ;
        RECT 34.950 631.950 37.050 632.400 ;
        RECT 199.950 631.950 202.050 632.400 ;
        RECT 349.950 631.950 352.050 632.400 ;
        RECT 460.950 633.600 463.050 634.050 ;
        RECT 508.950 633.600 511.050 634.050 ;
        RECT 460.950 632.400 511.050 633.600 ;
        RECT 460.950 631.950 463.050 632.400 ;
        RECT 508.950 631.950 511.050 632.400 ;
        RECT 169.950 630.600 172.050 631.050 ;
        RECT 205.950 630.600 208.050 631.050 ;
        RECT 169.950 629.400 208.050 630.600 ;
        RECT 169.950 628.950 172.050 629.400 ;
        RECT 205.950 628.950 208.050 629.400 ;
        RECT 262.950 630.600 265.050 631.050 ;
        RECT 322.950 630.600 325.050 631.050 ;
        RECT 262.950 629.400 325.050 630.600 ;
        RECT 262.950 628.950 265.050 629.400 ;
        RECT 322.950 628.950 325.050 629.400 ;
        RECT 625.950 630.600 628.050 631.050 ;
        RECT 796.950 630.600 799.050 631.050 ;
        RECT 823.950 630.600 826.050 631.050 ;
        RECT 625.950 629.400 826.050 630.600 ;
        RECT 625.950 628.950 628.050 629.400 ;
        RECT 796.950 628.950 799.050 629.400 ;
        RECT 823.950 628.950 826.050 629.400 ;
        RECT 838.950 630.600 841.050 631.050 ;
        RECT 856.950 630.600 859.050 631.050 ;
        RECT 838.950 629.400 859.050 630.600 ;
        RECT 838.950 628.950 841.050 629.400 ;
        RECT 856.950 628.950 859.050 629.400 ;
        RECT 208.950 627.600 211.050 628.050 ;
        RECT 250.950 627.600 253.050 628.050 ;
        RECT 208.950 626.400 253.050 627.600 ;
        RECT 208.950 625.950 211.050 626.400 ;
        RECT 250.950 625.950 253.050 626.400 ;
        RECT 643.950 627.600 646.050 628.050 ;
        RECT 724.950 627.600 727.050 628.050 ;
        RECT 757.950 627.600 760.050 628.050 ;
        RECT 643.950 626.400 760.050 627.600 ;
        RECT 643.950 625.950 646.050 626.400 ;
        RECT 724.950 625.950 727.050 626.400 ;
        RECT 757.950 625.950 760.050 626.400 ;
        RECT 418.950 624.600 421.050 625.050 ;
        RECT 644.400 624.600 645.600 625.950 ;
        RECT 418.950 623.400 645.600 624.600 ;
        RECT 688.950 624.600 691.050 625.050 ;
        RECT 697.950 624.600 700.050 625.050 ;
        RECT 688.950 623.400 700.050 624.600 ;
        RECT 418.950 622.950 421.050 623.400 ;
        RECT 688.950 622.950 691.050 623.400 ;
        RECT 697.950 622.950 700.050 623.400 ;
        RECT 130.950 621.600 133.050 622.050 ;
        RECT 211.950 621.600 214.050 622.050 ;
        RECT 130.950 620.400 214.050 621.600 ;
        RECT 130.950 619.950 133.050 620.400 ;
        RECT 211.950 619.950 214.050 620.400 ;
        RECT 526.950 621.600 529.050 622.050 ;
        RECT 535.800 621.600 537.900 622.050 ;
        RECT 526.950 620.400 537.900 621.600 ;
        RECT 526.950 619.950 529.050 620.400 ;
        RECT 535.800 619.950 537.900 620.400 ;
        RECT 538.950 621.600 541.050 622.050 ;
        RECT 553.950 621.600 556.050 622.050 ;
        RECT 538.950 620.400 556.050 621.600 ;
        RECT 538.950 619.950 541.050 620.400 ;
        RECT 553.950 619.950 556.050 620.400 ;
        RECT 631.950 621.600 634.050 622.050 ;
        RECT 718.950 621.600 721.050 622.050 ;
        RECT 631.950 620.400 721.050 621.600 ;
        RECT 631.950 619.950 634.050 620.400 ;
        RECT 718.950 619.950 721.050 620.400 ;
        RECT 808.950 621.600 811.050 622.050 ;
        RECT 865.950 621.600 868.050 622.050 ;
        RECT 808.950 620.400 868.050 621.600 ;
        RECT 808.950 619.950 811.050 620.400 ;
        RECT 865.950 619.950 868.050 620.400 ;
        RECT 277.950 618.600 280.050 619.050 ;
        RECT 343.950 618.600 346.050 619.050 ;
        RECT 277.950 617.400 346.050 618.600 ;
        RECT 277.950 616.950 280.050 617.400 ;
        RECT 343.950 616.950 346.050 617.400 ;
        RECT 523.950 618.600 526.050 619.050 ;
        RECT 568.950 618.600 571.050 619.050 ;
        RECT 583.950 618.600 586.050 619.050 ;
        RECT 523.950 617.400 586.050 618.600 ;
        RECT 523.950 616.950 526.050 617.400 ;
        RECT 568.950 616.950 571.050 617.400 ;
        RECT 583.950 616.950 586.050 617.400 ;
        RECT 589.950 618.600 592.050 619.050 ;
        RECT 802.950 618.600 805.050 619.050 ;
        RECT 811.950 618.600 814.050 619.050 ;
        RECT 835.950 618.600 838.050 619.050 ;
        RECT 589.950 617.400 838.050 618.600 ;
        RECT 589.950 616.950 592.050 617.400 ;
        RECT 802.950 616.950 805.050 617.400 ;
        RECT 811.950 616.950 814.050 617.400 ;
        RECT 835.950 616.950 838.050 617.400 ;
        RECT 541.950 615.600 544.050 616.050 ;
        RECT 559.950 615.600 562.050 616.050 ;
        RECT 541.950 614.400 562.050 615.600 ;
        RECT 541.950 613.950 544.050 614.400 ;
        RECT 559.950 613.950 562.050 614.400 ;
        RECT 616.950 615.600 619.050 616.050 ;
        RECT 643.950 615.600 646.050 616.050 ;
        RECT 616.950 614.400 646.050 615.600 ;
        RECT 616.950 613.950 619.050 614.400 ;
        RECT 643.950 613.950 646.050 614.400 ;
        RECT 52.950 612.600 55.050 613.050 ;
        RECT 58.950 612.600 61.050 613.050 ;
        RECT 52.950 611.400 61.050 612.600 ;
        RECT 52.950 610.950 55.050 611.400 ;
        RECT 58.950 610.950 61.050 611.400 ;
        RECT 94.950 612.600 97.050 613.050 ;
        RECT 127.950 612.600 130.050 613.050 ;
        RECT 136.950 612.600 139.050 613.050 ;
        RECT 94.950 611.400 123.600 612.600 ;
        RECT 94.950 610.950 97.050 611.400 ;
        RECT 122.400 609.600 123.600 611.400 ;
        RECT 127.950 611.400 139.050 612.600 ;
        RECT 127.950 610.950 130.050 611.400 ;
        RECT 136.950 610.950 139.050 611.400 ;
        RECT 154.950 612.600 157.050 613.050 ;
        RECT 166.950 612.600 169.050 612.900 ;
        RECT 154.950 611.400 169.050 612.600 ;
        RECT 154.950 610.950 157.050 611.400 ;
        RECT 166.950 610.800 169.050 611.400 ;
        RECT 184.950 612.600 187.050 613.050 ;
        RECT 208.950 612.600 211.050 613.050 ;
        RECT 184.950 611.400 211.050 612.600 ;
        RECT 184.950 610.950 187.050 611.400 ;
        RECT 208.950 610.950 211.050 611.400 ;
        RECT 289.950 612.600 292.050 613.050 ;
        RECT 319.950 612.600 322.050 613.050 ;
        RECT 289.950 611.400 322.050 612.600 ;
        RECT 289.950 610.950 292.050 611.400 ;
        RECT 319.950 610.950 322.050 611.400 ;
        RECT 376.950 612.600 379.050 613.050 ;
        RECT 382.950 612.600 385.050 613.050 ;
        RECT 391.950 612.600 394.050 613.050 ;
        RECT 376.950 611.400 394.050 612.600 ;
        RECT 376.950 610.950 379.050 611.400 ;
        RECT 382.950 610.950 385.050 611.400 ;
        RECT 391.950 610.950 394.050 611.400 ;
        RECT 520.950 612.600 523.050 613.050 ;
        RECT 538.950 612.600 541.050 612.900 ;
        RECT 520.950 611.400 541.050 612.600 ;
        RECT 520.950 610.950 523.050 611.400 ;
        RECT 538.950 610.800 541.050 611.400 ;
        RECT 550.950 612.600 553.050 613.050 ;
        RECT 574.950 612.600 577.050 613.050 ;
        RECT 550.950 611.400 577.050 612.600 ;
        RECT 550.950 610.950 553.050 611.400 ;
        RECT 574.950 610.950 577.050 611.400 ;
        RECT 658.950 612.600 661.050 613.050 ;
        RECT 706.950 612.600 709.050 613.050 ;
        RECT 736.950 612.600 739.050 613.050 ;
        RECT 745.950 612.600 748.050 613.050 ;
        RECT 658.950 611.400 748.050 612.600 ;
        RECT 658.950 610.950 661.050 611.400 ;
        RECT 706.950 610.950 709.050 611.400 ;
        RECT 736.950 610.950 739.050 611.400 ;
        RECT 745.950 610.950 748.050 611.400 ;
        RECT 757.950 612.600 760.050 613.050 ;
        RECT 778.950 612.600 781.050 613.050 ;
        RECT 790.950 612.600 793.050 613.050 ;
        RECT 757.950 611.400 793.050 612.600 ;
        RECT 757.950 610.950 760.050 611.400 ;
        RECT 778.950 610.950 781.050 611.400 ;
        RECT 790.950 610.950 793.050 611.400 ;
        RECT 844.950 612.600 847.050 613.050 ;
        RECT 853.950 612.600 856.050 613.050 ;
        RECT 844.950 611.400 856.050 612.600 ;
        RECT 844.950 610.950 847.050 611.400 ;
        RECT 853.950 610.950 856.050 611.400 ;
        RECT 877.950 612.600 880.050 613.050 ;
        RECT 889.950 612.600 892.050 613.050 ;
        RECT 877.950 611.400 892.050 612.600 ;
        RECT 877.950 610.950 880.050 611.400 ;
        RECT 889.950 610.950 892.050 611.400 ;
        RECT 148.950 609.600 151.050 610.050 ;
        RECT 122.400 608.400 151.050 609.600 ;
        RECT 148.950 607.950 151.050 608.400 ;
        RECT 304.950 609.600 307.050 610.050 ;
        RECT 331.950 609.600 334.050 610.050 ;
        RECT 304.950 608.400 334.050 609.600 ;
        RECT 304.950 607.950 307.050 608.400 ;
        RECT 331.950 607.950 334.050 608.400 ;
        RECT 541.950 609.600 544.050 609.900 ;
        RECT 553.950 609.600 556.050 610.050 ;
        RECT 577.950 609.600 580.050 610.050 ;
        RECT 541.950 608.400 580.050 609.600 ;
        RECT 541.950 607.800 544.050 608.400 ;
        RECT 553.950 607.950 556.050 608.400 ;
        RECT 577.950 607.950 580.050 608.400 ;
        RECT 583.950 609.600 586.050 610.050 ;
        RECT 604.950 609.600 607.050 610.050 ;
        RECT 583.950 608.400 607.050 609.600 ;
        RECT 583.950 607.950 586.050 608.400 ;
        RECT 604.950 607.950 607.050 608.400 ;
        RECT 610.950 609.600 613.050 610.050 ;
        RECT 619.950 609.600 622.050 610.050 ;
        RECT 610.950 608.400 622.050 609.600 ;
        RECT 610.950 607.950 613.050 608.400 ;
        RECT 619.950 607.950 622.050 608.400 ;
        RECT 841.950 609.600 844.050 610.050 ;
        RECT 859.950 609.600 862.050 610.050 ;
        RECT 841.950 608.400 862.050 609.600 ;
        RECT 841.950 607.950 844.050 608.400 ;
        RECT 859.950 607.950 862.050 608.400 ;
        RECT 37.950 606.600 40.050 607.050 ;
        RECT 43.950 606.600 46.050 607.200 ;
        RECT 37.950 605.400 46.050 606.600 ;
        RECT 37.950 604.950 40.050 605.400 ;
        RECT 43.950 605.100 46.050 605.400 ;
        RECT 64.950 606.600 67.050 607.050 ;
        RECT 73.950 606.600 76.050 607.200 ;
        RECT 64.950 605.400 76.050 606.600 ;
        RECT 64.950 604.950 67.050 605.400 ;
        RECT 73.950 605.100 76.050 605.400 ;
        RECT 97.950 606.750 100.050 607.200 ;
        RECT 103.950 606.750 106.050 607.200 ;
        RECT 97.950 605.550 106.050 606.750 ;
        RECT 97.950 605.100 100.050 605.550 ;
        RECT 103.950 605.100 106.050 605.550 ;
        RECT 118.950 605.100 121.050 607.200 ;
        RECT 130.950 606.600 133.050 607.050 ;
        RECT 142.950 606.600 145.050 607.200 ;
        RECT 160.950 606.600 163.050 607.200 ;
        RECT 130.950 605.400 141.600 606.600 ;
        RECT 109.950 603.600 112.050 604.050 ;
        RECT 119.400 603.600 120.600 605.100 ;
        RECT 130.950 604.950 133.050 605.400 ;
        RECT 109.950 602.400 120.600 603.600 ;
        RECT 109.950 601.950 112.050 602.400 ;
        RECT 140.400 600.900 141.600 605.400 ;
        RECT 142.950 605.400 163.050 606.600 ;
        RECT 142.950 605.100 145.050 605.400 ;
        RECT 160.950 605.100 163.050 605.400 ;
        RECT 190.950 606.600 193.050 607.200 ;
        RECT 214.950 606.600 217.050 607.050 ;
        RECT 226.950 606.600 229.050 607.200 ;
        RECT 190.950 605.400 229.050 606.600 ;
        RECT 190.950 605.100 193.050 605.400 ;
        RECT 214.950 604.950 217.050 605.400 ;
        RECT 226.950 605.100 229.050 605.400 ;
        RECT 238.950 606.750 241.050 607.200 ;
        RECT 247.950 606.750 250.050 607.200 ;
        RECT 238.950 605.550 250.050 606.750 ;
        RECT 238.950 605.100 241.050 605.550 ;
        RECT 247.950 605.100 250.050 605.550 ;
        RECT 280.950 604.950 283.050 607.050 ;
        RECT 298.950 606.600 301.050 607.200 ;
        RECT 325.950 606.600 328.050 607.200 ;
        RECT 343.950 606.600 346.050 607.200 ;
        RECT 298.950 605.400 328.050 606.600 ;
        RECT 298.950 605.100 301.050 605.400 ;
        RECT 325.950 605.100 328.050 605.400 ;
        RECT 329.400 605.400 346.050 606.600 ;
        RECT 262.950 603.600 265.050 604.050 ;
        RECT 254.400 602.400 265.050 603.600 ;
        RECT 139.950 598.800 142.050 600.900 ;
        RECT 172.950 600.600 175.050 601.050 ;
        RECT 181.950 600.600 184.050 600.900 ;
        RECT 172.950 599.400 184.050 600.600 ;
        RECT 172.950 598.950 175.050 599.400 ;
        RECT 181.950 598.800 184.050 599.400 ;
        RECT 208.950 600.450 211.050 600.900 ;
        RECT 214.950 600.450 217.050 600.900 ;
        RECT 208.950 599.250 217.050 600.450 ;
        RECT 208.950 598.800 211.050 599.250 ;
        RECT 214.950 598.800 217.050 599.250 ;
        RECT 229.950 600.600 232.050 600.900 ;
        RECT 254.400 600.600 255.600 602.400 ;
        RECT 262.950 601.950 265.050 602.400 ;
        RECT 229.950 599.400 255.600 600.600 ;
        RECT 268.950 600.600 271.050 600.900 ;
        RECT 281.400 600.600 282.600 604.950 ;
        RECT 326.400 603.600 327.600 605.100 ;
        RECT 320.400 602.400 327.600 603.600 ;
        RECT 320.400 601.050 321.600 602.400 ;
        RECT 268.950 599.400 282.600 600.600 ;
        RECT 286.950 600.600 289.050 601.050 ;
        RECT 295.950 600.600 298.050 600.900 ;
        RECT 286.950 599.400 298.050 600.600 ;
        RECT 229.950 598.800 232.050 599.400 ;
        RECT 268.950 598.800 271.050 599.400 ;
        RECT 286.950 598.950 289.050 599.400 ;
        RECT 295.950 598.800 298.050 599.400 ;
        RECT 316.950 599.400 321.600 601.050 ;
        RECT 322.950 600.600 325.050 600.900 ;
        RECT 329.400 600.600 330.600 605.400 ;
        RECT 343.950 605.100 346.050 605.400 ;
        RECT 385.950 606.750 388.050 607.200 ;
        RECT 400.950 606.750 403.050 607.200 ;
        RECT 385.950 605.550 403.050 606.750 ;
        RECT 385.950 605.100 388.050 605.550 ;
        RECT 400.950 605.100 403.050 605.550 ;
        RECT 430.950 606.600 433.050 607.200 ;
        RECT 445.950 606.600 448.050 607.200 ;
        RECT 430.950 605.400 448.050 606.600 ;
        RECT 430.950 605.100 433.050 605.400 ;
        RECT 445.950 605.100 448.050 605.400 ;
        RECT 451.950 606.750 454.050 607.200 ;
        RECT 457.950 606.750 460.050 607.200 ;
        RECT 451.950 605.550 460.050 606.750 ;
        RECT 451.950 605.100 454.050 605.550 ;
        RECT 457.950 605.100 460.050 605.550 ;
        RECT 493.950 606.600 496.050 607.200 ;
        RECT 517.950 606.600 520.050 607.200 ;
        RECT 493.950 605.400 520.050 606.600 ;
        RECT 493.950 605.100 496.050 605.400 ;
        RECT 517.950 605.100 520.050 605.400 ;
        RECT 535.950 604.950 538.050 607.050 ;
        RECT 586.950 606.600 589.050 607.200 ;
        RECT 595.950 606.600 598.050 607.050 ;
        RECT 586.950 605.400 598.050 606.600 ;
        RECT 586.950 605.100 589.050 605.400 ;
        RECT 595.950 604.950 598.050 605.400 ;
        RECT 655.950 605.100 658.050 607.200 ;
        RECT 661.950 606.750 664.050 607.200 ;
        RECT 667.950 606.750 670.050 607.050 ;
        RECT 661.950 605.550 670.050 606.750 ;
        RECT 661.950 605.100 664.050 605.550 ;
        RECT 346.950 600.600 349.050 600.900 ;
        RECT 322.950 599.400 330.600 600.600 ;
        RECT 341.400 600.000 349.050 600.600 ;
        RECT 340.950 599.400 349.050 600.000 ;
        RECT 316.950 598.950 321.000 599.400 ;
        RECT 322.950 598.800 325.050 599.400 ;
        RECT 94.950 597.600 97.050 598.050 ;
        RECT 115.950 597.600 118.050 598.050 ;
        RECT 94.950 596.400 118.050 597.600 ;
        RECT 94.950 595.950 97.050 596.400 ;
        RECT 115.950 595.950 118.050 596.400 ;
        RECT 148.950 597.600 151.050 598.050 ;
        RECT 157.950 597.600 160.050 598.050 ;
        RECT 148.950 596.400 160.050 597.600 ;
        RECT 148.950 595.950 151.050 596.400 ;
        RECT 157.950 595.950 160.050 596.400 ;
        RECT 223.950 597.600 226.050 598.050 ;
        RECT 238.950 597.600 241.050 598.050 ;
        RECT 280.950 597.600 283.050 598.050 ;
        RECT 319.950 597.600 322.050 598.050 ;
        RECT 223.950 596.400 322.050 597.600 ;
        RECT 223.950 595.950 226.050 596.400 ;
        RECT 238.950 595.950 241.050 596.400 ;
        RECT 280.950 595.950 283.050 596.400 ;
        RECT 319.950 595.950 322.050 596.400 ;
        RECT 328.950 597.600 331.050 598.050 ;
        RECT 334.950 597.600 337.050 598.050 ;
        RECT 328.950 596.400 337.050 597.600 ;
        RECT 328.950 595.950 331.050 596.400 ;
        RECT 334.950 595.950 337.050 596.400 ;
        RECT 340.950 595.950 343.050 599.400 ;
        RECT 346.950 598.800 349.050 599.400 ;
        RECT 364.950 600.600 367.050 600.900 ;
        RECT 376.950 600.600 379.050 601.050 ;
        RECT 364.950 599.400 379.050 600.600 ;
        RECT 364.950 598.800 367.050 599.400 ;
        RECT 376.950 598.950 379.050 599.400 ;
        RECT 409.950 600.600 412.050 600.900 ;
        RECT 421.950 600.600 424.050 601.050 ;
        RECT 427.950 600.600 430.050 600.900 ;
        RECT 409.950 599.400 430.050 600.600 ;
        RECT 409.950 598.800 412.050 599.400 ;
        RECT 421.950 598.950 424.050 599.400 ;
        RECT 427.950 598.800 430.050 599.400 ;
        RECT 454.950 600.600 457.050 600.900 ;
        RECT 460.950 600.600 463.050 601.050 ;
        RECT 454.950 599.400 463.050 600.600 ;
        RECT 454.950 598.800 457.050 599.400 ;
        RECT 460.950 598.950 463.050 599.400 ;
        RECT 514.950 600.600 517.050 600.900 ;
        RECT 523.950 600.600 526.050 601.050 ;
        RECT 514.950 599.400 526.050 600.600 ;
        RECT 536.400 600.600 537.600 604.950 ;
        RECT 656.400 603.600 657.600 605.100 ;
        RECT 667.950 604.950 670.050 605.550 ;
        RECT 676.950 605.100 679.050 607.200 ;
        RECT 712.950 606.600 715.050 607.200 ;
        RECT 730.950 606.750 733.050 607.200 ;
        RECT 742.950 606.750 745.050 607.200 ;
        RECT 730.950 606.600 745.050 606.750 ;
        RECT 712.950 605.550 745.050 606.600 ;
        RECT 712.950 605.400 733.050 605.550 ;
        RECT 712.950 605.100 715.050 605.400 ;
        RECT 730.950 605.100 733.050 605.400 ;
        RECT 742.950 605.100 745.050 605.550 ;
        RECT 763.950 606.750 766.050 607.200 ;
        RECT 769.950 606.750 772.050 607.200 ;
        RECT 763.950 605.550 772.050 606.750 ;
        RECT 763.950 605.100 766.050 605.550 ;
        RECT 769.950 605.100 772.050 605.550 ;
        RECT 784.950 606.750 787.050 607.200 ;
        RECT 793.950 606.750 796.050 607.200 ;
        RECT 784.950 606.600 796.050 606.750 ;
        RECT 808.950 606.600 811.050 607.200 ;
        RECT 784.950 605.550 811.050 606.600 ;
        RECT 784.950 605.100 787.050 605.550 ;
        RECT 793.950 605.400 811.050 605.550 ;
        RECT 793.950 605.100 796.050 605.400 ;
        RECT 808.950 605.100 811.050 605.400 ;
        RECT 853.950 605.100 856.050 607.200 ;
        RECT 862.950 606.600 865.050 607.050 ;
        RECT 868.950 606.600 871.050 607.050 ;
        RECT 862.950 605.400 871.050 606.600 ;
        RECT 667.950 603.600 670.050 603.900 ;
        RECT 677.400 603.600 678.600 605.100 ;
        RECT 656.400 602.400 678.600 603.600 ;
        RECT 667.950 601.800 670.050 602.400 ;
        RECT 547.800 600.600 549.900 601.050 ;
        RECT 536.400 599.400 549.900 600.600 ;
        RECT 514.950 598.800 517.050 599.400 ;
        RECT 523.950 598.950 526.050 599.400 ;
        RECT 547.800 598.950 549.900 599.400 ;
        RECT 550.950 600.450 553.050 600.900 ;
        RECT 556.950 600.450 559.050 600.900 ;
        RECT 550.950 599.250 559.050 600.450 ;
        RECT 550.950 598.800 553.050 599.250 ;
        RECT 556.950 598.800 559.050 599.250 ;
        RECT 574.950 600.450 577.050 600.900 ;
        RECT 607.950 600.450 610.050 600.900 ;
        RECT 574.950 599.250 610.050 600.450 ;
        RECT 574.950 598.800 577.050 599.250 ;
        RECT 607.950 598.800 610.050 599.250 ;
        RECT 613.950 600.600 616.050 600.900 ;
        RECT 622.950 600.600 625.050 601.050 ;
        RECT 613.950 599.400 625.050 600.600 ;
        RECT 613.950 598.800 616.050 599.400 ;
        RECT 622.950 598.950 625.050 599.400 ;
        RECT 634.950 600.600 637.050 600.900 ;
        RECT 652.950 600.600 655.050 600.900 ;
        RECT 634.950 599.400 655.050 600.600 ;
        RECT 634.950 598.800 637.050 599.400 ;
        RECT 652.950 598.800 655.050 599.400 ;
        RECT 697.950 600.600 700.050 601.050 ;
        RECT 703.950 600.600 706.050 600.900 ;
        RECT 697.950 599.400 706.050 600.600 ;
        RECT 697.950 598.950 700.050 599.400 ;
        RECT 703.950 598.800 706.050 599.400 ;
        RECT 718.950 600.600 721.050 601.050 ;
        RECT 727.950 600.600 730.050 600.900 ;
        RECT 718.950 599.400 730.050 600.600 ;
        RECT 718.950 598.950 721.050 599.400 ;
        RECT 727.950 598.800 730.050 599.400 ;
        RECT 742.950 600.600 745.050 601.050 ;
        RECT 754.950 600.600 757.050 600.900 ;
        RECT 742.950 599.400 757.050 600.600 ;
        RECT 742.950 598.950 745.050 599.400 ;
        RECT 754.950 598.800 757.050 599.400 ;
        RECT 760.950 600.450 763.050 600.900 ;
        RECT 775.950 600.450 778.050 600.900 ;
        RECT 760.950 599.250 778.050 600.450 ;
        RECT 760.950 598.800 763.050 599.250 ;
        RECT 775.950 598.800 778.050 599.250 ;
        RECT 823.950 600.450 826.050 600.900 ;
        RECT 829.950 600.450 832.050 600.900 ;
        RECT 823.950 599.250 832.050 600.450 ;
        RECT 823.950 598.800 826.050 599.250 ;
        RECT 829.950 598.800 832.050 599.250 ;
        RECT 847.950 600.600 850.050 601.050 ;
        RECT 854.400 600.600 855.600 605.100 ;
        RECT 862.950 604.950 865.050 605.400 ;
        RECT 868.950 604.950 871.050 605.400 ;
        RECT 877.950 605.100 880.050 607.200 ;
        RECT 883.950 606.600 886.050 607.200 ;
        RECT 892.950 606.600 895.050 607.050 ;
        RECT 883.950 605.400 895.050 606.600 ;
        RECT 883.950 605.100 886.050 605.400 ;
        RECT 847.950 599.400 855.600 600.600 ;
        RECT 847.950 598.950 850.050 599.400 ;
        RECT 878.400 598.050 879.600 605.100 ;
        RECT 892.950 604.950 895.050 605.400 ;
        RECT 481.950 597.600 484.050 598.050 ;
        RECT 508.950 597.600 511.050 598.050 ;
        RECT 481.950 596.400 511.050 597.600 ;
        RECT 481.950 595.950 484.050 596.400 ;
        RECT 508.950 595.950 511.050 596.400 ;
        RECT 538.950 597.600 541.050 598.050 ;
        RECT 568.950 597.600 571.050 598.050 ;
        RECT 538.950 596.400 571.050 597.600 ;
        RECT 538.950 595.950 541.050 596.400 ;
        RECT 568.950 595.950 571.050 596.400 ;
        RECT 877.950 595.950 880.050 598.050 ;
        RECT 883.950 597.600 886.050 598.050 ;
        RECT 898.950 597.600 901.050 598.050 ;
        RECT 883.950 596.400 901.050 597.600 ;
        RECT 883.950 595.950 886.050 596.400 ;
        RECT 898.950 595.950 901.050 596.400 ;
        RECT 118.950 594.600 121.050 595.050 ;
        RECT 127.950 594.600 130.050 595.050 ;
        RECT 118.950 593.400 130.050 594.600 ;
        RECT 118.950 592.950 121.050 593.400 ;
        RECT 127.950 592.950 130.050 593.400 ;
        RECT 175.950 594.600 178.050 595.050 ;
        RECT 187.950 594.600 190.050 595.050 ;
        RECT 175.950 593.400 190.050 594.600 ;
        RECT 175.950 592.950 178.050 593.400 ;
        RECT 187.950 592.950 190.050 593.400 ;
        RECT 274.950 594.600 277.050 595.050 ;
        RECT 292.950 594.600 295.050 595.050 ;
        RECT 274.950 593.400 295.050 594.600 ;
        RECT 274.950 592.950 277.050 593.400 ;
        RECT 292.950 592.950 295.050 593.400 ;
        RECT 337.950 594.600 340.050 595.050 ;
        RECT 343.950 594.600 346.050 595.050 ;
        RECT 337.950 593.400 346.050 594.600 ;
        RECT 337.950 592.950 340.050 593.400 ;
        RECT 343.950 592.950 346.050 593.400 ;
        RECT 502.950 594.600 505.050 595.050 ;
        RECT 532.950 594.600 535.050 595.050 ;
        RECT 502.950 593.400 535.050 594.600 ;
        RECT 502.950 592.950 505.050 593.400 ;
        RECT 532.950 592.950 535.050 593.400 ;
        RECT 667.950 594.600 670.050 595.050 ;
        RECT 706.950 594.600 709.050 595.050 ;
        RECT 781.950 594.600 784.050 595.050 ;
        RECT 667.950 593.400 784.050 594.600 ;
        RECT 667.950 592.950 670.050 593.400 ;
        RECT 706.950 592.950 709.050 593.400 ;
        RECT 781.950 592.950 784.050 593.400 ;
        RECT 787.950 594.600 790.050 595.050 ;
        RECT 811.950 594.600 814.050 595.050 ;
        RECT 850.950 594.600 853.050 595.050 ;
        RECT 787.950 593.400 853.050 594.600 ;
        RECT 787.950 592.950 790.050 593.400 ;
        RECT 811.950 592.950 814.050 593.400 ;
        RECT 850.950 592.950 853.050 593.400 ;
        RECT 139.950 591.600 142.050 592.050 ;
        RECT 163.950 591.600 166.050 592.050 ;
        RECT 139.950 590.400 166.050 591.600 ;
        RECT 139.950 589.950 142.050 590.400 ;
        RECT 163.950 589.950 166.050 590.400 ;
        RECT 250.950 591.600 253.050 592.050 ;
        RECT 289.950 591.600 292.050 592.050 ;
        RECT 301.950 591.600 304.050 592.050 ;
        RECT 250.950 590.400 304.050 591.600 ;
        RECT 250.950 589.950 253.050 590.400 ;
        RECT 289.950 589.950 292.050 590.400 ;
        RECT 301.950 589.950 304.050 590.400 ;
        RECT 388.950 591.600 391.050 592.050 ;
        RECT 448.950 591.600 451.050 592.050 ;
        RECT 388.950 590.400 451.050 591.600 ;
        RECT 388.950 589.950 391.050 590.400 ;
        RECT 448.950 589.950 451.050 590.400 ;
        RECT 472.950 591.600 475.050 592.050 ;
        RECT 490.950 591.600 493.050 592.050 ;
        RECT 472.950 590.400 493.050 591.600 ;
        RECT 472.950 589.950 475.050 590.400 ;
        RECT 490.950 589.950 493.050 590.400 ;
        RECT 562.950 591.600 565.050 592.050 ;
        RECT 583.950 591.600 586.050 592.050 ;
        RECT 682.950 591.600 685.050 592.050 ;
        RECT 562.950 590.400 685.050 591.600 ;
        RECT 562.950 589.950 565.050 590.400 ;
        RECT 583.950 589.950 586.050 590.400 ;
        RECT 682.950 589.950 685.050 590.400 ;
        RECT 709.950 591.600 712.050 592.050 ;
        RECT 733.950 591.600 736.050 592.050 ;
        RECT 805.950 591.600 808.050 592.050 ;
        RECT 709.950 590.400 808.050 591.600 ;
        RECT 709.950 589.950 712.050 590.400 ;
        RECT 733.950 589.950 736.050 590.400 ;
        RECT 805.950 589.950 808.050 590.400 ;
        RECT 856.950 591.600 859.050 592.050 ;
        RECT 880.950 591.600 883.050 592.050 ;
        RECT 856.950 590.400 883.050 591.600 ;
        RECT 856.950 589.950 859.050 590.400 ;
        RECT 880.950 589.950 883.050 590.400 ;
        RECT 25.950 588.600 28.050 589.050 ;
        RECT 37.950 588.600 40.050 589.050 ;
        RECT 25.950 587.400 40.050 588.600 ;
        RECT 25.950 586.950 28.050 587.400 ;
        RECT 37.950 586.950 40.050 587.400 ;
        RECT 151.950 588.600 154.050 589.050 ;
        RECT 169.950 588.600 172.050 589.050 ;
        RECT 151.950 587.400 172.050 588.600 ;
        RECT 151.950 586.950 154.050 587.400 ;
        RECT 169.950 586.950 172.050 587.400 ;
        RECT 244.950 588.600 247.050 589.050 ;
        RECT 253.950 588.600 256.050 589.050 ;
        RECT 244.950 587.400 256.050 588.600 ;
        RECT 244.950 586.950 247.050 587.400 ;
        RECT 253.950 586.950 256.050 587.400 ;
        RECT 505.950 588.600 508.050 589.050 ;
        RECT 571.950 588.600 574.050 589.050 ;
        RECT 505.950 587.400 574.050 588.600 ;
        RECT 505.950 586.950 508.050 587.400 ;
        RECT 571.950 586.950 574.050 587.400 ;
        RECT 784.950 588.600 787.050 589.050 ;
        RECT 793.950 588.600 796.050 589.050 ;
        RECT 784.950 587.400 796.050 588.600 ;
        RECT 784.950 586.950 787.050 587.400 ;
        RECT 793.950 586.950 796.050 587.400 ;
        RECT 808.950 588.600 811.050 589.050 ;
        RECT 820.950 588.600 823.050 589.050 ;
        RECT 808.950 587.400 823.050 588.600 ;
        RECT 808.950 586.950 811.050 587.400 ;
        RECT 820.950 586.950 823.050 587.400 ;
        RECT 76.950 585.600 79.050 586.050 ;
        RECT 103.950 585.600 106.050 586.050 ;
        RECT 190.950 585.600 193.050 586.050 ;
        RECT 76.950 584.400 193.050 585.600 ;
        RECT 76.950 583.950 79.050 584.400 ;
        RECT 103.950 583.950 106.050 584.400 ;
        RECT 190.950 583.950 193.050 584.400 ;
        RECT 319.950 585.600 322.050 586.050 ;
        RECT 382.950 585.600 385.050 586.050 ;
        RECT 445.950 585.600 448.050 586.050 ;
        RECT 319.950 584.400 448.050 585.600 ;
        RECT 319.950 583.950 322.050 584.400 ;
        RECT 382.950 583.950 385.050 584.400 ;
        RECT 445.950 583.950 448.050 584.400 ;
        RECT 490.950 585.600 493.050 586.050 ;
        RECT 523.950 585.600 526.050 586.050 ;
        RECT 490.950 584.400 526.050 585.600 ;
        RECT 490.950 583.950 493.050 584.400 ;
        RECT 523.950 583.950 526.050 584.400 ;
        RECT 658.950 585.600 661.050 586.050 ;
        RECT 679.950 585.600 682.050 586.050 ;
        RECT 658.950 584.400 682.050 585.600 ;
        RECT 658.950 583.950 661.050 584.400 ;
        RECT 679.950 583.950 682.050 584.400 ;
        RECT 760.950 585.600 763.050 586.050 ;
        RECT 769.950 585.600 772.050 586.050 ;
        RECT 799.950 585.600 802.050 586.050 ;
        RECT 760.950 584.400 802.050 585.600 ;
        RECT 760.950 583.950 763.050 584.400 ;
        RECT 769.950 583.950 772.050 584.400 ;
        RECT 799.950 583.950 802.050 584.400 ;
        RECT 835.950 585.600 838.050 586.050 ;
        RECT 844.950 585.600 847.050 586.050 ;
        RECT 835.950 584.400 847.050 585.600 ;
        RECT 835.950 583.950 838.050 584.400 ;
        RECT 844.950 583.950 847.050 584.400 ;
        RECT 37.950 582.600 40.050 583.050 ;
        RECT 82.950 582.600 85.050 583.050 ;
        RECT 37.950 581.400 85.050 582.600 ;
        RECT 37.950 580.950 40.050 581.400 ;
        RECT 82.950 580.950 85.050 581.400 ;
        RECT 127.950 582.600 130.050 583.050 ;
        RECT 133.950 582.600 136.050 583.050 ;
        RECT 127.950 581.400 136.050 582.600 ;
        RECT 127.950 580.950 130.050 581.400 ;
        RECT 133.950 580.950 136.050 581.400 ;
        RECT 244.950 582.600 247.050 583.050 ;
        RECT 283.950 582.600 286.050 583.050 ;
        RECT 244.950 581.400 286.050 582.600 ;
        RECT 244.950 580.950 247.050 581.400 ;
        RECT 283.950 580.950 286.050 581.400 ;
        RECT 550.950 582.600 553.050 583.050 ;
        RECT 568.950 582.600 571.050 583.050 ;
        RECT 550.950 581.400 571.050 582.600 ;
        RECT 550.950 580.950 553.050 581.400 ;
        RECT 568.950 580.950 571.050 581.400 ;
        RECT 826.950 582.600 829.050 583.050 ;
        RECT 868.950 582.600 871.050 583.050 ;
        RECT 826.950 581.400 871.050 582.600 ;
        RECT 826.950 580.950 829.050 581.400 ;
        RECT 868.950 580.950 871.050 581.400 ;
        RECT 874.950 582.600 877.050 583.050 ;
        RECT 898.950 582.600 901.050 583.050 ;
        RECT 874.950 581.400 901.050 582.600 ;
        RECT 874.950 580.950 877.050 581.400 ;
        RECT 898.950 580.950 901.050 581.400 ;
        RECT 19.950 579.600 22.050 580.050 ;
        RECT 157.950 579.600 160.050 580.050 ;
        RECT 19.950 578.400 160.050 579.600 ;
        RECT 19.950 577.950 22.050 578.400 ;
        RECT 157.950 577.950 160.050 578.400 ;
        RECT 337.950 579.600 340.050 580.050 ;
        RECT 385.950 579.600 388.050 580.050 ;
        RECT 337.950 578.400 388.050 579.600 ;
        RECT 337.950 577.950 340.050 578.400 ;
        RECT 385.950 577.950 388.050 578.400 ;
        RECT 577.950 579.600 580.050 580.050 ;
        RECT 604.950 579.600 607.050 580.050 ;
        RECT 577.950 578.400 607.050 579.600 ;
        RECT 577.950 577.950 580.050 578.400 ;
        RECT 604.950 577.950 607.050 578.400 ;
        RECT 643.950 579.600 646.050 580.050 ;
        RECT 658.950 579.600 661.050 580.050 ;
        RECT 643.950 578.400 661.050 579.600 ;
        RECT 643.950 577.950 646.050 578.400 ;
        RECT 658.950 577.950 661.050 578.400 ;
        RECT 679.950 579.600 682.050 580.050 ;
        RECT 730.950 579.600 733.050 580.050 ;
        RECT 739.950 579.600 742.050 580.050 ;
        RECT 772.950 579.600 775.050 580.050 ;
        RECT 679.950 578.400 775.050 579.600 ;
        RECT 679.950 577.950 682.050 578.400 ;
        RECT 730.950 577.950 733.050 578.400 ;
        RECT 739.950 577.950 742.050 578.400 ;
        RECT 772.950 577.950 775.050 578.400 ;
        RECT 832.950 579.600 835.050 580.050 ;
        RECT 844.950 579.600 847.050 580.050 ;
        RECT 832.950 578.400 847.050 579.600 ;
        RECT 832.950 577.950 835.050 578.400 ;
        RECT 844.950 577.950 847.050 578.400 ;
        RECT 850.950 579.600 853.050 580.050 ;
        RECT 856.950 579.600 859.050 580.050 ;
        RECT 850.950 578.400 859.050 579.600 ;
        RECT 850.950 577.950 853.050 578.400 ;
        RECT 856.950 577.950 859.050 578.400 ;
        RECT 64.950 576.600 67.050 577.050 ;
        RECT 70.950 576.600 73.050 577.050 ;
        RECT 64.950 575.400 73.050 576.600 ;
        RECT 64.950 574.950 67.050 575.400 ;
        RECT 70.950 574.950 73.050 575.400 ;
        RECT 76.950 576.600 79.050 577.050 ;
        RECT 109.950 576.600 112.050 577.050 ;
        RECT 121.950 576.600 124.050 577.050 ;
        RECT 76.950 575.400 124.050 576.600 ;
        RECT 76.950 574.950 79.050 575.400 ;
        RECT 109.950 574.950 112.050 575.400 ;
        RECT 121.950 574.950 124.050 575.400 ;
        RECT 292.950 576.600 295.050 577.050 ;
        RECT 338.400 576.600 339.600 577.950 ;
        RECT 292.950 575.400 339.600 576.600 ;
        RECT 346.950 576.600 349.050 577.050 ;
        RECT 364.950 576.600 367.050 577.050 ;
        RECT 346.950 575.400 367.050 576.600 ;
        RECT 292.950 574.950 295.050 575.400 ;
        RECT 346.950 574.950 349.050 575.400 ;
        RECT 364.950 574.950 367.050 575.400 ;
        RECT 532.950 576.600 535.050 577.050 ;
        RECT 556.950 576.600 559.050 577.050 ;
        RECT 532.950 575.400 559.050 576.600 ;
        RECT 532.950 574.950 535.050 575.400 ;
        RECT 556.950 574.950 559.050 575.400 ;
        RECT 562.950 576.600 565.050 577.050 ;
        RECT 574.950 576.600 577.050 577.050 ;
        RECT 562.950 575.400 577.050 576.600 ;
        RECT 562.950 574.950 565.050 575.400 ;
        RECT 574.950 574.950 577.050 575.400 ;
        RECT 787.950 576.600 790.050 577.050 ;
        RECT 796.950 576.600 799.050 577.050 ;
        RECT 787.950 575.400 799.050 576.600 ;
        RECT 787.950 574.950 790.050 575.400 ;
        RECT 796.950 574.950 799.050 575.400 ;
        RECT 133.950 573.750 136.050 574.200 ;
        RECT 139.950 573.750 142.050 574.200 ;
        RECT 133.950 572.550 142.050 573.750 ;
        RECT 133.950 572.100 136.050 572.550 ;
        RECT 139.950 572.100 142.050 572.550 ;
        RECT 226.950 573.750 229.050 574.200 ;
        RECT 229.950 573.750 232.050 574.050 ;
        RECT 232.950 573.750 235.050 574.200 ;
        RECT 226.950 572.550 235.050 573.750 ;
        RECT 226.950 572.100 229.050 572.550 ;
        RECT 229.950 571.950 232.050 572.550 ;
        RECT 232.950 572.100 235.050 572.550 ;
        RECT 253.950 573.750 256.050 574.200 ;
        RECT 265.950 573.750 268.050 574.200 ;
        RECT 253.950 572.550 268.050 573.750 ;
        RECT 253.950 572.100 256.050 572.550 ;
        RECT 265.950 572.100 268.050 572.550 ;
        RECT 271.950 573.600 274.050 574.200 ;
        RECT 286.950 573.600 289.050 574.050 ;
        RECT 304.950 573.600 307.050 574.050 ;
        RECT 271.950 572.400 307.050 573.600 ;
        RECT 271.950 572.100 274.050 572.400 ;
        RECT 286.950 571.950 289.050 572.400 ;
        RECT 304.950 571.950 307.050 572.400 ;
        RECT 391.950 573.750 394.050 574.200 ;
        RECT 415.950 573.750 418.050 574.200 ;
        RECT 391.950 572.550 418.050 573.750 ;
        RECT 391.950 572.100 394.050 572.550 ;
        RECT 415.950 572.100 418.050 572.550 ;
        RECT 445.950 573.750 448.050 574.200 ;
        RECT 472.950 573.750 475.050 574.200 ;
        RECT 445.950 573.600 475.050 573.750 ;
        RECT 502.950 573.600 505.050 574.050 ;
        RECT 445.950 572.550 505.050 573.600 ;
        RECT 445.950 572.100 448.050 572.550 ;
        RECT 472.950 572.400 505.050 572.550 ;
        RECT 472.950 572.100 475.050 572.400 ;
        RECT 502.950 571.950 505.050 572.400 ;
        RECT 508.950 573.750 511.050 574.200 ;
        RECT 514.950 573.750 517.050 574.200 ;
        RECT 508.950 572.550 517.050 573.750 ;
        RECT 508.950 572.100 511.050 572.550 ;
        RECT 514.950 572.100 517.050 572.550 ;
        RECT 211.950 570.600 214.050 571.050 ;
        RECT 349.950 570.600 352.050 571.050 ;
        RECT 529.950 570.600 532.050 574.050 ;
        RECT 538.950 573.600 541.050 574.200 ;
        RECT 553.950 573.600 556.050 574.050 ;
        RECT 538.950 572.400 556.050 573.600 ;
        RECT 538.950 572.100 541.050 572.400 ;
        RECT 553.950 571.950 556.050 572.400 ;
        RECT 577.950 573.600 582.000 574.050 ;
        RECT 610.950 573.600 613.050 574.200 ;
        RECT 577.950 571.950 582.600 573.600 ;
        RECT 211.950 569.400 225.600 570.600 ;
        RECT 211.950 568.950 214.050 569.400 ;
        RECT 52.950 567.600 55.050 567.900 ;
        RECT 58.950 567.600 61.050 568.050 ;
        RECT 52.950 566.400 61.050 567.600 ;
        RECT 52.950 565.800 55.050 566.400 ;
        RECT 58.950 565.950 61.050 566.400 ;
        RECT 100.950 567.600 103.050 567.900 ;
        RECT 130.950 567.600 133.050 567.900 ;
        RECT 100.950 566.400 133.050 567.600 ;
        RECT 100.950 565.800 103.050 566.400 ;
        RECT 130.950 565.800 133.050 566.400 ;
        RECT 139.950 567.600 142.050 568.050 ;
        RECT 151.950 567.600 154.050 567.900 ;
        RECT 139.950 566.400 154.050 567.600 ;
        RECT 139.950 565.950 142.050 566.400 ;
        RECT 151.950 565.800 154.050 566.400 ;
        RECT 205.950 567.600 208.050 567.900 ;
        RECT 214.950 567.600 217.050 568.050 ;
        RECT 205.950 566.400 217.050 567.600 ;
        RECT 224.400 567.600 225.600 569.400 ;
        RECT 335.400 569.400 352.050 570.600 ;
        RECT 335.400 567.900 336.600 569.400 ;
        RECT 349.950 568.950 352.050 569.400 ;
        RECT 527.400 570.000 532.050 570.600 ;
        RECT 527.400 569.400 531.600 570.000 ;
        RECT 241.950 567.600 244.050 567.900 ;
        RECT 224.400 566.400 244.050 567.600 ;
        RECT 205.950 565.800 208.050 566.400 ;
        RECT 214.950 565.950 217.050 566.400 ;
        RECT 241.950 565.800 244.050 566.400 ;
        RECT 268.950 565.800 271.050 567.900 ;
        RECT 274.950 567.600 277.050 567.900 ;
        RECT 298.950 567.600 301.050 567.900 ;
        RECT 313.950 567.600 316.050 567.900 ;
        RECT 274.950 566.400 316.050 567.600 ;
        RECT 274.950 565.800 277.050 566.400 ;
        RECT 298.950 565.800 301.050 566.400 ;
        RECT 313.950 565.800 316.050 566.400 ;
        RECT 334.950 565.800 337.050 567.900 ;
        RECT 409.950 567.600 412.050 567.900 ;
        RECT 415.950 567.600 418.050 568.050 ;
        RECT 409.950 566.400 418.050 567.600 ;
        RECT 409.950 565.800 412.050 566.400 ;
        RECT 415.950 565.950 418.050 566.400 ;
        RECT 433.950 567.600 436.050 567.900 ;
        RECT 451.950 567.600 454.050 567.900 ;
        RECT 433.950 566.400 454.050 567.600 ;
        RECT 433.950 565.800 436.050 566.400 ;
        RECT 451.950 565.800 454.050 566.400 ;
        RECT 457.950 567.450 460.050 567.900 ;
        RECT 469.950 567.450 472.050 567.900 ;
        RECT 457.950 566.250 472.050 567.450 ;
        RECT 457.950 565.800 460.050 566.250 ;
        RECT 469.950 565.800 472.050 566.250 ;
        RECT 517.950 567.600 520.050 567.900 ;
        RECT 527.400 567.600 528.600 569.400 ;
        RECT 517.950 566.400 528.600 567.600 ;
        RECT 529.950 567.450 532.050 567.900 ;
        RECT 541.950 567.600 544.050 567.900 ;
        RECT 553.950 567.600 556.050 568.050 ;
        RECT 581.400 567.900 582.600 571.950 ;
        RECT 602.400 572.400 613.050 573.600 ;
        RECT 602.400 568.050 603.600 572.400 ;
        RECT 610.950 572.100 613.050 572.400 ;
        RECT 622.950 573.750 625.050 574.200 ;
        RECT 631.950 573.750 634.050 574.200 ;
        RECT 622.950 572.550 634.050 573.750 ;
        RECT 622.950 572.100 625.050 572.550 ;
        RECT 631.950 572.100 634.050 572.550 ;
        RECT 697.950 573.600 700.050 574.050 ;
        RECT 712.950 573.600 715.050 574.200 ;
        RECT 697.950 572.400 715.050 573.600 ;
        RECT 697.950 571.950 700.050 572.400 ;
        RECT 712.950 572.100 715.050 572.400 ;
        RECT 718.950 573.600 721.050 574.050 ;
        RECT 751.950 573.600 754.050 574.200 ;
        RECT 718.950 572.400 754.050 573.600 ;
        RECT 718.950 571.950 721.050 572.400 ;
        RECT 751.950 572.100 754.050 572.400 ;
        RECT 763.950 573.600 766.050 574.050 ;
        RECT 769.950 573.600 772.050 574.200 ;
        RECT 763.950 572.400 772.050 573.600 ;
        RECT 763.950 571.950 766.050 572.400 ;
        RECT 769.950 572.100 772.050 572.400 ;
        RECT 775.950 572.100 778.050 574.200 ;
        RECT 811.950 573.750 814.050 574.200 ;
        RECT 820.950 573.750 823.050 574.200 ;
        RECT 811.950 572.550 823.050 573.750 ;
        RECT 811.950 572.100 814.050 572.550 ;
        RECT 820.950 572.100 823.050 572.550 ;
        RECT 826.950 573.600 829.050 574.200 ;
        RECT 847.950 573.600 850.050 577.050 ;
        RECT 862.950 573.600 865.050 574.050 ;
        RECT 871.950 573.600 874.050 574.200 ;
        RECT 826.950 572.400 846.600 573.600 ;
        RECT 847.950 573.000 852.600 573.600 ;
        RECT 848.400 572.400 852.600 573.000 ;
        RECT 826.950 572.100 829.050 572.400 ;
        RECT 541.950 567.450 556.050 567.600 ;
        RECT 529.950 566.400 556.050 567.450 ;
        RECT 517.950 565.800 520.050 566.400 ;
        RECT 529.950 566.250 544.050 566.400 ;
        RECT 529.950 565.800 532.050 566.250 ;
        RECT 541.950 565.800 544.050 566.250 ;
        RECT 553.950 565.950 556.050 566.400 ;
        RECT 565.950 567.450 568.050 567.900 ;
        RECT 571.950 567.450 574.050 567.900 ;
        RECT 580.950 567.600 583.050 567.900 ;
        RECT 565.950 566.250 574.050 567.450 ;
        RECT 565.950 565.800 568.050 566.250 ;
        RECT 571.950 565.800 574.050 566.250 ;
        RECT 575.400 566.400 583.050 567.600 ;
        RECT 190.950 564.600 193.050 565.050 ;
        RECT 223.950 564.600 226.050 565.050 ;
        RECT 190.950 563.400 226.050 564.600 ;
        RECT 269.400 564.600 270.600 565.800 ;
        RECT 280.950 564.600 283.050 565.050 ;
        RECT 269.400 563.400 283.050 564.600 ;
        RECT 190.950 562.950 193.050 563.400 ;
        RECT 223.950 562.950 226.050 563.400 ;
        RECT 280.950 562.950 283.050 563.400 ;
        RECT 304.950 564.600 307.050 565.050 ;
        RECT 340.950 564.600 343.050 565.050 ;
        RECT 575.400 564.600 576.600 566.400 ;
        RECT 580.950 565.800 583.050 566.400 ;
        RECT 601.950 565.950 604.050 568.050 ;
        RECT 613.950 567.600 616.050 567.900 ;
        RECT 622.950 567.600 625.050 568.050 ;
        RECT 613.950 566.400 625.050 567.600 ;
        RECT 613.950 565.800 616.050 566.400 ;
        RECT 622.950 565.950 625.050 566.400 ;
        RECT 709.950 567.600 712.050 567.900 ;
        RECT 727.950 567.600 730.050 567.900 ;
        RECT 709.950 566.400 730.050 567.600 ;
        RECT 709.950 565.800 712.050 566.400 ;
        RECT 727.950 565.800 730.050 566.400 ;
        RECT 739.950 567.450 742.050 567.900 ;
        RECT 754.950 567.450 757.050 567.900 ;
        RECT 739.950 566.250 757.050 567.450 ;
        RECT 776.400 567.600 777.600 572.100 ;
        RECT 781.950 567.600 784.050 568.050 ;
        RECT 776.400 566.400 784.050 567.600 ;
        RECT 739.950 565.800 742.050 566.250 ;
        RECT 754.950 565.800 757.050 566.250 ;
        RECT 781.950 565.950 784.050 566.400 ;
        RECT 787.950 567.450 790.050 567.900 ;
        RECT 796.950 567.450 799.050 567.900 ;
        RECT 787.950 566.250 799.050 567.450 ;
        RECT 787.950 565.800 790.050 566.250 ;
        RECT 796.950 565.800 799.050 566.250 ;
        RECT 823.950 567.450 826.050 567.900 ;
        RECT 835.950 567.450 838.050 567.900 ;
        RECT 823.950 566.250 838.050 567.450 ;
        RECT 845.400 567.600 846.600 572.400 ;
        RECT 851.400 570.600 852.600 572.400 ;
        RECT 862.950 572.400 874.050 573.600 ;
        RECT 862.950 571.950 865.050 572.400 ;
        RECT 871.950 572.100 874.050 572.400 ;
        RECT 877.950 572.100 880.050 574.200 ;
        RECT 851.400 569.400 855.600 570.600 ;
        RECT 854.400 567.900 855.600 569.400 ;
        RECT 847.950 567.600 850.050 567.900 ;
        RECT 845.400 566.400 850.050 567.600 ;
        RECT 823.950 565.800 826.050 566.250 ;
        RECT 835.950 565.800 838.050 566.250 ;
        RECT 847.950 565.800 850.050 566.400 ;
        RECT 853.950 565.800 856.050 567.900 ;
        RECT 865.950 567.600 868.050 568.050 ;
        RECT 878.400 567.600 879.600 572.100 ;
        RECT 865.950 566.400 879.600 567.600 ;
        RECT 865.950 565.950 868.050 566.400 ;
        RECT 304.950 563.400 343.050 564.600 ;
        RECT 304.950 562.950 307.050 563.400 ;
        RECT 340.950 562.950 343.050 563.400 ;
        RECT 545.400 563.400 576.600 564.600 ;
        RECT 670.950 564.600 673.050 565.050 ;
        RECT 703.950 564.600 706.050 565.050 ;
        RECT 670.950 563.400 706.050 564.600 ;
        RECT 247.950 561.600 250.050 562.050 ;
        RECT 274.950 561.600 277.050 562.050 ;
        RECT 247.950 560.400 277.050 561.600 ;
        RECT 247.950 559.950 250.050 560.400 ;
        RECT 274.950 559.950 277.050 560.400 ;
        RECT 319.950 561.600 322.050 562.050 ;
        RECT 385.950 561.600 388.050 562.050 ;
        RECT 418.950 561.600 421.050 562.050 ;
        RECT 319.950 560.400 384.600 561.600 ;
        RECT 319.950 559.950 322.050 560.400 ;
        RECT 383.400 559.050 384.600 560.400 ;
        RECT 385.950 560.400 421.050 561.600 ;
        RECT 385.950 559.950 388.050 560.400 ;
        RECT 418.950 559.950 421.050 560.400 ;
        RECT 469.950 561.600 472.050 562.050 ;
        RECT 499.950 561.600 502.050 562.050 ;
        RECT 505.950 561.600 508.050 562.050 ;
        RECT 469.950 560.400 508.050 561.600 ;
        RECT 469.950 559.950 472.050 560.400 ;
        RECT 499.950 559.950 502.050 560.400 ;
        RECT 505.950 559.950 508.050 560.400 ;
        RECT 523.950 561.600 526.050 562.050 ;
        RECT 545.400 561.600 546.600 563.400 ;
        RECT 670.950 562.950 673.050 563.400 ;
        RECT 703.950 562.950 706.050 563.400 ;
        RECT 772.950 564.600 775.050 565.050 ;
        RECT 788.400 564.600 789.600 565.800 ;
        RECT 772.950 563.400 789.600 564.600 ;
        RECT 874.950 564.600 877.050 565.050 ;
        RECT 898.950 564.600 901.050 565.050 ;
        RECT 874.950 563.400 901.050 564.600 ;
        RECT 772.950 562.950 775.050 563.400 ;
        RECT 874.950 562.950 877.050 563.400 ;
        RECT 898.950 562.950 901.050 563.400 ;
        RECT 523.950 560.400 546.600 561.600 ;
        RECT 547.950 561.600 550.050 562.050 ;
        RECT 559.950 561.600 562.050 562.050 ;
        RECT 565.950 561.600 568.050 562.050 ;
        RECT 547.950 560.400 568.050 561.600 ;
        RECT 523.950 559.950 526.050 560.400 ;
        RECT 547.950 559.950 550.050 560.400 ;
        RECT 559.950 559.950 562.050 560.400 ;
        RECT 565.950 559.950 568.050 560.400 ;
        RECT 571.950 561.600 574.050 562.050 ;
        RECT 634.950 561.600 637.050 562.050 ;
        RECT 571.950 560.400 637.050 561.600 ;
        RECT 571.950 559.950 574.050 560.400 ;
        RECT 634.950 559.950 637.050 560.400 ;
        RECT 748.950 561.600 751.050 562.050 ;
        RECT 763.950 561.600 766.050 562.050 ;
        RECT 748.950 560.400 766.050 561.600 ;
        RECT 748.950 559.950 751.050 560.400 ;
        RECT 763.950 559.950 766.050 560.400 ;
        RECT 781.950 561.600 784.050 562.050 ;
        RECT 835.950 561.600 838.050 562.050 ;
        RECT 868.950 561.600 871.050 562.050 ;
        RECT 781.950 560.400 804.600 561.600 ;
        RECT 781.950 559.950 784.050 560.400 ;
        RECT 803.400 559.050 804.600 560.400 ;
        RECT 835.950 560.400 871.050 561.600 ;
        RECT 835.950 559.950 838.050 560.400 ;
        RECT 868.950 559.950 871.050 560.400 ;
        RECT 40.950 558.600 43.050 559.050 ;
        RECT 73.950 558.600 76.050 559.050 ;
        RECT 40.950 557.400 76.050 558.600 ;
        RECT 40.950 556.950 43.050 557.400 ;
        RECT 73.950 556.950 76.050 557.400 ;
        RECT 322.950 558.600 325.050 559.050 ;
        RECT 373.950 558.600 376.050 559.050 ;
        RECT 322.950 557.400 376.050 558.600 ;
        RECT 322.950 556.950 325.050 557.400 ;
        RECT 373.950 556.950 376.050 557.400 ;
        RECT 382.950 558.600 385.050 559.050 ;
        RECT 433.950 558.600 436.050 559.050 ;
        RECT 382.950 557.400 436.050 558.600 ;
        RECT 382.950 556.950 385.050 557.400 ;
        RECT 433.950 556.950 436.050 557.400 ;
        RECT 466.950 558.600 469.050 559.050 ;
        RECT 532.950 558.600 535.050 559.050 ;
        RECT 466.950 557.400 535.050 558.600 ;
        RECT 466.950 556.950 469.050 557.400 ;
        RECT 532.950 556.950 535.050 557.400 ;
        RECT 757.950 558.600 760.050 559.050 ;
        RECT 778.950 558.600 781.050 559.050 ;
        RECT 757.950 557.400 781.050 558.600 ;
        RECT 757.950 556.950 760.050 557.400 ;
        RECT 778.950 556.950 781.050 557.400 ;
        RECT 802.950 558.600 805.050 559.050 ;
        RECT 832.950 558.600 835.050 559.050 ;
        RECT 802.950 557.400 835.050 558.600 ;
        RECT 802.950 556.950 805.050 557.400 ;
        RECT 832.950 556.950 835.050 557.400 ;
        RECT 172.950 555.600 175.050 556.050 ;
        RECT 241.950 555.600 244.050 556.050 ;
        RECT 490.950 555.600 493.050 556.050 ;
        RECT 508.950 555.600 511.050 556.050 ;
        RECT 541.950 555.600 544.050 556.050 ;
        RECT 172.950 554.400 544.050 555.600 ;
        RECT 172.950 553.950 175.050 554.400 ;
        RECT 241.950 553.950 244.050 554.400 ;
        RECT 490.950 553.950 493.050 554.400 ;
        RECT 508.950 553.950 511.050 554.400 ;
        RECT 541.950 553.950 544.050 554.400 ;
        RECT 553.950 555.600 556.050 556.050 ;
        RECT 628.950 555.600 631.050 556.050 ;
        RECT 553.950 554.400 631.050 555.600 ;
        RECT 553.950 553.950 556.050 554.400 ;
        RECT 628.950 553.950 631.050 554.400 ;
        RECT 838.950 555.600 841.050 556.050 ;
        RECT 892.950 555.600 895.050 556.050 ;
        RECT 838.950 554.400 895.050 555.600 ;
        RECT 838.950 553.950 841.050 554.400 ;
        RECT 892.950 553.950 895.050 554.400 ;
        RECT 355.950 552.600 358.050 553.050 ;
        RECT 388.950 552.600 391.050 553.050 ;
        RECT 355.950 551.400 391.050 552.600 ;
        RECT 355.950 550.950 358.050 551.400 ;
        RECT 388.950 550.950 391.050 551.400 ;
        RECT 421.950 552.600 424.050 553.050 ;
        RECT 481.950 552.600 484.050 553.050 ;
        RECT 421.950 551.400 484.050 552.600 ;
        RECT 421.950 550.950 424.050 551.400 ;
        RECT 481.950 550.950 484.050 551.400 ;
        RECT 733.950 552.600 736.050 553.050 ;
        RECT 853.950 552.600 856.050 553.050 ;
        RECT 733.950 551.400 856.050 552.600 ;
        RECT 733.950 550.950 736.050 551.400 ;
        RECT 853.950 550.950 856.050 551.400 ;
        RECT 865.950 552.600 868.050 553.050 ;
        RECT 874.950 552.600 877.050 553.050 ;
        RECT 865.950 551.400 877.050 552.600 ;
        RECT 865.950 550.950 868.050 551.400 ;
        RECT 874.950 550.950 877.050 551.400 ;
        RECT 88.950 549.600 91.050 550.050 ;
        RECT 109.950 549.600 112.050 550.050 ;
        RECT 184.950 549.600 187.050 550.050 ;
        RECT 199.950 549.600 202.050 550.050 ;
        RECT 88.950 548.400 202.050 549.600 ;
        RECT 88.950 547.950 91.050 548.400 ;
        RECT 109.950 547.950 112.050 548.400 ;
        RECT 184.950 547.950 187.050 548.400 ;
        RECT 199.950 547.950 202.050 548.400 ;
        RECT 403.950 549.600 406.050 550.050 ;
        RECT 517.950 549.600 520.050 550.050 ;
        RECT 403.950 548.400 520.050 549.600 ;
        RECT 403.950 547.950 406.050 548.400 ;
        RECT 517.950 547.950 520.050 548.400 ;
        RECT 388.950 546.600 391.050 547.050 ;
        RECT 466.950 546.600 469.050 547.050 ;
        RECT 388.950 545.400 469.050 546.600 ;
        RECT 388.950 544.950 391.050 545.400 ;
        RECT 466.950 544.950 469.050 545.400 ;
        RECT 640.950 546.600 643.050 547.050 ;
        RECT 718.950 546.600 721.050 547.050 ;
        RECT 640.950 545.400 721.050 546.600 ;
        RECT 640.950 544.950 643.050 545.400 ;
        RECT 718.950 544.950 721.050 545.400 ;
        RECT 760.950 546.600 763.050 547.050 ;
        RECT 862.950 546.600 865.050 547.050 ;
        RECT 760.950 545.400 865.050 546.600 ;
        RECT 760.950 544.950 763.050 545.400 ;
        RECT 862.950 544.950 865.050 545.400 ;
        RECT 232.950 543.600 235.050 544.050 ;
        RECT 259.950 543.600 262.050 544.050 ;
        RECT 232.950 542.400 262.050 543.600 ;
        RECT 232.950 541.950 235.050 542.400 ;
        RECT 259.950 541.950 262.050 542.400 ;
        RECT 310.950 543.600 313.050 544.050 ;
        RECT 385.950 543.600 388.050 544.050 ;
        RECT 310.950 542.400 388.050 543.600 ;
        RECT 310.950 541.950 313.050 542.400 ;
        RECT 385.950 541.950 388.050 542.400 ;
        RECT 430.950 543.600 433.050 544.050 ;
        RECT 445.950 543.600 448.050 544.050 ;
        RECT 430.950 542.400 448.050 543.600 ;
        RECT 430.950 541.950 433.050 542.400 ;
        RECT 445.950 541.950 448.050 542.400 ;
        RECT 454.950 543.600 457.050 544.050 ;
        RECT 514.950 543.600 517.050 544.050 ;
        RECT 454.950 542.400 517.050 543.600 ;
        RECT 454.950 541.950 457.050 542.400 ;
        RECT 514.950 541.950 517.050 542.400 ;
        RECT 793.950 543.600 796.050 544.050 ;
        RECT 832.950 543.600 835.050 544.050 ;
        RECT 838.950 543.600 841.050 544.050 ;
        RECT 793.950 542.400 841.050 543.600 ;
        RECT 793.950 541.950 796.050 542.400 ;
        RECT 832.950 541.950 835.050 542.400 ;
        RECT 838.950 541.950 841.050 542.400 ;
        RECT 226.950 540.600 229.050 541.050 ;
        RECT 301.950 540.600 304.050 541.050 ;
        RECT 226.950 539.400 304.050 540.600 ;
        RECT 226.950 538.950 229.050 539.400 ;
        RECT 301.950 538.950 304.050 539.400 ;
        RECT 445.950 540.600 448.050 540.900 ;
        RECT 517.950 540.600 520.050 541.050 ;
        RECT 445.950 539.400 520.050 540.600 ;
        RECT 445.950 538.800 448.050 539.400 ;
        RECT 517.950 538.950 520.050 539.400 ;
        RECT 544.950 540.600 547.050 541.050 ;
        RECT 601.950 540.600 604.050 541.050 ;
        RECT 544.950 539.400 604.050 540.600 ;
        RECT 544.950 538.950 547.050 539.400 ;
        RECT 601.950 538.950 604.050 539.400 ;
        RECT 628.950 540.600 631.050 541.050 ;
        RECT 655.950 540.600 658.050 541.050 ;
        RECT 628.950 539.400 658.050 540.600 ;
        RECT 628.950 538.950 631.050 539.400 ;
        RECT 655.950 538.950 658.050 539.400 ;
        RECT 880.950 540.600 883.050 541.050 ;
        RECT 889.950 540.600 892.050 541.050 ;
        RECT 880.950 539.400 892.050 540.600 ;
        RECT 880.950 538.950 883.050 539.400 ;
        RECT 889.950 538.950 892.050 539.400 ;
        RECT 121.950 537.600 124.050 538.050 ;
        RECT 133.950 537.600 136.050 538.050 ;
        RECT 160.950 537.600 163.050 538.050 ;
        RECT 121.950 536.400 163.050 537.600 ;
        RECT 121.950 535.950 124.050 536.400 ;
        RECT 133.950 535.950 136.050 536.400 ;
        RECT 160.950 535.950 163.050 536.400 ;
        RECT 520.950 537.600 523.050 538.050 ;
        RECT 538.800 537.600 540.900 538.050 ;
        RECT 520.950 536.400 540.900 537.600 ;
        RECT 520.950 535.950 523.050 536.400 ;
        RECT 538.800 535.950 540.900 536.400 ;
        RECT 541.950 537.600 544.050 538.050 ;
        RECT 577.950 537.600 580.050 538.050 ;
        RECT 541.950 536.400 580.050 537.600 ;
        RECT 541.950 535.950 544.050 536.400 ;
        RECT 577.950 535.950 580.050 536.400 ;
        RECT 616.950 537.600 619.050 538.050 ;
        RECT 697.950 537.600 700.050 538.050 ;
        RECT 616.950 536.400 700.050 537.600 ;
        RECT 616.950 535.950 619.050 536.400 ;
        RECT 697.950 535.950 700.050 536.400 ;
        RECT 112.950 534.600 115.050 535.050 ;
        RECT 86.400 533.400 115.050 534.600 ;
        RECT 79.950 531.600 82.050 532.050 ;
        RECT 86.400 531.600 87.600 533.400 ;
        RECT 112.950 532.950 115.050 533.400 ;
        RECT 457.950 534.600 460.050 535.050 ;
        RECT 487.950 534.600 490.050 535.050 ;
        RECT 502.950 534.600 505.050 535.050 ;
        RECT 457.950 533.400 505.050 534.600 ;
        RECT 457.950 532.950 460.050 533.400 ;
        RECT 487.950 532.950 490.050 533.400 ;
        RECT 502.950 532.950 505.050 533.400 ;
        RECT 517.950 534.600 520.050 535.050 ;
        RECT 544.950 534.600 547.050 535.050 ;
        RECT 517.950 533.400 547.050 534.600 ;
        RECT 517.950 532.950 520.050 533.400 ;
        RECT 544.950 532.950 547.050 533.400 ;
        RECT 715.950 534.600 718.050 535.050 ;
        RECT 778.950 534.600 781.050 535.050 ;
        RECT 715.950 533.400 781.050 534.600 ;
        RECT 715.950 532.950 718.050 533.400 ;
        RECT 778.950 532.950 781.050 533.400 ;
        RECT 841.950 534.600 844.050 535.050 ;
        RECT 856.950 534.600 859.050 535.050 ;
        RECT 886.950 534.600 889.050 535.050 ;
        RECT 841.950 533.400 889.050 534.600 ;
        RECT 841.950 532.950 844.050 533.400 ;
        RECT 856.950 532.950 859.050 533.400 ;
        RECT 886.950 532.950 889.050 533.400 ;
        RECT 79.950 530.400 87.600 531.600 ;
        RECT 121.950 531.600 124.050 532.050 ;
        RECT 178.950 531.600 181.050 532.050 ;
        RECT 121.950 530.400 181.050 531.600 ;
        RECT 79.950 529.950 82.050 530.400 ;
        RECT 121.950 529.950 124.050 530.400 ;
        RECT 178.950 529.950 181.050 530.400 ;
        RECT 364.950 531.600 367.050 532.050 ;
        RECT 394.950 531.600 397.050 532.050 ;
        RECT 364.950 530.400 397.050 531.600 ;
        RECT 364.950 529.950 367.050 530.400 ;
        RECT 394.950 529.950 397.050 530.400 ;
        RECT 661.950 531.600 664.050 531.900 ;
        RECT 667.950 531.600 670.050 532.050 ;
        RECT 661.950 530.400 670.050 531.600 ;
        RECT 661.950 529.800 664.050 530.400 ;
        RECT 667.950 529.950 670.050 530.400 ;
        RECT 697.950 531.600 700.050 532.050 ;
        RECT 703.950 531.600 706.050 532.050 ;
        RECT 745.950 531.600 748.050 532.050 ;
        RECT 697.950 530.400 748.050 531.600 ;
        RECT 697.950 529.950 700.050 530.400 ;
        RECT 703.950 529.950 706.050 530.400 ;
        RECT 745.950 529.950 748.050 530.400 ;
        RECT 784.950 529.950 787.050 532.050 ;
        RECT 862.950 531.600 865.050 532.050 ;
        RECT 877.950 531.600 880.050 532.050 ;
        RECT 862.950 530.400 880.050 531.600 ;
        RECT 862.950 529.950 865.050 530.400 ;
        RECT 877.950 529.950 880.050 530.400 ;
        RECT 43.950 528.600 46.050 529.200 ;
        RECT 52.950 528.600 55.050 529.200 ;
        RECT 88.950 528.600 91.050 529.200 ;
        RECT 43.950 527.400 51.600 528.600 ;
        RECT 43.950 527.100 46.050 527.400 ;
        RECT 50.400 525.600 51.600 527.400 ;
        RECT 52.950 527.400 91.050 528.600 ;
        RECT 52.950 527.100 55.050 527.400 ;
        RECT 88.950 527.100 91.050 527.400 ;
        RECT 139.950 528.750 142.050 529.200 ;
        RECT 145.950 528.750 148.050 529.200 ;
        RECT 139.950 528.600 148.050 528.750 ;
        RECT 154.950 528.600 157.050 529.200 ;
        RECT 139.950 527.550 157.050 528.600 ;
        RECT 139.950 527.100 142.050 527.550 ;
        RECT 145.950 527.400 157.050 527.550 ;
        RECT 145.950 527.100 148.050 527.400 ;
        RECT 154.950 527.100 157.050 527.400 ;
        RECT 259.950 528.600 262.050 529.200 ;
        RECT 268.950 528.600 271.050 529.050 ;
        RECT 259.950 527.400 271.050 528.600 ;
        RECT 259.950 527.100 262.050 527.400 ;
        RECT 268.950 526.950 271.050 527.400 ;
        RECT 277.950 528.600 280.050 529.200 ;
        RECT 295.950 528.600 298.050 529.200 ;
        RECT 322.950 528.600 325.050 529.200 ;
        RECT 277.950 527.400 325.050 528.600 ;
        RECT 277.950 527.100 280.050 527.400 ;
        RECT 295.950 527.100 298.050 527.400 ;
        RECT 322.950 527.100 325.050 527.400 ;
        RECT 334.950 528.750 337.050 529.200 ;
        RECT 343.950 528.750 346.050 529.200 ;
        RECT 334.950 527.550 346.050 528.750 ;
        RECT 334.950 527.100 337.050 527.550 ;
        RECT 343.950 527.100 346.050 527.550 ;
        RECT 349.950 528.750 352.050 529.200 ;
        RECT 355.950 528.750 358.050 529.200 ;
        RECT 349.950 527.550 358.050 528.750 ;
        RECT 349.950 527.100 352.050 527.550 ;
        RECT 355.950 527.100 358.050 527.550 ;
        RECT 364.950 527.100 367.050 529.200 ;
        RECT 370.950 528.750 373.050 529.200 ;
        RECT 379.800 528.750 381.900 529.200 ;
        RECT 370.950 527.550 381.900 528.750 ;
        RECT 370.950 527.100 373.050 527.550 ;
        RECT 379.800 527.100 381.900 527.550 ;
        RECT 382.950 528.750 385.050 529.200 ;
        RECT 388.950 528.750 391.050 529.200 ;
        RECT 382.950 527.550 391.050 528.750 ;
        RECT 382.950 527.100 385.050 527.550 ;
        RECT 388.950 527.100 391.050 527.550 ;
        RECT 406.950 528.750 409.050 529.200 ;
        RECT 415.950 528.750 418.050 529.200 ;
        RECT 406.950 528.600 418.050 528.750 ;
        RECT 439.950 528.600 442.050 529.200 ;
        RECT 406.950 527.550 442.050 528.600 ;
        RECT 406.950 527.100 409.050 527.550 ;
        RECT 415.950 527.400 442.050 527.550 ;
        RECT 415.950 527.100 418.050 527.400 ;
        RECT 439.950 527.100 442.050 527.400 ;
        RECT 50.400 524.400 63.600 525.600 ;
        RECT 62.400 522.900 63.600 524.400 ;
        RECT 365.400 523.050 366.600 527.100 ;
        RECT 448.950 526.950 451.050 529.050 ;
        RECT 463.950 528.600 466.050 529.200 ;
        RECT 455.400 527.400 466.050 528.600 ;
        RECT 19.950 522.600 22.050 522.900 ;
        RECT 25.950 522.600 28.050 522.900 ;
        RECT 19.950 521.400 28.050 522.600 ;
        RECT 19.950 520.800 22.050 521.400 ;
        RECT 25.950 520.800 28.050 521.400 ;
        RECT 61.950 520.800 64.050 522.900 ;
        RECT 115.950 522.450 118.050 522.900 ;
        RECT 121.950 522.450 124.050 522.900 ;
        RECT 115.950 521.250 124.050 522.450 ;
        RECT 115.950 520.800 118.050 521.250 ;
        RECT 121.950 520.800 124.050 521.250 ;
        RECT 136.950 522.600 139.050 522.900 ;
        RECT 157.950 522.600 160.050 522.900 ;
        RECT 136.950 521.400 160.050 522.600 ;
        RECT 136.950 520.800 139.050 521.400 ;
        RECT 157.950 520.800 160.050 521.400 ;
        RECT 163.950 522.600 166.050 522.900 ;
        RECT 181.950 522.600 184.050 522.900 ;
        RECT 163.950 521.400 184.050 522.600 ;
        RECT 163.950 520.800 166.050 521.400 ;
        RECT 181.950 520.800 184.050 521.400 ;
        RECT 268.950 522.450 271.050 522.900 ;
        RECT 274.950 522.450 277.050 522.900 ;
        RECT 268.950 521.250 277.050 522.450 ;
        RECT 268.950 520.800 271.050 521.250 ;
        RECT 274.950 520.800 277.050 521.250 ;
        RECT 304.950 522.450 307.050 522.900 ;
        RECT 310.950 522.450 313.050 522.900 ;
        RECT 304.950 521.250 313.050 522.450 ;
        RECT 304.950 520.800 307.050 521.250 ;
        RECT 310.950 520.800 313.050 521.250 ;
        RECT 361.950 521.400 366.600 523.050 ;
        RECT 379.950 522.450 382.050 522.900 ;
        RECT 391.950 522.450 394.050 522.900 ;
        RECT 361.950 520.950 366.000 521.400 ;
        RECT 379.950 521.250 394.050 522.450 ;
        RECT 379.950 520.800 382.050 521.250 ;
        RECT 391.950 520.800 394.050 521.250 ;
        RECT 397.950 522.600 400.050 522.900 ;
        RECT 406.950 522.600 409.050 523.050 ;
        RECT 397.950 521.400 409.050 522.600 ;
        RECT 397.950 520.800 400.050 521.400 ;
        RECT 406.950 520.950 409.050 521.400 ;
        RECT 412.950 522.600 415.050 522.900 ;
        RECT 436.950 522.600 439.050 522.900 ;
        RECT 412.950 521.400 439.050 522.600 ;
        RECT 412.950 520.800 415.050 521.400 ;
        RECT 436.950 520.800 439.050 521.400 ;
        RECT 442.950 522.600 445.050 522.900 ;
        RECT 449.400 522.600 450.600 526.950 ;
        RECT 455.400 526.050 456.600 527.400 ;
        RECT 463.950 527.100 466.050 527.400 ;
        RECT 469.950 528.600 472.050 529.050 ;
        RECT 478.950 528.600 481.050 529.050 ;
        RECT 511.950 528.600 514.050 529.200 ;
        RECT 469.950 527.400 481.050 528.600 ;
        RECT 469.950 526.950 472.050 527.400 ;
        RECT 478.950 526.950 481.050 527.400 ;
        RECT 500.400 527.400 514.050 528.600 ;
        RECT 451.950 524.400 456.600 526.050 ;
        RECT 451.950 523.950 456.000 524.400 ;
        RECT 500.400 523.050 501.600 527.400 ;
        RECT 511.950 527.100 514.050 527.400 ;
        RECT 538.950 528.600 541.050 529.200 ;
        RECT 553.950 528.600 556.050 529.200 ;
        RECT 538.950 527.400 556.050 528.600 ;
        RECT 538.950 527.100 541.050 527.400 ;
        RECT 553.950 527.100 556.050 527.400 ;
        RECT 565.950 526.950 568.050 529.050 ;
        RECT 571.950 528.750 574.050 529.200 ;
        RECT 598.950 528.750 601.050 529.200 ;
        RECT 571.950 527.550 601.050 528.750 ;
        RECT 571.950 527.100 574.050 527.550 ;
        RECT 598.950 527.100 601.050 527.550 ;
        RECT 604.950 527.100 607.050 529.200 ;
        RECT 613.950 528.750 616.050 529.200 ;
        RECT 622.950 528.750 625.050 529.200 ;
        RECT 613.950 527.550 625.050 528.750 ;
        RECT 613.950 527.100 616.050 527.550 ;
        RECT 622.950 527.100 625.050 527.550 ;
        RECT 643.950 528.750 646.050 529.200 ;
        RECT 652.950 528.750 655.050 529.200 ;
        RECT 643.950 527.550 655.050 528.750 ;
        RECT 673.950 528.600 676.050 529.200 ;
        RECT 688.950 528.600 691.050 529.200 ;
        RECT 643.950 527.100 646.050 527.550 ;
        RECT 652.950 527.100 655.050 527.550 ;
        RECT 668.400 527.400 691.050 528.600 ;
        RECT 442.950 521.400 450.600 522.600 ;
        RECT 472.950 522.600 475.050 522.900 ;
        RECT 490.950 522.600 493.050 522.900 ;
        RECT 472.950 521.400 493.050 522.600 ;
        RECT 442.950 520.800 445.050 521.400 ;
        RECT 472.950 520.800 475.050 521.400 ;
        RECT 490.950 520.800 493.050 521.400 ;
        RECT 499.950 520.950 502.050 523.050 ;
        RECT 520.950 522.600 523.050 522.900 ;
        RECT 550.950 522.600 553.050 523.050 ;
        RECT 520.950 521.400 553.050 522.600 ;
        RECT 520.950 520.800 523.050 521.400 ;
        RECT 550.950 520.950 553.050 521.400 ;
        RECT 220.950 519.600 223.050 520.050 ;
        RECT 298.950 519.600 301.050 520.050 ;
        RECT 334.950 519.600 337.050 520.050 ;
        RECT 349.950 519.600 352.050 520.050 ;
        RECT 220.950 518.400 352.050 519.600 ;
        RECT 220.950 517.950 223.050 518.400 ;
        RECT 298.950 517.950 301.050 518.400 ;
        RECT 334.950 517.950 337.050 518.400 ;
        RECT 349.950 517.950 352.050 518.400 ;
        RECT 427.950 519.600 430.050 520.050 ;
        RECT 457.950 519.600 460.050 520.050 ;
        RECT 427.950 518.400 460.050 519.600 ;
        RECT 427.950 517.950 430.050 518.400 ;
        RECT 457.950 517.950 460.050 518.400 ;
        RECT 502.950 519.600 505.050 520.050 ;
        RECT 532.950 519.600 535.050 520.050 ;
        RECT 541.950 519.600 544.050 520.050 ;
        RECT 502.950 518.400 531.600 519.600 ;
        RECT 502.950 517.950 505.050 518.400 ;
        RECT 109.950 516.600 112.050 517.050 ;
        RECT 130.950 516.600 133.050 517.050 ;
        RECT 109.950 515.400 133.050 516.600 ;
        RECT 109.950 514.950 112.050 515.400 ;
        RECT 130.950 514.950 133.050 515.400 ;
        RECT 346.950 516.600 349.050 517.050 ;
        RECT 367.950 516.600 370.050 517.050 ;
        RECT 382.950 516.600 385.050 517.050 ;
        RECT 346.950 515.400 385.050 516.600 ;
        RECT 346.950 514.950 349.050 515.400 ;
        RECT 367.950 514.950 370.050 515.400 ;
        RECT 382.950 514.950 385.050 515.400 ;
        RECT 418.950 516.600 421.050 517.050 ;
        RECT 454.950 516.600 457.050 517.050 ;
        RECT 418.950 515.400 457.050 516.600 ;
        RECT 530.400 516.600 531.600 518.400 ;
        RECT 532.950 518.400 544.050 519.600 ;
        RECT 532.950 517.950 535.050 518.400 ;
        RECT 541.950 517.950 544.050 518.400 ;
        RECT 553.950 519.600 556.050 520.050 ;
        RECT 566.400 519.600 567.600 526.950 ;
        RECT 568.950 525.600 571.050 526.050 ;
        RECT 605.400 525.600 606.600 527.100 ;
        RECT 668.400 525.600 669.600 527.400 ;
        RECT 673.950 527.100 676.050 527.400 ;
        RECT 688.950 527.100 691.050 527.400 ;
        RECT 721.950 528.750 724.050 529.200 ;
        RECT 727.950 528.750 730.050 529.200 ;
        RECT 721.950 528.600 730.050 528.750 ;
        RECT 739.950 528.600 742.050 529.200 ;
        RECT 721.950 527.550 742.050 528.600 ;
        RECT 721.950 527.100 724.050 527.550 ;
        RECT 727.950 527.400 742.050 527.550 ;
        RECT 727.950 527.100 730.050 527.400 ;
        RECT 739.950 527.100 742.050 527.400 ;
        RECT 745.950 528.600 748.050 529.200 ;
        RECT 772.950 528.600 775.050 529.200 ;
        RECT 745.950 527.400 775.050 528.600 ;
        RECT 745.950 527.100 748.050 527.400 ;
        RECT 772.950 527.100 775.050 527.400 ;
        RECT 785.400 525.600 786.600 529.950 ;
        RECT 799.950 528.750 802.050 529.200 ;
        RECT 805.950 528.750 808.050 529.200 ;
        RECT 799.950 528.600 808.050 528.750 ;
        RECT 817.950 528.600 820.050 529.200 ;
        RECT 799.950 527.550 820.050 528.600 ;
        RECT 799.950 527.100 802.050 527.550 ;
        RECT 805.950 527.400 820.050 527.550 ;
        RECT 805.950 527.100 808.050 527.400 ;
        RECT 817.950 527.100 820.050 527.400 ;
        RECT 823.950 527.100 826.050 529.200 ;
        RECT 829.950 528.750 832.050 529.200 ;
        RECT 841.950 528.750 844.050 529.200 ;
        RECT 829.950 527.550 844.050 528.750 ;
        RECT 829.950 527.100 832.050 527.550 ;
        RECT 841.950 527.100 844.050 527.550 ;
        RECT 568.950 524.400 669.600 525.600 ;
        RECT 782.400 524.400 786.600 525.600 ;
        RECT 568.950 523.950 571.050 524.400 ;
        RECT 782.400 523.050 783.600 524.400 ;
        RECT 580.950 522.600 583.050 522.900 ;
        RECT 631.950 522.600 634.050 522.900 ;
        RECT 580.950 521.400 634.050 522.600 ;
        RECT 580.950 520.800 583.050 521.400 ;
        RECT 631.950 520.800 634.050 521.400 ;
        RECT 670.950 522.600 673.050 522.900 ;
        RECT 712.950 522.600 715.050 522.900 ;
        RECT 733.950 522.600 736.050 523.050 ;
        RECT 670.950 521.400 736.050 522.600 ;
        RECT 670.950 520.800 673.050 521.400 ;
        RECT 712.950 520.800 715.050 521.400 ;
        RECT 733.950 520.950 736.050 521.400 ;
        RECT 748.950 522.600 751.050 522.900 ;
        RECT 757.800 522.600 759.900 523.050 ;
        RECT 748.950 521.400 759.900 522.600 ;
        RECT 748.950 520.800 751.050 521.400 ;
        RECT 757.800 520.950 759.900 521.400 ;
        RECT 760.950 522.450 763.050 522.900 ;
        RECT 769.950 522.450 772.050 522.900 ;
        RECT 760.950 521.250 772.050 522.450 ;
        RECT 760.950 520.800 763.050 521.250 ;
        RECT 769.950 520.800 772.050 521.250 ;
        RECT 778.950 521.400 783.600 523.050 ;
        RECT 784.950 522.600 787.050 523.050 ;
        RECT 790.950 522.600 793.050 522.900 ;
        RECT 784.950 521.400 793.050 522.600 ;
        RECT 778.950 520.950 783.000 521.400 ;
        RECT 784.950 520.950 787.050 521.400 ;
        RECT 790.950 520.800 793.050 521.400 ;
        RECT 796.950 522.600 799.050 522.900 ;
        RECT 824.400 522.600 825.600 527.100 ;
        RECT 859.950 526.950 862.050 529.050 ;
        RECT 860.400 523.050 861.600 526.950 ;
        RECT 874.950 525.600 877.050 529.050 ;
        RECT 892.950 527.100 895.050 529.200 ;
        RECT 872.400 525.000 877.050 525.600 ;
        RECT 872.400 524.400 876.600 525.000 ;
        RECT 838.950 522.600 841.050 522.900 ;
        RECT 796.950 521.400 841.050 522.600 ;
        RECT 796.950 520.800 799.050 521.400 ;
        RECT 838.950 520.800 841.050 521.400 ;
        RECT 859.950 520.950 862.050 523.050 ;
        RECT 872.400 522.900 873.600 524.400 ;
        RECT 871.950 520.800 874.050 522.900 ;
        RECT 877.950 522.600 880.050 523.050 ;
        RECT 889.950 522.600 892.050 522.900 ;
        RECT 877.950 521.400 892.050 522.600 ;
        RECT 877.950 520.950 880.050 521.400 ;
        RECT 889.950 520.800 892.050 521.400 ;
        RECT 553.950 518.400 567.600 519.600 ;
        RECT 595.950 519.600 598.050 520.050 ;
        RECT 613.950 519.600 616.050 520.050 ;
        RECT 595.950 518.400 616.050 519.600 ;
        RECT 553.950 517.950 556.050 518.400 ;
        RECT 595.950 517.950 598.050 518.400 ;
        RECT 613.950 517.950 616.050 518.400 ;
        RECT 742.950 519.600 745.050 520.050 ;
        RECT 761.400 519.600 762.600 520.800 ;
        RECT 893.400 520.050 894.600 527.100 ;
        RECT 898.950 526.950 901.050 529.050 ;
        RECT 899.400 523.050 900.600 526.950 ;
        RECT 898.950 520.950 901.050 523.050 ;
        RECT 742.950 518.400 762.600 519.600 ;
        RECT 775.950 519.600 778.050 520.050 ;
        RECT 805.950 519.600 808.050 520.050 ;
        RECT 775.950 518.400 808.050 519.600 ;
        RECT 742.950 517.950 745.050 518.400 ;
        RECT 775.950 517.950 778.050 518.400 ;
        RECT 805.950 517.950 808.050 518.400 ;
        RECT 820.950 519.600 823.050 520.050 ;
        RECT 832.950 519.600 835.050 520.050 ;
        RECT 820.950 518.400 835.050 519.600 ;
        RECT 820.950 517.950 823.050 518.400 ;
        RECT 832.950 517.950 835.050 518.400 ;
        RECT 892.950 517.950 895.050 520.050 ;
        RECT 535.950 516.600 538.050 517.050 ;
        RECT 530.400 515.400 538.050 516.600 ;
        RECT 418.950 514.950 421.050 515.400 ;
        RECT 454.950 514.950 457.050 515.400 ;
        RECT 535.950 514.950 538.050 515.400 ;
        RECT 550.950 516.600 553.050 517.050 ;
        RECT 556.950 516.600 559.050 517.050 ;
        RECT 571.950 516.600 574.050 517.050 ;
        RECT 550.950 515.400 574.050 516.600 ;
        RECT 550.950 514.950 553.050 515.400 ;
        RECT 556.950 514.950 559.050 515.400 ;
        RECT 571.950 514.950 574.050 515.400 ;
        RECT 601.950 516.600 604.050 517.050 ;
        RECT 646.950 516.600 649.050 517.050 ;
        RECT 601.950 515.400 649.050 516.600 ;
        RECT 601.950 514.950 604.050 515.400 ;
        RECT 646.950 514.950 649.050 515.400 ;
        RECT 301.950 513.600 304.050 514.050 ;
        RECT 379.950 513.600 382.050 514.050 ;
        RECT 301.950 512.400 382.050 513.600 ;
        RECT 301.950 511.950 304.050 512.400 ;
        RECT 379.950 511.950 382.050 512.400 ;
        RECT 430.950 513.600 433.050 514.050 ;
        RECT 448.950 513.600 451.050 514.050 ;
        RECT 430.950 512.400 451.050 513.600 ;
        RECT 430.950 511.950 433.050 512.400 ;
        RECT 448.950 511.950 451.050 512.400 ;
        RECT 505.950 513.600 508.050 514.050 ;
        RECT 625.950 513.600 628.050 514.050 ;
        RECT 505.950 512.400 628.050 513.600 ;
        RECT 505.950 511.950 508.050 512.400 ;
        RECT 625.950 511.950 628.050 512.400 ;
        RECT 874.950 513.600 877.050 514.050 ;
        RECT 895.950 513.600 898.050 514.050 ;
        RECT 874.950 512.400 898.050 513.600 ;
        RECT 874.950 511.950 877.050 512.400 ;
        RECT 895.950 511.950 898.050 512.400 ;
        RECT 325.950 510.600 328.050 511.050 ;
        RECT 427.950 510.600 430.050 511.050 ;
        RECT 325.950 509.400 430.050 510.600 ;
        RECT 325.950 508.950 328.050 509.400 ;
        RECT 427.950 508.950 430.050 509.400 ;
        RECT 496.950 510.600 499.050 511.050 ;
        RECT 661.950 510.600 664.050 511.050 ;
        RECT 694.950 510.600 697.050 511.050 ;
        RECT 496.950 509.400 697.050 510.600 ;
        RECT 496.950 508.950 499.050 509.400 ;
        RECT 661.950 508.950 664.050 509.400 ;
        RECT 694.950 508.950 697.050 509.400 ;
        RECT 829.950 510.600 832.050 511.050 ;
        RECT 877.950 510.600 880.050 511.050 ;
        RECT 829.950 509.400 880.050 510.600 ;
        RECT 829.950 508.950 832.050 509.400 ;
        RECT 877.950 508.950 880.050 509.400 ;
        RECT 34.950 507.600 37.050 508.050 ;
        RECT 88.950 507.600 91.050 508.050 ;
        RECT 34.950 506.400 91.050 507.600 ;
        RECT 34.950 505.950 37.050 506.400 ;
        RECT 88.950 505.950 91.050 506.400 ;
        RECT 334.950 507.600 337.050 508.050 ;
        RECT 391.950 507.600 394.050 508.050 ;
        RECT 334.950 506.400 394.050 507.600 ;
        RECT 334.950 505.950 337.050 506.400 ;
        RECT 391.950 505.950 394.050 506.400 ;
        RECT 478.950 507.600 481.050 508.050 ;
        RECT 499.950 507.600 502.050 508.050 ;
        RECT 478.950 506.400 502.050 507.600 ;
        RECT 478.950 505.950 481.050 506.400 ;
        RECT 499.950 505.950 502.050 506.400 ;
        RECT 550.950 507.600 553.050 508.050 ;
        RECT 559.950 507.600 562.050 508.050 ;
        RECT 550.950 506.400 562.050 507.600 ;
        RECT 550.950 505.950 553.050 506.400 ;
        RECT 559.950 505.950 562.050 506.400 ;
        RECT 703.950 507.600 706.050 508.050 ;
        RECT 709.950 507.600 712.050 508.050 ;
        RECT 703.950 506.400 712.050 507.600 ;
        RECT 703.950 505.950 706.050 506.400 ;
        RECT 709.950 505.950 712.050 506.400 ;
        RECT 727.950 507.600 730.050 508.050 ;
        RECT 754.950 507.600 757.050 508.050 ;
        RECT 814.950 507.600 817.050 508.050 ;
        RECT 727.950 506.400 817.050 507.600 ;
        RECT 727.950 505.950 730.050 506.400 ;
        RECT 754.950 505.950 757.050 506.400 ;
        RECT 814.950 505.950 817.050 506.400 ;
        RECT 139.950 504.600 142.050 505.050 ;
        RECT 145.950 504.600 148.050 505.050 ;
        RECT 139.950 503.400 148.050 504.600 ;
        RECT 139.950 502.950 142.050 503.400 ;
        RECT 145.950 502.950 148.050 503.400 ;
        RECT 202.950 504.600 205.050 505.050 ;
        RECT 268.950 504.600 271.050 505.050 ;
        RECT 280.950 504.600 283.050 505.050 ;
        RECT 202.950 503.400 283.050 504.600 ;
        RECT 202.950 502.950 205.050 503.400 ;
        RECT 268.950 502.950 271.050 503.400 ;
        RECT 280.950 502.950 283.050 503.400 ;
        RECT 361.950 504.600 364.050 505.050 ;
        RECT 409.950 504.600 412.050 505.050 ;
        RECT 433.950 504.600 436.050 505.050 ;
        RECT 361.950 503.400 412.050 504.600 ;
        RECT 361.950 502.950 364.050 503.400 ;
        RECT 409.950 502.950 412.050 503.400 ;
        RECT 419.400 503.400 436.050 504.600 ;
        RECT 355.950 501.600 358.050 502.050 ;
        RECT 367.950 501.600 370.050 502.050 ;
        RECT 355.950 500.400 370.050 501.600 ;
        RECT 355.950 499.950 358.050 500.400 ;
        RECT 367.950 499.950 370.050 500.400 ;
        RECT 373.950 501.600 376.050 502.050 ;
        RECT 419.400 501.600 420.600 503.400 ;
        RECT 433.950 502.950 436.050 503.400 ;
        RECT 442.950 504.600 445.050 505.050 ;
        RECT 454.950 504.600 457.050 505.050 ;
        RECT 442.950 503.400 457.050 504.600 ;
        RECT 442.950 502.950 445.050 503.400 ;
        RECT 454.950 502.950 457.050 503.400 ;
        RECT 622.950 504.600 625.050 505.050 ;
        RECT 631.950 504.600 634.050 505.050 ;
        RECT 622.950 503.400 634.050 504.600 ;
        RECT 622.950 502.950 625.050 503.400 ;
        RECT 631.950 502.950 634.050 503.400 ;
        RECT 796.950 504.600 799.050 505.050 ;
        RECT 850.950 504.600 853.050 505.050 ;
        RECT 796.950 503.400 853.050 504.600 ;
        RECT 796.950 502.950 799.050 503.400 ;
        RECT 850.950 502.950 853.050 503.400 ;
        RECT 373.950 500.400 420.600 501.600 ;
        RECT 421.950 501.600 424.050 502.050 ;
        RECT 430.950 501.600 433.050 502.050 ;
        RECT 421.950 500.400 433.050 501.600 ;
        RECT 373.950 499.950 376.050 500.400 ;
        RECT 421.950 499.950 424.050 500.400 ;
        RECT 430.950 499.950 433.050 500.400 ;
        RECT 436.950 501.600 439.050 502.050 ;
        RECT 451.950 501.600 454.050 502.050 ;
        RECT 469.950 501.600 472.050 502.050 ;
        RECT 478.800 501.600 480.900 502.050 ;
        RECT 436.950 500.400 480.900 501.600 ;
        RECT 436.950 499.950 439.050 500.400 ;
        RECT 451.950 499.950 454.050 500.400 ;
        RECT 469.950 499.950 472.050 500.400 ;
        RECT 478.800 499.950 480.900 500.400 ;
        RECT 529.950 501.600 532.050 502.050 ;
        RECT 544.950 501.600 547.050 502.050 ;
        RECT 529.950 500.400 547.050 501.600 ;
        RECT 529.950 499.950 532.050 500.400 ;
        RECT 544.950 499.950 547.050 500.400 ;
        RECT 613.950 501.600 616.050 502.050 ;
        RECT 670.950 501.600 673.050 502.050 ;
        RECT 613.950 500.400 673.050 501.600 ;
        RECT 613.950 499.950 616.050 500.400 ;
        RECT 670.950 499.950 673.050 500.400 ;
        RECT 703.950 501.600 706.050 502.050 ;
        RECT 742.950 501.600 745.050 502.050 ;
        RECT 703.950 500.400 745.050 501.600 ;
        RECT 703.950 499.950 706.050 500.400 ;
        RECT 742.950 499.950 745.050 500.400 ;
        RECT 322.950 498.600 325.050 499.050 ;
        RECT 331.950 498.600 334.050 499.050 ;
        RECT 322.950 497.400 334.050 498.600 ;
        RECT 322.950 496.950 325.050 497.400 ;
        RECT 331.950 496.950 334.050 497.400 ;
        RECT 340.950 498.600 343.050 499.050 ;
        RECT 370.950 498.600 373.050 499.050 ;
        RECT 340.950 497.400 373.050 498.600 ;
        RECT 340.950 496.950 343.050 497.400 ;
        RECT 370.950 496.950 373.050 497.400 ;
        RECT 403.950 498.600 406.050 499.050 ;
        RECT 412.950 498.600 415.050 499.050 ;
        RECT 403.950 497.400 415.050 498.600 ;
        RECT 403.950 496.950 406.050 497.400 ;
        RECT 412.950 496.950 415.050 497.400 ;
        RECT 433.950 498.600 436.050 499.050 ;
        RECT 466.950 498.600 469.050 499.050 ;
        RECT 511.950 498.600 514.050 499.050 ;
        RECT 433.950 497.400 514.050 498.600 ;
        RECT 433.950 496.950 436.050 497.400 ;
        RECT 466.950 496.950 469.050 497.400 ;
        RECT 511.950 496.950 514.050 497.400 ;
        RECT 541.950 498.600 544.050 499.050 ;
        RECT 640.950 498.600 643.050 499.050 ;
        RECT 655.950 498.600 658.050 499.050 ;
        RECT 541.950 497.400 606.600 498.600 ;
        RECT 541.950 496.950 544.050 497.400 ;
        RECT 19.950 495.600 22.050 496.200 ;
        RECT 25.950 495.600 28.050 496.200 ;
        RECT 19.950 494.400 28.050 495.600 ;
        RECT 19.950 494.100 22.050 494.400 ;
        RECT 25.950 494.100 28.050 494.400 ;
        RECT 73.950 495.600 76.050 496.200 ;
        RECT 91.950 495.600 94.050 496.050 ;
        RECT 73.950 494.400 94.050 495.600 ;
        RECT 73.950 494.100 76.050 494.400 ;
        RECT 91.950 493.950 94.050 494.400 ;
        RECT 106.950 495.600 109.050 496.200 ;
        RECT 115.950 495.600 118.050 496.050 ;
        RECT 121.950 495.600 124.050 496.200 ;
        RECT 106.950 494.400 124.050 495.600 ;
        RECT 106.950 494.100 109.050 494.400 ;
        RECT 115.950 493.950 118.050 494.400 ;
        RECT 121.950 494.100 124.050 494.400 ;
        RECT 145.950 494.100 148.050 496.200 ;
        RECT 235.950 495.600 238.050 496.200 ;
        RECT 244.950 495.600 247.050 496.050 ;
        RECT 235.950 494.400 247.050 495.600 ;
        RECT 235.950 494.100 238.050 494.400 ;
        RECT 146.400 492.600 147.600 494.100 ;
        RECT 244.950 493.950 247.050 494.400 ;
        RECT 250.950 495.600 253.050 496.050 ;
        RECT 274.950 495.600 277.050 496.200 ;
        RECT 250.950 494.400 277.050 495.600 ;
        RECT 250.950 493.950 253.050 494.400 ;
        RECT 274.950 494.100 277.050 494.400 ;
        RECT 280.950 495.600 283.050 496.200 ;
        RECT 334.950 495.600 337.050 496.050 ;
        RECT 280.950 494.400 337.050 495.600 ;
        RECT 280.950 494.100 283.050 494.400 ;
        RECT 334.950 493.950 337.050 494.400 ;
        RECT 391.950 495.600 394.050 496.200 ;
        RECT 421.950 495.600 424.050 496.050 ;
        RECT 391.950 494.400 424.050 495.600 ;
        RECT 391.950 494.100 394.050 494.400 ;
        RECT 421.950 493.950 424.050 494.400 ;
        RECT 445.950 495.600 448.050 496.050 ;
        RECT 460.950 495.600 463.050 496.200 ;
        RECT 445.950 494.400 463.050 495.600 ;
        RECT 445.950 493.950 448.050 494.400 ;
        RECT 460.950 494.100 463.050 494.400 ;
        RECT 475.950 495.750 478.050 496.200 ;
        RECT 487.950 495.750 490.050 496.200 ;
        RECT 475.950 494.550 490.050 495.750 ;
        RECT 475.950 494.100 478.050 494.550 ;
        RECT 487.950 494.100 490.050 494.550 ;
        RECT 520.950 495.600 523.050 496.050 ;
        RECT 526.950 495.600 529.050 496.050 ;
        RECT 520.950 494.400 529.050 495.600 ;
        RECT 520.950 493.950 523.050 494.400 ;
        RECT 526.950 493.950 529.050 494.400 ;
        RECT 535.950 494.100 538.050 496.200 ;
        RECT 559.950 495.600 562.050 496.200 ;
        RECT 539.400 494.400 562.050 495.600 ;
        RECT 154.950 492.600 157.050 493.050 ;
        RECT 146.400 491.400 157.050 492.600 ;
        RECT 154.950 490.950 157.050 491.400 ;
        RECT 310.950 492.600 313.050 493.050 ;
        RECT 442.950 492.600 445.050 493.050 ;
        RECT 310.950 491.400 445.050 492.600 ;
        RECT 310.950 490.950 313.050 491.400 ;
        RECT 442.950 490.950 445.050 491.400 ;
        RECT 526.950 492.600 529.050 492.900 ;
        RECT 536.400 492.600 537.600 494.100 ;
        RECT 526.950 491.400 537.600 492.600 ;
        RECT 526.950 490.800 529.050 491.400 ;
        RECT 37.950 489.600 40.050 490.050 ;
        RECT 43.950 489.600 46.050 489.900 ;
        RECT 37.950 488.400 46.050 489.600 ;
        RECT 37.950 487.950 40.050 488.400 ;
        RECT 43.950 487.800 46.050 488.400 ;
        RECT 82.950 489.450 85.050 489.900 ;
        RECT 88.950 489.600 91.050 489.900 ;
        RECT 97.950 489.600 100.050 489.900 ;
        RECT 88.950 489.450 100.050 489.600 ;
        RECT 82.950 488.400 100.050 489.450 ;
        RECT 82.950 488.250 91.050 488.400 ;
        RECT 82.950 487.800 85.050 488.250 ;
        RECT 88.950 487.800 91.050 488.250 ;
        RECT 97.950 487.800 100.050 488.400 ;
        RECT 124.950 489.600 127.050 489.900 ;
        RECT 142.950 489.600 145.050 489.900 ;
        RECT 124.950 488.400 145.050 489.600 ;
        RECT 124.950 487.800 127.050 488.400 ;
        RECT 142.950 487.800 145.050 488.400 ;
        RECT 268.950 489.600 271.050 490.050 ;
        RECT 277.950 489.600 280.050 489.900 ;
        RECT 268.950 488.400 280.050 489.600 ;
        RECT 268.950 487.950 271.050 488.400 ;
        RECT 277.950 487.800 280.050 488.400 ;
        RECT 304.950 489.600 307.050 489.900 ;
        RECT 337.950 489.600 340.050 489.900 ;
        RECT 304.950 488.400 340.050 489.600 ;
        RECT 304.950 487.800 307.050 488.400 ;
        RECT 337.950 487.800 340.050 488.400 ;
        RECT 343.950 489.450 346.050 489.900 ;
        RECT 349.950 489.450 352.050 489.900 ;
        RECT 394.950 489.600 397.050 489.900 ;
        RECT 343.950 488.250 352.050 489.450 ;
        RECT 343.950 487.800 346.050 488.250 ;
        RECT 349.950 487.800 352.050 488.250 ;
        RECT 380.400 488.400 397.050 489.600 ;
        RECT 145.950 486.600 148.050 487.050 ;
        RECT 157.950 486.600 160.050 487.050 ;
        RECT 145.950 485.400 160.050 486.600 ;
        RECT 145.950 484.950 148.050 485.400 ;
        RECT 157.950 484.950 160.050 485.400 ;
        RECT 370.950 486.600 373.050 487.050 ;
        RECT 380.400 486.600 381.600 488.400 ;
        RECT 394.950 487.800 397.050 488.400 ;
        RECT 412.950 489.600 415.050 489.900 ;
        RECT 418.800 489.600 420.900 490.050 ;
        RECT 412.950 488.400 420.900 489.600 ;
        RECT 412.950 487.800 415.050 488.400 ;
        RECT 418.800 487.950 420.900 488.400 ;
        RECT 421.950 489.450 424.050 489.900 ;
        RECT 427.950 489.450 430.050 489.900 ;
        RECT 421.950 488.250 430.050 489.450 ;
        RECT 421.950 487.800 424.050 488.250 ;
        RECT 427.950 487.800 430.050 488.250 ;
        RECT 463.950 489.450 466.050 489.900 ;
        RECT 469.950 489.450 472.050 489.900 ;
        RECT 463.950 488.250 472.050 489.450 ;
        RECT 463.950 487.800 466.050 488.250 ;
        RECT 469.950 487.800 472.050 488.250 ;
        RECT 517.950 489.600 520.050 489.900 ;
        RECT 523.950 489.600 526.050 490.050 ;
        RECT 532.950 489.600 535.050 489.900 ;
        RECT 539.400 489.600 540.600 494.400 ;
        RECT 559.950 494.100 562.050 494.400 ;
        RECT 565.950 495.600 568.050 496.200 ;
        RECT 598.950 495.600 601.050 496.050 ;
        RECT 565.950 494.400 601.050 495.600 ;
        RECT 565.950 494.100 568.050 494.400 ;
        RECT 598.950 493.950 601.050 494.400 ;
        RECT 605.400 495.600 606.600 497.400 ;
        RECT 640.950 497.400 658.050 498.600 ;
        RECT 640.950 496.950 643.050 497.400 ;
        RECT 655.950 496.950 658.050 497.400 ;
        RECT 691.950 498.600 694.050 499.050 ;
        RECT 697.950 498.600 700.050 499.050 ;
        RECT 691.950 497.400 700.050 498.600 ;
        RECT 691.950 496.950 694.050 497.400 ;
        RECT 697.950 496.950 700.050 497.400 ;
        RECT 760.950 498.600 763.050 499.050 ;
        RECT 769.950 498.600 772.050 499.050 ;
        RECT 760.950 497.400 772.050 498.600 ;
        RECT 760.950 496.950 763.050 497.400 ;
        RECT 769.950 496.950 772.050 497.400 ;
        RECT 892.950 496.950 895.050 499.050 ;
        RECT 607.950 495.600 610.050 496.200 ;
        RECT 605.400 494.400 610.050 495.600 ;
        RECT 517.950 488.400 535.050 489.600 ;
        RECT 536.400 489.000 540.600 489.600 ;
        RECT 517.950 487.800 520.050 488.400 ;
        RECT 523.950 487.950 526.050 488.400 ;
        RECT 532.950 487.800 535.050 488.400 ;
        RECT 535.950 488.400 540.600 489.000 ;
        RECT 568.950 489.450 571.050 489.900 ;
        RECT 574.950 489.450 577.050 489.900 ;
        RECT 370.950 485.400 381.600 486.600 ;
        RECT 370.950 484.950 373.050 485.400 ;
        RECT 535.950 484.950 538.050 488.400 ;
        RECT 568.950 488.250 577.050 489.450 ;
        RECT 568.950 487.800 571.050 488.250 ;
        RECT 574.950 487.800 577.050 488.250 ;
        RECT 586.950 489.600 589.050 489.900 ;
        RECT 605.400 489.600 606.600 494.400 ;
        RECT 607.950 494.100 610.050 494.400 ;
        RECT 637.950 495.600 640.050 496.200 ;
        RECT 708.000 495.600 712.050 496.050 ;
        RECT 637.950 494.400 663.600 495.600 ;
        RECT 637.950 494.100 640.050 494.400 ;
        RECT 662.400 493.050 663.600 494.400 ;
        RECT 707.400 493.950 712.050 495.600 ;
        RECT 721.950 495.750 724.050 496.200 ;
        RECT 745.950 495.750 748.050 496.200 ;
        RECT 721.950 495.600 748.050 495.750 ;
        RECT 784.800 495.600 786.900 496.050 ;
        RECT 721.950 494.550 786.900 495.600 ;
        RECT 721.950 494.100 724.050 494.550 ;
        RECT 745.950 494.400 786.900 494.550 ;
        RECT 745.950 494.100 748.050 494.400 ;
        RECT 784.800 493.950 786.900 494.400 ;
        RECT 787.950 495.600 790.050 496.050 ;
        RECT 796.950 495.600 799.050 496.200 ;
        RECT 787.950 494.400 799.050 495.600 ;
        RECT 787.950 493.950 790.050 494.400 ;
        RECT 796.950 494.100 799.050 494.400 ;
        RECT 808.950 495.750 811.050 496.200 ;
        RECT 817.950 495.750 820.050 496.200 ;
        RECT 808.950 494.550 820.050 495.750 ;
        RECT 808.950 494.100 811.050 494.550 ;
        RECT 817.950 494.100 820.050 494.550 ;
        RECT 823.950 494.100 826.050 496.200 ;
        RECT 835.950 495.750 838.050 496.200 ;
        RECT 844.950 495.750 847.050 496.200 ;
        RECT 835.950 494.550 847.050 495.750 ;
        RECT 835.950 494.100 838.050 494.550 ;
        RECT 844.950 494.100 847.050 494.550 ;
        RECT 856.950 495.750 859.050 496.200 ;
        RECT 865.950 495.750 868.050 496.200 ;
        RECT 856.950 494.550 868.050 495.750 ;
        RECT 856.950 494.100 859.050 494.550 ;
        RECT 865.950 494.100 868.050 494.550 ;
        RECT 662.400 491.400 667.050 493.050 ;
        RECT 663.000 490.950 667.050 491.400 ;
        RECT 670.950 492.600 673.050 493.050 ;
        RECT 691.950 492.600 694.050 493.050 ;
        RECT 670.950 491.400 694.050 492.600 ;
        RECT 670.950 490.950 673.050 491.400 ;
        RECT 691.950 490.950 694.050 491.400 ;
        RECT 707.400 489.900 708.600 493.950 ;
        RECT 586.950 488.400 606.600 489.600 ;
        RECT 622.950 489.450 625.050 489.900 ;
        RECT 628.950 489.450 631.050 489.900 ;
        RECT 586.950 487.800 589.050 488.400 ;
        RECT 622.950 488.250 631.050 489.450 ;
        RECT 622.950 487.800 625.050 488.250 ;
        RECT 628.950 487.800 631.050 488.250 ;
        RECT 706.950 487.800 709.050 489.900 ;
        RECT 742.950 489.600 745.050 489.900 ;
        RECT 772.950 489.600 775.050 489.900 ;
        RECT 742.950 488.400 775.050 489.600 ;
        RECT 742.950 487.800 745.050 488.400 ;
        RECT 772.950 487.800 775.050 488.400 ;
        RECT 784.950 489.450 787.050 489.900 ;
        RECT 793.950 489.600 796.050 489.900 ;
        RECT 814.950 489.600 817.050 489.900 ;
        RECT 793.950 489.450 817.050 489.600 ;
        RECT 784.950 488.400 817.050 489.450 ;
        RECT 824.400 489.600 825.600 494.100 ;
        RECT 871.950 493.950 874.050 496.050 ;
        RECT 886.950 495.600 889.050 496.200 ;
        RECT 884.400 494.400 889.050 495.600 ;
        RECT 872.400 490.050 873.600 493.950 ;
        RECT 829.950 489.600 832.050 490.050 ;
        RECT 824.400 488.400 832.050 489.600 ;
        RECT 784.950 488.250 796.050 488.400 ;
        RECT 784.950 487.800 787.050 488.250 ;
        RECT 793.950 487.800 796.050 488.250 ;
        RECT 814.950 487.800 817.050 488.400 ;
        RECT 829.950 487.950 832.050 488.400 ;
        RECT 871.950 487.950 874.050 490.050 ;
        RECT 884.400 487.050 885.600 494.400 ;
        RECT 886.950 494.100 889.050 494.400 ;
        RECT 889.950 489.450 892.050 489.900 ;
        RECT 893.400 489.450 894.600 496.950 ;
        RECT 895.950 489.450 898.050 489.900 ;
        RECT 889.950 488.250 898.050 489.450 ;
        RECT 889.950 487.800 892.050 488.250 ;
        RECT 895.950 487.800 898.050 488.250 ;
        RECT 544.950 486.600 547.050 487.050 ;
        RECT 553.950 486.600 556.050 487.050 ;
        RECT 562.950 486.600 565.050 487.050 ;
        RECT 544.950 485.400 565.050 486.600 ;
        RECT 544.950 484.950 547.050 485.400 ;
        RECT 553.950 484.950 556.050 485.400 ;
        RECT 562.950 484.950 565.050 485.400 ;
        RECT 595.950 486.600 598.050 487.050 ;
        RECT 610.950 486.600 613.050 487.050 ;
        RECT 796.950 486.600 799.050 487.050 ;
        RECT 595.950 485.400 613.050 486.600 ;
        RECT 595.950 484.950 598.050 485.400 ;
        RECT 610.950 484.950 613.050 485.400 ;
        RECT 752.400 485.400 799.050 486.600 ;
        RECT 752.400 484.050 753.600 485.400 ;
        RECT 796.950 484.950 799.050 485.400 ;
        RECT 847.950 486.600 850.050 487.050 ;
        RECT 868.950 486.600 871.050 487.050 ;
        RECT 847.950 485.400 871.050 486.600 ;
        RECT 847.950 484.950 850.050 485.400 ;
        RECT 868.950 484.950 871.050 485.400 ;
        RECT 883.950 484.950 886.050 487.050 ;
        RECT 244.950 483.600 247.050 484.050 ;
        RECT 283.950 483.600 286.050 484.050 ;
        RECT 298.950 483.600 301.050 484.050 ;
        RECT 310.950 483.600 313.050 484.050 ;
        RECT 244.950 482.400 313.050 483.600 ;
        RECT 244.950 481.950 247.050 482.400 ;
        RECT 283.950 481.950 286.050 482.400 ;
        RECT 298.950 481.950 301.050 482.400 ;
        RECT 310.950 481.950 313.050 482.400 ;
        RECT 394.950 483.600 397.050 484.050 ;
        RECT 433.950 483.600 436.050 484.050 ;
        RECT 475.950 483.600 478.050 484.050 ;
        RECT 394.950 482.400 478.050 483.600 ;
        RECT 394.950 481.950 397.050 482.400 ;
        RECT 433.950 481.950 436.050 482.400 ;
        RECT 475.950 481.950 478.050 482.400 ;
        RECT 565.950 483.600 568.050 484.050 ;
        RECT 598.950 483.600 601.050 484.050 ;
        RECT 565.950 482.400 601.050 483.600 ;
        RECT 565.950 481.950 568.050 482.400 ;
        RECT 598.950 481.950 601.050 482.400 ;
        RECT 664.950 483.600 667.050 484.050 ;
        RECT 751.950 483.600 754.050 484.050 ;
        RECT 664.950 482.400 754.050 483.600 ;
        RECT 869.400 483.600 870.600 484.950 ;
        RECT 880.950 483.600 883.050 484.050 ;
        RECT 869.400 482.400 883.050 483.600 ;
        RECT 664.950 481.950 667.050 482.400 ;
        RECT 751.950 481.950 754.050 482.400 ;
        RECT 880.950 481.950 883.050 482.400 ;
        RECT 412.950 480.600 415.050 481.050 ;
        RECT 424.950 480.600 427.050 481.050 ;
        RECT 457.950 480.600 460.050 481.050 ;
        RECT 412.950 479.400 460.050 480.600 ;
        RECT 412.950 478.950 415.050 479.400 ;
        RECT 424.950 478.950 427.050 479.400 ;
        RECT 457.950 478.950 460.050 479.400 ;
        RECT 472.950 480.600 475.050 481.050 ;
        RECT 544.950 480.600 547.050 481.050 ;
        RECT 472.950 479.400 547.050 480.600 ;
        RECT 472.950 478.950 475.050 479.400 ;
        RECT 544.950 478.950 547.050 479.400 ;
        RECT 574.950 480.600 577.050 481.050 ;
        RECT 649.950 480.600 652.050 481.050 ;
        RECT 574.950 479.400 652.050 480.600 ;
        RECT 574.950 478.950 577.050 479.400 ;
        RECT 649.950 478.950 652.050 479.400 ;
        RECT 826.950 480.600 829.050 481.050 ;
        RECT 883.950 480.600 886.050 481.050 ;
        RECT 826.950 479.400 886.050 480.600 ;
        RECT 826.950 478.950 829.050 479.400 ;
        RECT 883.950 478.950 886.050 479.400 ;
        RECT 277.950 477.600 280.050 478.050 ;
        RECT 361.950 477.600 364.050 478.050 ;
        RECT 277.950 476.400 364.050 477.600 ;
        RECT 277.950 475.950 280.050 476.400 ;
        RECT 361.950 475.950 364.050 476.400 ;
        RECT 388.950 477.600 391.050 478.050 ;
        RECT 403.950 477.600 406.050 478.050 ;
        RECT 388.950 476.400 406.050 477.600 ;
        RECT 388.950 475.950 391.050 476.400 ;
        RECT 403.950 475.950 406.050 476.400 ;
        RECT 571.950 477.600 574.050 478.050 ;
        RECT 658.950 477.600 661.050 478.050 ;
        RECT 673.950 477.600 676.050 478.050 ;
        RECT 571.950 476.400 676.050 477.600 ;
        RECT 571.950 475.950 574.050 476.400 ;
        RECT 658.950 475.950 661.050 476.400 ;
        RECT 673.950 475.950 676.050 476.400 ;
        RECT 754.950 477.600 757.050 478.050 ;
        RECT 760.950 477.600 763.050 478.050 ;
        RECT 827.400 477.600 828.600 478.950 ;
        RECT 754.950 476.400 828.600 477.600 ;
        RECT 832.950 477.600 835.050 478.050 ;
        RECT 871.950 477.600 874.050 478.050 ;
        RECT 832.950 476.400 874.050 477.600 ;
        RECT 754.950 475.950 757.050 476.400 ;
        RECT 760.950 475.950 763.050 476.400 ;
        RECT 832.950 475.950 835.050 476.400 ;
        RECT 871.950 475.950 874.050 476.400 ;
        RECT 418.950 474.600 421.050 475.050 ;
        RECT 448.950 474.600 451.050 475.050 ;
        RECT 418.950 473.400 451.050 474.600 ;
        RECT 418.950 472.950 421.050 473.400 ;
        RECT 448.950 472.950 451.050 473.400 ;
        RECT 562.950 474.600 565.050 475.050 ;
        RECT 634.950 474.600 637.050 475.050 ;
        RECT 562.950 473.400 637.050 474.600 ;
        RECT 562.950 472.950 565.050 473.400 ;
        RECT 634.950 472.950 637.050 473.400 ;
        RECT 301.950 471.600 304.050 472.050 ;
        RECT 331.950 471.600 334.050 472.050 ;
        RECT 472.950 471.600 475.050 472.050 ;
        RECT 301.950 470.400 475.050 471.600 ;
        RECT 301.950 469.950 304.050 470.400 ;
        RECT 331.950 469.950 334.050 470.400 ;
        RECT 472.950 469.950 475.050 470.400 ;
        RECT 799.950 471.600 802.050 472.050 ;
        RECT 805.950 471.600 808.050 472.050 ;
        RECT 799.950 470.400 808.050 471.600 ;
        RECT 799.950 469.950 802.050 470.400 ;
        RECT 805.950 469.950 808.050 470.400 ;
        RECT 91.950 468.600 94.050 469.050 ;
        RECT 106.950 468.600 109.050 469.050 ;
        RECT 154.950 468.600 157.050 469.050 ;
        RECT 91.950 467.400 157.050 468.600 ;
        RECT 91.950 466.950 94.050 467.400 ;
        RECT 106.950 466.950 109.050 467.400 ;
        RECT 154.950 466.950 157.050 467.400 ;
        RECT 379.950 468.600 382.050 469.050 ;
        RECT 412.950 468.600 415.050 469.050 ;
        RECT 379.950 467.400 415.050 468.600 ;
        RECT 379.950 466.950 382.050 467.400 ;
        RECT 412.950 466.950 415.050 467.400 ;
        RECT 421.950 468.600 424.050 469.050 ;
        RECT 475.950 468.600 478.050 469.050 ;
        RECT 493.950 468.600 496.050 469.050 ;
        RECT 421.950 467.400 496.050 468.600 ;
        RECT 421.950 466.950 424.050 467.400 ;
        RECT 475.950 466.950 478.050 467.400 ;
        RECT 493.950 466.950 496.050 467.400 ;
        RECT 823.950 468.600 826.050 469.050 ;
        RECT 859.950 468.600 862.050 469.050 ;
        RECT 823.950 467.400 862.050 468.600 ;
        RECT 823.950 466.950 826.050 467.400 ;
        RECT 859.950 466.950 862.050 467.400 ;
        RECT 820.950 465.600 823.050 466.050 ;
        RECT 898.950 465.600 901.050 466.050 ;
        RECT 820.950 464.400 901.050 465.600 ;
        RECT 820.950 463.950 823.050 464.400 ;
        RECT 898.950 463.950 901.050 464.400 ;
        RECT 55.950 462.600 58.050 463.050 ;
        RECT 76.950 462.600 79.050 463.050 ;
        RECT 91.950 462.600 94.050 463.050 ;
        RECT 169.950 462.600 172.050 463.050 ;
        RECT 55.950 461.400 172.050 462.600 ;
        RECT 55.950 460.950 58.050 461.400 ;
        RECT 76.950 460.950 79.050 461.400 ;
        RECT 91.950 460.950 94.050 461.400 ;
        RECT 169.950 460.950 172.050 461.400 ;
        RECT 286.950 462.600 289.050 463.050 ;
        RECT 304.950 462.600 307.050 463.050 ;
        RECT 286.950 461.400 307.050 462.600 ;
        RECT 286.950 460.950 289.050 461.400 ;
        RECT 304.950 460.950 307.050 461.400 ;
        RECT 802.950 462.600 805.050 463.050 ;
        RECT 841.950 462.600 844.050 463.050 ;
        RECT 802.950 461.400 844.050 462.600 ;
        RECT 802.950 460.950 805.050 461.400 ;
        RECT 841.950 460.950 844.050 461.400 ;
        RECT 259.950 459.600 262.050 460.050 ;
        RECT 268.950 459.600 271.050 460.050 ;
        RECT 394.950 459.600 397.050 460.050 ;
        RECT 259.950 458.400 271.050 459.600 ;
        RECT 259.950 457.950 262.050 458.400 ;
        RECT 268.950 457.950 271.050 458.400 ;
        RECT 380.400 458.400 397.050 459.600 ;
        RECT 380.400 457.050 381.600 458.400 ;
        RECT 394.950 457.950 397.050 458.400 ;
        RECT 442.950 459.600 445.050 460.050 ;
        RECT 460.950 459.600 463.050 460.050 ;
        RECT 505.950 459.600 508.050 460.050 ;
        RECT 442.950 458.400 508.050 459.600 ;
        RECT 442.950 457.950 445.050 458.400 ;
        RECT 460.950 457.950 463.050 458.400 ;
        RECT 505.950 457.950 508.050 458.400 ;
        RECT 598.950 459.600 601.050 460.050 ;
        RECT 619.950 459.600 622.050 460.050 ;
        RECT 598.950 458.400 622.050 459.600 ;
        RECT 598.950 457.950 601.050 458.400 ;
        RECT 619.950 457.950 622.050 458.400 ;
        RECT 634.950 459.600 637.050 460.050 ;
        RECT 646.950 459.600 649.050 460.050 ;
        RECT 634.950 458.400 649.050 459.600 ;
        RECT 634.950 457.950 637.050 458.400 ;
        RECT 646.950 457.950 649.050 458.400 ;
        RECT 868.950 459.600 871.050 460.050 ;
        RECT 898.950 459.600 901.050 460.050 ;
        RECT 868.950 458.400 901.050 459.600 ;
        RECT 868.950 457.950 871.050 458.400 ;
        RECT 898.950 457.950 901.050 458.400 ;
        RECT 115.950 456.600 118.050 457.050 ;
        RECT 124.950 456.600 127.050 457.050 ;
        RECT 160.950 456.600 163.050 457.050 ;
        RECT 115.950 455.400 163.050 456.600 ;
        RECT 115.950 454.950 118.050 455.400 ;
        RECT 124.950 454.950 127.050 455.400 ;
        RECT 160.950 454.950 163.050 455.400 ;
        RECT 202.950 456.600 205.050 457.050 ;
        RECT 211.950 456.600 214.050 457.050 ;
        RECT 202.950 455.400 214.050 456.600 ;
        RECT 202.950 454.950 205.050 455.400 ;
        RECT 211.950 454.950 214.050 455.400 ;
        RECT 346.950 456.600 349.050 457.050 ;
        RECT 379.950 456.600 382.050 457.050 ;
        RECT 346.950 455.400 382.050 456.600 ;
        RECT 346.950 454.950 349.050 455.400 ;
        RECT 379.950 454.950 382.050 455.400 ;
        RECT 409.950 456.600 412.050 457.050 ;
        RECT 430.950 456.600 433.050 457.050 ;
        RECT 409.950 455.400 433.050 456.600 ;
        RECT 409.950 454.950 412.050 455.400 ;
        RECT 430.950 454.950 433.050 455.400 ;
        RECT 436.950 456.600 439.050 457.050 ;
        RECT 472.950 456.600 475.050 457.050 ;
        RECT 538.950 456.600 541.050 457.050 ;
        RECT 436.950 455.400 541.050 456.600 ;
        RECT 436.950 454.950 439.050 455.400 ;
        RECT 472.950 454.950 475.050 455.400 ;
        RECT 538.950 454.950 541.050 455.400 ;
        RECT 706.950 456.600 709.050 457.050 ;
        RECT 718.950 456.600 721.050 457.050 ;
        RECT 706.950 455.400 721.050 456.600 ;
        RECT 706.950 454.950 709.050 455.400 ;
        RECT 718.950 454.950 721.050 455.400 ;
        RECT 742.950 456.600 745.050 457.050 ;
        RECT 748.950 456.600 751.050 457.050 ;
        RECT 742.950 455.400 751.050 456.600 ;
        RECT 742.950 454.950 745.050 455.400 ;
        RECT 748.950 454.950 751.050 455.400 ;
        RECT 766.950 456.600 769.050 457.050 ;
        RECT 772.950 456.600 775.050 457.050 ;
        RECT 781.950 456.600 784.050 457.050 ;
        RECT 829.950 456.600 832.050 457.050 ;
        RECT 766.950 455.400 832.050 456.600 ;
        RECT 766.950 454.950 769.050 455.400 ;
        RECT 772.950 454.950 775.050 455.400 ;
        RECT 781.950 454.950 784.050 455.400 ;
        RECT 829.950 454.950 832.050 455.400 ;
        RECT 847.950 456.600 850.050 457.050 ;
        RECT 865.950 456.600 868.050 457.050 ;
        RECT 847.950 455.400 868.050 456.600 ;
        RECT 847.950 454.950 850.050 455.400 ;
        RECT 865.950 454.950 868.050 455.400 ;
        RECT 385.950 453.600 388.050 454.050 ;
        RECT 403.950 453.600 406.050 454.050 ;
        RECT 385.950 452.400 406.050 453.600 ;
        RECT 385.950 451.950 388.050 452.400 ;
        RECT 403.950 451.950 406.050 452.400 ;
        RECT 625.950 453.600 628.050 454.050 ;
        RECT 643.800 453.600 645.900 454.050 ;
        RECT 625.950 452.400 645.900 453.600 ;
        RECT 625.950 451.950 628.050 452.400 ;
        RECT 643.800 451.950 645.900 452.400 ;
        RECT 646.950 453.600 649.050 454.050 ;
        RECT 661.950 453.600 664.050 454.050 ;
        RECT 646.950 452.400 664.050 453.600 ;
        RECT 646.950 451.950 649.050 452.400 ;
        RECT 661.950 451.950 664.050 452.400 ;
        RECT 667.950 451.950 673.050 454.050 ;
        RECT 763.950 453.600 766.050 454.050 ;
        RECT 752.400 452.400 766.050 453.600 ;
        RECT 115.950 450.600 118.050 451.200 ;
        RECT 133.950 450.600 136.050 451.200 ;
        RECT 115.950 449.400 136.050 450.600 ;
        RECT 115.950 449.100 118.050 449.400 ;
        RECT 133.950 449.100 136.050 449.400 ;
        RECT 139.950 449.100 142.050 451.200 ;
        RECT 349.950 450.750 352.050 451.200 ;
        RECT 355.950 450.750 358.050 451.200 ;
        RECT 349.950 449.550 358.050 450.750 ;
        RECT 400.950 450.600 403.050 451.050 ;
        RECT 349.950 449.100 352.050 449.550 ;
        RECT 355.950 449.100 358.050 449.550 ;
        RECT 392.400 449.400 403.050 450.600 ;
        RECT 22.950 444.600 25.050 444.900 ;
        RECT 28.950 444.600 31.050 444.900 ;
        RECT 22.950 443.400 31.050 444.600 ;
        RECT 22.950 442.800 25.050 443.400 ;
        RECT 28.950 442.800 31.050 443.400 ;
        RECT 106.950 444.450 109.050 444.900 ;
        RECT 112.950 444.450 115.050 444.900 ;
        RECT 106.950 443.250 115.050 444.450 ;
        RECT 106.950 442.800 109.050 443.250 ;
        RECT 112.950 442.800 115.050 443.250 ;
        RECT 124.950 444.450 127.050 444.900 ;
        RECT 130.950 444.450 133.050 444.900 ;
        RECT 124.950 443.250 133.050 444.450 ;
        RECT 124.950 442.800 127.050 443.250 ;
        RECT 130.950 442.800 133.050 443.250 ;
        RECT 140.400 441.600 141.600 449.100 ;
        RECT 244.950 444.450 247.050 444.900 ;
        RECT 253.950 444.450 256.050 444.900 ;
        RECT 244.950 443.250 256.050 444.450 ;
        RECT 244.950 442.800 247.050 443.250 ;
        RECT 253.950 442.800 256.050 443.250 ;
        RECT 346.950 444.600 349.050 445.050 ;
        RECT 358.950 444.600 361.050 444.900 ;
        RECT 346.950 443.400 361.050 444.600 ;
        RECT 346.950 442.950 349.050 443.400 ;
        RECT 358.950 442.800 361.050 443.400 ;
        RECT 388.950 444.600 391.050 444.900 ;
        RECT 392.400 444.600 393.600 449.400 ;
        RECT 400.950 448.950 403.050 449.400 ;
        RECT 424.950 448.950 427.050 451.050 ;
        RECT 430.950 450.600 433.050 451.200 ;
        RECT 454.950 450.600 457.050 451.200 ;
        RECT 430.950 449.400 457.050 450.600 ;
        RECT 430.950 449.100 433.050 449.400 ;
        RECT 454.950 449.100 457.050 449.400 ;
        RECT 472.950 450.600 475.050 451.050 ;
        RECT 472.950 449.400 480.600 450.600 ;
        RECT 472.950 448.950 475.050 449.400 ;
        RECT 425.400 445.050 426.600 448.950 ;
        RECT 388.950 443.400 393.600 444.600 ;
        RECT 394.950 444.450 397.050 444.900 ;
        RECT 406.950 444.450 409.050 444.900 ;
        RECT 388.950 442.800 391.050 443.400 ;
        RECT 394.950 443.250 409.050 444.450 ;
        RECT 394.950 442.800 397.050 443.250 ;
        RECT 406.950 442.800 409.050 443.250 ;
        RECT 424.800 442.950 426.900 445.050 ;
        RECT 427.950 444.600 430.050 444.900 ;
        RECT 451.950 444.600 454.050 444.900 ;
        RECT 427.950 443.400 454.050 444.600 ;
        RECT 427.950 442.800 430.050 443.400 ;
        RECT 451.950 442.800 454.050 443.400 ;
        RECT 457.950 444.600 460.050 444.900 ;
        RECT 466.950 444.600 469.050 445.050 ;
        RECT 479.400 444.900 480.600 449.400 ;
        RECT 481.950 448.950 484.050 451.050 ;
        RECT 490.950 450.750 493.050 451.050 ;
        RECT 499.950 450.750 502.050 451.200 ;
        RECT 490.950 449.550 502.050 450.750 ;
        RECT 490.950 448.950 493.050 449.550 ;
        RECT 499.950 449.100 502.050 449.550 ;
        RECT 514.950 450.600 517.050 451.050 ;
        RECT 529.950 450.600 532.050 451.050 ;
        RECT 514.950 449.400 532.050 450.600 ;
        RECT 514.950 448.950 517.050 449.400 ;
        RECT 529.950 448.950 532.050 449.400 ;
        RECT 550.950 450.600 553.050 451.200 ;
        RECT 559.950 450.750 562.050 451.200 ;
        RECT 565.950 450.750 568.050 451.200 ;
        RECT 559.950 450.600 568.050 450.750 ;
        RECT 550.950 449.550 568.050 450.600 ;
        RECT 550.950 449.400 562.050 449.550 ;
        RECT 550.950 449.100 553.050 449.400 ;
        RECT 559.950 449.100 562.050 449.400 ;
        RECT 565.950 449.100 568.050 449.550 ;
        RECT 592.950 450.600 595.050 451.050 ;
        RECT 604.950 450.600 607.050 451.050 ;
        RECT 592.950 449.400 607.050 450.600 ;
        RECT 592.950 448.950 595.050 449.400 ;
        RECT 604.950 448.950 607.050 449.400 ;
        RECT 619.950 450.750 622.050 451.200 ;
        RECT 658.950 450.750 661.050 451.200 ;
        RECT 619.950 449.550 661.050 450.750 ;
        RECT 619.950 449.100 622.050 449.550 ;
        RECT 658.950 449.100 661.050 449.550 ;
        RECT 676.950 449.100 679.050 451.200 ;
        RECT 682.950 450.600 685.050 451.050 ;
        RECT 694.950 450.600 697.050 451.200 ;
        RECT 682.950 449.400 697.050 450.600 ;
        RECT 457.950 443.400 469.050 444.600 ;
        RECT 457.950 442.800 460.050 443.400 ;
        RECT 466.950 442.950 469.050 443.400 ;
        RECT 478.950 442.800 481.050 444.900 ;
        RECT 148.950 441.600 151.050 441.900 ;
        RECT 163.950 441.600 166.050 442.050 ;
        RECT 181.950 441.600 184.050 442.050 ;
        RECT 140.400 440.400 184.050 441.600 ;
        RECT 148.950 439.800 151.050 440.400 ;
        RECT 163.950 439.950 166.050 440.400 ;
        RECT 181.950 439.950 184.050 440.400 ;
        RECT 136.950 438.600 139.050 439.050 ;
        RECT 145.950 438.600 148.050 439.050 ;
        RECT 136.950 437.400 148.050 438.600 ;
        RECT 136.950 436.950 139.050 437.400 ;
        RECT 145.950 436.950 148.050 437.400 ;
        RECT 157.950 438.600 160.050 439.050 ;
        RECT 169.950 438.600 172.050 439.050 ;
        RECT 157.950 437.400 172.050 438.600 ;
        RECT 157.950 436.950 160.050 437.400 ;
        RECT 169.950 436.950 172.050 437.400 ;
        RECT 316.950 438.600 319.050 439.050 ;
        RECT 391.950 438.600 394.050 439.050 ;
        RECT 424.950 438.600 427.050 439.050 ;
        RECT 316.950 437.400 427.050 438.600 ;
        RECT 316.950 436.950 319.050 437.400 ;
        RECT 391.950 436.950 394.050 437.400 ;
        RECT 424.950 436.950 427.050 437.400 ;
        RECT 466.950 438.600 469.050 439.050 ;
        RECT 482.400 438.600 483.600 448.950 ;
        RECT 661.950 447.600 664.050 448.050 ;
        RECT 677.400 447.600 678.600 449.100 ;
        RECT 682.950 448.950 685.050 449.400 ;
        RECT 694.950 449.100 697.050 449.400 ;
        RECT 700.950 450.600 703.050 451.200 ;
        RECT 718.950 450.600 721.050 451.200 ;
        RECT 700.950 449.400 721.050 450.600 ;
        RECT 700.950 449.100 703.050 449.400 ;
        RECT 718.950 449.100 721.050 449.400 ;
        RECT 742.950 450.600 745.050 451.200 ;
        RECT 752.400 450.600 753.600 452.400 ;
        RECT 763.950 451.950 766.050 452.400 ;
        RECT 811.950 453.600 814.050 454.050 ;
        RECT 841.950 453.600 844.050 454.050 ;
        RECT 856.950 453.600 859.050 454.050 ;
        RECT 811.950 452.400 859.050 453.600 ;
        RECT 811.950 451.950 814.050 452.400 ;
        RECT 841.950 451.950 844.050 452.400 ;
        RECT 856.950 451.950 859.050 452.400 ;
        RECT 742.950 449.400 753.600 450.600 ;
        RECT 817.950 450.600 820.050 451.200 ;
        RECT 835.950 450.600 838.050 451.200 ;
        RECT 817.950 449.400 838.050 450.600 ;
        RECT 742.950 449.100 745.050 449.400 ;
        RECT 817.950 449.100 820.050 449.400 ;
        RECT 835.950 449.100 838.050 449.400 ;
        RECT 859.950 450.600 862.050 451.200 ;
        RECT 883.950 450.600 886.050 451.200 ;
        RECT 859.950 449.400 886.050 450.600 ;
        RECT 859.950 449.100 862.050 449.400 ;
        RECT 883.950 449.100 886.050 449.400 ;
        RECT 661.950 446.400 678.600 447.600 ;
        RECT 719.400 447.600 720.600 449.100 ;
        RECT 730.950 447.600 733.050 448.050 ;
        RECT 754.950 447.600 757.050 448.050 ;
        RECT 719.400 446.400 733.050 447.600 ;
        RECT 661.950 445.950 664.050 446.400 ;
        RECT 730.950 445.950 733.050 446.400 ;
        RECT 746.400 446.400 757.050 447.600 ;
        RECT 484.950 444.600 487.050 444.900 ;
        RECT 502.950 444.600 505.050 444.900 ;
        RECT 484.950 443.400 505.050 444.600 ;
        RECT 484.950 442.800 487.050 443.400 ;
        RECT 502.950 442.800 505.050 443.400 ;
        RECT 535.950 444.450 538.050 444.900 ;
        RECT 541.950 444.450 544.050 444.900 ;
        RECT 535.950 443.250 544.050 444.450 ;
        RECT 535.950 442.800 538.050 443.250 ;
        RECT 541.950 442.800 544.050 443.250 ;
        RECT 547.950 444.600 550.050 444.900 ;
        RECT 568.950 444.600 571.050 444.900 ;
        RECT 610.950 444.600 613.050 445.050 ;
        RECT 746.400 444.900 747.600 446.400 ;
        RECT 754.950 445.950 757.050 446.400 ;
        RECT 547.950 444.000 555.600 444.600 ;
        RECT 547.950 443.400 556.050 444.000 ;
        RECT 547.950 442.800 550.050 443.400 ;
        RECT 553.950 439.950 556.050 443.400 ;
        RECT 568.950 443.400 613.050 444.600 ;
        RECT 568.950 442.800 571.050 443.400 ;
        RECT 610.950 442.950 613.050 443.400 ;
        RECT 622.950 444.450 625.050 444.900 ;
        RECT 628.950 444.450 631.050 444.900 ;
        RECT 622.950 443.250 631.050 444.450 ;
        RECT 622.950 442.800 625.050 443.250 ;
        RECT 628.950 442.800 631.050 443.250 ;
        RECT 745.950 442.800 748.050 444.900 ;
        RECT 790.950 444.600 793.050 444.900 ;
        RECT 808.950 444.600 811.050 444.900 ;
        RECT 790.950 443.400 811.050 444.600 ;
        RECT 790.950 442.800 793.050 443.400 ;
        RECT 808.950 442.800 811.050 443.400 ;
        RECT 826.950 444.600 829.050 445.050 ;
        RECT 832.950 444.600 835.050 444.900 ;
        RECT 826.950 443.400 835.050 444.600 ;
        RECT 826.950 442.950 829.050 443.400 ;
        RECT 832.950 442.800 835.050 443.400 ;
        RECT 850.950 444.600 853.050 445.050 ;
        RECT 856.950 444.600 859.050 444.900 ;
        RECT 850.950 443.400 859.050 444.600 ;
        RECT 850.950 442.950 853.050 443.400 ;
        RECT 856.950 442.800 859.050 443.400 ;
        RECT 604.950 441.600 607.050 442.050 ;
        RECT 643.950 441.600 646.050 442.050 ;
        RECT 604.950 440.400 646.050 441.600 ;
        RECT 604.950 439.950 607.050 440.400 ;
        RECT 643.950 439.950 646.050 440.400 ;
        RECT 658.950 441.600 661.050 442.050 ;
        RECT 667.950 441.600 670.050 442.050 ;
        RECT 658.950 440.400 670.050 441.600 ;
        RECT 658.950 439.950 661.050 440.400 ;
        RECT 667.950 439.950 670.050 440.400 ;
        RECT 706.950 441.600 709.050 442.050 ;
        RECT 721.950 441.600 724.050 442.050 ;
        RECT 706.950 440.400 724.050 441.600 ;
        RECT 860.400 441.600 861.600 449.100 ;
        RECT 895.950 448.950 898.050 451.050 ;
        RECT 877.950 444.450 880.050 444.900 ;
        RECT 886.950 444.450 889.050 444.900 ;
        RECT 877.950 443.250 889.050 444.450 ;
        RECT 877.950 442.800 880.050 443.250 ;
        RECT 886.950 442.800 889.050 443.250 ;
        RECT 892.950 444.600 895.050 444.900 ;
        RECT 896.400 444.600 897.600 448.950 ;
        RECT 892.950 443.400 897.600 444.600 ;
        RECT 892.950 442.800 895.050 443.400 ;
        RECT 865.950 441.600 868.050 442.050 ;
        RECT 860.400 440.400 868.050 441.600 ;
        RECT 706.950 439.950 709.050 440.400 ;
        RECT 721.950 439.950 724.050 440.400 ;
        RECT 865.950 439.950 868.050 440.400 ;
        RECT 466.950 437.400 483.600 438.600 ;
        RECT 559.950 438.600 562.050 439.050 ;
        RECT 571.950 438.600 574.050 439.050 ;
        RECT 559.950 437.400 574.050 438.600 ;
        RECT 466.950 436.950 469.050 437.400 ;
        RECT 559.950 436.950 562.050 437.400 ;
        RECT 571.950 436.950 574.050 437.400 ;
        RECT 589.950 438.600 592.050 439.050 ;
        RECT 604.950 438.600 607.050 438.900 ;
        RECT 589.950 437.400 607.050 438.600 ;
        RECT 589.950 436.950 592.050 437.400 ;
        RECT 604.950 436.800 607.050 437.400 ;
        RECT 649.950 438.600 652.050 439.050 ;
        RECT 673.950 438.600 676.050 439.050 ;
        RECT 700.950 438.600 703.050 439.050 ;
        RECT 649.950 437.400 703.050 438.600 ;
        RECT 649.950 436.950 652.050 437.400 ;
        RECT 673.950 436.950 676.050 437.400 ;
        RECT 700.950 436.950 703.050 437.400 ;
        RECT 802.950 438.600 805.050 439.050 ;
        RECT 808.950 438.600 811.050 439.050 ;
        RECT 814.950 438.600 817.050 439.050 ;
        RECT 826.950 438.600 829.050 439.050 ;
        RECT 838.950 438.600 841.050 439.050 ;
        RECT 802.950 437.400 841.050 438.600 ;
        RECT 802.950 436.950 805.050 437.400 ;
        RECT 808.950 436.950 811.050 437.400 ;
        RECT 814.950 436.950 817.050 437.400 ;
        RECT 826.950 436.950 829.050 437.400 ;
        RECT 838.950 436.950 841.050 437.400 ;
        RECT 862.950 435.600 865.050 436.050 ;
        RECT 877.950 435.600 880.050 436.050 ;
        RECT 862.950 434.400 880.050 435.600 ;
        RECT 862.950 433.950 865.050 434.400 ;
        RECT 877.950 433.950 880.050 434.400 ;
        RECT 364.950 432.600 367.050 433.050 ;
        RECT 397.950 432.600 400.050 433.050 ;
        RECT 364.950 431.400 400.050 432.600 ;
        RECT 364.950 430.950 367.050 431.400 ;
        RECT 397.950 430.950 400.050 431.400 ;
        RECT 412.950 432.600 415.050 433.050 ;
        RECT 466.950 432.600 469.050 433.050 ;
        RECT 412.950 431.400 469.050 432.600 ;
        RECT 412.950 430.950 415.050 431.400 ;
        RECT 466.950 430.950 469.050 431.400 ;
        RECT 478.950 432.600 481.050 433.050 ;
        RECT 493.950 432.600 496.050 433.050 ;
        RECT 478.950 431.400 496.050 432.600 ;
        RECT 478.950 430.950 481.050 431.400 ;
        RECT 493.950 430.950 496.050 431.400 ;
        RECT 508.950 432.600 511.050 433.050 ;
        RECT 550.950 432.600 553.050 433.050 ;
        RECT 586.950 432.600 589.050 433.050 ;
        RECT 508.950 431.400 589.050 432.600 ;
        RECT 508.950 430.950 511.050 431.400 ;
        RECT 550.950 430.950 553.050 431.400 ;
        RECT 586.950 430.950 589.050 431.400 ;
        RECT 697.950 432.600 700.050 433.050 ;
        RECT 724.950 432.600 727.050 433.050 ;
        RECT 733.950 432.600 736.050 433.050 ;
        RECT 775.950 432.600 778.050 433.050 ;
        RECT 697.950 431.400 778.050 432.600 ;
        RECT 697.950 430.950 700.050 431.400 ;
        RECT 724.950 430.950 727.050 431.400 ;
        RECT 733.950 430.950 736.050 431.400 ;
        RECT 775.950 430.950 778.050 431.400 ;
        RECT 841.950 432.600 844.050 433.050 ;
        RECT 859.950 432.600 862.050 433.050 ;
        RECT 841.950 431.400 862.050 432.600 ;
        RECT 841.950 430.950 844.050 431.400 ;
        RECT 859.950 430.950 862.050 431.400 ;
        RECT 292.950 429.600 295.050 430.050 ;
        RECT 382.950 429.600 385.050 430.050 ;
        RECT 400.950 429.600 403.050 430.050 ;
        RECT 292.950 428.400 403.050 429.600 ;
        RECT 292.950 427.950 295.050 428.400 ;
        RECT 382.950 427.950 385.050 428.400 ;
        RECT 400.950 427.950 403.050 428.400 ;
        RECT 421.950 429.600 424.050 430.050 ;
        RECT 436.950 429.600 439.050 430.050 ;
        RECT 421.950 428.400 439.050 429.600 ;
        RECT 421.950 427.950 424.050 428.400 ;
        RECT 436.950 427.950 439.050 428.400 ;
        RECT 634.950 429.600 637.050 430.050 ;
        RECT 652.950 429.600 655.050 430.050 ;
        RECT 634.950 428.400 655.050 429.600 ;
        RECT 634.950 427.950 637.050 428.400 ;
        RECT 652.950 427.950 655.050 428.400 ;
        RECT 40.950 426.600 43.050 427.050 ;
        RECT 64.950 426.600 67.050 427.050 ;
        RECT 40.950 425.400 67.050 426.600 ;
        RECT 40.950 424.950 43.050 425.400 ;
        RECT 64.950 424.950 67.050 425.400 ;
        RECT 268.950 426.600 271.050 427.050 ;
        RECT 403.950 426.600 406.050 427.050 ;
        RECT 418.950 426.600 421.050 427.050 ;
        RECT 268.950 425.400 421.050 426.600 ;
        RECT 268.950 424.950 271.050 425.400 ;
        RECT 403.950 424.950 406.050 425.400 ;
        RECT 418.950 424.950 421.050 425.400 ;
        RECT 577.950 426.600 580.050 427.050 ;
        RECT 646.950 426.600 649.050 427.050 ;
        RECT 577.950 425.400 649.050 426.600 ;
        RECT 577.950 424.950 580.050 425.400 ;
        RECT 646.950 424.950 649.050 425.400 ;
        RECT 820.950 426.600 823.050 427.050 ;
        RECT 847.950 426.600 850.050 427.050 ;
        RECT 820.950 425.400 850.050 426.600 ;
        RECT 820.950 424.950 823.050 425.400 ;
        RECT 847.950 424.950 850.050 425.400 ;
        RECT 859.950 426.600 862.050 427.050 ;
        RECT 874.950 426.600 877.050 427.050 ;
        RECT 859.950 425.400 877.050 426.600 ;
        RECT 859.950 424.950 862.050 425.400 ;
        RECT 874.950 424.950 877.050 425.400 ;
        RECT 265.950 423.600 268.050 424.050 ;
        RECT 277.950 423.600 280.050 424.050 ;
        RECT 265.950 422.400 280.050 423.600 ;
        RECT 265.950 421.950 268.050 422.400 ;
        RECT 277.950 421.950 280.050 422.400 ;
        RECT 337.950 423.600 340.050 424.050 ;
        RECT 370.950 423.600 373.050 424.050 ;
        RECT 382.950 423.600 385.050 424.050 ;
        RECT 337.950 422.400 385.050 423.600 ;
        RECT 337.950 421.950 340.050 422.400 ;
        RECT 370.950 421.950 373.050 422.400 ;
        RECT 382.950 421.950 385.050 422.400 ;
        RECT 457.950 423.600 460.050 424.050 ;
        RECT 484.950 423.600 487.050 424.050 ;
        RECT 490.950 423.600 493.050 424.050 ;
        RECT 457.950 422.400 493.050 423.600 ;
        RECT 457.950 421.950 460.050 422.400 ;
        RECT 484.950 421.950 487.050 422.400 ;
        RECT 490.950 421.950 493.050 422.400 ;
        RECT 679.950 423.600 682.050 424.050 ;
        RECT 694.950 423.600 697.050 424.050 ;
        RECT 742.950 423.600 745.050 424.050 ;
        RECT 679.950 422.400 745.050 423.600 ;
        RECT 679.950 421.950 682.050 422.400 ;
        RECT 694.950 421.950 697.050 422.400 ;
        RECT 742.950 421.950 745.050 422.400 ;
        RECT 61.950 420.600 64.050 421.050 ;
        RECT 103.950 420.600 106.050 421.050 ;
        RECT 61.950 419.400 106.050 420.600 ;
        RECT 61.950 418.950 64.050 419.400 ;
        RECT 103.950 418.950 106.050 419.400 ;
        RECT 262.950 420.600 265.050 421.050 ;
        RECT 286.950 420.600 289.050 421.050 ;
        RECT 262.950 419.400 289.050 420.600 ;
        RECT 262.950 418.950 265.050 419.400 ;
        RECT 286.950 418.950 289.050 419.400 ;
        RECT 409.950 420.600 412.050 421.050 ;
        RECT 427.950 420.600 430.050 421.050 ;
        RECT 409.950 419.400 430.050 420.600 ;
        RECT 409.950 418.950 412.050 419.400 ;
        RECT 427.950 418.950 430.050 419.400 ;
        RECT 433.950 420.600 436.050 421.050 ;
        RECT 451.950 420.600 454.050 421.050 ;
        RECT 433.950 419.400 450.600 420.600 ;
        RECT 433.950 418.950 436.050 419.400 ;
        RECT 19.950 417.600 22.050 418.200 ;
        RECT 67.950 417.600 70.050 418.200 ;
        RECT 19.950 416.400 70.050 417.600 ;
        RECT 19.950 416.100 22.050 416.400 ;
        RECT 67.950 416.100 70.050 416.400 ;
        RECT 253.950 417.750 256.050 418.200 ;
        RECT 262.950 417.750 265.050 418.200 ;
        RECT 253.950 416.550 265.050 417.750 ;
        RECT 253.950 416.100 256.050 416.550 ;
        RECT 262.950 416.100 265.050 416.550 ;
        RECT 364.950 417.600 367.050 418.200 ;
        RECT 376.950 417.600 379.050 418.050 ;
        RECT 364.950 416.400 379.050 417.600 ;
        RECT 364.950 416.100 367.050 416.400 ;
        RECT 376.950 415.950 379.050 416.400 ;
        RECT 430.950 416.100 433.050 418.200 ;
        RECT 449.400 417.600 450.600 419.400 ;
        RECT 451.950 419.400 489.600 420.600 ;
        RECT 451.950 418.950 454.050 419.400 ;
        RECT 449.400 416.400 456.600 417.600 ;
        RECT 431.400 414.600 432.600 416.100 ;
        RECT 416.400 413.400 432.600 414.600 ;
        RECT 142.950 411.600 145.050 412.050 ;
        RECT 151.950 411.600 154.050 411.900 ;
        RECT 142.950 410.400 154.050 411.600 ;
        RECT 142.950 409.950 145.050 410.400 ;
        RECT 151.950 409.800 154.050 410.400 ;
        RECT 280.950 411.450 283.050 412.050 ;
        RECT 310.950 411.450 313.050 412.050 ;
        RECT 313.950 411.450 316.050 411.900 ;
        RECT 280.950 410.250 316.050 411.450 ;
        RECT 280.950 409.950 283.050 410.250 ;
        RECT 310.950 409.950 313.050 410.250 ;
        RECT 313.950 409.800 316.050 410.250 ;
        RECT 406.950 411.600 409.050 411.900 ;
        RECT 416.400 411.600 417.600 413.400 ;
        RECT 455.400 411.900 456.600 416.400 ;
        RECT 466.950 414.600 469.050 415.050 ;
        RECT 488.400 414.600 489.600 419.400 ;
        RECT 721.950 418.950 724.050 421.050 ;
        RECT 802.950 420.600 805.050 421.050 ;
        RECT 814.950 420.600 817.050 421.050 ;
        RECT 802.950 419.400 817.050 420.600 ;
        RECT 802.950 418.950 805.050 419.400 ;
        RECT 814.950 418.950 817.050 419.400 ;
        RECT 502.950 417.600 505.050 418.200 ;
        RECT 547.950 417.600 550.050 418.050 ;
        RECT 502.950 416.400 550.050 417.600 ;
        RECT 502.950 416.100 505.050 416.400 ;
        RECT 547.950 415.950 550.050 416.400 ;
        RECT 610.950 417.600 613.050 418.200 ;
        RECT 622.950 417.750 625.050 418.200 ;
        RECT 634.950 417.750 637.050 418.200 ;
        RECT 622.950 417.600 637.050 417.750 ;
        RECT 652.950 417.600 655.050 418.200 ;
        RECT 610.950 416.550 637.050 417.600 ;
        RECT 610.950 416.400 625.050 416.550 ;
        RECT 610.950 416.100 613.050 416.400 ;
        RECT 622.950 416.100 625.050 416.400 ;
        RECT 634.950 416.100 637.050 416.550 ;
        RECT 638.400 416.400 655.050 417.600 ;
        RECT 466.950 413.400 483.600 414.600 ;
        RECT 488.400 413.400 507.600 414.600 ;
        RECT 466.950 412.950 469.050 413.400 ;
        RECT 482.400 411.900 483.600 413.400 ;
        RECT 506.400 411.900 507.600 413.400 ;
        RECT 638.400 411.900 639.600 416.400 ;
        RECT 652.950 416.100 655.050 416.400 ;
        RECT 673.950 417.600 676.050 418.200 ;
        RECT 706.950 417.600 709.050 418.050 ;
        RECT 718.950 417.600 721.050 418.200 ;
        RECT 673.950 416.400 684.600 417.600 ;
        RECT 673.950 416.100 676.050 416.400 ;
        RECT 683.400 412.050 684.600 416.400 ;
        RECT 706.950 416.400 721.050 417.600 ;
        RECT 706.950 415.950 709.050 416.400 ;
        RECT 718.950 416.100 721.050 416.400 ;
        RECT 722.400 414.600 723.600 418.950 ;
        RECT 748.950 417.600 751.050 418.200 ;
        RECT 760.950 417.750 763.050 418.200 ;
        RECT 769.950 417.750 772.050 418.200 ;
        RECT 760.950 417.600 772.050 417.750 ;
        RECT 748.950 416.550 772.050 417.600 ;
        RECT 748.950 416.400 763.050 416.550 ;
        RECT 748.950 416.100 751.050 416.400 ;
        RECT 760.950 416.100 763.050 416.400 ;
        RECT 769.950 416.100 772.050 416.550 ;
        RECT 793.950 417.750 796.050 418.200 ;
        RECT 820.950 417.750 823.050 418.200 ;
        RECT 793.950 416.550 823.050 417.750 ;
        RECT 793.950 416.100 796.050 416.550 ;
        RECT 820.950 416.100 823.050 416.550 ;
        RECT 835.950 416.100 838.050 418.200 ;
        RECT 880.950 417.750 883.050 418.200 ;
        RECT 895.950 417.750 898.050 418.200 ;
        RECT 880.950 416.550 898.050 417.750 ;
        RECT 880.950 416.100 883.050 416.550 ;
        RECT 895.950 416.100 898.050 416.550 ;
        RECT 704.400 413.400 723.600 414.600 ;
        RECT 406.950 410.400 417.600 411.600 ;
        RECT 418.950 411.450 421.050 411.900 ;
        RECT 427.950 411.450 430.050 411.900 ;
        RECT 406.950 409.800 409.050 410.400 ;
        RECT 418.950 410.250 430.050 411.450 ;
        RECT 418.950 409.800 421.050 410.250 ;
        RECT 427.950 409.800 430.050 410.250 ;
        RECT 454.950 409.800 457.050 411.900 ;
        RECT 481.950 409.800 484.050 411.900 ;
        RECT 490.950 411.450 493.050 411.900 ;
        RECT 499.950 411.450 502.050 411.900 ;
        RECT 490.950 410.250 502.050 411.450 ;
        RECT 490.950 409.800 493.050 410.250 ;
        RECT 499.950 409.800 502.050 410.250 ;
        RECT 505.950 409.800 508.050 411.900 ;
        RECT 550.950 411.450 553.050 411.900 ;
        RECT 556.950 411.450 559.050 411.900 ;
        RECT 550.950 410.250 559.050 411.450 ;
        RECT 550.950 409.800 553.050 410.250 ;
        RECT 556.950 409.800 559.050 410.250 ;
        RECT 565.950 411.450 568.050 411.900 ;
        RECT 580.950 411.450 583.050 411.900 ;
        RECT 565.950 410.250 583.050 411.450 ;
        RECT 565.950 409.800 568.050 410.250 ;
        RECT 580.950 409.800 583.050 410.250 ;
        RECT 613.950 411.600 616.050 411.900 ;
        RECT 631.950 411.600 634.050 411.900 ;
        RECT 613.950 410.400 634.050 411.600 ;
        RECT 613.950 409.800 616.050 410.400 ;
        RECT 631.950 409.800 634.050 410.400 ;
        RECT 637.950 409.800 640.050 411.900 ;
        RECT 655.950 411.600 658.050 411.900 ;
        RECT 661.950 411.600 664.050 412.050 ;
        RECT 655.950 410.400 664.050 411.600 ;
        RECT 655.950 409.800 658.050 410.400 ;
        RECT 661.950 409.950 664.050 410.400 ;
        RECT 682.950 409.950 685.050 412.050 ;
        RECT 704.400 411.900 705.600 413.400 ;
        RECT 722.400 411.900 723.600 413.400 ;
        RECT 703.950 409.800 706.050 411.900 ;
        RECT 721.950 409.800 724.050 411.900 ;
        RECT 727.950 411.600 730.050 411.900 ;
        RECT 733.950 411.600 736.050 412.050 ;
        RECT 727.950 410.400 736.050 411.600 ;
        RECT 727.950 409.800 730.050 410.400 ;
        RECT 733.950 409.950 736.050 410.400 ;
        RECT 751.950 411.600 754.050 411.900 ;
        RECT 772.950 411.600 775.050 411.900 ;
        RECT 751.950 410.400 775.050 411.600 ;
        RECT 751.950 409.800 754.050 410.400 ;
        RECT 772.950 409.800 775.050 410.400 ;
        RECT 790.950 411.600 793.050 411.900 ;
        RECT 802.950 411.600 805.050 412.050 ;
        RECT 790.950 410.400 805.050 411.600 ;
        RECT 790.950 409.800 793.050 410.400 ;
        RECT 802.950 409.950 805.050 410.400 ;
        RECT 820.950 411.600 823.050 412.050 ;
        RECT 836.400 411.600 837.600 416.100 ;
        RECT 820.950 410.400 837.600 411.600 ;
        RECT 820.950 409.950 823.050 410.400 ;
        RECT 346.950 408.600 349.050 409.050 ;
        RECT 361.950 408.600 364.050 409.050 ;
        RECT 346.950 407.400 364.050 408.600 ;
        RECT 346.950 406.950 349.050 407.400 ;
        RECT 361.950 406.950 364.050 407.400 ;
        RECT 376.950 408.600 379.050 409.050 ;
        RECT 400.950 408.600 403.050 409.050 ;
        RECT 376.950 407.400 403.050 408.600 ;
        RECT 376.950 406.950 379.050 407.400 ;
        RECT 400.950 406.950 403.050 407.400 ;
        RECT 511.950 408.600 514.050 409.050 ;
        RECT 538.950 408.600 541.050 409.050 ;
        RECT 511.950 407.400 541.050 408.600 ;
        RECT 511.950 406.950 514.050 407.400 ;
        RECT 538.950 406.950 541.050 407.400 ;
        RECT 547.950 408.600 550.050 409.050 ;
        RECT 559.950 408.600 562.050 409.050 ;
        RECT 547.950 407.400 562.050 408.600 ;
        RECT 547.950 406.950 550.050 407.400 ;
        RECT 559.950 406.950 562.050 407.400 ;
        RECT 607.950 408.600 610.050 409.050 ;
        RECT 637.950 408.600 640.050 409.050 ;
        RECT 607.950 407.400 640.050 408.600 ;
        RECT 607.950 406.950 610.050 407.400 ;
        RECT 637.950 406.950 640.050 407.400 ;
        RECT 670.950 408.600 673.050 409.050 ;
        RECT 688.950 408.600 691.050 409.050 ;
        RECT 670.950 407.400 691.050 408.600 ;
        RECT 670.950 406.950 673.050 407.400 ;
        RECT 688.950 406.950 691.050 407.400 ;
        RECT 811.950 408.600 814.050 409.050 ;
        RECT 829.950 408.600 832.050 409.050 ;
        RECT 811.950 407.400 832.050 408.600 ;
        RECT 811.950 406.950 814.050 407.400 ;
        RECT 829.950 406.950 832.050 407.400 ;
        RECT 871.950 408.600 874.050 409.050 ;
        RECT 883.950 408.600 886.050 409.050 ;
        RECT 871.950 407.400 886.050 408.600 ;
        RECT 871.950 406.950 874.050 407.400 ;
        RECT 883.950 406.950 886.050 407.400 ;
        RECT 442.950 405.600 445.050 406.050 ;
        RECT 472.950 405.600 475.050 406.050 ;
        RECT 442.950 404.400 475.050 405.600 ;
        RECT 442.950 403.950 445.050 404.400 ;
        RECT 472.950 403.950 475.050 404.400 ;
        RECT 505.950 405.600 508.050 406.050 ;
        RECT 565.950 405.600 568.050 406.050 ;
        RECT 505.950 404.400 568.050 405.600 ;
        RECT 505.950 403.950 508.050 404.400 ;
        RECT 565.950 403.950 568.050 404.400 ;
        RECT 721.950 405.600 724.050 406.050 ;
        RECT 745.950 405.600 748.050 406.050 ;
        RECT 721.950 404.400 748.050 405.600 ;
        RECT 721.950 403.950 724.050 404.400 ;
        RECT 745.950 403.950 748.050 404.400 ;
        RECT 802.950 405.600 805.050 406.050 ;
        RECT 838.950 405.600 841.050 406.050 ;
        RECT 802.950 404.400 841.050 405.600 ;
        RECT 802.950 403.950 805.050 404.400 ;
        RECT 838.950 403.950 841.050 404.400 ;
        RECT 94.950 402.600 97.050 403.050 ;
        RECT 145.950 402.600 148.050 403.050 ;
        RECT 169.950 402.600 172.050 403.050 ;
        RECT 94.950 401.400 172.050 402.600 ;
        RECT 94.950 400.950 97.050 401.400 ;
        RECT 145.950 400.950 148.050 401.400 ;
        RECT 169.950 400.950 172.050 401.400 ;
        RECT 400.950 402.600 403.050 403.050 ;
        RECT 433.950 402.600 436.050 403.050 ;
        RECT 457.950 402.600 460.050 403.050 ;
        RECT 400.950 401.400 460.050 402.600 ;
        RECT 400.950 400.950 403.050 401.400 ;
        RECT 433.950 400.950 436.050 401.400 ;
        RECT 457.950 400.950 460.050 401.400 ;
        RECT 571.950 402.600 574.050 403.050 ;
        RECT 583.950 402.600 586.050 403.050 ;
        RECT 571.950 401.400 586.050 402.600 ;
        RECT 571.950 400.950 574.050 401.400 ;
        RECT 583.950 400.950 586.050 401.400 ;
        RECT 637.950 402.600 640.050 403.050 ;
        RECT 655.950 402.600 658.050 403.050 ;
        RECT 883.950 402.600 886.050 403.050 ;
        RECT 637.950 401.400 658.050 402.600 ;
        RECT 637.950 400.950 640.050 401.400 ;
        RECT 655.950 400.950 658.050 401.400 ;
        RECT 842.400 401.400 886.050 402.600 ;
        RECT 842.400 400.050 843.600 401.400 ;
        RECT 883.950 400.950 886.050 401.400 ;
        RECT 205.950 399.600 208.050 400.050 ;
        RECT 265.950 399.600 268.050 400.050 ;
        RECT 289.950 399.600 292.050 400.050 ;
        RECT 205.950 398.400 292.050 399.600 ;
        RECT 205.950 397.950 208.050 398.400 ;
        RECT 265.950 397.950 268.050 398.400 ;
        RECT 289.950 397.950 292.050 398.400 ;
        RECT 295.950 399.600 298.050 400.050 ;
        RECT 322.950 399.600 325.050 400.050 ;
        RECT 367.950 399.600 370.050 400.050 ;
        RECT 403.950 399.600 406.050 400.050 ;
        RECT 295.950 398.400 406.050 399.600 ;
        RECT 295.950 397.950 298.050 398.400 ;
        RECT 322.950 397.950 325.050 398.400 ;
        RECT 367.950 397.950 370.050 398.400 ;
        RECT 403.950 397.950 406.050 398.400 ;
        RECT 445.950 399.600 448.050 400.050 ;
        RECT 460.950 399.600 463.050 400.050 ;
        RECT 445.950 398.400 463.050 399.600 ;
        RECT 445.950 397.950 448.050 398.400 ;
        RECT 460.950 397.950 463.050 398.400 ;
        RECT 538.950 399.600 541.050 400.050 ;
        RECT 565.950 399.600 568.050 400.050 ;
        RECT 538.950 398.400 568.050 399.600 ;
        RECT 538.950 397.950 541.050 398.400 ;
        RECT 565.950 397.950 568.050 398.400 ;
        RECT 622.950 399.600 625.050 400.050 ;
        RECT 634.950 399.600 637.050 400.050 ;
        RECT 688.950 399.600 691.050 400.050 ;
        RECT 622.950 398.400 691.050 399.600 ;
        RECT 622.950 397.950 625.050 398.400 ;
        RECT 634.950 397.950 637.050 398.400 ;
        RECT 688.950 397.950 691.050 398.400 ;
        RECT 766.950 399.600 769.050 400.050 ;
        RECT 796.950 399.600 799.050 400.050 ;
        RECT 766.950 398.400 799.050 399.600 ;
        RECT 766.950 397.950 769.050 398.400 ;
        RECT 796.950 397.950 799.050 398.400 ;
        RECT 817.950 399.600 820.050 400.050 ;
        RECT 841.950 399.600 844.050 400.050 ;
        RECT 817.950 398.400 844.050 399.600 ;
        RECT 817.950 397.950 820.050 398.400 ;
        RECT 841.950 397.950 844.050 398.400 ;
        RECT 523.950 396.600 526.050 397.050 ;
        RECT 535.950 396.600 538.050 397.050 ;
        RECT 523.950 395.400 538.050 396.600 ;
        RECT 523.950 394.950 526.050 395.400 ;
        RECT 535.950 394.950 538.050 395.400 ;
        RECT 799.950 396.600 802.050 397.050 ;
        RECT 856.950 396.600 859.050 397.050 ;
        RECT 892.950 396.600 895.050 397.050 ;
        RECT 799.950 395.400 895.050 396.600 ;
        RECT 799.950 394.950 802.050 395.400 ;
        RECT 856.950 394.950 859.050 395.400 ;
        RECT 892.950 394.950 895.050 395.400 ;
        RECT 88.950 393.600 91.050 394.050 ;
        RECT 130.950 393.600 133.050 394.050 ;
        RECT 88.950 392.400 133.050 393.600 ;
        RECT 88.950 391.950 91.050 392.400 ;
        RECT 130.950 391.950 133.050 392.400 ;
        RECT 379.950 393.600 382.050 394.050 ;
        RECT 439.950 393.600 442.050 394.050 ;
        RECT 379.950 392.400 442.050 393.600 ;
        RECT 379.950 391.950 382.050 392.400 ;
        RECT 439.950 391.950 442.050 392.400 ;
        RECT 448.950 393.600 451.050 394.050 ;
        RECT 511.950 393.600 514.050 394.050 ;
        RECT 448.950 392.400 514.050 393.600 ;
        RECT 448.950 391.950 451.050 392.400 ;
        RECT 511.950 391.950 514.050 392.400 ;
        RECT 631.950 393.600 634.050 394.050 ;
        RECT 649.950 393.600 652.050 394.050 ;
        RECT 682.950 393.600 685.050 394.050 ;
        RECT 631.950 392.400 685.050 393.600 ;
        RECT 631.950 391.950 634.050 392.400 ;
        RECT 649.950 391.950 652.050 392.400 ;
        RECT 682.950 391.950 685.050 392.400 ;
        RECT 688.950 393.600 691.050 394.050 ;
        RECT 712.950 393.600 715.050 394.050 ;
        RECT 688.950 392.400 715.050 393.600 ;
        RECT 688.950 391.950 691.050 392.400 ;
        RECT 712.950 391.950 715.050 392.400 ;
        RECT 760.950 393.600 763.050 394.050 ;
        RECT 766.950 393.600 769.050 394.050 ;
        RECT 760.950 392.400 769.050 393.600 ;
        RECT 760.950 391.950 763.050 392.400 ;
        RECT 766.950 391.950 769.050 392.400 ;
        RECT 244.950 390.600 247.050 391.050 ;
        RECT 316.950 390.600 319.050 391.050 ;
        RECT 244.950 389.400 319.050 390.600 ;
        RECT 244.950 388.950 247.050 389.400 ;
        RECT 316.950 388.950 319.050 389.400 ;
        RECT 325.950 390.600 328.050 391.050 ;
        RECT 442.950 390.600 445.050 391.050 ;
        RECT 325.950 389.400 445.050 390.600 ;
        RECT 325.950 388.950 328.050 389.400 ;
        RECT 442.950 388.950 445.050 389.400 ;
        RECT 526.950 390.600 529.050 391.050 ;
        RECT 532.950 390.600 535.050 391.050 ;
        RECT 526.950 389.400 535.050 390.600 ;
        RECT 526.950 388.950 529.050 389.400 ;
        RECT 532.950 388.950 535.050 389.400 ;
        RECT 745.950 390.600 748.050 391.050 ;
        RECT 751.950 390.600 754.050 391.050 ;
        RECT 745.950 389.400 754.050 390.600 ;
        RECT 745.950 388.950 748.050 389.400 ;
        RECT 751.950 388.950 754.050 389.400 ;
        RECT 370.950 387.600 373.050 388.050 ;
        RECT 379.950 387.600 382.050 388.050 ;
        RECT 370.950 386.400 382.050 387.600 ;
        RECT 370.950 385.950 373.050 386.400 ;
        RECT 379.950 385.950 382.050 386.400 ;
        RECT 511.950 387.600 514.050 388.050 ;
        RECT 544.950 387.600 547.050 388.050 ;
        RECT 511.950 386.400 547.050 387.600 ;
        RECT 511.950 385.950 514.050 386.400 ;
        RECT 544.950 385.950 547.050 386.400 ;
        RECT 661.950 387.600 664.050 388.050 ;
        RECT 673.950 387.600 676.050 388.050 ;
        RECT 661.950 386.400 676.050 387.600 ;
        RECT 661.950 385.950 664.050 386.400 ;
        RECT 673.950 385.950 676.050 386.400 ;
        RECT 682.950 387.600 685.050 388.050 ;
        RECT 706.950 387.600 709.050 388.050 ;
        RECT 682.950 386.400 709.050 387.600 ;
        RECT 682.950 385.950 685.050 386.400 ;
        RECT 706.950 385.950 709.050 386.400 ;
        RECT 826.950 387.600 829.050 388.050 ;
        RECT 838.950 387.600 841.050 388.050 ;
        RECT 826.950 386.400 841.050 387.600 ;
        RECT 826.950 385.950 829.050 386.400 ;
        RECT 838.950 385.950 841.050 386.400 ;
        RECT 862.950 387.600 865.050 388.050 ;
        RECT 898.950 387.600 901.050 388.050 ;
        RECT 862.950 386.400 901.050 387.600 ;
        RECT 862.950 385.950 865.050 386.400 ;
        RECT 898.950 385.950 901.050 386.400 ;
        RECT 409.950 384.600 412.050 385.050 ;
        RECT 454.950 384.600 457.050 385.050 ;
        RECT 409.950 383.400 457.050 384.600 ;
        RECT 409.950 382.950 412.050 383.400 ;
        RECT 454.950 382.950 457.050 383.400 ;
        RECT 574.950 384.600 577.050 385.050 ;
        RECT 631.950 384.600 634.050 385.050 ;
        RECT 574.950 383.400 634.050 384.600 ;
        RECT 574.950 382.950 577.050 383.400 ;
        RECT 631.950 382.950 634.050 383.400 ;
        RECT 640.950 384.600 643.050 385.050 ;
        RECT 661.950 384.600 664.050 384.900 ;
        RECT 640.950 383.400 664.050 384.600 ;
        RECT 640.950 382.950 643.050 383.400 ;
        RECT 661.950 382.800 664.050 383.400 ;
        RECT 316.950 381.600 319.050 382.050 ;
        RECT 370.950 381.600 373.050 382.050 ;
        RECT 397.950 381.600 400.050 382.050 ;
        RECT 316.950 380.400 373.050 381.600 ;
        RECT 316.950 379.950 319.050 380.400 ;
        RECT 370.950 379.950 373.050 380.400 ;
        RECT 380.400 380.400 400.050 381.600 ;
        RECT 52.950 378.600 55.050 379.050 ;
        RECT 76.950 378.600 79.050 379.050 ;
        RECT 88.950 378.600 91.050 379.050 ;
        RECT 52.950 377.400 91.050 378.600 ;
        RECT 52.950 376.950 55.050 377.400 ;
        RECT 76.950 376.950 79.050 377.400 ;
        RECT 88.950 376.950 91.050 377.400 ;
        RECT 196.950 378.600 199.050 379.050 ;
        RECT 205.950 378.600 208.050 379.050 ;
        RECT 196.950 377.400 208.050 378.600 ;
        RECT 196.950 376.950 199.050 377.400 ;
        RECT 205.950 376.950 208.050 377.400 ;
        RECT 265.950 378.600 268.050 379.050 ;
        RECT 283.950 378.600 286.050 379.050 ;
        RECT 265.950 377.400 286.050 378.600 ;
        RECT 265.950 376.950 268.050 377.400 ;
        RECT 283.950 376.950 286.050 377.400 ;
        RECT 373.950 378.600 376.050 379.050 ;
        RECT 380.400 378.600 381.600 380.400 ;
        RECT 397.950 379.950 400.050 380.400 ;
        RECT 589.950 381.600 592.050 382.050 ;
        RECT 694.950 381.600 697.050 382.050 ;
        RECT 706.950 381.600 709.050 382.050 ;
        RECT 730.950 381.600 733.050 382.050 ;
        RECT 589.950 380.400 733.050 381.600 ;
        RECT 589.950 379.950 592.050 380.400 ;
        RECT 694.950 379.950 697.050 380.400 ;
        RECT 706.950 379.950 709.050 380.400 ;
        RECT 730.950 379.950 733.050 380.400 ;
        RECT 736.950 381.600 739.050 382.050 ;
        RECT 742.950 381.600 745.050 382.050 ;
        RECT 754.950 381.600 757.050 382.050 ;
        RECT 736.950 380.400 757.050 381.600 ;
        RECT 736.950 379.950 739.050 380.400 ;
        RECT 742.950 379.950 745.050 380.400 ;
        RECT 754.950 379.950 757.050 380.400 ;
        RECT 373.950 377.400 381.600 378.600 ;
        RECT 595.950 378.600 598.050 379.050 ;
        RECT 622.950 378.600 625.050 379.050 ;
        RECT 595.950 377.400 625.050 378.600 ;
        RECT 373.950 376.950 376.050 377.400 ;
        RECT 595.950 376.950 598.050 377.400 ;
        RECT 622.950 376.950 625.050 377.400 ;
        RECT 826.950 378.600 829.050 379.050 ;
        RECT 877.950 378.600 880.050 379.050 ;
        RECT 826.950 377.400 880.050 378.600 ;
        RECT 826.950 376.950 829.050 377.400 ;
        RECT 877.950 376.950 880.050 377.400 ;
        RECT 421.950 375.600 424.050 376.050 ;
        RECT 448.950 375.600 451.050 376.050 ;
        RECT 421.950 374.400 451.050 375.600 ;
        RECT 421.950 373.950 424.050 374.400 ;
        RECT 448.950 373.950 451.050 374.400 ;
        RECT 526.950 375.600 529.050 376.050 ;
        RECT 562.950 375.600 565.050 376.050 ;
        RECT 526.950 374.400 565.050 375.600 ;
        RECT 526.950 373.950 529.050 374.400 ;
        RECT 562.950 373.950 565.050 374.400 ;
        RECT 43.950 372.600 46.050 373.200 ;
        RECT 79.950 372.750 82.050 373.200 ;
        RECT 94.950 372.750 97.050 373.200 ;
        RECT 43.950 371.400 63.600 372.600 ;
        RECT 43.950 371.100 46.050 371.400 ;
        RECT 62.400 366.900 63.600 371.400 ;
        RECT 79.950 371.550 97.050 372.750 ;
        RECT 79.950 371.100 82.050 371.550 ;
        RECT 94.950 371.100 97.050 371.550 ;
        RECT 121.950 372.750 124.050 373.200 ;
        RECT 130.950 372.750 133.050 373.200 ;
        RECT 121.950 371.550 133.050 372.750 ;
        RECT 121.950 371.100 124.050 371.550 ;
        RECT 130.950 371.100 133.050 371.550 ;
        RECT 136.950 371.100 139.050 373.200 ;
        RECT 154.950 371.100 157.050 373.200 ;
        RECT 178.950 372.600 181.050 373.200 ;
        RECT 184.800 372.600 186.900 373.050 ;
        RECT 178.950 371.400 186.900 372.600 ;
        RECT 178.950 371.100 181.050 371.400 ;
        RECT 137.400 369.600 138.600 371.100 ;
        RECT 148.950 369.600 151.050 370.050 ;
        RECT 137.400 368.400 151.050 369.600 ;
        RECT 155.400 369.600 156.600 371.100 ;
        RECT 184.800 370.950 186.900 371.400 ;
        RECT 187.950 372.750 190.050 373.200 ;
        RECT 202.950 372.750 205.050 373.200 ;
        RECT 187.950 371.550 205.050 372.750 ;
        RECT 187.950 371.100 190.050 371.550 ;
        RECT 202.950 371.100 205.050 371.550 ;
        RECT 238.950 371.100 241.050 373.200 ;
        RECT 271.950 372.600 274.050 373.200 ;
        RECT 286.950 372.600 289.050 373.200 ;
        RECT 271.950 371.400 289.050 372.600 ;
        RECT 271.950 371.100 274.050 371.400 ;
        RECT 286.950 371.100 289.050 371.400 ;
        RECT 295.950 372.600 298.050 373.200 ;
        RECT 331.950 372.600 334.050 373.050 ;
        RECT 295.950 371.400 334.050 372.600 ;
        RECT 295.950 371.100 298.050 371.400 ;
        RECT 166.950 369.600 169.050 370.050 ;
        RECT 155.400 368.400 169.050 369.600 ;
        RECT 148.950 367.950 151.050 368.400 ;
        RECT 166.950 367.950 169.050 368.400 ;
        RECT 208.950 369.600 211.050 370.050 ;
        RECT 239.400 369.600 240.600 371.100 ;
        RECT 287.400 369.600 288.600 371.100 ;
        RECT 331.950 370.950 334.050 371.400 ;
        RECT 337.950 372.600 340.050 373.200 ;
        RECT 373.950 372.600 376.050 373.200 ;
        RECT 337.950 371.400 376.050 372.600 ;
        RECT 337.950 371.100 340.050 371.400 ;
        RECT 373.950 371.100 376.050 371.400 ;
        RECT 385.950 372.600 388.050 373.050 ;
        RECT 418.950 372.600 421.050 373.200 ;
        RECT 385.950 371.400 421.050 372.600 ;
        RECT 385.950 370.950 388.050 371.400 ;
        RECT 418.950 371.100 421.050 371.400 ;
        RECT 472.950 372.600 475.050 373.200 ;
        RECT 517.950 372.600 520.050 373.200 ;
        RECT 472.950 371.400 520.050 372.600 ;
        RECT 472.950 371.100 475.050 371.400 ;
        RECT 517.950 371.100 520.050 371.400 ;
        RECT 523.950 370.950 526.050 373.050 ;
        RECT 556.950 372.750 559.050 373.200 ;
        RECT 580.950 372.750 583.050 373.200 ;
        RECT 556.950 371.550 583.050 372.750 ;
        RECT 556.950 371.100 559.050 371.550 ;
        RECT 580.950 371.100 583.050 371.550 ;
        RECT 601.950 372.600 604.050 373.200 ;
        RECT 610.950 372.600 613.050 373.050 ;
        RECT 616.950 372.600 619.050 373.200 ;
        RECT 601.950 371.400 619.050 372.600 ;
        RECT 601.950 371.100 604.050 371.400 ;
        RECT 610.950 370.950 613.050 371.400 ;
        RECT 616.950 371.100 619.050 371.400 ;
        RECT 634.950 372.600 639.000 373.050 ;
        RECT 634.950 370.950 639.600 372.600 ;
        RECT 712.950 371.100 715.050 373.200 ;
        RECT 367.950 369.600 370.050 370.050 ;
        RECT 208.950 368.400 370.050 369.600 ;
        RECT 208.950 367.950 211.050 368.400 ;
        RECT 367.950 367.950 370.050 368.400 ;
        RECT 505.950 369.600 508.050 370.050 ;
        RECT 524.400 369.600 525.600 370.950 ;
        RECT 505.950 368.400 525.600 369.600 ;
        RECT 505.950 367.950 508.050 368.400 ;
        RECT 19.950 366.600 22.050 366.900 ;
        RECT 25.950 366.600 28.050 366.900 ;
        RECT 19.950 365.400 28.050 366.600 ;
        RECT 19.950 364.800 22.050 365.400 ;
        RECT 25.950 364.800 28.050 365.400 ;
        RECT 61.950 364.800 64.050 366.900 ;
        RECT 109.950 366.600 112.050 366.900 ;
        RECT 121.950 366.600 124.050 367.050 ;
        RECT 109.950 365.400 124.050 366.600 ;
        RECT 109.950 364.800 112.050 365.400 ;
        RECT 121.950 364.950 124.050 365.400 ;
        RECT 139.950 366.600 142.050 366.900 ;
        RECT 157.950 366.600 160.050 366.900 ;
        RECT 139.950 365.400 160.050 366.600 ;
        RECT 139.950 364.800 142.050 365.400 ;
        RECT 157.950 364.800 160.050 365.400 ;
        RECT 184.950 366.450 187.050 366.900 ;
        RECT 193.950 366.450 196.050 366.900 ;
        RECT 184.950 365.250 196.050 366.450 ;
        RECT 184.950 364.800 187.050 365.250 ;
        RECT 193.950 364.800 196.050 365.250 ;
        RECT 391.950 366.450 394.050 366.900 ;
        RECT 439.950 366.450 442.050 366.900 ;
        RECT 391.950 365.250 442.050 366.450 ;
        RECT 391.950 364.800 394.050 365.250 ;
        RECT 439.950 364.800 442.050 365.250 ;
        RECT 457.950 366.450 460.050 366.900 ;
        RECT 469.950 366.450 472.050 366.900 ;
        RECT 457.950 365.250 472.050 366.450 ;
        RECT 457.950 364.800 460.050 365.250 ;
        RECT 469.950 364.800 472.050 365.250 ;
        RECT 562.950 366.450 565.050 366.900 ;
        RECT 571.950 366.450 574.050 366.900 ;
        RECT 562.950 365.250 574.050 366.450 ;
        RECT 562.950 364.800 565.050 365.250 ;
        RECT 571.950 364.800 574.050 365.250 ;
        RECT 580.950 366.600 583.050 367.050 ;
        RECT 638.400 366.900 639.600 370.950 ;
        RECT 713.400 367.050 714.600 371.100 ;
        RECT 724.950 370.950 727.050 373.050 ;
        RECT 736.950 371.100 739.050 373.200 ;
        RECT 760.950 372.600 763.050 373.200 ;
        RECT 769.950 372.750 772.050 373.200 ;
        RECT 775.950 372.750 778.050 373.200 ;
        RECT 769.950 372.600 778.050 372.750 ;
        RECT 760.950 371.550 778.050 372.600 ;
        RECT 760.950 371.400 772.050 371.550 ;
        RECT 760.950 371.100 763.050 371.400 ;
        RECT 769.950 371.100 772.050 371.400 ;
        RECT 775.950 371.100 778.050 371.550 ;
        RECT 781.950 371.100 784.050 373.200 ;
        RECT 793.950 372.750 796.050 373.200 ;
        RECT 805.950 372.750 808.050 373.200 ;
        RECT 793.950 371.550 808.050 372.750 ;
        RECT 793.950 371.100 796.050 371.550 ;
        RECT 805.950 371.100 808.050 371.550 ;
        RECT 811.950 372.750 814.050 373.200 ;
        RECT 817.950 372.750 820.050 373.200 ;
        RECT 811.950 371.550 820.050 372.750 ;
        RECT 829.950 372.600 832.050 376.050 ;
        RECT 874.950 373.950 877.050 376.050 ;
        RECT 811.950 371.100 814.050 371.550 ;
        RECT 817.950 371.100 820.050 371.550 ;
        RECT 827.400 372.000 832.050 372.600 ;
        RECT 832.950 372.600 835.050 373.200 ;
        RECT 850.950 372.600 853.050 373.200 ;
        RECT 827.400 371.400 831.600 372.000 ;
        RECT 832.950 371.400 853.050 372.600 ;
        RECT 598.950 366.600 601.050 366.900 ;
        RECT 580.950 365.400 601.050 366.600 ;
        RECT 580.950 364.950 583.050 365.400 ;
        RECT 598.950 364.800 601.050 365.400 ;
        RECT 637.950 364.800 640.050 366.900 ;
        RECT 649.950 366.450 652.050 366.900 ;
        RECT 658.950 366.450 661.050 366.900 ;
        RECT 649.950 365.250 661.050 366.450 ;
        RECT 649.950 364.800 652.050 365.250 ;
        RECT 658.950 364.800 661.050 365.250 ;
        RECT 673.950 366.450 676.050 366.900 ;
        RECT 679.950 366.450 682.050 366.900 ;
        RECT 673.950 365.250 682.050 366.450 ;
        RECT 673.950 364.800 676.050 365.250 ;
        RECT 679.950 364.800 682.050 365.250 ;
        RECT 697.950 366.600 700.050 367.050 ;
        RECT 703.950 366.600 706.050 366.900 ;
        RECT 697.950 365.400 706.050 366.600 ;
        RECT 713.400 365.400 718.050 367.050 ;
        RECT 725.400 366.600 726.600 370.950 ;
        RECT 737.400 367.050 738.600 371.100 ;
        RECT 727.950 366.600 730.050 366.900 ;
        RECT 725.400 365.400 730.050 366.600 ;
        RECT 737.400 365.400 742.050 367.050 ;
        RECT 697.950 364.950 700.050 365.400 ;
        RECT 703.950 364.800 706.050 365.400 ;
        RECT 714.000 364.950 718.050 365.400 ;
        RECT 727.950 364.800 730.050 365.400 ;
        RECT 738.000 364.950 742.050 365.400 ;
        RECT 745.950 366.600 748.050 367.050 ;
        RECT 751.950 366.600 754.050 366.900 ;
        RECT 745.950 365.400 754.050 366.600 ;
        RECT 745.950 364.950 748.050 365.400 ;
        RECT 751.950 364.800 754.050 365.400 ;
        RECT 757.950 366.600 760.050 366.900 ;
        RECT 772.950 366.600 775.050 366.900 ;
        RECT 757.950 366.450 775.050 366.600 ;
        RECT 778.950 366.450 781.050 366.900 ;
        RECT 757.950 365.400 781.050 366.450 ;
        RECT 757.950 364.800 760.050 365.400 ;
        RECT 772.950 365.250 781.050 365.400 ;
        RECT 772.950 364.800 775.050 365.250 ;
        RECT 778.950 364.800 781.050 365.250 ;
        RECT 166.950 363.600 169.050 364.050 ;
        RECT 175.950 363.600 178.050 364.050 ;
        RECT 208.950 363.600 211.050 364.050 ;
        RECT 166.950 362.400 211.050 363.600 ;
        RECT 166.950 361.950 169.050 362.400 ;
        RECT 175.950 361.950 178.050 362.400 ;
        RECT 208.950 361.950 211.050 362.400 ;
        RECT 313.950 363.600 316.050 364.050 ;
        RECT 325.950 363.600 328.050 364.050 ;
        RECT 313.950 362.400 328.050 363.600 ;
        RECT 313.950 361.950 316.050 362.400 ;
        RECT 325.950 361.950 328.050 362.400 ;
        RECT 367.950 363.600 370.050 364.050 ;
        RECT 385.950 363.600 388.050 364.050 ;
        RECT 367.950 362.400 388.050 363.600 ;
        RECT 367.950 361.950 370.050 362.400 ;
        RECT 385.950 361.950 388.050 362.400 ;
        RECT 496.950 363.600 499.050 364.050 ;
        RECT 511.950 363.600 514.050 364.050 ;
        RECT 496.950 362.400 514.050 363.600 ;
        RECT 496.950 361.950 499.050 362.400 ;
        RECT 511.950 361.950 514.050 362.400 ;
        RECT 418.950 360.600 421.050 361.050 ;
        RECT 442.950 360.600 445.050 361.050 ;
        RECT 418.950 359.400 445.050 360.600 ;
        RECT 418.950 358.950 421.050 359.400 ;
        RECT 442.950 358.950 445.050 359.400 ;
        RECT 454.950 360.600 457.050 361.050 ;
        RECT 493.950 360.600 496.050 361.050 ;
        RECT 454.950 359.400 496.050 360.600 ;
        RECT 454.950 358.950 457.050 359.400 ;
        RECT 493.950 358.950 496.050 359.400 ;
        RECT 532.950 360.600 535.050 361.050 ;
        RECT 547.950 360.600 550.050 361.050 ;
        RECT 532.950 359.400 550.050 360.600 ;
        RECT 532.950 358.950 535.050 359.400 ;
        RECT 547.950 358.950 550.050 359.400 ;
        RECT 592.950 360.600 595.050 361.050 ;
        RECT 619.950 360.600 622.050 361.050 ;
        RECT 592.950 359.400 622.050 360.600 ;
        RECT 592.950 358.950 595.050 359.400 ;
        RECT 619.950 358.950 622.050 359.400 ;
        RECT 631.950 360.600 634.050 361.050 ;
        RECT 721.950 360.600 724.050 361.050 ;
        RECT 631.950 359.400 724.050 360.600 ;
        RECT 782.400 360.600 783.600 371.100 ;
        RECT 784.950 366.600 787.050 366.900 ;
        RECT 793.950 366.600 796.050 367.050 ;
        RECT 784.950 365.400 796.050 366.600 ;
        RECT 827.400 366.600 828.600 371.400 ;
        RECT 832.950 371.100 835.050 371.400 ;
        RECT 850.950 371.100 853.050 371.400 ;
        RECT 875.400 366.900 876.600 373.950 ;
        RECT 877.950 372.750 880.050 373.200 ;
        RECT 898.950 372.750 901.050 373.200 ;
        RECT 877.950 371.550 901.050 372.750 ;
        RECT 877.950 371.100 880.050 371.550 ;
        RECT 898.950 371.100 901.050 371.550 ;
        RECT 829.950 366.600 832.050 366.900 ;
        RECT 827.400 365.400 832.050 366.600 ;
        RECT 784.950 364.800 787.050 365.400 ;
        RECT 793.950 364.950 796.050 365.400 ;
        RECT 829.950 364.800 832.050 365.400 ;
        RECT 874.950 364.800 877.050 366.900 ;
        RECT 796.950 363.600 799.050 364.050 ;
        RECT 802.950 363.600 805.050 364.050 ;
        RECT 796.950 362.400 805.050 363.600 ;
        RECT 796.950 361.950 799.050 362.400 ;
        RECT 802.950 361.950 805.050 362.400 ;
        RECT 877.950 363.600 880.050 364.050 ;
        RECT 883.950 363.600 886.050 364.050 ;
        RECT 877.950 362.400 886.050 363.600 ;
        RECT 877.950 361.950 880.050 362.400 ;
        RECT 883.950 361.950 886.050 362.400 ;
        RECT 787.950 360.600 790.050 361.050 ;
        RECT 782.400 359.400 790.050 360.600 ;
        RECT 631.950 358.950 634.050 359.400 ;
        RECT 721.950 358.950 724.050 359.400 ;
        RECT 787.950 358.950 790.050 359.400 ;
        RECT 793.950 360.600 796.050 361.050 ;
        RECT 817.950 360.600 820.050 361.050 ;
        RECT 793.950 359.400 820.050 360.600 ;
        RECT 793.950 358.950 796.050 359.400 ;
        RECT 817.950 358.950 820.050 359.400 ;
        RECT 868.950 360.600 871.050 361.050 ;
        RECT 895.950 360.600 898.050 361.050 ;
        RECT 868.950 359.400 898.050 360.600 ;
        RECT 868.950 358.950 871.050 359.400 ;
        RECT 895.950 358.950 898.050 359.400 ;
        RECT 127.950 357.600 130.050 358.050 ;
        RECT 175.950 357.600 178.050 358.050 ;
        RECT 187.950 357.600 190.050 358.050 ;
        RECT 220.950 357.600 223.050 358.050 ;
        RECT 127.950 356.400 223.050 357.600 ;
        RECT 127.950 355.950 130.050 356.400 ;
        RECT 175.950 355.950 178.050 356.400 ;
        RECT 187.950 355.950 190.050 356.400 ;
        RECT 220.950 355.950 223.050 356.400 ;
        RECT 94.950 354.600 97.050 355.050 ;
        RECT 409.950 354.600 412.050 355.050 ;
        RECT 94.950 353.400 412.050 354.600 ;
        RECT 94.950 352.950 97.050 353.400 ;
        RECT 409.950 352.950 412.050 353.400 ;
        RECT 445.950 354.600 448.050 355.050 ;
        RECT 463.950 354.600 466.050 355.050 ;
        RECT 445.950 353.400 466.050 354.600 ;
        RECT 445.950 352.950 448.050 353.400 ;
        RECT 463.950 352.950 466.050 353.400 ;
        RECT 517.950 354.600 520.050 355.050 ;
        RECT 535.950 354.600 538.050 355.050 ;
        RECT 517.950 353.400 538.050 354.600 ;
        RECT 517.950 352.950 520.050 353.400 ;
        RECT 535.950 352.950 538.050 353.400 ;
        RECT 715.950 354.600 718.050 355.050 ;
        RECT 721.950 354.600 724.050 355.050 ;
        RECT 739.950 354.600 742.050 355.050 ;
        RECT 793.950 354.600 796.050 355.050 ;
        RECT 715.950 353.400 796.050 354.600 ;
        RECT 715.950 352.950 718.050 353.400 ;
        RECT 721.950 352.950 724.050 353.400 ;
        RECT 739.950 352.950 742.050 353.400 ;
        RECT 793.950 352.950 796.050 353.400 ;
        RECT 298.950 351.600 301.050 352.050 ;
        RECT 340.950 351.600 343.050 352.050 ;
        RECT 298.950 350.400 343.050 351.600 ;
        RECT 298.950 349.950 301.050 350.400 ;
        RECT 340.950 349.950 343.050 350.400 ;
        RECT 433.950 351.600 436.050 352.050 ;
        RECT 472.950 351.600 475.050 352.050 ;
        RECT 433.950 350.400 475.050 351.600 ;
        RECT 433.950 349.950 436.050 350.400 ;
        RECT 472.950 349.950 475.050 350.400 ;
        RECT 850.950 351.600 853.050 352.050 ;
        RECT 886.950 351.600 889.050 352.050 ;
        RECT 850.950 350.400 889.050 351.600 ;
        RECT 850.950 349.950 853.050 350.400 ;
        RECT 886.950 349.950 889.050 350.400 ;
        RECT 97.950 348.600 100.050 349.050 ;
        RECT 112.950 348.600 115.050 349.050 ;
        RECT 97.950 347.400 115.050 348.600 ;
        RECT 97.950 346.950 100.050 347.400 ;
        RECT 112.950 346.950 115.050 347.400 ;
        RECT 286.950 348.600 289.050 349.050 ;
        RECT 376.950 348.600 379.050 349.050 ;
        RECT 391.950 348.600 394.050 349.050 ;
        RECT 286.950 347.400 394.050 348.600 ;
        RECT 286.950 346.950 289.050 347.400 ;
        RECT 376.950 346.950 379.050 347.400 ;
        RECT 391.950 346.950 394.050 347.400 ;
        RECT 400.950 348.600 403.050 349.050 ;
        RECT 418.950 348.600 421.050 349.050 ;
        RECT 400.950 347.400 421.050 348.600 ;
        RECT 400.950 346.950 403.050 347.400 ;
        RECT 418.950 346.950 421.050 347.400 ;
        RECT 484.950 348.600 487.050 349.050 ;
        RECT 592.950 348.600 595.050 349.050 ;
        RECT 484.950 347.400 595.050 348.600 ;
        RECT 484.950 346.950 487.050 347.400 ;
        RECT 592.950 346.950 595.050 347.400 ;
        RECT 697.950 348.600 700.050 349.050 ;
        RECT 709.950 348.600 712.050 349.050 ;
        RECT 733.950 348.600 736.050 349.050 ;
        RECT 739.950 348.600 742.050 349.050 ;
        RECT 697.950 347.400 742.050 348.600 ;
        RECT 697.950 346.950 700.050 347.400 ;
        RECT 709.950 346.950 712.050 347.400 ;
        RECT 733.950 346.950 736.050 347.400 ;
        RECT 739.950 346.950 742.050 347.400 ;
        RECT 811.950 348.600 814.050 349.050 ;
        RECT 841.950 348.600 844.050 349.050 ;
        RECT 811.950 347.400 844.050 348.600 ;
        RECT 811.950 346.950 814.050 347.400 ;
        RECT 841.950 346.950 844.050 347.400 ;
        RECT 874.950 348.600 877.050 349.050 ;
        RECT 889.950 348.600 892.050 349.050 ;
        RECT 874.950 347.400 892.050 348.600 ;
        RECT 874.950 346.950 877.050 347.400 ;
        RECT 889.950 346.950 892.050 347.400 ;
        RECT 148.950 345.600 151.050 346.050 ;
        RECT 181.950 345.600 184.050 346.050 ;
        RECT 148.950 344.400 184.050 345.600 ;
        RECT 148.950 343.950 151.050 344.400 ;
        RECT 181.950 343.950 184.050 344.400 ;
        RECT 199.950 345.600 202.050 346.050 ;
        RECT 217.800 345.600 219.900 346.050 ;
        RECT 199.950 344.400 219.900 345.600 ;
        RECT 199.950 343.950 202.050 344.400 ;
        RECT 217.800 343.950 219.900 344.400 ;
        RECT 334.950 345.600 337.050 346.050 ;
        RECT 358.950 345.600 361.050 346.050 ;
        RECT 334.950 344.400 361.050 345.600 ;
        RECT 334.950 343.950 337.050 344.400 ;
        RECT 358.950 343.950 361.050 344.400 ;
        RECT 397.950 345.600 400.050 346.050 ;
        RECT 427.950 345.600 430.050 346.050 ;
        RECT 451.950 345.600 454.050 346.050 ;
        RECT 397.950 344.400 454.050 345.600 ;
        RECT 397.950 343.950 400.050 344.400 ;
        RECT 427.950 343.950 430.050 344.400 ;
        RECT 451.950 343.950 454.050 344.400 ;
        RECT 673.950 345.600 676.050 346.050 ;
        RECT 688.950 345.600 691.050 346.050 ;
        RECT 673.950 344.400 691.050 345.600 ;
        RECT 673.950 343.950 676.050 344.400 ;
        RECT 688.950 343.950 691.050 344.400 ;
        RECT 22.950 342.600 25.050 343.050 ;
        RECT 103.950 342.600 106.050 343.050 ;
        RECT 22.950 341.400 106.050 342.600 ;
        RECT 22.950 340.950 25.050 341.400 ;
        RECT 103.950 340.950 106.050 341.400 ;
        RECT 121.950 342.600 124.050 343.050 ;
        RECT 169.950 342.600 172.050 343.050 ;
        RECT 121.950 341.400 172.050 342.600 ;
        RECT 121.950 340.950 124.050 341.400 ;
        RECT 169.950 340.950 172.050 341.400 ;
        RECT 472.950 342.600 475.050 343.050 ;
        RECT 499.950 342.600 502.050 343.050 ;
        RECT 472.950 341.400 502.050 342.600 ;
        RECT 472.950 340.950 475.050 341.400 ;
        RECT 499.950 340.950 502.050 341.400 ;
        RECT 514.950 342.600 517.050 343.050 ;
        RECT 526.950 342.600 529.050 343.050 ;
        RECT 514.950 341.400 529.050 342.600 ;
        RECT 514.950 340.950 517.050 341.400 ;
        RECT 526.950 340.950 529.050 341.400 ;
        RECT 541.950 342.600 544.050 343.050 ;
        RECT 556.950 342.600 559.050 343.050 ;
        RECT 541.950 341.400 559.050 342.600 ;
        RECT 541.950 340.950 544.050 341.400 ;
        RECT 556.950 340.950 559.050 341.400 ;
        RECT 694.950 340.950 697.050 343.050 ;
        RECT 741.000 342.600 745.050 343.050 ;
        RECT 740.400 340.950 745.050 342.600 ;
        RECT 754.950 342.600 757.050 343.050 ;
        RECT 760.950 342.600 763.050 343.050 ;
        RECT 754.950 341.400 763.050 342.600 ;
        RECT 754.950 340.950 757.050 341.400 ;
        RECT 760.950 340.950 763.050 341.400 ;
        RECT 802.950 342.600 805.050 343.050 ;
        RECT 808.950 342.600 811.050 343.050 ;
        RECT 837.000 342.600 841.050 343.050 ;
        RECT 802.950 341.400 811.050 342.600 ;
        RECT 802.950 340.950 805.050 341.400 ;
        RECT 808.950 340.950 811.050 341.400 ;
        RECT 836.400 340.950 841.050 342.600 ;
        RECT 43.950 339.600 46.050 340.200 ;
        RECT 49.950 339.600 52.050 340.200 ;
        RECT 205.950 339.600 208.050 340.200 ;
        RECT 43.950 338.400 52.050 339.600 ;
        RECT 43.950 338.100 46.050 338.400 ;
        RECT 49.950 338.100 52.050 338.400 ;
        RECT 185.400 338.400 208.050 339.600 ;
        RECT 185.400 333.900 186.600 338.400 ;
        RECT 205.950 338.100 208.050 338.400 ;
        RECT 223.950 339.600 226.050 340.050 ;
        RECT 232.950 339.600 235.050 340.200 ;
        RECT 223.950 338.400 235.050 339.600 ;
        RECT 223.950 337.950 226.050 338.400 ;
        RECT 232.950 338.100 235.050 338.400 ;
        RECT 256.950 339.600 259.050 340.200 ;
        RECT 268.950 339.600 271.050 340.050 ;
        RECT 274.950 339.600 277.050 340.200 ;
        RECT 256.950 338.400 277.050 339.600 ;
        RECT 256.950 338.100 259.050 338.400 ;
        RECT 268.950 337.950 271.050 338.400 ;
        RECT 274.950 338.100 277.050 338.400 ;
        RECT 298.950 339.600 301.050 340.200 ;
        RECT 310.950 339.600 313.050 340.050 ;
        RECT 298.950 338.400 313.050 339.600 ;
        RECT 298.950 338.100 301.050 338.400 ;
        RECT 310.950 337.950 313.050 338.400 ;
        RECT 337.950 339.600 340.050 340.050 ;
        RECT 346.950 339.600 349.050 340.050 ;
        RECT 337.950 338.400 349.050 339.600 ;
        RECT 337.950 337.950 340.050 338.400 ;
        RECT 346.950 337.950 349.050 338.400 ;
        RECT 355.950 339.750 358.050 340.200 ;
        RECT 367.950 339.750 370.050 340.200 ;
        RECT 355.950 338.550 370.050 339.750 ;
        RECT 355.950 338.100 358.050 338.550 ;
        RECT 367.950 338.100 370.050 338.550 ;
        RECT 394.950 339.750 397.050 340.200 ;
        RECT 400.950 339.750 403.050 340.200 ;
        RECT 394.950 338.550 403.050 339.750 ;
        RECT 394.950 338.100 397.050 338.550 ;
        RECT 400.950 338.100 403.050 338.550 ;
        RECT 406.950 339.600 409.050 340.200 ;
        RECT 439.950 339.600 442.050 340.050 ;
        RECT 406.950 338.400 442.050 339.600 ;
        RECT 406.950 338.100 409.050 338.400 ;
        RECT 439.950 337.950 442.050 338.400 ;
        RECT 457.950 339.600 460.050 340.200 ;
        RECT 466.950 339.600 469.050 340.050 ;
        RECT 478.950 339.600 481.050 340.200 ;
        RECT 457.950 338.400 469.050 339.600 ;
        RECT 457.950 338.100 460.050 338.400 ;
        RECT 466.950 337.950 469.050 338.400 ;
        RECT 476.400 338.400 481.050 339.600 ;
        RECT 476.400 336.600 477.600 338.400 ;
        RECT 478.950 338.100 481.050 338.400 ;
        RECT 490.950 339.750 493.050 340.200 ;
        RECT 529.950 339.750 532.050 340.200 ;
        RECT 490.950 338.550 532.050 339.750 ;
        RECT 490.950 338.100 493.050 338.550 ;
        RECT 529.950 338.100 532.050 338.550 ;
        RECT 550.950 338.100 553.050 340.200 ;
        RECT 562.950 339.600 565.050 340.050 ;
        RECT 577.950 339.600 580.050 340.200 ;
        RECT 562.950 338.400 580.050 339.600 ;
        RECT 470.400 336.000 477.600 336.600 ;
        RECT 469.950 335.400 477.600 336.000 ;
        RECT 184.950 331.800 187.050 333.900 ;
        RECT 190.950 333.600 193.050 333.900 ;
        RECT 202.950 333.600 205.050 333.900 ;
        RECT 190.950 333.450 205.050 333.600 ;
        RECT 223.950 333.450 226.050 333.900 ;
        RECT 190.950 332.400 226.050 333.450 ;
        RECT 190.950 331.800 193.050 332.400 ;
        RECT 202.950 332.250 226.050 332.400 ;
        RECT 202.950 331.800 205.050 332.250 ;
        RECT 223.950 331.800 226.050 332.250 ;
        RECT 277.950 333.600 280.050 333.900 ;
        RECT 286.950 333.600 289.050 334.050 ;
        RECT 277.950 332.400 289.050 333.600 ;
        RECT 277.950 331.800 280.050 332.400 ;
        RECT 286.950 331.950 289.050 332.400 ;
        RECT 301.950 333.450 304.050 333.900 ;
        RECT 307.950 333.600 310.050 333.900 ;
        RECT 316.950 333.600 319.050 333.900 ;
        RECT 307.950 333.450 319.050 333.600 ;
        RECT 301.950 332.400 319.050 333.450 ;
        RECT 301.950 332.250 310.050 332.400 ;
        RECT 301.950 331.800 304.050 332.250 ;
        RECT 307.950 331.800 310.050 332.250 ;
        RECT 316.950 331.800 319.050 332.400 ;
        RECT 391.950 333.450 394.050 333.900 ;
        RECT 403.950 333.450 406.050 333.900 ;
        RECT 391.950 332.250 406.050 333.450 ;
        RECT 391.950 331.800 394.050 332.250 ;
        RECT 403.950 331.800 406.050 332.250 ;
        RECT 418.950 333.450 421.050 333.900 ;
        RECT 424.950 333.600 427.050 333.900 ;
        RECT 454.950 333.600 457.050 333.900 ;
        RECT 424.950 333.450 457.050 333.600 ;
        RECT 418.950 332.400 457.050 333.450 ;
        RECT 418.950 332.250 427.050 332.400 ;
        RECT 418.950 331.800 421.050 332.250 ;
        RECT 424.950 331.800 427.050 332.250 ;
        RECT 454.950 331.800 457.050 332.400 ;
        RECT 469.950 331.950 472.050 335.400 ;
        RECT 481.950 333.450 484.050 333.900 ;
        RECT 490.950 333.450 493.050 333.900 ;
        RECT 481.950 332.250 493.050 333.450 ;
        RECT 481.950 331.800 484.050 332.250 ;
        RECT 490.950 331.800 493.050 332.250 ;
        RECT 496.950 333.450 499.050 333.900 ;
        RECT 526.950 333.600 529.050 333.900 ;
        RECT 551.400 333.600 552.600 338.100 ;
        RECT 562.950 337.950 565.050 338.400 ;
        RECT 577.950 338.100 580.050 338.400 ;
        RECT 583.950 339.600 586.050 340.200 ;
        RECT 589.950 339.600 592.050 340.050 ;
        RECT 601.950 339.600 604.050 340.200 ;
        RECT 583.950 338.400 604.050 339.600 ;
        RECT 583.950 338.100 586.050 338.400 ;
        RECT 589.950 337.950 592.050 338.400 ;
        RECT 601.950 338.100 604.050 338.400 ;
        RECT 625.950 339.750 628.050 340.200 ;
        RECT 637.950 339.750 640.050 340.200 ;
        RECT 625.950 338.550 640.050 339.750 ;
        RECT 625.950 338.100 628.050 338.550 ;
        RECT 637.950 338.100 640.050 338.550 ;
        RECT 526.950 333.450 552.600 333.600 ;
        RECT 496.950 332.400 552.600 333.450 ;
        RECT 553.950 333.450 556.050 333.900 ;
        RECT 562.950 333.450 565.050 333.900 ;
        RECT 496.950 332.250 529.050 332.400 ;
        RECT 496.950 331.800 499.050 332.250 ;
        RECT 526.950 331.800 529.050 332.250 ;
        RECT 553.950 332.250 565.050 333.450 ;
        RECT 553.950 331.800 556.050 332.250 ;
        RECT 562.950 331.800 565.050 332.250 ;
        RECT 637.950 333.600 640.050 334.050 ;
        RECT 695.400 333.900 696.600 340.950 ;
        RECT 703.950 339.600 706.050 340.200 ;
        RECT 727.950 339.600 730.050 340.050 ;
        RECT 740.400 339.600 741.600 340.950 ;
        RECT 703.950 338.400 730.050 339.600 ;
        RECT 703.950 338.100 706.050 338.400 ;
        RECT 727.950 337.950 730.050 338.400 ;
        RECT 737.400 338.400 741.600 339.600 ;
        RECT 745.950 339.750 748.050 340.200 ;
        RECT 751.950 339.750 754.050 340.200 ;
        RECT 745.950 338.550 754.050 339.750 ;
        RECT 737.400 333.900 738.600 338.400 ;
        RECT 745.950 338.100 748.050 338.550 ;
        RECT 751.950 338.100 754.050 338.550 ;
        RECT 775.950 339.600 778.050 340.050 ;
        RECT 787.950 339.600 790.050 340.200 ;
        RECT 775.950 338.400 790.050 339.600 ;
        RECT 775.950 337.950 778.050 338.400 ;
        RECT 787.950 338.100 790.050 338.400 ;
        RECT 823.950 339.600 826.050 340.050 ;
        RECT 832.950 339.600 835.050 340.200 ;
        RECT 823.950 338.400 835.050 339.600 ;
        RECT 823.950 337.950 826.050 338.400 ;
        RECT 832.950 338.100 835.050 338.400 ;
        RECT 836.400 336.600 837.600 340.950 ;
        RECT 850.950 337.950 853.050 340.050 ;
        RECT 830.400 335.400 837.600 336.600 ;
        RECT 830.400 333.900 831.600 335.400 ;
        RECT 851.400 334.050 852.600 337.950 ;
        RECT 865.950 336.600 868.050 340.050 ;
        RECT 865.950 336.000 870.600 336.600 ;
        RECT 866.400 335.400 870.600 336.000 ;
        RECT 652.950 333.600 655.050 333.900 ;
        RECT 637.950 332.400 655.050 333.600 ;
        RECT 637.950 331.950 640.050 332.400 ;
        RECT 652.950 331.800 655.050 332.400 ;
        RECT 694.950 331.800 697.050 333.900 ;
        RECT 700.950 333.600 703.050 333.900 ;
        RECT 718.950 333.600 721.050 333.900 ;
        RECT 700.950 332.400 721.050 333.600 ;
        RECT 700.950 331.800 703.050 332.400 ;
        RECT 718.950 331.800 721.050 332.400 ;
        RECT 736.950 331.800 739.050 333.900 ;
        RECT 751.950 333.450 754.050 333.900 ;
        RECT 763.950 333.450 766.050 333.900 ;
        RECT 751.950 332.250 766.050 333.450 ;
        RECT 751.950 331.800 754.050 332.250 ;
        RECT 763.950 331.800 766.050 332.250 ;
        RECT 769.950 333.450 772.050 333.900 ;
        RECT 775.950 333.450 778.050 333.900 ;
        RECT 769.950 332.250 778.050 333.450 ;
        RECT 769.950 331.800 772.050 332.250 ;
        RECT 775.950 331.800 778.050 332.250 ;
        RECT 829.950 331.800 832.050 333.900 ;
        RECT 850.950 331.950 853.050 334.050 ;
        RECT 869.400 333.600 870.600 335.400 ;
        RECT 874.950 333.600 877.050 334.050 ;
        RECT 869.400 332.400 877.050 333.600 ;
        RECT 874.950 331.950 877.050 332.400 ;
        RECT 76.950 330.600 79.050 331.050 ;
        RECT 85.950 330.600 88.050 331.050 ;
        RECT 130.950 330.600 133.050 331.050 ;
        RECT 145.950 330.600 148.050 331.050 ;
        RECT 76.950 329.400 148.050 330.600 ;
        RECT 76.950 328.950 79.050 329.400 ;
        RECT 85.950 328.950 88.050 329.400 ;
        RECT 130.950 328.950 133.050 329.400 ;
        RECT 145.950 328.950 148.050 329.400 ;
        RECT 430.950 330.600 433.050 331.050 ;
        RECT 448.950 330.600 451.050 331.050 ;
        RECT 430.950 329.400 451.050 330.600 ;
        RECT 430.950 328.950 433.050 329.400 ;
        RECT 448.950 328.950 451.050 329.400 ;
        RECT 493.950 330.600 496.050 330.900 ;
        RECT 502.950 330.600 505.050 331.050 ;
        RECT 493.950 329.400 505.050 330.600 ;
        RECT 493.950 328.800 496.050 329.400 ;
        RECT 502.950 328.950 505.050 329.400 ;
        RECT 643.950 330.600 646.050 331.050 ;
        RECT 649.950 330.600 652.050 331.050 ;
        RECT 643.950 329.400 652.050 330.600 ;
        RECT 643.950 328.950 646.050 329.400 ;
        RECT 649.950 328.950 652.050 329.400 ;
        RECT 349.950 327.600 352.050 328.050 ;
        RECT 388.950 327.600 391.050 328.050 ;
        RECT 349.950 326.400 391.050 327.600 ;
        RECT 349.950 325.950 352.050 326.400 ;
        RECT 388.950 325.950 391.050 326.400 ;
        RECT 466.950 327.600 469.050 328.050 ;
        RECT 532.950 327.600 535.050 328.050 ;
        RECT 547.950 327.600 550.050 328.050 ;
        RECT 466.950 326.400 550.050 327.600 ;
        RECT 466.950 325.950 469.050 326.400 ;
        RECT 532.950 325.950 535.050 326.400 ;
        RECT 547.950 325.950 550.050 326.400 ;
        RECT 556.950 327.600 559.050 328.050 ;
        RECT 592.950 327.600 595.050 328.050 ;
        RECT 622.950 327.600 625.050 328.050 ;
        RECT 556.950 326.400 625.050 327.600 ;
        RECT 556.950 325.950 559.050 326.400 ;
        RECT 592.950 325.950 595.050 326.400 ;
        RECT 622.950 325.950 625.050 326.400 ;
        RECT 652.950 327.600 655.050 328.050 ;
        RECT 670.950 327.600 673.050 328.050 ;
        RECT 652.950 326.400 673.050 327.600 ;
        RECT 652.950 325.950 655.050 326.400 ;
        RECT 670.950 325.950 673.050 326.400 ;
        RECT 835.950 327.600 838.050 328.050 ;
        RECT 856.950 327.600 859.050 328.050 ;
        RECT 835.950 326.400 859.050 327.600 ;
        RECT 835.950 325.950 838.050 326.400 ;
        RECT 856.950 325.950 859.050 326.400 ;
        RECT 322.950 324.600 325.050 325.050 ;
        RECT 337.950 324.600 340.050 325.050 ;
        RECT 373.950 324.600 376.050 325.050 ;
        RECT 394.950 324.600 397.050 325.050 ;
        RECT 403.950 324.600 406.050 325.050 ;
        RECT 322.950 323.400 406.050 324.600 ;
        RECT 322.950 322.950 325.050 323.400 ;
        RECT 337.950 322.950 340.050 323.400 ;
        RECT 373.950 322.950 376.050 323.400 ;
        RECT 394.950 322.950 397.050 323.400 ;
        RECT 403.950 322.950 406.050 323.400 ;
        RECT 439.950 324.600 442.050 325.050 ;
        RECT 496.950 324.600 499.050 325.050 ;
        RECT 439.950 323.400 499.050 324.600 ;
        RECT 439.950 322.950 442.050 323.400 ;
        RECT 496.950 322.950 499.050 323.400 ;
        RECT 862.950 324.600 865.050 325.050 ;
        RECT 886.950 324.600 889.050 325.050 ;
        RECT 892.950 324.600 895.050 325.050 ;
        RECT 862.950 323.400 895.050 324.600 ;
        RECT 862.950 322.950 865.050 323.400 ;
        RECT 886.950 322.950 889.050 323.400 ;
        RECT 892.950 322.950 895.050 323.400 ;
        RECT 112.950 321.600 115.050 322.050 ;
        RECT 190.950 321.600 193.050 322.050 ;
        RECT 112.950 320.400 193.050 321.600 ;
        RECT 112.950 319.950 115.050 320.400 ;
        RECT 190.950 319.950 193.050 320.400 ;
        RECT 382.950 321.600 385.050 322.050 ;
        RECT 475.950 321.600 478.050 322.050 ;
        RECT 493.950 321.600 496.050 322.050 ;
        RECT 382.950 320.400 496.050 321.600 ;
        RECT 382.950 319.950 385.050 320.400 ;
        RECT 475.950 319.950 478.050 320.400 ;
        RECT 493.950 319.950 496.050 320.400 ;
        RECT 502.950 321.600 505.050 322.050 ;
        RECT 517.950 321.600 520.050 322.050 ;
        RECT 610.950 321.600 613.050 322.050 ;
        RECT 688.950 321.600 691.050 322.050 ;
        RECT 502.950 320.400 691.050 321.600 ;
        RECT 502.950 319.950 505.050 320.400 ;
        RECT 517.950 319.950 520.050 320.400 ;
        RECT 610.950 319.950 613.050 320.400 ;
        RECT 688.950 319.950 691.050 320.400 ;
        RECT 772.950 321.600 775.050 322.050 ;
        RECT 778.950 321.600 781.050 322.050 ;
        RECT 790.950 321.600 793.050 322.050 ;
        RECT 772.950 320.400 793.050 321.600 ;
        RECT 772.950 319.950 775.050 320.400 ;
        RECT 778.950 319.950 781.050 320.400 ;
        RECT 790.950 319.950 793.050 320.400 ;
        RECT 211.950 318.600 214.050 319.050 ;
        RECT 343.950 318.600 346.050 319.050 ;
        RECT 211.950 317.400 346.050 318.600 ;
        RECT 211.950 316.950 214.050 317.400 ;
        RECT 343.950 316.950 346.050 317.400 ;
        RECT 355.950 318.600 358.050 319.050 ;
        RECT 394.950 318.600 397.050 319.050 ;
        RECT 409.950 318.600 412.050 319.050 ;
        RECT 355.950 317.400 412.050 318.600 ;
        RECT 355.950 316.950 358.050 317.400 ;
        RECT 394.950 316.950 397.050 317.400 ;
        RECT 409.950 316.950 412.050 317.400 ;
        RECT 580.950 318.600 583.050 319.050 ;
        RECT 619.950 318.600 622.050 319.050 ;
        RECT 580.950 317.400 622.050 318.600 ;
        RECT 580.950 316.950 583.050 317.400 ;
        RECT 619.950 316.950 622.050 317.400 ;
        RECT 841.950 318.600 844.050 319.050 ;
        RECT 847.950 318.600 850.050 319.050 ;
        RECT 841.950 317.400 850.050 318.600 ;
        RECT 841.950 316.950 844.050 317.400 ;
        RECT 847.950 316.950 850.050 317.400 ;
        RECT 508.950 315.600 511.050 316.050 ;
        RECT 553.950 315.600 556.050 316.050 ;
        RECT 508.950 314.400 556.050 315.600 ;
        RECT 508.950 313.950 511.050 314.400 ;
        RECT 553.950 313.950 556.050 314.400 ;
        RECT 343.950 312.600 346.050 313.050 ;
        RECT 439.950 312.600 442.050 313.050 ;
        RECT 343.950 311.400 442.050 312.600 ;
        RECT 343.950 310.950 346.050 311.400 ;
        RECT 439.950 310.950 442.050 311.400 ;
        RECT 829.950 312.600 832.050 313.050 ;
        RECT 847.950 312.600 850.050 313.050 ;
        RECT 829.950 311.400 850.050 312.600 ;
        RECT 829.950 310.950 832.050 311.400 ;
        RECT 847.950 310.950 850.050 311.400 ;
        RECT 490.950 309.600 493.050 310.050 ;
        RECT 526.950 309.600 529.050 310.050 ;
        RECT 490.950 308.400 529.050 309.600 ;
        RECT 490.950 307.950 493.050 308.400 ;
        RECT 526.950 307.950 529.050 308.400 ;
        RECT 601.950 309.600 604.050 310.050 ;
        RECT 616.950 309.600 619.050 310.050 ;
        RECT 601.950 308.400 619.050 309.600 ;
        RECT 601.950 307.950 604.050 308.400 ;
        RECT 616.950 307.950 619.050 308.400 ;
        RECT 823.950 309.600 826.050 310.050 ;
        RECT 871.950 309.600 874.050 310.050 ;
        RECT 823.950 308.400 874.050 309.600 ;
        RECT 823.950 307.950 826.050 308.400 ;
        RECT 871.950 307.950 874.050 308.400 ;
        RECT 10.950 306.600 13.050 307.050 ;
        RECT 46.950 306.600 49.050 307.050 ;
        RECT 136.950 306.600 139.050 307.050 ;
        RECT 10.950 305.400 139.050 306.600 ;
        RECT 10.950 304.950 13.050 305.400 ;
        RECT 46.950 304.950 49.050 305.400 ;
        RECT 136.950 304.950 139.050 305.400 ;
        RECT 232.950 306.600 235.050 307.050 ;
        RECT 241.950 306.600 244.050 307.050 ;
        RECT 250.950 306.600 253.050 307.050 ;
        RECT 232.950 305.400 253.050 306.600 ;
        RECT 232.950 304.950 235.050 305.400 ;
        RECT 241.950 304.950 244.050 305.400 ;
        RECT 250.950 304.950 253.050 305.400 ;
        RECT 298.950 306.600 301.050 307.050 ;
        RECT 340.950 306.600 343.050 307.050 ;
        RECT 298.950 305.400 343.050 306.600 ;
        RECT 298.950 304.950 301.050 305.400 ;
        RECT 340.950 304.950 343.050 305.400 ;
        RECT 532.950 306.600 535.050 307.050 ;
        RECT 556.950 306.600 559.050 307.050 ;
        RECT 532.950 305.400 559.050 306.600 ;
        RECT 532.950 304.950 535.050 305.400 ;
        RECT 556.950 304.950 559.050 305.400 ;
        RECT 571.950 306.600 574.050 307.050 ;
        RECT 583.950 306.600 586.050 307.050 ;
        RECT 571.950 305.400 586.050 306.600 ;
        RECT 571.950 304.950 574.050 305.400 ;
        RECT 583.950 304.950 586.050 305.400 ;
        RECT 589.950 306.600 592.050 307.050 ;
        RECT 706.950 306.600 709.050 307.050 ;
        RECT 589.950 305.400 709.050 306.600 ;
        RECT 589.950 304.950 592.050 305.400 ;
        RECT 706.950 304.950 709.050 305.400 ;
        RECT 778.950 306.600 781.050 307.050 ;
        RECT 793.950 306.600 796.050 307.050 ;
        RECT 778.950 305.400 796.050 306.600 ;
        RECT 778.950 304.950 781.050 305.400 ;
        RECT 793.950 304.950 796.050 305.400 ;
        RECT 178.950 303.600 181.050 304.050 ;
        RECT 196.950 303.600 199.050 304.050 ;
        RECT 178.950 302.400 199.050 303.600 ;
        RECT 178.950 301.950 181.050 302.400 ;
        RECT 196.950 301.950 199.050 302.400 ;
        RECT 289.950 303.600 292.050 304.050 ;
        RECT 304.950 303.600 307.050 304.050 ;
        RECT 289.950 302.400 307.050 303.600 ;
        RECT 289.950 301.950 292.050 302.400 ;
        RECT 304.950 301.950 307.050 302.400 ;
        RECT 343.950 303.600 346.050 304.050 ;
        RECT 349.950 303.600 352.050 304.050 ;
        RECT 358.950 303.600 361.050 304.050 ;
        RECT 379.950 303.600 382.050 304.050 ;
        RECT 343.950 302.400 382.050 303.600 ;
        RECT 343.950 301.950 346.050 302.400 ;
        RECT 349.950 301.950 352.050 302.400 ;
        RECT 358.950 301.950 361.050 302.400 ;
        RECT 379.950 301.950 382.050 302.400 ;
        RECT 52.950 300.600 55.050 301.050 ;
        RECT 133.950 300.600 136.050 301.050 ;
        RECT 52.950 299.400 136.050 300.600 ;
        RECT 52.950 298.950 55.050 299.400 ;
        RECT 133.950 298.950 136.050 299.400 ;
        RECT 151.950 300.600 154.050 301.050 ;
        RECT 178.950 300.600 181.050 300.900 ;
        RECT 151.950 299.400 181.050 300.600 ;
        RECT 151.950 298.950 154.050 299.400 ;
        RECT 178.950 298.800 181.050 299.400 ;
        RECT 208.950 300.600 211.050 301.050 ;
        RECT 241.950 300.600 244.050 301.050 ;
        RECT 289.950 300.600 292.050 300.900 ;
        RECT 208.950 299.400 292.050 300.600 ;
        RECT 208.950 298.950 211.050 299.400 ;
        RECT 241.950 298.950 244.050 299.400 ;
        RECT 289.950 298.800 292.050 299.400 ;
        RECT 310.950 300.600 313.050 301.050 ;
        RECT 322.950 300.600 325.050 301.050 ;
        RECT 310.950 299.400 325.050 300.600 ;
        RECT 310.950 298.950 313.050 299.400 ;
        RECT 322.950 298.950 325.050 299.400 ;
        RECT 454.950 300.600 457.050 301.050 ;
        RECT 484.950 300.600 487.050 301.050 ;
        RECT 514.950 300.600 517.050 301.050 ;
        RECT 454.950 299.400 517.050 300.600 ;
        RECT 454.950 298.950 457.050 299.400 ;
        RECT 484.950 298.950 487.050 299.400 ;
        RECT 514.950 298.950 517.050 299.400 ;
        RECT 520.950 300.600 523.050 301.050 ;
        RECT 550.950 300.600 553.050 301.050 ;
        RECT 520.950 299.400 553.050 300.600 ;
        RECT 520.950 298.950 523.050 299.400 ;
        RECT 550.950 298.950 553.050 299.400 ;
        RECT 559.950 300.600 562.050 301.050 ;
        RECT 637.950 300.600 640.050 301.050 ;
        RECT 559.950 299.400 640.050 300.600 ;
        RECT 559.950 298.950 562.050 299.400 ;
        RECT 637.950 298.950 640.050 299.400 ;
        RECT 664.950 300.600 667.050 301.050 ;
        RECT 673.950 300.600 676.050 301.050 ;
        RECT 664.950 299.400 676.050 300.600 ;
        RECT 664.950 298.950 667.050 299.400 ;
        RECT 673.950 298.950 676.050 299.400 ;
        RECT 769.950 300.600 772.050 301.050 ;
        RECT 784.950 300.600 787.050 301.050 ;
        RECT 769.950 299.400 787.050 300.600 ;
        RECT 769.950 298.950 772.050 299.400 ;
        RECT 784.950 298.950 787.050 299.400 ;
        RECT 856.800 298.950 858.900 301.050 ;
        RECT 253.950 297.600 256.050 298.050 ;
        RECT 262.950 297.600 265.050 298.050 ;
        RECT 253.950 296.400 265.050 297.600 ;
        RECT 253.950 295.950 256.050 296.400 ;
        RECT 262.950 295.950 265.050 296.400 ;
        RECT 331.950 297.600 334.050 298.050 ;
        RECT 355.950 297.600 358.050 298.050 ;
        RECT 373.950 297.600 376.050 298.050 ;
        RECT 331.950 296.400 376.050 297.600 ;
        RECT 331.950 295.950 334.050 296.400 ;
        RECT 355.950 295.950 358.050 296.400 ;
        RECT 373.950 295.950 376.050 296.400 ;
        RECT 463.950 297.600 466.050 298.050 ;
        RECT 469.950 297.600 472.050 297.900 ;
        RECT 463.950 296.400 472.050 297.600 ;
        RECT 463.950 295.950 466.050 296.400 ;
        RECT 469.950 295.800 472.050 296.400 ;
        RECT 487.950 297.600 490.050 298.050 ;
        RECT 538.950 297.600 541.050 298.050 ;
        RECT 544.950 297.600 547.050 298.050 ;
        RECT 487.950 296.400 547.050 297.600 ;
        RECT 487.950 295.950 490.050 296.400 ;
        RECT 538.950 295.950 541.050 296.400 ;
        RECT 544.950 295.950 547.050 296.400 ;
        RECT 676.950 297.600 679.050 298.050 ;
        RECT 685.950 297.600 688.050 298.050 ;
        RECT 676.950 296.400 688.050 297.600 ;
        RECT 676.950 295.950 679.050 296.400 ;
        RECT 685.950 295.950 688.050 296.400 ;
        RECT 796.950 297.600 799.050 298.050 ;
        RECT 802.950 297.600 805.050 298.050 ;
        RECT 796.950 296.400 805.050 297.600 ;
        RECT 796.950 295.950 799.050 296.400 ;
        RECT 802.950 295.950 805.050 296.400 ;
        RECT 811.950 297.600 814.050 298.050 ;
        RECT 829.950 297.600 832.050 298.050 ;
        RECT 811.950 296.400 832.050 297.600 ;
        RECT 811.950 295.950 814.050 296.400 ;
        RECT 829.950 295.950 832.050 296.400 ;
        RECT 857.250 297.600 858.450 298.950 ;
        RECT 874.950 297.600 877.050 298.050 ;
        RECT 857.250 296.400 877.050 297.600 ;
        RECT 28.950 294.600 31.050 295.200 ;
        RECT 52.950 294.600 55.050 295.200 ;
        RECT 28.950 293.400 55.050 294.600 ;
        RECT 28.950 293.100 31.050 293.400 ;
        RECT 52.950 293.100 55.050 293.400 ;
        RECT 70.950 294.750 73.050 295.200 ;
        RECT 76.950 294.750 79.050 295.200 ;
        RECT 70.950 293.550 79.050 294.750 ;
        RECT 70.950 293.100 73.050 293.550 ;
        RECT 76.950 293.100 79.050 293.550 ;
        RECT 94.950 294.750 97.050 295.200 ;
        RECT 103.950 294.750 106.050 295.200 ;
        RECT 94.950 293.550 106.050 294.750 ;
        RECT 109.950 294.600 112.050 295.200 ;
        RECT 151.950 294.600 154.050 295.200 ;
        RECT 94.950 293.100 97.050 293.550 ;
        RECT 103.950 293.100 106.050 293.550 ;
        RECT 107.400 293.400 154.050 294.600 ;
        RECT 97.950 291.600 100.050 292.050 ;
        RECT 107.400 291.600 108.600 293.400 ;
        RECT 109.950 293.100 112.050 293.400 ;
        RECT 151.950 293.100 154.050 293.400 ;
        RECT 172.950 293.100 175.050 295.200 ;
        RECT 202.950 294.750 205.050 295.200 ;
        RECT 208.950 294.750 211.050 295.200 ;
        RECT 202.950 294.600 211.050 294.750 ;
        RECT 179.400 293.550 211.050 294.600 ;
        RECT 179.400 293.400 205.050 293.550 ;
        RECT 97.950 290.400 108.600 291.600 ;
        RECT 163.950 291.600 166.050 292.050 ;
        RECT 173.400 291.600 174.600 293.100 ;
        RECT 179.400 291.600 180.600 293.400 ;
        RECT 202.950 293.100 205.050 293.400 ;
        RECT 208.950 293.100 211.050 293.550 ;
        RECT 277.950 294.750 280.050 295.200 ;
        RECT 283.950 294.750 286.050 295.200 ;
        RECT 277.950 293.550 286.050 294.750 ;
        RECT 277.950 293.100 280.050 293.550 ;
        RECT 283.950 293.100 286.050 293.550 ;
        RECT 313.950 294.600 316.050 295.200 ;
        RECT 340.950 294.600 343.050 295.050 ;
        RECT 409.950 294.750 412.050 295.200 ;
        RECT 418.950 294.750 421.050 295.200 ;
        RECT 313.950 293.400 354.600 294.600 ;
        RECT 313.950 293.100 316.050 293.400 ;
        RECT 340.950 292.950 343.050 293.400 ;
        RECT 163.950 290.400 180.600 291.600 ;
        RECT 353.400 291.600 354.600 293.400 ;
        RECT 409.950 293.550 421.050 294.750 ;
        RECT 409.950 293.100 412.050 293.550 ;
        RECT 418.950 293.100 421.050 293.550 ;
        RECT 463.950 294.600 466.050 294.900 ;
        RECT 481.950 294.600 484.050 295.050 ;
        RECT 463.950 293.400 484.050 294.600 ;
        RECT 463.950 292.800 466.050 293.400 ;
        RECT 481.950 292.950 484.050 293.400 ;
        RECT 496.950 293.100 499.050 295.200 ;
        RECT 508.950 294.750 511.050 295.200 ;
        RECT 520.950 294.750 523.050 295.200 ;
        RECT 508.950 293.550 523.050 294.750 ;
        RECT 508.950 293.100 511.050 293.550 ;
        RECT 520.950 293.100 523.050 293.550 ;
        RECT 547.950 293.100 550.050 295.200 ;
        RECT 592.950 294.600 595.050 295.200 ;
        RECT 664.950 294.600 667.050 295.200 ;
        RECT 669.000 294.600 673.050 295.050 ;
        RECT 587.400 293.400 595.050 294.600 ;
        RECT 353.400 290.400 372.600 291.600 ;
        RECT 97.950 289.950 100.050 290.400 ;
        RECT 163.950 289.950 166.050 290.400 ;
        RECT 58.950 288.450 61.050 288.900 ;
        RECT 67.950 288.450 70.050 288.900 ;
        RECT 58.950 287.250 70.050 288.450 ;
        RECT 58.950 286.800 61.050 287.250 ;
        RECT 67.950 286.800 70.050 287.250 ;
        RECT 106.950 288.600 109.050 288.900 ;
        RECT 121.950 288.600 124.050 289.050 ;
        RECT 106.950 287.400 124.050 288.600 ;
        RECT 106.950 286.800 109.050 287.400 ;
        RECT 121.950 286.950 124.050 287.400 ;
        RECT 169.950 288.450 172.050 288.900 ;
        RECT 187.950 288.450 190.050 288.900 ;
        RECT 169.950 287.250 190.050 288.450 ;
        RECT 169.950 286.800 172.050 287.250 ;
        RECT 187.950 286.800 190.050 287.250 ;
        RECT 250.950 288.450 253.050 288.900 ;
        RECT 259.950 288.450 262.050 288.900 ;
        RECT 250.950 287.250 262.050 288.450 ;
        RECT 250.950 286.800 253.050 287.250 ;
        RECT 259.950 286.800 262.050 287.250 ;
        RECT 265.950 288.450 268.050 288.900 ;
        RECT 271.950 288.450 274.050 288.900 ;
        RECT 265.950 287.250 274.050 288.450 ;
        RECT 265.950 286.800 268.050 287.250 ;
        RECT 271.950 286.800 274.050 287.250 ;
        RECT 304.950 288.450 307.050 288.900 ;
        RECT 307.950 288.450 310.050 289.050 ;
        RECT 310.950 288.450 313.050 288.900 ;
        RECT 304.950 287.250 313.050 288.450 ;
        RECT 304.950 286.800 307.050 287.250 ;
        RECT 307.950 286.950 310.050 287.250 ;
        RECT 310.950 286.800 313.050 287.250 ;
        RECT 322.950 288.450 325.050 288.900 ;
        RECT 328.950 288.450 331.050 288.900 ;
        RECT 322.950 287.250 331.050 288.450 ;
        RECT 371.400 288.600 372.600 290.400 ;
        RECT 376.950 288.600 379.050 288.900 ;
        RECT 371.400 287.400 379.050 288.600 ;
        RECT 322.950 286.800 325.050 287.250 ;
        RECT 328.950 286.800 331.050 287.250 ;
        RECT 376.950 286.800 379.050 287.400 ;
        RECT 394.950 288.450 397.050 288.900 ;
        RECT 400.950 288.600 403.050 288.900 ;
        RECT 424.950 288.600 427.050 288.900 ;
        RECT 400.950 288.450 427.050 288.600 ;
        RECT 394.950 287.400 427.050 288.450 ;
        RECT 394.950 287.250 403.050 287.400 ;
        RECT 394.950 286.800 397.050 287.250 ;
        RECT 400.950 286.800 403.050 287.250 ;
        RECT 424.950 286.800 427.050 287.400 ;
        RECT 497.400 286.050 498.600 293.100 ;
        RECT 499.950 288.600 502.050 288.900 ;
        RECT 508.950 288.600 511.050 289.050 ;
        RECT 499.950 287.400 511.050 288.600 ;
        RECT 499.950 286.800 502.050 287.400 ;
        RECT 508.950 286.950 511.050 287.400 ;
        RECT 514.950 288.450 517.050 288.900 ;
        RECT 529.950 288.600 532.050 288.900 ;
        RECT 548.400 288.600 549.600 293.100 ;
        RECT 587.400 291.600 588.600 293.400 ;
        RECT 592.950 293.100 595.050 293.400 ;
        RECT 659.400 293.400 667.050 294.600 ;
        RECT 572.400 290.400 588.600 291.600 ;
        RECT 529.950 288.450 549.600 288.600 ;
        RECT 514.950 287.400 549.600 288.450 ;
        RECT 550.950 288.600 553.050 288.900 ;
        RECT 556.950 288.600 559.050 289.050 ;
        RECT 572.400 288.900 573.600 290.400 ;
        RECT 550.950 287.400 559.050 288.600 ;
        RECT 514.950 287.250 532.050 287.400 ;
        RECT 514.950 286.800 517.050 287.250 ;
        RECT 529.950 286.800 532.050 287.250 ;
        RECT 550.950 286.800 553.050 287.400 ;
        RECT 556.950 286.950 559.050 287.400 ;
        RECT 571.950 286.800 574.050 288.900 ;
        RECT 586.950 288.450 589.050 288.900 ;
        RECT 595.950 288.450 598.050 288.900 ;
        RECT 586.950 287.250 598.050 288.450 ;
        RECT 586.950 286.800 589.050 287.250 ;
        RECT 595.950 286.800 598.050 287.250 ;
        RECT 616.950 288.450 619.050 288.900 ;
        RECT 622.950 288.450 625.050 288.900 ;
        RECT 616.950 287.250 625.050 288.450 ;
        RECT 616.950 286.800 619.050 287.250 ;
        RECT 622.950 286.800 625.050 287.250 ;
        RECT 634.950 288.600 637.050 289.050 ;
        RECT 640.950 288.600 643.050 288.900 ;
        RECT 659.400 288.600 660.600 293.400 ;
        RECT 664.950 293.100 667.050 293.400 ;
        RECT 668.400 292.950 673.050 294.600 ;
        RECT 697.950 294.750 700.050 295.200 ;
        RECT 712.950 294.750 715.050 295.200 ;
        RECT 697.950 293.550 715.050 294.750 ;
        RECT 697.950 293.100 700.050 293.550 ;
        RECT 712.950 293.100 715.050 293.550 ;
        RECT 724.950 294.750 727.050 295.200 ;
        RECT 733.950 294.750 736.050 295.200 ;
        RECT 724.950 293.550 736.050 294.750 ;
        RECT 724.950 293.100 727.050 293.550 ;
        RECT 733.950 293.100 736.050 293.550 ;
        RECT 739.950 293.100 742.050 295.200 ;
        RECT 757.950 293.100 760.050 295.200 ;
        RECT 763.950 294.600 766.050 295.200 ;
        RECT 784.950 294.600 787.050 295.200 ;
        RECT 763.950 293.400 787.050 294.600 ;
        RECT 763.950 293.100 766.050 293.400 ;
        RECT 784.950 293.100 787.050 293.400 ;
        RECT 805.950 294.750 808.050 295.200 ;
        RECT 820.950 294.750 823.050 295.200 ;
        RECT 805.950 293.550 823.050 294.750 ;
        RECT 805.950 293.100 808.050 293.550 ;
        RECT 820.950 293.100 823.050 293.550 ;
        RECT 857.250 294.600 858.450 296.400 ;
        RECT 874.950 295.950 877.050 296.400 ;
        RECT 857.250 293.400 861.600 294.600 ;
        RECT 668.400 291.600 669.600 292.950 ;
        RECT 662.400 290.400 669.600 291.600 ;
        RECT 662.400 288.900 663.600 290.400 ;
        RECT 740.400 289.050 741.600 293.100 ;
        RECT 748.950 291.600 751.050 292.050 ;
        RECT 758.400 291.600 759.600 293.100 ;
        RECT 748.950 290.400 759.600 291.600 ;
        RECT 785.400 291.600 786.600 293.100 ;
        RECT 841.950 291.600 844.050 292.050 ;
        RECT 785.400 290.400 792.600 291.600 ;
        RECT 748.950 289.950 751.050 290.400 ;
        RECT 634.950 287.400 660.600 288.600 ;
        RECT 634.950 286.950 637.050 287.400 ;
        RECT 640.950 286.800 643.050 287.400 ;
        RECT 661.950 286.800 664.050 288.900 ;
        RECT 691.950 288.600 694.050 288.900 ;
        RECT 697.950 288.600 700.050 289.050 ;
        RECT 691.950 287.400 700.050 288.600 ;
        RECT 740.400 287.400 745.050 289.050 ;
        RECT 691.950 286.800 694.050 287.400 ;
        RECT 697.950 286.950 700.050 287.400 ;
        RECT 741.000 286.950 745.050 287.400 ;
        RECT 769.950 288.600 772.050 289.050 ;
        RECT 787.950 288.600 790.050 288.900 ;
        RECT 769.950 287.400 790.050 288.600 ;
        RECT 791.400 288.600 792.600 290.400 ;
        RECT 812.400 290.400 844.050 291.600 ;
        RECT 860.400 291.600 861.600 293.400 ;
        RECT 865.950 291.600 868.050 295.050 ;
        RECT 860.400 290.400 864.600 291.600 ;
        RECT 865.950 291.000 870.600 291.600 ;
        RECT 866.400 290.400 870.600 291.000 ;
        RECT 802.950 288.600 805.050 288.900 ;
        RECT 791.400 287.400 805.050 288.600 ;
        RECT 769.950 286.950 772.050 287.400 ;
        RECT 787.950 286.800 790.050 287.400 ;
        RECT 802.950 286.800 805.050 287.400 ;
        RECT 808.950 288.600 811.050 288.900 ;
        RECT 812.400 288.600 813.600 290.400 ;
        RECT 841.950 289.950 844.050 290.400 ;
        RECT 863.400 288.900 864.600 290.400 ;
        RECT 808.950 287.400 813.600 288.600 ;
        RECT 808.950 286.800 811.050 287.400 ;
        RECT 862.950 286.800 865.050 288.900 ;
        RECT 869.400 288.600 870.600 290.400 ;
        RECT 877.950 288.600 880.050 288.900 ;
        RECT 869.400 287.400 880.050 288.600 ;
        RECT 877.950 286.800 880.050 287.400 ;
        RECT 292.950 285.600 295.050 286.050 ;
        RECT 298.950 285.600 301.050 286.050 ;
        RECT 292.950 284.400 301.050 285.600 ;
        RECT 292.950 283.950 295.050 284.400 ;
        RECT 298.950 283.950 301.050 284.400 ;
        RECT 340.950 285.600 343.050 286.050 ;
        RECT 352.950 285.600 355.050 286.050 ;
        RECT 340.950 284.400 355.050 285.600 ;
        RECT 340.950 283.950 343.050 284.400 ;
        RECT 352.950 283.950 355.050 284.400 ;
        RECT 472.950 285.600 475.050 286.050 ;
        RECT 487.950 285.600 490.050 286.050 ;
        RECT 472.950 284.400 490.050 285.600 ;
        RECT 472.950 283.950 475.050 284.400 ;
        RECT 487.950 283.950 490.050 284.400 ;
        RECT 496.950 283.950 499.050 286.050 ;
        RECT 538.950 285.600 541.050 286.050 ;
        RECT 580.950 285.600 583.050 286.050 ;
        RECT 538.950 284.400 583.050 285.600 ;
        RECT 538.950 283.950 541.050 284.400 ;
        RECT 580.950 283.950 583.050 284.400 ;
        RECT 151.950 282.600 154.050 283.050 ;
        RECT 211.950 282.600 214.050 283.050 ;
        RECT 151.950 281.400 214.050 282.600 ;
        RECT 151.950 280.950 154.050 281.400 ;
        RECT 211.950 280.950 214.050 281.400 ;
        RECT 523.950 282.600 526.050 283.050 ;
        RECT 535.950 282.600 538.050 283.050 ;
        RECT 523.950 281.400 538.050 282.600 ;
        RECT 523.950 280.950 526.050 281.400 ;
        RECT 535.950 280.950 538.050 281.400 ;
        RECT 547.950 282.600 550.050 283.050 ;
        RECT 571.950 282.600 574.050 283.050 ;
        RECT 547.950 281.400 574.050 282.600 ;
        RECT 547.950 280.950 550.050 281.400 ;
        RECT 571.950 280.950 574.050 281.400 ;
        RECT 130.950 279.600 133.050 280.050 ;
        RECT 199.950 279.600 202.050 280.050 ;
        RECT 130.950 278.400 202.050 279.600 ;
        RECT 130.950 277.950 133.050 278.400 ;
        RECT 199.950 277.950 202.050 278.400 ;
        RECT 214.950 279.600 217.050 280.050 ;
        RECT 220.950 279.600 223.050 280.050 ;
        RECT 214.950 278.400 223.050 279.600 ;
        RECT 214.950 277.950 217.050 278.400 ;
        RECT 220.950 277.950 223.050 278.400 ;
        RECT 358.950 279.600 361.050 280.050 ;
        RECT 373.950 279.600 376.050 280.050 ;
        RECT 358.950 278.400 376.050 279.600 ;
        RECT 358.950 277.950 361.050 278.400 ;
        RECT 373.950 277.950 376.050 278.400 ;
        RECT 571.950 279.600 574.050 279.900 ;
        RECT 601.950 279.600 604.050 280.050 ;
        RECT 571.950 278.400 604.050 279.600 ;
        RECT 571.950 277.800 574.050 278.400 ;
        RECT 601.950 277.950 604.050 278.400 ;
        RECT 667.950 279.600 670.050 280.050 ;
        RECT 709.950 279.600 712.050 280.050 ;
        RECT 667.950 278.400 712.050 279.600 ;
        RECT 667.950 277.950 670.050 278.400 ;
        RECT 709.950 277.950 712.050 278.400 ;
        RECT 736.950 279.600 739.050 280.050 ;
        RECT 748.950 279.600 751.050 280.050 ;
        RECT 736.950 278.400 751.050 279.600 ;
        RECT 736.950 277.950 739.050 278.400 ;
        RECT 748.950 277.950 751.050 278.400 ;
        RECT 760.950 279.600 763.050 280.050 ;
        RECT 793.950 279.600 796.050 280.050 ;
        RECT 829.950 279.600 832.050 280.050 ;
        RECT 760.950 278.400 832.050 279.600 ;
        RECT 760.950 277.950 763.050 278.400 ;
        RECT 793.950 277.950 796.050 278.400 ;
        RECT 829.950 277.950 832.050 278.400 ;
        RECT 166.950 276.600 169.050 277.050 ;
        RECT 172.950 276.600 175.050 277.050 ;
        RECT 166.950 275.400 175.050 276.600 ;
        RECT 166.950 274.950 169.050 275.400 ;
        RECT 172.950 274.950 175.050 275.400 ;
        RECT 253.950 276.600 256.050 277.050 ;
        RECT 277.950 276.600 280.050 277.050 ;
        RECT 301.950 276.600 304.050 277.050 ;
        RECT 253.950 275.400 304.050 276.600 ;
        RECT 253.950 274.950 256.050 275.400 ;
        RECT 277.950 274.950 280.050 275.400 ;
        RECT 301.950 274.950 304.050 275.400 ;
        RECT 475.950 276.600 478.050 277.050 ;
        RECT 493.950 276.600 496.050 277.050 ;
        RECT 475.950 275.400 496.050 276.600 ;
        RECT 475.950 274.950 478.050 275.400 ;
        RECT 493.950 274.950 496.050 275.400 ;
        RECT 541.950 276.600 544.050 277.050 ;
        RECT 565.950 276.600 568.050 277.050 ;
        RECT 634.950 276.600 637.050 277.050 ;
        RECT 541.950 275.400 637.050 276.600 ;
        RECT 541.950 274.950 544.050 275.400 ;
        RECT 565.950 274.950 568.050 275.400 ;
        RECT 634.950 274.950 637.050 275.400 ;
        RECT 715.950 276.600 718.050 277.050 ;
        RECT 727.950 276.600 730.050 276.900 ;
        RECT 751.950 276.600 754.050 277.050 ;
        RECT 715.950 275.400 754.050 276.600 ;
        RECT 715.950 274.950 718.050 275.400 ;
        RECT 727.950 274.800 730.050 275.400 ;
        RECT 751.950 274.950 754.050 275.400 ;
        RECT 772.950 276.600 775.050 277.050 ;
        RECT 787.950 276.600 790.050 277.050 ;
        RECT 772.950 275.400 790.050 276.600 ;
        RECT 772.950 274.950 775.050 275.400 ;
        RECT 787.950 274.950 790.050 275.400 ;
        RECT 853.950 276.600 856.050 277.050 ;
        RECT 898.950 276.600 901.050 277.050 ;
        RECT 853.950 275.400 901.050 276.600 ;
        RECT 853.950 274.950 856.050 275.400 ;
        RECT 898.950 274.950 901.050 275.400 ;
        RECT 22.950 273.600 25.050 274.050 ;
        RECT 34.950 273.600 37.050 274.050 ;
        RECT 22.950 272.400 37.050 273.600 ;
        RECT 22.950 271.950 25.050 272.400 ;
        RECT 34.950 271.950 37.050 272.400 ;
        RECT 142.950 273.600 145.050 274.050 ;
        RECT 154.950 273.600 157.050 274.050 ;
        RECT 142.950 272.400 157.050 273.600 ;
        RECT 142.950 271.950 145.050 272.400 ;
        RECT 154.950 271.950 157.050 272.400 ;
        RECT 190.950 273.600 193.050 274.050 ;
        RECT 199.950 273.600 202.050 274.050 ;
        RECT 214.950 273.600 217.050 274.050 ;
        RECT 190.950 272.400 217.050 273.600 ;
        RECT 190.950 271.950 193.050 272.400 ;
        RECT 199.950 271.950 202.050 272.400 ;
        RECT 214.950 271.950 217.050 272.400 ;
        RECT 478.950 273.600 481.050 274.050 ;
        RECT 487.950 273.600 490.050 274.050 ;
        RECT 478.950 272.400 490.050 273.600 ;
        RECT 478.950 271.950 481.050 272.400 ;
        RECT 487.950 271.950 490.050 272.400 ;
        RECT 106.950 270.600 109.050 271.050 ;
        RECT 115.950 270.600 118.050 271.050 ;
        RECT 106.950 269.400 118.050 270.600 ;
        RECT 106.950 268.950 109.050 269.400 ;
        RECT 115.950 268.950 118.050 269.400 ;
        RECT 205.950 270.600 208.050 271.050 ;
        RECT 241.950 270.600 244.050 271.050 ;
        RECT 472.950 270.600 475.050 271.050 ;
        RECT 493.950 270.600 496.050 271.050 ;
        RECT 205.950 269.400 496.050 270.600 ;
        RECT 205.950 268.950 208.050 269.400 ;
        RECT 241.950 268.950 244.050 269.400 ;
        RECT 472.950 268.950 475.050 269.400 ;
        RECT 493.950 268.950 496.050 269.400 ;
        RECT 577.950 270.600 580.050 271.050 ;
        RECT 718.950 270.600 721.050 271.050 ;
        RECT 742.950 270.600 745.050 271.050 ;
        RECT 577.950 269.400 745.050 270.600 ;
        RECT 577.950 268.950 580.050 269.400 ;
        RECT 718.950 268.950 721.050 269.400 ;
        RECT 742.950 268.950 745.050 269.400 ;
        RECT 799.950 270.600 802.050 271.050 ;
        RECT 850.950 270.600 853.050 271.050 ;
        RECT 799.950 269.400 853.050 270.600 ;
        RECT 799.950 268.950 802.050 269.400 ;
        RECT 850.950 268.950 853.050 269.400 ;
        RECT 19.950 267.600 22.050 268.050 ;
        RECT 28.950 267.600 31.050 268.050 ;
        RECT 19.950 266.400 31.050 267.600 ;
        RECT 19.950 265.950 22.050 266.400 ;
        RECT 28.950 265.950 31.050 266.400 ;
        RECT 52.950 267.600 55.050 268.050 ;
        RECT 58.950 267.600 61.050 268.050 ;
        RECT 94.950 267.600 97.050 268.050 ;
        RECT 52.950 266.400 97.050 267.600 ;
        RECT 52.950 265.950 55.050 266.400 ;
        RECT 58.950 265.950 61.050 266.400 ;
        RECT 94.950 265.950 97.050 266.400 ;
        RECT 187.950 267.600 190.050 268.050 ;
        RECT 202.950 267.600 205.050 268.050 ;
        RECT 187.950 266.400 205.050 267.600 ;
        RECT 187.950 265.950 190.050 266.400 ;
        RECT 202.950 265.950 205.050 266.400 ;
        RECT 208.950 267.600 211.050 268.050 ;
        RECT 232.950 267.600 235.050 268.050 ;
        RECT 208.950 266.400 235.050 267.600 ;
        RECT 208.950 265.950 211.050 266.400 ;
        RECT 232.950 265.950 235.050 266.400 ;
        RECT 382.950 267.600 385.050 268.050 ;
        RECT 397.950 267.600 400.050 268.050 ;
        RECT 382.950 266.400 400.050 267.600 ;
        RECT 382.950 265.950 385.050 266.400 ;
        RECT 397.950 265.950 400.050 266.400 ;
        RECT 454.950 267.600 457.050 268.050 ;
        RECT 466.950 267.600 469.050 268.050 ;
        RECT 454.950 266.400 469.050 267.600 ;
        RECT 454.950 265.950 457.050 266.400 ;
        RECT 466.950 265.950 469.050 266.400 ;
        RECT 664.950 267.600 667.050 268.050 ;
        RECT 673.800 267.600 675.900 268.050 ;
        RECT 664.950 266.400 675.900 267.600 ;
        RECT 664.950 265.950 667.050 266.400 ;
        RECT 673.800 265.950 675.900 266.400 ;
        RECT 676.950 267.600 679.050 268.050 ;
        RECT 688.950 267.600 691.050 268.050 ;
        RECT 676.950 266.400 691.050 267.600 ;
        RECT 676.950 265.950 679.050 266.400 ;
        RECT 688.950 265.950 691.050 266.400 ;
        RECT 748.950 267.600 751.050 268.050 ;
        RECT 781.950 267.600 784.050 268.050 ;
        RECT 820.950 267.600 823.050 268.050 ;
        RECT 748.950 266.400 823.050 267.600 ;
        RECT 748.950 265.950 751.050 266.400 ;
        RECT 781.950 265.950 784.050 266.400 ;
        RECT 820.950 265.950 823.050 266.400 ;
        RECT 877.950 267.600 880.050 268.050 ;
        RECT 889.950 267.600 892.050 268.050 ;
        RECT 877.950 266.400 892.050 267.600 ;
        RECT 877.950 265.950 880.050 266.400 ;
        RECT 889.950 265.950 892.050 266.400 ;
        RECT 31.950 264.600 34.050 265.050 ;
        RECT 40.950 264.600 43.050 265.050 ;
        RECT 97.950 264.600 100.050 265.050 ;
        RECT 31.950 263.400 100.050 264.600 ;
        RECT 31.950 262.950 34.050 263.400 ;
        RECT 40.950 262.950 43.050 263.400 ;
        RECT 97.950 262.950 100.050 263.400 ;
        RECT 286.950 264.600 289.050 264.900 ;
        RECT 322.950 264.600 325.050 265.050 ;
        RECT 286.950 263.400 325.050 264.600 ;
        RECT 286.950 262.800 289.050 263.400 ;
        RECT 322.950 262.950 325.050 263.400 ;
        RECT 442.950 264.600 445.050 265.050 ;
        RECT 448.950 264.600 451.050 265.050 ;
        RECT 469.950 264.600 472.050 265.050 ;
        RECT 484.950 264.600 487.050 265.050 ;
        RECT 490.950 264.600 493.050 264.900 ;
        RECT 442.950 263.400 465.600 264.600 ;
        RECT 442.950 262.950 445.050 263.400 ;
        RECT 448.950 262.950 451.050 263.400 ;
        RECT 64.950 260.100 67.050 262.200 ;
        RECT 112.950 261.600 115.050 262.200 ;
        RECT 193.950 261.600 196.050 262.200 ;
        RECT 208.950 261.600 211.050 262.200 ;
        RECT 112.950 260.400 117.600 261.600 ;
        RECT 112.950 260.100 115.050 260.400 ;
        RECT 25.950 255.450 28.050 255.900 ;
        RECT 31.950 255.450 34.050 256.050 ;
        RECT 25.950 254.250 34.050 255.450 ;
        RECT 25.950 253.800 28.050 254.250 ;
        RECT 31.950 253.950 34.050 254.250 ;
        RECT 43.950 255.600 46.050 255.900 ;
        RECT 61.950 255.600 64.050 255.900 ;
        RECT 43.950 254.400 64.050 255.600 ;
        RECT 43.950 253.800 46.050 254.400 ;
        RECT 61.950 253.800 64.050 254.400 ;
        RECT 65.400 253.050 66.600 260.100 ;
        RECT 97.950 258.600 100.050 259.050 ;
        RECT 97.950 257.400 111.600 258.600 ;
        RECT 97.950 256.950 100.050 257.400 ;
        RECT 70.950 255.600 73.050 256.050 ;
        RECT 110.400 255.900 111.600 257.400 ;
        RECT 116.400 256.050 117.600 260.400 ;
        RECT 193.950 260.400 211.050 261.600 ;
        RECT 193.950 260.100 196.050 260.400 ;
        RECT 208.950 260.100 211.050 260.400 ;
        RECT 232.950 260.100 235.050 262.200 ;
        RECT 292.950 261.600 295.050 262.050 ;
        RECT 307.950 261.600 310.050 262.200 ;
        RECT 292.950 260.400 310.050 261.600 ;
        RECT 233.400 258.600 234.600 260.100 ;
        RECT 292.950 259.950 295.050 260.400 ;
        RECT 307.950 260.100 310.050 260.400 ;
        RECT 313.950 261.600 316.050 262.200 ;
        RECT 337.950 261.600 340.050 262.200 ;
        RECT 346.950 261.600 349.050 262.050 ;
        RECT 313.950 260.400 324.600 261.600 ;
        RECT 313.950 260.100 316.050 260.400 ;
        RECT 218.400 257.400 234.600 258.600 ;
        RECT 323.400 259.050 324.600 260.400 ;
        RECT 337.950 260.400 349.050 261.600 ;
        RECT 337.950 260.100 340.050 260.400 ;
        RECT 346.950 259.950 349.050 260.400 ;
        RECT 376.950 261.750 379.050 262.200 ;
        RECT 385.950 261.750 388.050 262.200 ;
        RECT 376.950 260.550 388.050 261.750 ;
        RECT 376.950 260.100 379.050 260.550 ;
        RECT 385.950 260.100 388.050 260.550 ;
        RECT 391.950 261.600 394.050 262.200 ;
        RECT 400.950 261.600 403.050 262.050 ;
        RECT 391.950 260.400 403.050 261.600 ;
        RECT 391.950 260.100 394.050 260.400 ;
        RECT 400.950 259.950 403.050 260.400 ;
        RECT 406.950 261.600 409.050 262.200 ;
        RECT 418.950 261.600 421.050 262.050 ;
        RECT 406.950 260.400 421.050 261.600 ;
        RECT 406.950 260.100 409.050 260.400 ;
        RECT 418.950 259.950 421.050 260.400 ;
        RECT 460.950 260.100 463.050 262.200 ;
        RECT 464.400 261.600 465.600 263.400 ;
        RECT 469.950 263.400 480.600 264.600 ;
        RECT 469.950 262.950 472.050 263.400 ;
        RECT 475.950 261.600 478.050 262.200 ;
        RECT 464.400 260.400 478.050 261.600 ;
        RECT 479.400 261.600 480.600 263.400 ;
        RECT 484.950 263.400 493.050 264.600 ;
        RECT 484.950 262.950 487.050 263.400 ;
        RECT 490.950 262.800 493.050 263.400 ;
        RECT 505.950 264.600 508.050 265.050 ;
        RECT 529.950 264.600 532.050 265.050 ;
        RECT 505.950 263.400 532.050 264.600 ;
        RECT 505.950 262.950 508.050 263.400 ;
        RECT 529.950 262.950 532.050 263.400 ;
        RECT 589.950 264.600 592.050 265.050 ;
        RECT 646.950 264.600 649.050 265.050 ;
        RECT 589.950 263.400 649.050 264.600 ;
        RECT 589.950 262.950 592.050 263.400 ;
        RECT 646.950 262.950 649.050 263.400 ;
        RECT 784.950 264.600 787.050 265.050 ;
        RECT 805.950 264.600 808.050 265.050 ;
        RECT 856.950 264.600 859.050 265.050 ;
        RECT 784.950 263.400 816.600 264.600 ;
        RECT 784.950 262.950 787.050 263.400 ;
        RECT 805.950 262.950 808.050 263.400 ;
        RECT 481.950 261.600 484.050 262.200 ;
        RECT 479.400 260.400 484.050 261.600 ;
        RECT 475.950 260.100 478.050 260.400 ;
        RECT 481.950 260.100 484.050 260.400 ;
        RECT 499.950 261.750 502.050 262.200 ;
        RECT 517.950 261.750 520.050 262.200 ;
        RECT 499.950 260.550 520.050 261.750 ;
        RECT 499.950 260.100 502.050 260.550 ;
        RECT 517.950 260.100 520.050 260.550 ;
        RECT 538.950 261.600 541.050 262.050 ;
        RECT 547.950 261.600 550.050 262.200 ;
        RECT 538.950 260.400 550.050 261.600 ;
        RECT 323.400 257.400 328.050 259.050 ;
        RECT 461.400 258.600 462.600 260.100 ;
        RECT 538.950 259.950 541.050 260.400 ;
        RECT 547.950 260.100 550.050 260.400 ;
        RECT 577.950 261.600 580.050 262.050 ;
        RECT 583.950 261.600 586.050 262.050 ;
        RECT 577.950 260.400 586.050 261.600 ;
        RECT 577.950 259.950 580.050 260.400 ;
        RECT 583.950 259.950 586.050 260.400 ;
        RECT 613.950 261.600 616.050 262.200 ;
        RECT 643.950 261.750 646.050 262.200 ;
        RECT 658.950 261.750 661.050 262.200 ;
        RECT 613.950 260.400 621.600 261.600 ;
        RECT 613.950 260.100 616.050 260.400 ;
        RECT 461.400 258.000 474.600 258.600 ;
        RECT 461.400 257.400 475.050 258.000 ;
        RECT 85.950 255.600 88.050 255.900 ;
        RECT 70.950 254.400 88.050 255.600 ;
        RECT 70.950 253.950 73.050 254.400 ;
        RECT 85.950 253.800 88.050 254.400 ;
        RECT 109.950 253.800 112.050 255.900 ;
        RECT 115.950 253.950 118.050 256.050 ;
        RECT 145.950 255.450 148.050 255.900 ;
        RECT 154.950 255.600 157.050 255.900 ;
        RECT 163.950 255.600 166.050 256.050 ;
        RECT 154.950 255.450 166.050 255.600 ;
        RECT 145.950 254.400 166.050 255.450 ;
        RECT 145.950 254.250 157.050 254.400 ;
        RECT 145.950 253.800 148.050 254.250 ;
        RECT 154.950 253.800 157.050 254.250 ;
        RECT 163.950 253.950 166.050 254.400 ;
        RECT 190.950 255.450 193.050 255.900 ;
        RECT 199.950 255.450 202.050 255.900 ;
        RECT 190.950 254.250 202.050 255.450 ;
        RECT 190.950 253.800 193.050 254.250 ;
        RECT 199.950 253.800 202.050 254.250 ;
        RECT 211.950 255.600 214.050 255.900 ;
        RECT 218.400 255.600 219.600 257.400 ;
        RECT 324.000 256.950 328.050 257.400 ;
        RECT 211.950 254.400 219.600 255.600 ;
        RECT 241.950 255.600 244.050 256.050 ;
        RECT 250.950 255.600 253.050 255.900 ;
        RECT 241.950 254.400 253.050 255.600 ;
        RECT 211.950 253.800 214.050 254.400 ;
        RECT 241.950 253.950 244.050 254.400 ;
        RECT 250.950 253.800 253.050 254.400 ;
        RECT 280.950 255.450 283.050 255.900 ;
        RECT 292.950 255.450 295.050 255.900 ;
        RECT 280.950 254.250 295.050 255.450 ;
        RECT 280.950 253.800 283.050 254.250 ;
        RECT 292.950 253.800 295.050 254.250 ;
        RECT 301.950 255.450 304.050 255.900 ;
        RECT 310.950 255.450 313.050 255.900 ;
        RECT 301.950 254.250 313.050 255.450 ;
        RECT 301.950 253.800 304.050 254.250 ;
        RECT 310.950 253.800 313.050 254.250 ;
        RECT 316.950 255.450 319.050 255.900 ;
        RECT 322.950 255.450 325.050 255.900 ;
        RECT 316.950 254.250 325.050 255.450 ;
        RECT 316.950 253.800 319.050 254.250 ;
        RECT 322.950 253.800 325.050 254.250 ;
        RECT 439.950 255.450 442.050 255.900 ;
        RECT 451.950 255.600 454.050 255.900 ;
        RECT 451.950 255.450 471.600 255.600 ;
        RECT 439.950 254.400 471.600 255.450 ;
        RECT 439.950 254.250 454.050 254.400 ;
        RECT 439.950 253.800 442.050 254.250 ;
        RECT 451.950 253.800 454.050 254.250 ;
        RECT 65.400 251.400 70.050 253.050 ;
        RECT 66.000 250.950 70.050 251.400 ;
        RECT 19.950 249.600 22.050 250.050 ;
        RECT 52.950 249.600 55.050 250.050 ;
        RECT 19.950 248.400 55.050 249.600 ;
        RECT 136.950 249.600 139.050 253.050 ;
        RECT 184.950 252.600 187.050 253.050 ;
        RECT 220.950 252.600 223.050 253.050 ;
        RECT 232.950 252.600 235.050 253.050 ;
        RECT 184.950 251.400 235.050 252.600 ;
        RECT 293.400 252.600 294.600 253.800 ;
        RECT 334.950 252.600 337.050 253.050 ;
        RECT 293.400 251.400 337.050 252.600 ;
        RECT 470.400 252.600 471.600 254.400 ;
        RECT 472.950 253.950 475.050 257.400 ;
        RECT 620.400 256.050 621.600 260.400 ;
        RECT 643.950 260.550 661.050 261.750 ;
        RECT 673.950 261.600 676.050 262.200 ;
        RECT 643.950 260.100 646.050 260.550 ;
        RECT 658.950 260.100 661.050 260.550 ;
        RECT 662.400 260.400 676.050 261.600 ;
        RECT 662.400 258.600 663.600 260.400 ;
        RECT 673.950 260.100 676.050 260.400 ;
        RECT 679.950 261.600 682.050 262.200 ;
        RECT 697.950 261.600 700.050 262.200 ;
        RECT 679.950 260.400 700.050 261.600 ;
        RECT 679.950 260.100 682.050 260.400 ;
        RECT 697.950 260.100 700.050 260.400 ;
        RECT 703.950 261.750 706.050 262.200 ;
        RECT 712.950 261.750 715.050 262.200 ;
        RECT 703.950 260.550 715.050 261.750 ;
        RECT 703.950 260.100 706.050 260.550 ;
        RECT 712.950 260.100 715.050 260.550 ;
        RECT 757.950 261.600 760.050 262.200 ;
        RECT 781.950 261.600 784.050 262.200 ;
        RECT 757.950 260.400 784.050 261.600 ;
        RECT 757.950 260.100 760.050 260.400 ;
        RECT 781.950 260.100 784.050 260.400 ;
        RECT 799.950 261.600 802.050 262.050 ;
        RECT 799.950 260.400 810.600 261.600 ;
        RECT 799.950 259.950 802.050 260.400 ;
        RECT 632.400 257.400 663.600 258.600 ;
        RECT 484.950 255.450 487.050 255.900 ;
        RECT 490.950 255.450 493.050 255.900 ;
        RECT 484.950 254.250 493.050 255.450 ;
        RECT 484.950 253.800 487.050 254.250 ;
        RECT 490.950 253.800 493.050 254.250 ;
        RECT 550.950 255.450 553.050 255.900 ;
        RECT 559.950 255.450 562.050 255.900 ;
        RECT 550.950 254.250 562.050 255.450 ;
        RECT 550.950 253.800 553.050 254.250 ;
        RECT 559.950 253.800 562.050 254.250 ;
        RECT 580.950 255.450 583.050 255.900 ;
        RECT 586.950 255.450 589.050 255.900 ;
        RECT 580.950 254.250 589.050 255.450 ;
        RECT 580.950 253.800 583.050 254.250 ;
        RECT 586.950 253.800 589.050 254.250 ;
        RECT 619.950 253.950 622.050 256.050 ;
        RECT 632.400 255.900 633.600 257.400 ;
        RECT 809.400 255.900 810.600 260.400 ;
        RECT 811.950 260.100 814.050 262.200 ;
        RECT 815.400 261.600 816.600 263.400 ;
        RECT 842.400 263.400 859.050 264.600 ;
        RECT 842.400 262.200 843.600 263.400 ;
        RECT 856.950 262.950 859.050 263.400 ;
        RECT 826.950 261.600 829.050 262.200 ;
        RECT 815.400 260.400 829.050 261.600 ;
        RECT 826.950 260.100 829.050 260.400 ;
        RECT 832.950 261.750 835.050 262.200 ;
        RECT 841.950 261.750 844.050 262.200 ;
        RECT 832.950 260.550 844.050 261.750 ;
        RECT 877.950 261.600 880.050 262.200 ;
        RECT 832.950 260.100 835.050 260.550 ;
        RECT 841.950 260.100 844.050 260.550 ;
        RECT 854.400 260.400 880.050 261.600 ;
        RECT 812.400 258.600 813.600 260.100 ;
        RECT 812.400 257.400 846.600 258.600 ;
        RECT 631.950 253.800 634.050 255.900 ;
        RECT 637.950 255.450 640.050 255.900 ;
        RECT 643.950 255.450 646.050 255.900 ;
        RECT 637.950 254.250 646.050 255.450 ;
        RECT 637.950 253.800 640.050 254.250 ;
        RECT 643.950 253.800 646.050 254.250 ;
        RECT 682.950 255.450 685.050 255.900 ;
        RECT 688.950 255.450 691.050 255.900 ;
        RECT 682.950 254.250 691.050 255.450 ;
        RECT 682.950 253.800 685.050 254.250 ;
        RECT 688.950 253.800 691.050 254.250 ;
        RECT 721.950 255.600 724.050 255.900 ;
        RECT 748.950 255.600 751.050 255.900 ;
        RECT 721.950 254.400 751.050 255.600 ;
        RECT 721.950 253.800 724.050 254.400 ;
        RECT 748.950 253.800 751.050 254.400 ;
        RECT 760.950 255.600 763.050 255.900 ;
        RECT 778.950 255.600 781.050 255.900 ;
        RECT 760.950 254.400 781.050 255.600 ;
        RECT 760.950 253.800 763.050 254.400 ;
        RECT 778.950 253.800 781.050 254.400 ;
        RECT 808.950 253.800 811.050 255.900 ;
        RECT 478.950 252.600 481.050 253.050 ;
        RECT 470.400 251.400 481.050 252.600 ;
        RECT 184.950 250.950 187.050 251.400 ;
        RECT 220.950 250.950 223.050 251.400 ;
        RECT 232.950 250.950 235.050 251.400 ;
        RECT 334.950 250.950 337.050 251.400 ;
        RECT 478.950 250.950 481.050 251.400 ;
        RECT 649.950 252.600 652.050 253.050 ;
        RECT 682.950 252.600 685.050 252.750 ;
        RECT 706.950 252.600 709.050 253.050 ;
        RECT 649.950 251.400 709.050 252.600 ;
        RECT 649.950 250.950 652.050 251.400 ;
        RECT 682.950 250.650 685.050 251.400 ;
        RECT 706.950 250.950 709.050 251.400 ;
        RECT 757.950 252.600 760.050 253.050 ;
        RECT 784.950 252.600 787.050 253.050 ;
        RECT 802.950 252.600 805.050 253.050 ;
        RECT 845.400 252.900 846.600 257.400 ;
        RECT 854.400 255.900 855.600 260.400 ;
        RECT 877.950 260.100 880.050 260.400 ;
        RECT 853.950 253.800 856.050 255.900 ;
        RECT 868.950 255.450 871.050 255.900 ;
        RECT 874.950 255.450 877.050 255.900 ;
        RECT 868.950 254.250 877.050 255.450 ;
        RECT 868.950 253.800 871.050 254.250 ;
        RECT 874.950 253.800 877.050 254.250 ;
        RECT 757.950 251.400 805.050 252.600 ;
        RECT 757.950 250.950 760.050 251.400 ;
        RECT 784.950 250.950 787.050 251.400 ;
        RECT 802.950 250.950 805.050 251.400 ;
        RECT 844.950 250.800 847.050 252.900 ;
        RECT 157.950 249.600 160.050 250.050 ;
        RECT 136.950 249.000 160.050 249.600 ;
        RECT 137.400 248.400 160.050 249.000 ;
        RECT 19.950 247.950 22.050 248.400 ;
        RECT 52.950 247.950 55.050 248.400 ;
        RECT 157.950 247.950 160.050 248.400 ;
        RECT 202.950 249.600 205.050 250.050 ;
        RECT 268.950 249.600 271.050 250.050 ;
        RECT 202.950 248.400 271.050 249.600 ;
        RECT 202.950 247.950 205.050 248.400 ;
        RECT 268.950 247.950 271.050 248.400 ;
        RECT 382.950 249.600 385.050 250.050 ;
        RECT 397.950 249.600 400.050 250.050 ;
        RECT 403.950 249.600 406.050 250.050 ;
        RECT 382.950 248.400 406.050 249.600 ;
        RECT 382.950 247.950 385.050 248.400 ;
        RECT 397.950 247.950 400.050 248.400 ;
        RECT 403.950 247.950 406.050 248.400 ;
        RECT 424.950 249.600 427.050 250.050 ;
        RECT 448.950 249.600 451.050 250.050 ;
        RECT 508.950 249.600 511.050 250.050 ;
        RECT 520.950 249.600 523.050 250.050 ;
        RECT 424.950 248.400 523.050 249.600 ;
        RECT 424.950 247.950 427.050 248.400 ;
        RECT 448.950 247.950 451.050 248.400 ;
        RECT 508.950 247.950 511.050 248.400 ;
        RECT 520.950 247.950 523.050 248.400 ;
        RECT 553.950 249.600 556.050 250.050 ;
        RECT 586.950 249.600 589.050 250.050 ;
        RECT 592.950 249.600 595.050 250.050 ;
        RECT 553.950 248.400 595.050 249.600 ;
        RECT 553.950 247.950 556.050 248.400 ;
        RECT 586.950 247.950 589.050 248.400 ;
        RECT 592.950 247.950 595.050 248.400 ;
        RECT 610.950 249.600 613.050 250.050 ;
        RECT 637.950 249.600 640.050 250.050 ;
        RECT 610.950 248.400 640.050 249.600 ;
        RECT 610.950 247.950 613.050 248.400 ;
        RECT 637.950 247.950 640.050 248.400 ;
        RECT 742.950 249.600 745.050 250.050 ;
        RECT 754.950 249.600 757.050 250.050 ;
        RECT 742.950 248.400 757.050 249.600 ;
        RECT 742.950 247.950 745.050 248.400 ;
        RECT 754.950 247.950 757.050 248.400 ;
        RECT 829.950 249.600 832.050 250.050 ;
        RECT 853.950 249.600 856.050 250.050 ;
        RECT 829.950 248.400 856.050 249.600 ;
        RECT 829.950 247.950 832.050 248.400 ;
        RECT 853.950 247.950 856.050 248.400 ;
        RECT 388.950 246.600 391.050 247.050 ;
        RECT 502.950 246.600 505.050 247.050 ;
        RECT 388.950 245.400 505.050 246.600 ;
        RECT 388.950 244.950 391.050 245.400 ;
        RECT 502.950 244.950 505.050 245.400 ;
        RECT 694.950 243.600 697.050 244.050 ;
        RECT 715.950 243.600 718.050 244.050 ;
        RECT 724.950 243.600 727.050 244.050 ;
        RECT 694.950 242.400 727.050 243.600 ;
        RECT 694.950 241.950 697.050 242.400 ;
        RECT 715.950 241.950 718.050 242.400 ;
        RECT 724.950 241.950 727.050 242.400 ;
        RECT 400.950 240.600 403.050 241.050 ;
        RECT 472.950 240.600 475.050 241.050 ;
        RECT 517.950 240.600 520.050 241.050 ;
        RECT 400.950 239.400 420.600 240.600 ;
        RECT 400.950 238.950 403.050 239.400 ;
        RECT 151.950 237.600 154.050 238.050 ;
        RECT 166.950 237.600 169.050 238.050 ;
        RECT 151.950 236.400 169.050 237.600 ;
        RECT 419.400 237.600 420.600 239.400 ;
        RECT 472.950 239.400 520.050 240.600 ;
        RECT 472.950 238.950 475.050 239.400 ;
        RECT 517.950 238.950 520.050 239.400 ;
        RECT 559.950 240.600 562.050 241.050 ;
        RECT 823.950 240.600 826.050 241.050 ;
        RECT 559.950 239.400 826.050 240.600 ;
        RECT 559.950 238.950 562.050 239.400 ;
        RECT 823.950 238.950 826.050 239.400 ;
        RECT 838.950 240.600 841.050 241.050 ;
        RECT 859.950 240.600 862.050 241.050 ;
        RECT 838.950 239.400 862.050 240.600 ;
        RECT 838.950 238.950 841.050 239.400 ;
        RECT 859.950 238.950 862.050 239.400 ;
        RECT 454.950 237.600 457.050 238.050 ;
        RECT 419.400 236.400 457.050 237.600 ;
        RECT 151.950 235.950 154.050 236.400 ;
        RECT 166.950 235.950 169.050 236.400 ;
        RECT 454.950 235.950 457.050 236.400 ;
        RECT 487.950 237.600 490.050 238.050 ;
        RECT 553.950 237.600 556.050 238.050 ;
        RECT 487.950 236.400 556.050 237.600 ;
        RECT 487.950 235.950 490.050 236.400 ;
        RECT 553.950 235.950 556.050 236.400 ;
        RECT 361.950 234.600 364.050 235.050 ;
        RECT 370.950 234.600 373.050 235.050 ;
        RECT 361.950 233.400 373.050 234.600 ;
        RECT 361.950 232.950 364.050 233.400 ;
        RECT 370.950 232.950 373.050 233.400 ;
        RECT 382.950 234.600 385.050 235.050 ;
        RECT 388.950 234.600 391.050 235.050 ;
        RECT 382.950 233.400 391.050 234.600 ;
        RECT 382.950 232.950 385.050 233.400 ;
        RECT 388.950 232.950 391.050 233.400 ;
        RECT 412.950 234.600 415.050 235.050 ;
        RECT 460.950 234.600 463.050 235.050 ;
        RECT 412.950 233.400 463.050 234.600 ;
        RECT 412.950 232.950 415.050 233.400 ;
        RECT 460.950 232.950 463.050 233.400 ;
        RECT 715.950 234.600 718.050 235.050 ;
        RECT 751.950 234.600 754.050 235.050 ;
        RECT 715.950 233.400 754.050 234.600 ;
        RECT 715.950 232.950 718.050 233.400 ;
        RECT 751.950 232.950 754.050 233.400 ;
        RECT 778.950 234.600 781.050 235.050 ;
        RECT 841.950 234.600 844.050 235.050 ;
        RECT 778.950 233.400 844.050 234.600 ;
        RECT 778.950 232.950 781.050 233.400 ;
        RECT 841.950 232.950 844.050 233.400 ;
        RECT 271.950 231.600 274.050 232.050 ;
        RECT 325.950 231.600 328.050 232.050 ;
        RECT 376.950 231.600 379.050 232.050 ;
        RECT 409.950 231.600 412.050 232.050 ;
        RECT 271.950 230.400 324.600 231.600 ;
        RECT 271.950 229.950 274.050 230.400 ;
        RECT 211.950 228.600 214.050 229.050 ;
        RECT 223.950 228.600 226.050 229.050 ;
        RECT 211.950 227.400 226.050 228.600 ;
        RECT 211.950 226.950 214.050 227.400 ;
        RECT 223.950 226.950 226.050 227.400 ;
        RECT 295.950 228.600 298.050 229.050 ;
        RECT 310.950 228.600 313.050 229.050 ;
        RECT 295.950 227.400 313.050 228.600 ;
        RECT 323.400 228.600 324.600 230.400 ;
        RECT 325.950 230.400 412.050 231.600 ;
        RECT 325.950 229.950 328.050 230.400 ;
        RECT 376.950 229.950 379.050 230.400 ;
        RECT 409.950 229.950 412.050 230.400 ;
        RECT 469.950 231.600 472.050 232.050 ;
        RECT 526.950 231.600 529.050 232.050 ;
        RECT 469.950 230.400 529.050 231.600 ;
        RECT 469.950 229.950 472.050 230.400 ;
        RECT 526.950 229.950 529.050 230.400 ;
        RECT 550.950 231.600 553.050 232.050 ;
        RECT 577.950 231.600 580.050 232.050 ;
        RECT 550.950 230.400 580.050 231.600 ;
        RECT 550.950 229.950 553.050 230.400 ;
        RECT 577.950 229.950 580.050 230.400 ;
        RECT 667.950 231.600 670.050 232.050 ;
        RECT 766.950 231.600 769.050 232.050 ;
        RECT 667.950 230.400 769.050 231.600 ;
        RECT 667.950 229.950 670.050 230.400 ;
        RECT 766.950 229.950 769.050 230.400 ;
        RECT 364.950 228.600 367.050 229.050 ;
        RECT 388.950 228.600 391.050 229.050 ;
        RECT 439.950 228.600 442.050 229.050 ;
        RECT 323.400 227.400 391.050 228.600 ;
        RECT 295.950 226.950 298.050 227.400 ;
        RECT 310.950 226.950 313.050 227.400 ;
        RECT 364.950 226.950 367.050 227.400 ;
        RECT 388.950 226.950 391.050 227.400 ;
        RECT 398.400 227.400 442.050 228.600 ;
        RECT 67.950 225.600 70.050 226.050 ;
        RECT 109.950 225.600 112.050 226.050 ;
        RECT 124.950 225.600 127.050 226.050 ;
        RECT 67.950 224.400 127.050 225.600 ;
        RECT 67.950 223.950 70.050 224.400 ;
        RECT 109.950 223.950 112.050 224.400 ;
        RECT 124.950 223.950 127.050 224.400 ;
        RECT 379.950 225.600 382.050 226.050 ;
        RECT 398.400 225.600 399.600 227.400 ;
        RECT 439.950 226.950 442.050 227.400 ;
        RECT 676.950 228.600 679.050 229.050 ;
        RECT 676.950 227.400 693.600 228.600 ;
        RECT 676.950 226.950 679.050 227.400 ;
        RECT 379.950 224.400 399.600 225.600 ;
        RECT 637.950 225.600 640.050 226.050 ;
        RECT 646.950 225.600 649.050 226.050 ;
        RECT 637.950 224.400 649.050 225.600 ;
        RECT 692.400 225.600 693.600 227.400 ;
        RECT 742.950 225.600 745.050 226.050 ;
        RECT 692.400 224.400 745.050 225.600 ;
        RECT 379.950 223.950 382.050 224.400 ;
        RECT 637.950 223.950 640.050 224.400 ;
        RECT 646.950 223.950 649.050 224.400 ;
        RECT 742.950 223.950 745.050 224.400 ;
        RECT 178.950 222.600 181.050 223.050 ;
        RECT 184.950 222.600 187.050 223.050 ;
        RECT 178.950 221.400 187.050 222.600 ;
        RECT 178.950 220.950 181.050 221.400 ;
        RECT 184.950 220.950 187.050 221.400 ;
        RECT 202.950 222.600 205.050 223.050 ;
        RECT 208.950 222.600 211.050 223.050 ;
        RECT 220.950 222.600 223.050 223.050 ;
        RECT 271.950 222.600 274.050 223.050 ;
        RECT 202.950 221.400 223.050 222.600 ;
        RECT 202.950 220.950 205.050 221.400 ;
        RECT 208.950 220.950 211.050 221.400 ;
        RECT 220.950 220.950 223.050 221.400 ;
        RECT 251.400 221.400 274.050 222.600 ;
        RECT 251.400 220.050 252.600 221.400 ;
        RECT 271.950 220.950 274.050 221.400 ;
        RECT 415.950 222.600 418.050 223.050 ;
        RECT 433.950 222.600 436.050 223.050 ;
        RECT 415.950 221.400 436.050 222.600 ;
        RECT 415.950 220.950 418.050 221.400 ;
        RECT 433.950 220.950 436.050 221.400 ;
        RECT 466.950 222.600 469.050 223.050 ;
        RECT 478.950 222.600 481.050 223.050 ;
        RECT 466.950 221.400 481.050 222.600 ;
        RECT 466.950 220.950 469.050 221.400 ;
        RECT 478.950 220.950 481.050 221.400 ;
        RECT 487.950 222.600 490.050 223.050 ;
        RECT 508.950 222.600 511.050 223.050 ;
        RECT 487.950 221.400 511.050 222.600 ;
        RECT 487.950 220.950 490.050 221.400 ;
        RECT 508.950 220.950 511.050 221.400 ;
        RECT 514.950 222.600 517.050 223.050 ;
        RECT 529.950 222.600 532.050 223.050 ;
        RECT 514.950 221.400 532.050 222.600 ;
        RECT 514.950 220.950 517.050 221.400 ;
        RECT 529.950 220.950 532.050 221.400 ;
        RECT 535.950 222.600 538.050 223.050 ;
        RECT 541.950 222.600 544.050 223.050 ;
        RECT 535.950 221.400 544.050 222.600 ;
        RECT 535.950 220.950 538.050 221.400 ;
        RECT 541.950 220.950 544.050 221.400 ;
        RECT 556.950 222.600 559.050 223.050 ;
        RECT 601.950 222.600 604.050 223.050 ;
        RECT 556.950 221.400 604.050 222.600 ;
        RECT 556.950 220.950 559.050 221.400 ;
        RECT 601.950 220.950 604.050 221.400 ;
        RECT 670.950 222.600 673.050 223.050 ;
        RECT 688.950 222.600 691.050 223.050 ;
        RECT 700.950 222.600 703.050 223.050 ;
        RECT 718.950 222.600 721.050 223.050 ;
        RECT 670.950 221.400 721.050 222.600 ;
        RECT 670.950 220.950 673.050 221.400 ;
        RECT 688.950 220.950 691.050 221.400 ;
        RECT 700.950 220.950 703.050 221.400 ;
        RECT 718.950 220.950 721.050 221.400 ;
        RECT 751.950 222.600 754.050 223.050 ;
        RECT 784.950 222.600 787.050 223.050 ;
        RECT 751.950 221.400 787.050 222.600 ;
        RECT 751.950 220.950 754.050 221.400 ;
        RECT 784.950 220.950 787.050 221.400 ;
        RECT 799.950 222.600 802.050 223.050 ;
        RECT 805.950 222.600 808.050 223.050 ;
        RECT 799.950 221.400 808.050 222.600 ;
        RECT 799.950 220.950 802.050 221.400 ;
        RECT 805.950 220.950 808.050 221.400 ;
        RECT 817.950 222.600 820.050 223.050 ;
        RECT 859.950 222.600 862.050 223.050 ;
        RECT 877.950 222.600 880.050 223.050 ;
        RECT 817.950 221.400 880.050 222.600 ;
        RECT 817.950 220.950 820.050 221.400 ;
        RECT 859.950 220.950 862.050 221.400 ;
        RECT 877.950 220.950 880.050 221.400 ;
        RECT 235.950 219.600 238.050 220.050 ;
        RECT 250.950 219.600 253.050 220.050 ;
        RECT 235.950 218.400 253.050 219.600 ;
        RECT 235.950 217.950 238.050 218.400 ;
        RECT 250.950 217.950 253.050 218.400 ;
        RECT 298.950 219.600 301.050 220.050 ;
        RECT 319.950 219.600 322.050 220.050 ;
        RECT 298.950 218.400 322.050 219.600 ;
        RECT 298.950 217.950 301.050 218.400 ;
        RECT 319.950 217.950 322.050 218.400 ;
        RECT 490.950 219.600 493.050 220.050 ;
        RECT 505.950 219.600 508.050 220.050 ;
        RECT 568.950 219.600 571.050 220.050 ;
        RECT 583.950 219.600 586.050 220.050 ;
        RECT 490.950 218.400 516.600 219.600 ;
        RECT 490.950 217.950 493.050 218.400 ;
        RECT 505.950 217.950 508.050 218.400 ;
        RECT 28.950 216.750 31.050 217.200 ;
        RECT 34.800 216.750 36.900 217.200 ;
        RECT 28.950 215.550 36.900 216.750 ;
        RECT 28.950 215.100 31.050 215.550 ;
        RECT 34.800 215.100 36.900 215.550 ;
        RECT 37.950 216.750 40.050 217.200 ;
        RECT 43.950 216.750 46.050 217.200 ;
        RECT 37.950 215.550 46.050 216.750 ;
        RECT 37.950 215.100 40.050 215.550 ;
        RECT 43.950 215.100 46.050 215.550 ;
        RECT 88.950 216.750 91.050 217.200 ;
        RECT 97.950 216.750 100.050 217.200 ;
        RECT 88.950 215.550 100.050 216.750 ;
        RECT 88.950 215.100 91.050 215.550 ;
        RECT 97.950 215.100 100.050 215.550 ;
        RECT 103.950 216.750 106.050 217.200 ;
        RECT 115.950 216.750 118.050 217.200 ;
        RECT 103.950 215.550 118.050 216.750 ;
        RECT 103.950 215.100 106.050 215.550 ;
        RECT 115.950 215.100 118.050 215.550 ;
        RECT 130.950 216.750 133.050 217.200 ;
        RECT 139.950 216.750 142.050 217.200 ;
        RECT 130.950 215.550 142.050 216.750 ;
        RECT 130.950 215.100 133.050 215.550 ;
        RECT 139.950 215.100 142.050 215.550 ;
        RECT 172.950 216.600 175.050 217.200 ;
        RECT 193.950 216.600 196.050 217.200 ;
        RECT 172.950 215.400 196.050 216.600 ;
        RECT 172.950 215.100 175.050 215.400 ;
        RECT 193.950 215.100 196.050 215.400 ;
        RECT 199.950 215.100 202.050 217.200 ;
        RECT 259.950 216.750 262.050 217.200 ;
        RECT 265.950 216.750 268.050 217.200 ;
        RECT 259.950 215.550 268.050 216.750 ;
        RECT 259.950 215.100 262.050 215.550 ;
        RECT 265.950 215.100 268.050 215.550 ;
        RECT 283.950 216.750 286.050 217.200 ;
        RECT 298.950 216.750 301.050 217.200 ;
        RECT 283.950 215.550 301.050 216.750 ;
        RECT 283.950 215.100 286.050 215.550 ;
        RECT 298.950 215.100 301.050 215.550 ;
        RECT 325.950 216.750 328.050 217.200 ;
        RECT 334.950 216.750 337.050 217.200 ;
        RECT 325.950 215.550 337.050 216.750 ;
        RECT 340.950 216.600 343.050 217.200 ;
        RECT 325.950 215.100 328.050 215.550 ;
        RECT 334.950 215.100 337.050 215.550 ;
        RECT 338.400 215.400 343.050 216.600 ;
        RECT 200.400 213.600 201.600 215.100 ;
        RECT 200.400 212.400 225.600 213.600 ;
        RECT 82.950 210.600 85.050 211.050 ;
        RECT 224.400 210.900 225.600 212.400 ;
        RECT 338.400 211.050 339.600 215.400 ;
        RECT 340.950 215.100 343.050 215.400 ;
        RECT 370.950 216.600 373.050 217.050 ;
        RECT 382.950 216.600 385.050 217.050 ;
        RECT 370.950 215.400 385.050 216.600 ;
        RECT 370.950 214.950 373.050 215.400 ;
        RECT 382.950 214.950 385.050 215.400 ;
        RECT 400.950 216.750 403.050 217.200 ;
        RECT 415.950 216.750 418.050 217.200 ;
        RECT 400.950 215.550 418.050 216.750 ;
        RECT 400.950 215.100 403.050 215.550 ;
        RECT 415.950 215.100 418.050 215.550 ;
        RECT 427.950 216.600 430.050 217.050 ;
        RECT 457.950 216.600 460.050 217.050 ;
        RECT 427.950 215.400 460.050 216.600 ;
        RECT 427.950 214.950 430.050 215.400 ;
        RECT 457.950 214.950 460.050 215.400 ;
        RECT 493.950 216.750 496.050 217.200 ;
        RECT 499.950 216.750 502.050 217.200 ;
        RECT 493.950 215.550 502.050 216.750 ;
        RECT 493.950 215.100 496.050 215.550 ;
        RECT 499.950 215.100 502.050 215.550 ;
        RECT 515.400 216.600 516.600 218.400 ;
        RECT 568.950 218.400 586.050 219.600 ;
        RECT 602.400 219.600 603.600 220.950 ;
        RECT 637.950 219.600 640.050 220.050 ;
        RECT 602.400 218.400 640.050 219.600 ;
        RECT 568.950 217.950 571.050 218.400 ;
        RECT 583.950 217.950 586.050 218.400 ;
        RECT 637.950 217.950 640.050 218.400 ;
        RECT 655.950 219.600 658.050 220.050 ;
        RECT 664.950 219.600 667.050 220.050 ;
        RECT 655.950 218.400 667.050 219.600 ;
        RECT 655.950 217.950 658.050 218.400 ;
        RECT 664.950 217.950 667.050 218.400 ;
        RECT 790.950 219.600 793.050 220.050 ;
        RECT 796.950 219.600 799.050 220.050 ;
        RECT 808.950 219.600 811.050 219.900 ;
        RECT 790.950 218.400 811.050 219.600 ;
        RECT 790.950 217.950 793.050 218.400 ;
        RECT 796.950 217.950 799.050 218.400 ;
        RECT 808.950 217.800 811.050 218.400 ;
        RECT 826.950 219.600 829.050 220.050 ;
        RECT 832.950 219.600 835.050 220.050 ;
        RECT 826.950 218.400 835.050 219.600 ;
        RECT 826.950 217.950 829.050 218.400 ;
        RECT 832.950 217.950 835.050 218.400 ;
        RECT 517.950 216.600 520.050 217.200 ;
        RECT 535.950 216.600 538.050 217.200 ;
        RECT 515.400 215.400 520.050 216.600 ;
        RECT 517.950 215.100 520.050 215.400 ;
        RECT 521.400 215.400 538.050 216.600 ;
        RECT 475.950 213.600 478.050 214.050 ;
        RECT 521.400 213.600 522.600 215.400 ;
        RECT 535.950 215.100 538.050 215.400 ;
        RECT 592.950 216.600 595.050 217.200 ;
        RECT 622.950 216.750 625.050 217.200 ;
        RECT 628.950 216.750 631.050 217.200 ;
        RECT 592.950 215.400 612.600 216.600 ;
        RECT 592.950 215.100 595.050 215.400 ;
        RECT 475.950 212.400 522.600 213.600 ;
        RECT 475.950 211.950 478.050 212.400 ;
        RECT 94.950 210.600 97.050 210.900 ;
        RECT 82.950 209.400 97.050 210.600 ;
        RECT 82.950 208.950 85.050 209.400 ;
        RECT 94.950 208.800 97.050 209.400 ;
        RECT 121.950 210.600 124.050 210.900 ;
        RECT 154.950 210.600 157.050 210.900 ;
        RECT 121.950 209.400 157.050 210.600 ;
        RECT 121.950 208.800 124.050 209.400 ;
        RECT 154.950 208.800 157.050 209.400 ;
        RECT 175.950 210.450 178.050 210.900 ;
        RECT 184.950 210.600 187.050 210.900 ;
        RECT 196.950 210.600 199.050 210.900 ;
        RECT 184.950 210.450 199.050 210.600 ;
        RECT 175.950 209.400 199.050 210.450 ;
        RECT 175.950 209.250 187.050 209.400 ;
        RECT 175.950 208.800 178.050 209.250 ;
        RECT 184.950 208.800 187.050 209.250 ;
        RECT 196.950 208.800 199.050 209.400 ;
        RECT 223.950 208.800 226.050 210.900 ;
        RECT 274.950 210.600 277.050 210.900 ;
        RECT 283.950 210.600 286.050 211.050 ;
        RECT 274.950 209.400 286.050 210.600 ;
        RECT 274.950 208.800 277.050 209.400 ;
        RECT 283.950 208.950 286.050 209.400 ;
        RECT 310.950 210.450 313.050 210.900 ;
        RECT 322.950 210.450 325.050 210.900 ;
        RECT 310.950 209.250 325.050 210.450 ;
        RECT 310.950 208.800 313.050 209.250 ;
        RECT 322.950 208.800 325.050 209.250 ;
        RECT 337.950 208.950 340.050 211.050 ;
        RECT 343.950 210.450 346.050 210.900 ;
        RECT 352.950 210.450 355.050 210.900 ;
        RECT 343.950 209.250 355.050 210.450 ;
        RECT 343.950 208.800 346.050 209.250 ;
        RECT 352.950 208.800 355.050 209.250 ;
        RECT 376.950 210.450 379.050 210.900 ;
        RECT 385.950 210.450 388.050 210.900 ;
        RECT 376.950 209.250 388.050 210.450 ;
        RECT 376.950 208.800 379.050 209.250 ;
        RECT 385.950 208.800 388.050 209.250 ;
        RECT 418.950 210.600 421.050 210.900 ;
        RECT 424.950 210.600 427.050 211.050 ;
        RECT 436.950 210.600 439.050 210.900 ;
        RECT 418.950 209.400 439.050 210.600 ;
        RECT 418.950 208.800 421.050 209.400 ;
        RECT 424.950 208.950 427.050 209.400 ;
        RECT 436.950 208.800 439.050 209.400 ;
        RECT 454.950 210.450 457.050 210.900 ;
        RECT 463.950 210.450 466.050 210.900 ;
        RECT 454.950 209.250 466.050 210.450 ;
        RECT 454.950 208.800 457.050 209.250 ;
        RECT 463.950 208.800 466.050 209.250 ;
        RECT 484.950 210.600 487.050 210.900 ;
        RECT 502.950 210.600 505.050 211.050 ;
        RECT 484.950 209.400 505.050 210.600 ;
        RECT 484.950 208.800 487.050 209.400 ;
        RECT 502.950 208.950 505.050 209.400 ;
        RECT 511.950 210.450 514.050 210.900 ;
        RECT 520.950 210.450 523.050 210.900 ;
        RECT 511.950 209.250 523.050 210.450 ;
        RECT 511.950 208.800 514.050 209.250 ;
        RECT 520.950 208.800 523.050 209.250 ;
        RECT 526.950 210.450 529.050 210.900 ;
        RECT 538.950 210.450 541.050 210.900 ;
        RECT 526.950 209.250 541.050 210.450 ;
        RECT 526.950 208.800 529.050 209.250 ;
        RECT 538.950 208.800 541.050 209.250 ;
        RECT 544.950 210.600 547.050 210.900 ;
        RECT 559.950 210.600 562.050 211.050 ;
        RECT 611.400 210.900 612.600 215.400 ;
        RECT 622.950 215.550 631.050 216.750 ;
        RECT 666.000 216.600 670.050 217.050 ;
        RECT 622.950 215.100 625.050 215.550 ;
        RECT 628.950 215.100 631.050 215.550 ;
        RECT 665.400 214.950 670.050 216.600 ;
        RECT 673.950 216.600 676.050 217.050 ;
        RECT 682.950 216.600 685.050 217.200 ;
        RECT 673.950 215.400 685.050 216.600 ;
        RECT 673.950 214.950 676.050 215.400 ;
        RECT 682.950 215.100 685.050 215.400 ;
        RECT 697.950 216.600 700.050 217.050 ;
        RECT 706.950 216.600 709.050 217.200 ;
        RECT 697.950 215.400 709.050 216.600 ;
        RECT 697.950 214.950 700.050 215.400 ;
        RECT 706.950 215.100 709.050 215.400 ;
        RECT 718.950 216.600 723.000 217.050 ;
        RECT 730.950 216.750 733.050 217.200 ;
        RECT 739.950 216.750 742.050 217.200 ;
        RECT 718.950 214.950 723.600 216.600 ;
        RECT 730.950 215.550 742.050 216.750 ;
        RECT 730.950 215.100 733.050 215.550 ;
        RECT 739.950 215.100 742.050 215.550 ;
        RECT 757.950 216.750 760.050 217.200 ;
        RECT 763.950 216.750 766.050 217.200 ;
        RECT 757.950 215.550 766.050 216.750 ;
        RECT 757.950 215.100 760.050 215.550 ;
        RECT 763.950 215.100 766.050 215.550 ;
        RECT 772.950 216.750 775.050 217.200 ;
        RECT 778.950 216.750 781.050 217.200 ;
        RECT 772.950 215.550 781.050 216.750 ;
        RECT 772.950 215.100 775.050 215.550 ;
        RECT 778.950 215.100 781.050 215.550 ;
        RECT 802.950 215.100 805.050 217.200 ;
        RECT 820.950 216.600 825.000 217.050 ;
        RECT 844.950 216.600 847.050 217.050 ;
        RECT 544.950 209.400 562.050 210.600 ;
        RECT 544.950 208.800 547.050 209.400 ;
        RECT 559.950 208.950 562.050 209.400 ;
        RECT 568.950 210.600 571.050 210.900 ;
        RECT 574.950 210.600 577.050 210.900 ;
        RECT 568.950 209.400 577.050 210.600 ;
        RECT 568.950 208.800 571.050 209.400 ;
        RECT 574.950 208.800 577.050 209.400 ;
        RECT 610.950 208.800 613.050 210.900 ;
        RECT 643.950 210.600 646.050 211.050 ;
        RECT 665.400 210.900 666.600 214.950 ;
        RECT 658.950 210.600 661.050 210.900 ;
        RECT 643.950 209.400 661.050 210.600 ;
        RECT 643.950 208.950 646.050 209.400 ;
        RECT 658.950 208.800 661.050 209.400 ;
        RECT 664.950 208.800 667.050 210.900 ;
        RECT 691.950 210.600 694.050 211.050 ;
        RECT 718.950 210.600 721.050 211.050 ;
        RECT 691.950 209.400 721.050 210.600 ;
        RECT 722.400 210.600 723.600 214.950 ;
        RECT 727.950 210.600 730.050 210.900 ;
        RECT 722.400 209.400 730.050 210.600 ;
        RECT 691.950 208.950 694.050 209.400 ;
        RECT 718.950 208.950 721.050 209.400 ;
        RECT 727.950 208.800 730.050 209.400 ;
        RECT 742.950 210.600 745.050 211.050 ;
        RECT 748.950 210.600 751.050 210.900 ;
        RECT 742.950 209.400 751.050 210.600 ;
        RECT 742.950 208.950 745.050 209.400 ;
        RECT 748.950 208.800 751.050 209.400 ;
        RECT 754.950 210.450 757.050 210.900 ;
        RECT 760.950 210.450 763.050 210.900 ;
        RECT 754.950 209.250 763.050 210.450 ;
        RECT 754.950 208.800 757.050 209.250 ;
        RECT 760.950 208.800 763.050 209.250 ;
        RECT 766.950 210.600 769.050 211.050 ;
        RECT 775.950 210.600 778.050 210.900 ;
        RECT 766.950 209.400 778.050 210.600 ;
        RECT 766.950 208.950 769.050 209.400 ;
        RECT 775.950 208.800 778.050 209.400 ;
        RECT 796.950 210.600 799.050 211.050 ;
        RECT 803.400 210.600 804.600 215.100 ;
        RECT 820.950 214.950 825.600 216.600 ;
        RECT 839.400 216.000 847.050 216.600 ;
        RECT 796.950 209.400 804.600 210.600 ;
        RECT 805.950 210.600 808.050 210.900 ;
        RECT 814.950 210.600 817.050 211.050 ;
        RECT 824.400 210.900 825.600 214.950 ;
        RECT 838.950 215.400 847.050 216.000 ;
        RECT 838.950 211.950 841.050 215.400 ;
        RECT 844.950 214.950 847.050 215.400 ;
        RECT 805.950 209.400 817.050 210.600 ;
        RECT 796.950 208.950 799.050 209.400 ;
        RECT 805.950 208.800 808.050 209.400 ;
        RECT 814.950 208.950 817.050 209.400 ;
        RECT 823.950 208.800 826.050 210.900 ;
        RECT 46.950 207.600 49.050 208.050 ;
        RECT 88.950 207.600 91.050 208.050 ;
        RECT 46.950 206.400 91.050 207.600 ;
        RECT 46.950 205.950 49.050 206.400 ;
        RECT 88.950 205.950 91.050 206.400 ;
        RECT 361.950 207.600 364.050 208.050 ;
        RECT 377.400 207.600 378.600 208.800 ;
        RECT 361.950 206.400 378.600 207.600 ;
        RECT 487.950 207.600 490.050 208.050 ;
        RECT 499.950 207.600 502.050 208.050 ;
        RECT 487.950 206.400 502.050 207.600 ;
        RECT 361.950 205.950 364.050 206.400 ;
        RECT 487.950 205.950 490.050 206.400 ;
        RECT 499.950 205.950 502.050 206.400 ;
        RECT 673.950 207.600 676.050 208.050 ;
        RECT 703.950 207.600 706.050 208.050 ;
        RECT 673.950 206.400 706.050 207.600 ;
        RECT 673.950 205.950 676.050 206.400 ;
        RECT 703.950 205.950 706.050 206.400 ;
        RECT 769.950 207.600 772.050 208.050 ;
        RECT 781.950 207.600 784.050 208.050 ;
        RECT 793.950 207.600 796.050 208.050 ;
        RECT 769.950 206.400 796.050 207.600 ;
        RECT 769.950 205.950 772.050 206.400 ;
        RECT 781.950 205.950 784.050 206.400 ;
        RECT 793.950 205.950 796.050 206.400 ;
        RECT 847.950 207.600 850.050 208.050 ;
        RECT 859.950 207.600 862.050 208.050 ;
        RECT 847.950 206.400 862.050 207.600 ;
        RECT 847.950 205.950 850.050 206.400 ;
        RECT 859.950 205.950 862.050 206.400 ;
        RECT 19.950 204.600 22.050 205.050 ;
        RECT 61.950 204.600 64.050 205.050 ;
        RECT 19.950 203.400 64.050 204.600 ;
        RECT 19.950 202.950 22.050 203.400 ;
        RECT 61.950 202.950 64.050 203.400 ;
        RECT 76.950 204.600 79.050 205.050 ;
        RECT 82.950 204.600 85.050 205.050 ;
        RECT 76.950 203.400 85.050 204.600 ;
        RECT 89.400 204.600 90.600 205.950 ;
        RECT 130.950 204.600 133.050 205.050 ;
        RECT 89.400 203.400 133.050 204.600 ;
        RECT 76.950 202.950 79.050 203.400 ;
        RECT 82.950 202.950 85.050 203.400 ;
        RECT 130.950 202.950 133.050 203.400 ;
        RECT 199.950 204.600 202.050 205.050 ;
        RECT 211.950 204.600 214.050 205.050 ;
        RECT 217.950 204.600 220.050 205.050 ;
        RECT 199.950 203.400 220.050 204.600 ;
        RECT 199.950 202.950 202.050 203.400 ;
        RECT 211.950 202.950 214.050 203.400 ;
        RECT 217.950 202.950 220.050 203.400 ;
        RECT 232.950 204.600 235.050 205.050 ;
        RECT 247.950 204.600 250.050 205.050 ;
        RECT 268.950 204.600 271.050 205.050 ;
        RECT 232.950 203.400 271.050 204.600 ;
        RECT 232.950 202.950 235.050 203.400 ;
        RECT 247.950 202.950 250.050 203.400 ;
        RECT 268.950 202.950 271.050 203.400 ;
        RECT 403.950 204.600 406.050 205.050 ;
        RECT 412.950 204.600 415.050 205.050 ;
        RECT 403.950 203.400 415.050 204.600 ;
        RECT 403.950 202.950 406.050 203.400 ;
        RECT 412.950 202.950 415.050 203.400 ;
        RECT 430.950 204.600 433.050 205.050 ;
        RECT 475.950 204.600 478.050 205.050 ;
        RECT 430.950 203.400 478.050 204.600 ;
        RECT 430.950 202.950 433.050 203.400 ;
        RECT 475.950 202.950 478.050 203.400 ;
        RECT 646.950 204.600 649.050 205.050 ;
        RECT 658.950 204.600 661.050 205.050 ;
        RECT 646.950 203.400 661.050 204.600 ;
        RECT 646.950 202.950 649.050 203.400 ;
        RECT 658.950 202.950 661.050 203.400 ;
        RECT 721.950 204.600 724.050 205.050 ;
        RECT 727.950 204.600 730.050 205.050 ;
        RECT 721.950 203.400 730.050 204.600 ;
        RECT 721.950 202.950 724.050 203.400 ;
        RECT 727.950 202.950 730.050 203.400 ;
        RECT 736.950 204.600 739.050 205.050 ;
        RECT 763.950 204.600 766.050 205.050 ;
        RECT 736.950 203.400 766.050 204.600 ;
        RECT 736.950 202.950 739.050 203.400 ;
        RECT 763.950 202.950 766.050 203.400 ;
        RECT 841.950 204.600 844.050 205.050 ;
        RECT 874.950 204.600 877.050 205.050 ;
        RECT 841.950 203.400 877.050 204.600 ;
        RECT 841.950 202.950 844.050 203.400 ;
        RECT 874.950 202.950 877.050 203.400 ;
        RECT 100.950 201.600 103.050 202.050 ;
        RECT 109.950 201.600 112.050 202.050 ;
        RECT 100.950 200.400 112.050 201.600 ;
        RECT 100.950 199.950 103.050 200.400 ;
        RECT 109.950 199.950 112.050 200.400 ;
        RECT 295.950 201.600 298.050 202.050 ;
        RECT 310.950 201.600 313.050 202.050 ;
        RECT 295.950 200.400 313.050 201.600 ;
        RECT 295.950 199.950 298.050 200.400 ;
        RECT 310.950 199.950 313.050 200.400 ;
        RECT 367.950 201.600 370.050 202.050 ;
        RECT 379.950 201.600 382.050 202.050 ;
        RECT 367.950 200.400 382.050 201.600 ;
        RECT 367.950 199.950 370.050 200.400 ;
        RECT 379.950 199.950 382.050 200.400 ;
        RECT 412.950 201.600 415.050 201.900 ;
        RECT 427.950 201.600 430.050 202.050 ;
        RECT 412.950 200.400 430.050 201.600 ;
        RECT 412.950 199.800 415.050 200.400 ;
        RECT 427.950 199.950 430.050 200.400 ;
        RECT 478.950 201.600 481.050 202.050 ;
        RECT 490.950 201.600 493.050 202.050 ;
        RECT 496.950 201.600 499.050 202.050 ;
        RECT 478.950 200.400 499.050 201.600 ;
        RECT 478.950 199.950 481.050 200.400 ;
        RECT 490.950 199.950 493.050 200.400 ;
        RECT 496.950 199.950 499.050 200.400 ;
        RECT 733.950 201.600 736.050 202.050 ;
        RECT 769.950 201.600 772.050 202.050 ;
        RECT 796.950 201.600 799.050 202.050 ;
        RECT 733.950 200.400 799.050 201.600 ;
        RECT 733.950 199.950 736.050 200.400 ;
        RECT 769.950 199.950 772.050 200.400 ;
        RECT 796.950 199.950 799.050 200.400 ;
        RECT 16.950 198.600 19.050 199.050 ;
        RECT 37.950 198.600 40.050 199.050 ;
        RECT 16.950 197.400 40.050 198.600 ;
        RECT 16.950 196.950 19.050 197.400 ;
        RECT 37.950 196.950 40.050 197.400 ;
        RECT 151.950 198.600 154.050 199.050 ;
        RECT 157.950 198.600 160.050 199.050 ;
        RECT 151.950 197.400 160.050 198.600 ;
        RECT 151.950 196.950 154.050 197.400 ;
        RECT 157.950 196.950 160.050 197.400 ;
        RECT 211.950 198.600 214.050 199.050 ;
        RECT 259.950 198.600 262.050 199.050 ;
        RECT 211.950 197.400 262.050 198.600 ;
        RECT 211.950 196.950 214.050 197.400 ;
        RECT 259.950 196.950 262.050 197.400 ;
        RECT 601.950 198.600 604.050 199.050 ;
        RECT 619.950 198.600 622.050 199.050 ;
        RECT 601.950 197.400 622.050 198.600 ;
        RECT 601.950 196.950 604.050 197.400 ;
        RECT 619.950 196.950 622.050 197.400 ;
        RECT 631.950 198.600 634.050 199.050 ;
        RECT 673.950 198.600 676.050 199.050 ;
        RECT 631.950 197.400 676.050 198.600 ;
        RECT 631.950 196.950 634.050 197.400 ;
        RECT 673.950 196.950 676.050 197.400 ;
        RECT 748.950 198.600 751.050 199.050 ;
        RECT 775.950 198.600 778.050 199.050 ;
        RECT 748.950 197.400 778.050 198.600 ;
        RECT 748.950 196.950 751.050 197.400 ;
        RECT 775.950 196.950 778.050 197.400 ;
        RECT 400.950 195.600 403.050 196.050 ;
        RECT 481.950 195.600 484.050 196.050 ;
        RECT 505.950 195.600 508.050 196.050 ;
        RECT 400.950 194.400 417.600 195.600 ;
        RECT 400.950 193.950 403.050 194.400 ;
        RECT 46.950 192.600 49.050 193.050 ;
        RECT 103.950 192.600 106.050 193.050 ;
        RECT 46.950 191.400 106.050 192.600 ;
        RECT 46.950 190.950 49.050 191.400 ;
        RECT 103.950 190.950 106.050 191.400 ;
        RECT 112.950 192.600 115.050 193.050 ;
        RECT 148.950 192.600 151.050 193.050 ;
        RECT 112.950 191.400 151.050 192.600 ;
        RECT 112.950 190.950 115.050 191.400 ;
        RECT 148.950 190.950 151.050 191.400 ;
        RECT 190.950 192.600 193.050 193.050 ;
        RECT 217.950 192.600 220.050 193.050 ;
        RECT 238.950 192.600 241.050 193.050 ;
        RECT 190.950 191.400 241.050 192.600 ;
        RECT 416.400 192.600 417.600 194.400 ;
        RECT 481.950 194.400 508.050 195.600 ;
        RECT 481.950 193.950 484.050 194.400 ;
        RECT 505.950 193.950 508.050 194.400 ;
        RECT 529.950 195.600 532.050 196.050 ;
        RECT 721.950 195.600 724.050 196.050 ;
        RECT 529.950 194.400 724.050 195.600 ;
        RECT 529.950 193.950 532.050 194.400 ;
        RECT 721.950 193.950 724.050 194.400 ;
        RECT 730.950 195.600 733.050 196.050 ;
        RECT 739.950 195.600 742.050 196.050 ;
        RECT 730.950 194.400 742.050 195.600 ;
        RECT 730.950 193.950 733.050 194.400 ;
        RECT 739.950 193.950 742.050 194.400 ;
        RECT 745.950 195.600 748.050 196.050 ;
        RECT 793.950 195.600 796.050 196.050 ;
        RECT 799.950 195.600 802.050 196.050 ;
        RECT 745.950 194.400 792.600 195.600 ;
        RECT 745.950 193.950 748.050 194.400 ;
        RECT 436.950 192.600 439.050 193.050 ;
        RECT 416.400 191.400 439.050 192.600 ;
        RECT 190.950 190.950 193.050 191.400 ;
        RECT 217.950 190.950 220.050 191.400 ;
        RECT 238.950 190.950 241.050 191.400 ;
        RECT 436.950 190.950 439.050 191.400 ;
        RECT 586.950 192.600 589.050 193.050 ;
        RECT 742.950 192.600 745.050 193.050 ;
        RECT 586.950 191.400 745.050 192.600 ;
        RECT 791.400 192.600 792.600 194.400 ;
        RECT 793.950 194.400 802.050 195.600 ;
        RECT 793.950 193.950 796.050 194.400 ;
        RECT 799.950 193.950 802.050 194.400 ;
        RECT 805.950 192.600 808.050 193.050 ;
        RECT 791.400 191.400 808.050 192.600 ;
        RECT 586.950 190.950 589.050 191.400 ;
        RECT 742.950 190.950 745.050 191.400 ;
        RECT 805.950 190.950 808.050 191.400 ;
        RECT 193.950 189.600 196.050 190.050 ;
        RECT 202.950 189.600 205.050 190.050 ;
        RECT 193.950 188.400 205.050 189.600 ;
        RECT 193.950 187.950 196.050 188.400 ;
        RECT 202.950 187.950 205.050 188.400 ;
        RECT 298.950 189.600 301.050 190.050 ;
        RECT 316.950 189.600 319.050 190.050 ;
        RECT 298.950 188.400 319.050 189.600 ;
        RECT 298.950 187.950 301.050 188.400 ;
        RECT 316.950 187.950 319.050 188.400 ;
        RECT 391.950 189.600 394.050 190.050 ;
        RECT 412.950 189.600 415.050 190.050 ;
        RECT 391.950 188.400 415.050 189.600 ;
        RECT 391.950 187.950 394.050 188.400 ;
        RECT 412.950 187.950 415.050 188.400 ;
        RECT 469.950 189.600 472.050 190.050 ;
        RECT 511.950 189.600 514.050 190.050 ;
        RECT 469.950 188.400 514.050 189.600 ;
        RECT 469.950 187.950 472.050 188.400 ;
        RECT 511.950 187.950 514.050 188.400 ;
        RECT 532.950 189.600 535.050 190.050 ;
        RECT 583.950 189.600 586.050 190.050 ;
        RECT 532.950 188.400 586.050 189.600 ;
        RECT 532.950 187.950 535.050 188.400 ;
        RECT 583.950 187.950 586.050 188.400 ;
        RECT 640.950 189.600 643.050 190.050 ;
        RECT 670.950 189.600 673.050 190.050 ;
        RECT 640.950 188.400 673.050 189.600 ;
        RECT 640.950 187.950 643.050 188.400 ;
        RECT 670.950 187.950 673.050 188.400 ;
        RECT 697.950 189.600 700.050 190.050 ;
        RECT 709.950 189.600 712.050 190.050 ;
        RECT 697.950 188.400 712.050 189.600 ;
        RECT 697.950 187.950 700.050 188.400 ;
        RECT 709.950 187.950 712.050 188.400 ;
        RECT 718.950 189.600 721.050 190.050 ;
        RECT 730.950 189.600 733.050 190.050 ;
        RECT 718.950 188.400 733.050 189.600 ;
        RECT 718.950 187.950 721.050 188.400 ;
        RECT 730.950 187.950 733.050 188.400 ;
        RECT 736.950 189.600 739.050 190.050 ;
        RECT 766.950 189.600 769.050 190.050 ;
        RECT 736.950 188.400 769.050 189.600 ;
        RECT 736.950 187.950 739.050 188.400 ;
        RECT 766.950 187.950 769.050 188.400 ;
        RECT 820.950 189.600 823.050 190.050 ;
        RECT 847.950 189.600 850.050 190.050 ;
        RECT 820.950 188.400 850.050 189.600 ;
        RECT 820.950 187.950 823.050 188.400 ;
        RECT 847.950 187.950 850.050 188.400 ;
        RECT 856.950 189.600 859.050 190.050 ;
        RECT 871.950 189.600 874.050 190.050 ;
        RECT 856.950 188.400 874.050 189.600 ;
        RECT 856.950 187.950 859.050 188.400 ;
        RECT 871.950 187.950 874.050 188.400 ;
        RECT 37.950 186.600 40.050 187.050 ;
        RECT 43.950 186.600 46.050 187.050 ;
        RECT 70.950 186.600 73.050 187.050 ;
        RECT 37.950 185.400 73.050 186.600 ;
        RECT 37.950 184.950 40.050 185.400 ;
        RECT 43.950 184.950 46.050 185.400 ;
        RECT 70.950 184.950 73.050 185.400 ;
        RECT 85.950 186.600 88.050 187.050 ;
        RECT 124.950 186.600 127.050 187.050 ;
        RECT 85.950 185.400 127.050 186.600 ;
        RECT 85.950 184.950 88.050 185.400 ;
        RECT 124.950 184.950 127.050 185.400 ;
        RECT 178.950 186.600 181.050 187.050 ;
        RECT 208.950 186.600 211.050 187.050 ;
        RECT 178.950 185.400 211.050 186.600 ;
        RECT 178.950 184.950 181.050 185.400 ;
        RECT 208.950 184.950 211.050 185.400 ;
        RECT 235.950 186.600 238.050 187.050 ;
        RECT 241.950 186.600 244.050 187.050 ;
        RECT 235.950 185.400 244.050 186.600 ;
        RECT 235.950 184.950 238.050 185.400 ;
        RECT 241.950 184.950 244.050 185.400 ;
        RECT 259.950 186.600 262.050 187.050 ;
        RECT 268.950 186.600 271.050 187.050 ;
        RECT 259.950 185.400 271.050 186.600 ;
        RECT 259.950 184.950 262.050 185.400 ;
        RECT 268.950 184.950 271.050 185.400 ;
        RECT 322.950 186.600 325.050 187.050 ;
        RECT 337.950 186.600 340.050 187.050 ;
        RECT 322.950 185.400 340.050 186.600 ;
        RECT 322.950 184.950 325.050 185.400 ;
        RECT 337.950 184.950 340.050 185.400 ;
        RECT 415.950 186.600 418.050 187.050 ;
        RECT 448.950 186.600 451.050 187.050 ;
        RECT 415.950 185.400 451.050 186.600 ;
        RECT 415.950 184.950 418.050 185.400 ;
        RECT 448.950 184.950 451.050 185.400 ;
        RECT 466.950 186.600 469.050 187.050 ;
        RECT 481.950 186.600 484.050 187.050 ;
        RECT 466.950 185.400 484.050 186.600 ;
        RECT 466.950 184.950 469.050 185.400 ;
        RECT 481.950 184.950 484.050 185.400 ;
        RECT 502.950 186.600 505.050 187.050 ;
        RECT 508.950 186.600 511.050 187.050 ;
        RECT 502.950 185.400 511.050 186.600 ;
        RECT 502.950 184.950 505.050 185.400 ;
        RECT 508.950 184.950 511.050 185.400 ;
        RECT 523.950 186.600 526.050 187.050 ;
        RECT 550.950 186.600 553.050 187.050 ;
        RECT 556.950 186.600 559.050 187.050 ;
        RECT 523.950 185.400 559.050 186.600 ;
        RECT 523.950 184.950 526.050 185.400 ;
        RECT 550.950 184.950 553.050 185.400 ;
        RECT 556.950 184.950 559.050 185.400 ;
        RECT 685.950 186.600 688.050 187.050 ;
        RECT 712.950 186.600 715.050 187.050 ;
        RECT 685.950 185.400 720.600 186.600 ;
        RECT 685.950 184.950 688.050 185.400 ;
        RECT 712.950 184.950 715.050 185.400 ;
        RECT 55.950 183.600 58.050 184.200 ;
        RECT 67.950 183.600 70.050 184.050 ;
        RECT 55.950 182.400 70.050 183.600 ;
        RECT 55.950 182.100 58.050 182.400 ;
        RECT 67.950 181.950 70.050 182.400 ;
        RECT 88.950 183.600 91.050 184.050 ;
        RECT 97.950 183.600 100.050 184.200 ;
        RECT 88.950 182.400 100.050 183.600 ;
        RECT 88.950 181.950 91.050 182.400 ;
        RECT 97.950 182.100 100.050 182.400 ;
        RECT 130.950 183.750 133.050 184.200 ;
        RECT 142.950 183.750 145.050 184.200 ;
        RECT 130.950 182.550 145.050 183.750 ;
        RECT 130.950 182.100 133.050 182.550 ;
        RECT 142.950 182.100 145.050 182.550 ;
        RECT 184.950 183.600 187.050 184.200 ;
        RECT 199.950 183.600 202.050 184.200 ;
        RECT 184.950 182.400 202.050 183.600 ;
        RECT 184.950 182.100 187.050 182.400 ;
        RECT 199.950 182.100 202.050 182.400 ;
        RECT 223.950 183.600 226.050 184.200 ;
        RECT 232.950 183.600 235.050 184.050 ;
        RECT 223.950 182.400 235.050 183.600 ;
        RECT 223.950 182.100 226.050 182.400 ;
        RECT 232.950 181.950 235.050 182.400 ;
        RECT 247.950 183.600 250.050 184.200 ;
        RECT 256.950 183.600 259.050 184.050 ;
        RECT 247.950 182.400 259.050 183.600 ;
        RECT 247.950 182.100 250.050 182.400 ;
        RECT 256.950 181.950 259.050 182.400 ;
        RECT 274.950 183.600 277.050 184.050 ;
        RECT 283.950 183.600 286.050 184.200 ;
        RECT 274.950 182.400 286.050 183.600 ;
        RECT 274.950 181.950 277.050 182.400 ;
        RECT 283.950 182.100 286.050 182.400 ;
        RECT 289.950 183.600 292.050 184.200 ;
        RECT 301.950 183.750 304.050 184.200 ;
        RECT 310.950 183.750 313.050 184.200 ;
        RECT 301.950 183.600 313.050 183.750 ;
        RECT 289.950 182.550 313.050 183.600 ;
        RECT 289.950 182.400 304.050 182.550 ;
        RECT 289.950 182.100 292.050 182.400 ;
        RECT 301.950 182.100 304.050 182.400 ;
        RECT 310.950 182.100 313.050 182.550 ;
        RECT 316.950 183.600 319.050 184.200 ;
        RECT 325.950 183.600 328.050 184.050 ;
        RECT 316.950 182.400 328.050 183.600 ;
        RECT 316.950 182.100 319.050 182.400 ;
        RECT 325.950 181.950 328.050 182.400 ;
        RECT 358.950 183.750 361.050 184.200 ;
        RECT 364.950 183.750 367.050 184.200 ;
        RECT 358.950 183.600 367.050 183.750 ;
        RECT 388.950 183.600 391.050 184.200 ;
        RECT 358.950 182.550 391.050 183.600 ;
        RECT 358.950 182.100 361.050 182.550 ;
        RECT 364.950 182.400 391.050 182.550 ;
        RECT 364.950 182.100 367.050 182.400 ;
        RECT 388.950 182.100 391.050 182.400 ;
        RECT 394.950 183.600 397.050 184.200 ;
        RECT 400.800 183.600 402.900 184.050 ;
        RECT 394.950 182.400 402.900 183.600 ;
        RECT 394.950 182.100 397.050 182.400 ;
        RECT 400.800 181.950 402.900 182.400 ;
        RECT 403.950 183.750 406.050 184.200 ;
        RECT 409.950 183.750 412.050 184.200 ;
        RECT 403.950 182.550 412.050 183.750 ;
        RECT 403.950 182.100 406.050 182.550 ;
        RECT 409.950 182.100 412.050 182.550 ;
        RECT 445.950 183.600 448.050 184.050 ;
        RECT 457.950 183.600 460.050 184.200 ;
        RECT 484.950 183.600 487.050 184.050 ;
        RECT 517.950 183.600 520.050 184.200 ;
        RECT 445.950 182.400 487.050 183.600 ;
        RECT 445.950 181.950 448.050 182.400 ;
        RECT 457.950 182.100 460.050 182.400 ;
        RECT 484.950 181.950 487.050 182.400 ;
        RECT 512.400 182.400 520.050 183.600 ;
        RECT 85.950 180.600 88.050 181.050 ;
        RECT 322.950 180.600 325.050 181.050 ;
        RECT 512.400 180.600 513.600 182.400 ;
        RECT 517.950 182.100 520.050 182.400 ;
        RECT 538.950 183.750 541.050 184.200 ;
        RECT 544.950 183.750 547.050 184.200 ;
        RECT 538.950 183.600 547.050 183.750 ;
        RECT 562.950 183.600 565.050 184.200 ;
        RECT 538.950 182.550 565.050 183.600 ;
        RECT 538.950 182.100 541.050 182.550 ;
        RECT 544.950 182.400 565.050 182.550 ;
        RECT 544.950 182.100 547.050 182.400 ;
        RECT 562.950 182.100 565.050 182.400 ;
        RECT 592.950 183.600 595.050 184.200 ;
        RECT 598.950 183.600 601.050 184.050 ;
        RECT 604.950 183.600 607.050 184.050 ;
        RECT 592.950 182.400 607.050 183.600 ;
        RECT 592.950 182.100 595.050 182.400 ;
        RECT 598.950 181.950 601.050 182.400 ;
        RECT 604.950 181.950 607.050 182.400 ;
        RECT 646.950 183.600 649.050 184.200 ;
        RECT 664.950 183.600 667.050 184.050 ;
        RECT 646.950 182.400 667.050 183.600 ;
        RECT 646.950 182.100 649.050 182.400 ;
        RECT 664.950 181.950 667.050 182.400 ;
        RECT 703.950 183.600 706.050 184.200 ;
        RECT 719.400 183.600 720.600 185.400 ;
        RECT 751.950 183.600 754.050 184.200 ;
        RECT 703.950 182.400 711.600 183.600 ;
        RECT 719.400 182.400 754.050 183.600 ;
        RECT 703.950 182.100 706.050 182.400 ;
        RECT 59.400 179.400 88.050 180.600 ;
        RECT 19.950 177.450 22.050 177.900 ;
        RECT 28.950 177.450 31.050 177.900 ;
        RECT 19.950 176.250 31.050 177.450 ;
        RECT 19.950 175.800 22.050 176.250 ;
        RECT 28.950 175.800 31.050 176.250 ;
        RECT 34.950 177.600 37.050 177.900 ;
        RECT 46.950 177.600 49.050 178.050 ;
        RECT 59.400 177.900 60.600 179.400 ;
        RECT 85.950 178.950 88.050 179.400 ;
        RECT 293.400 179.400 325.050 180.600 ;
        RECT 506.400 180.000 513.600 180.600 ;
        RECT 34.950 176.400 49.050 177.600 ;
        RECT 34.950 175.800 37.050 176.400 ;
        RECT 46.950 175.950 49.050 176.400 ;
        RECT 58.950 175.800 61.050 177.900 ;
        RECT 67.950 177.450 70.050 177.900 ;
        RECT 73.950 177.450 76.050 177.900 ;
        RECT 67.950 176.250 76.050 177.450 ;
        RECT 67.950 175.800 70.050 176.250 ;
        RECT 73.950 175.800 76.050 176.250 ;
        RECT 106.950 177.450 109.050 177.900 ;
        RECT 118.950 177.450 121.050 177.900 ;
        RECT 106.950 176.250 121.050 177.450 ;
        RECT 106.950 175.800 109.050 176.250 ;
        RECT 118.950 175.800 121.050 176.250 ;
        RECT 160.950 175.800 163.050 177.900 ;
        RECT 181.950 177.600 184.050 177.900 ;
        RECT 190.950 177.600 193.050 178.050 ;
        RECT 181.950 176.400 193.050 177.600 ;
        RECT 181.950 175.800 184.050 176.400 ;
        RECT 190.950 175.950 193.050 176.400 ;
        RECT 202.950 177.600 205.050 177.900 ;
        RECT 208.950 177.600 211.050 178.050 ;
        RECT 202.950 176.400 211.050 177.600 ;
        RECT 202.950 175.800 205.050 176.400 ;
        RECT 208.950 175.950 211.050 176.400 ;
        RECT 235.950 177.450 238.050 177.900 ;
        RECT 244.950 177.450 247.050 177.900 ;
        RECT 235.950 176.250 247.050 177.450 ;
        RECT 235.950 175.800 238.050 176.250 ;
        RECT 244.950 175.800 247.050 176.250 ;
        RECT 265.950 177.600 268.050 177.900 ;
        RECT 277.950 177.600 280.050 178.050 ;
        RECT 293.400 177.900 294.600 179.400 ;
        RECT 314.400 177.900 315.600 179.400 ;
        RECT 322.950 178.950 325.050 179.400 ;
        RECT 505.950 179.400 513.600 180.000 ;
        RECT 265.950 176.400 280.050 177.600 ;
        RECT 265.950 175.800 268.050 176.400 ;
        RECT 277.950 175.950 280.050 176.400 ;
        RECT 292.950 175.800 295.050 177.900 ;
        RECT 313.950 175.800 316.050 177.900 ;
        RECT 343.950 177.600 346.050 177.900 ;
        RECT 358.950 177.600 361.050 178.050 ;
        RECT 343.950 176.400 361.050 177.600 ;
        RECT 343.950 175.800 346.050 176.400 ;
        RECT 358.950 175.950 361.050 176.400 ;
        RECT 412.950 177.600 415.050 177.900 ;
        RECT 433.950 177.600 436.050 177.900 ;
        RECT 412.950 176.400 436.050 177.600 ;
        RECT 412.950 175.800 415.050 176.400 ;
        RECT 433.950 175.800 436.050 176.400 ;
        RECT 439.950 177.450 442.050 177.900 ;
        RECT 445.950 177.450 448.050 177.900 ;
        RECT 439.950 176.250 448.050 177.450 ;
        RECT 439.950 175.800 442.050 176.250 ;
        RECT 445.950 175.800 448.050 176.250 ;
        RECT 478.950 177.600 481.050 177.900 ;
        RECT 487.950 177.600 490.050 178.050 ;
        RECT 493.950 177.600 496.050 177.900 ;
        RECT 478.950 176.400 496.050 177.600 ;
        RECT 478.950 175.800 481.050 176.400 ;
        RECT 487.950 175.950 490.050 176.400 ;
        RECT 493.950 175.800 496.050 176.400 ;
        RECT 505.950 175.950 508.050 179.400 ;
        RECT 710.400 178.050 711.600 182.400 ;
        RECT 751.950 182.100 754.050 182.400 ;
        RECT 757.950 182.100 760.050 184.200 ;
        RECT 781.950 183.600 784.050 184.200 ;
        RECT 767.400 182.400 784.050 183.600 ;
        RECT 758.400 180.600 759.600 182.100 ;
        RECT 767.400 180.600 768.600 182.400 ;
        RECT 781.950 182.100 784.050 182.400 ;
        RECT 799.950 183.600 802.050 184.200 ;
        RECT 805.950 183.600 808.050 184.200 ;
        RECT 817.950 183.600 820.050 184.050 ;
        RECT 799.950 182.400 804.600 183.600 ;
        RECT 799.950 182.100 802.050 182.400 ;
        RECT 758.400 179.400 768.600 180.600 ;
        RECT 803.400 180.600 804.600 182.400 ;
        RECT 805.950 182.400 820.050 183.600 ;
        RECT 805.950 182.100 808.050 182.400 ;
        RECT 817.950 181.950 820.050 182.400 ;
        RECT 826.950 183.600 829.050 184.200 ;
        RECT 832.950 183.600 835.050 187.050 ;
        RECT 826.950 183.000 835.050 183.600 ;
        RECT 859.950 183.600 862.050 184.050 ;
        RECT 898.950 183.600 901.050 184.050 ;
        RECT 826.950 182.400 834.600 183.000 ;
        RECT 859.950 182.400 901.050 183.600 ;
        RECT 826.950 182.100 829.050 182.400 ;
        RECT 859.950 181.950 862.050 182.400 ;
        RECT 898.950 181.950 901.050 182.400 ;
        RECT 856.950 180.600 859.050 180.900 ;
        RECT 803.400 179.400 859.050 180.600 ;
        RECT 526.950 177.450 529.050 177.900 ;
        RECT 532.950 177.450 535.050 177.900 ;
        RECT 526.950 176.250 535.050 177.450 ;
        RECT 526.950 175.800 529.050 176.250 ;
        RECT 532.950 175.800 535.050 176.250 ;
        RECT 631.950 177.450 634.050 177.900 ;
        RECT 637.950 177.450 640.050 177.900 ;
        RECT 631.950 176.250 640.050 177.450 ;
        RECT 631.950 175.800 634.050 176.250 ;
        RECT 637.950 175.800 640.050 176.250 ;
        RECT 643.950 177.600 646.050 177.900 ;
        RECT 667.950 177.600 670.050 177.900 ;
        RECT 643.950 176.400 670.050 177.600 ;
        RECT 710.400 176.400 715.050 178.050 ;
        RECT 643.950 175.800 646.050 176.400 ;
        RECT 667.950 175.800 670.050 176.400 ;
        RECT 711.000 175.950 715.050 176.400 ;
        RECT 724.950 177.450 727.050 177.900 ;
        RECT 730.950 177.450 733.050 177.900 ;
        RECT 724.950 176.250 733.050 177.450 ;
        RECT 724.950 175.800 727.050 176.250 ;
        RECT 730.950 175.800 733.050 176.250 ;
        RECT 736.950 177.600 739.050 177.900 ;
        RECT 758.400 177.600 759.600 179.400 ;
        RECT 856.950 178.800 859.050 179.400 ;
        RECT 736.950 176.400 759.600 177.600 ;
        RECT 769.950 177.600 772.050 178.050 ;
        RECT 787.950 177.600 790.050 178.050 ;
        RECT 769.950 176.400 790.050 177.600 ;
        RECT 736.950 175.800 739.050 176.400 ;
        RECT 769.950 175.950 772.050 176.400 ;
        RECT 787.950 175.950 790.050 176.400 ;
        RECT 817.950 177.450 820.050 177.900 ;
        RECT 829.950 177.450 832.050 177.900 ;
        RECT 817.950 176.250 832.050 177.450 ;
        RECT 817.950 175.800 820.050 176.250 ;
        RECT 829.950 175.800 832.050 176.250 ;
        RECT 127.950 171.600 130.050 172.050 ;
        RECT 161.400 171.600 162.600 175.800 ;
        RECT 220.950 174.600 223.050 175.050 ;
        RECT 236.400 174.600 237.600 175.800 ;
        RECT 220.950 173.400 237.600 174.600 ;
        RECT 556.950 174.600 559.050 175.050 ;
        RECT 583.950 174.600 586.050 175.050 ;
        RECT 556.950 173.400 586.050 174.600 ;
        RECT 220.950 172.950 223.050 173.400 ;
        RECT 556.950 172.950 559.050 173.400 ;
        RECT 583.950 172.950 586.050 173.400 ;
        RECT 589.950 174.600 592.050 175.050 ;
        RECT 601.950 174.600 604.050 175.050 ;
        RECT 589.950 173.400 604.050 174.600 ;
        RECT 589.950 172.950 592.050 173.400 ;
        RECT 601.950 172.950 604.050 173.400 ;
        RECT 760.950 174.600 763.050 175.050 ;
        RECT 778.950 174.600 781.050 175.050 ;
        RECT 790.950 174.600 793.050 175.050 ;
        RECT 760.950 173.400 793.050 174.600 ;
        RECT 760.950 172.950 763.050 173.400 ;
        RECT 778.950 172.950 781.050 173.400 ;
        RECT 790.950 172.950 793.050 173.400 ;
        RECT 199.950 171.600 202.050 172.050 ;
        RECT 127.950 170.400 202.050 171.600 ;
        RECT 127.950 169.950 130.050 170.400 ;
        RECT 199.950 169.950 202.050 170.400 ;
        RECT 370.950 171.600 373.050 172.050 ;
        RECT 385.950 171.600 388.050 172.050 ;
        RECT 403.950 171.600 406.050 172.050 ;
        RECT 460.950 171.600 463.050 172.050 ;
        RECT 370.950 170.400 463.050 171.600 ;
        RECT 370.950 169.950 373.050 170.400 ;
        RECT 385.950 169.950 388.050 170.400 ;
        RECT 403.950 169.950 406.050 170.400 ;
        RECT 460.950 169.950 463.050 170.400 ;
        RECT 520.950 171.600 523.050 172.050 ;
        RECT 565.950 171.600 568.050 172.050 ;
        RECT 520.950 170.400 568.050 171.600 ;
        RECT 520.950 169.950 523.050 170.400 ;
        RECT 565.950 169.950 568.050 170.400 ;
        RECT 694.950 171.600 697.050 172.050 ;
        RECT 724.950 171.600 727.050 172.050 ;
        RECT 694.950 170.400 727.050 171.600 ;
        RECT 694.950 169.950 697.050 170.400 ;
        RECT 724.950 169.950 727.050 170.400 ;
        RECT 730.950 171.600 733.050 172.050 ;
        RECT 745.950 171.600 748.050 172.050 ;
        RECT 730.950 170.400 748.050 171.600 ;
        RECT 730.950 169.950 733.050 170.400 ;
        RECT 745.950 169.950 748.050 170.400 ;
        RECT 226.950 168.600 229.050 169.050 ;
        RECT 259.950 168.600 262.050 169.050 ;
        RECT 328.950 168.600 331.050 169.050 ;
        RECT 361.950 168.600 364.050 169.050 ;
        RECT 226.950 167.400 364.050 168.600 ;
        RECT 226.950 166.950 229.050 167.400 ;
        RECT 259.950 166.950 262.050 167.400 ;
        RECT 328.950 166.950 331.050 167.400 ;
        RECT 361.950 166.950 364.050 167.400 ;
        RECT 607.950 168.600 610.050 169.050 ;
        RECT 625.950 168.600 628.050 169.050 ;
        RECT 607.950 167.400 628.050 168.600 ;
        RECT 607.950 166.950 610.050 167.400 ;
        RECT 625.950 166.950 628.050 167.400 ;
        RECT 844.950 168.600 847.050 169.050 ;
        RECT 859.950 168.600 862.050 169.050 ;
        RECT 844.950 167.400 862.050 168.600 ;
        RECT 844.950 166.950 847.050 167.400 ;
        RECT 859.950 166.950 862.050 167.400 ;
        RECT 232.950 165.600 235.050 166.050 ;
        RECT 286.950 165.600 289.050 166.050 ;
        RECT 307.950 165.600 310.050 166.050 ;
        RECT 232.950 164.400 310.050 165.600 ;
        RECT 232.950 163.950 235.050 164.400 ;
        RECT 286.950 163.950 289.050 164.400 ;
        RECT 307.950 163.950 310.050 164.400 ;
        RECT 508.950 165.600 511.050 166.050 ;
        RECT 730.950 165.600 733.050 166.050 ;
        RECT 508.950 164.400 733.050 165.600 ;
        RECT 508.950 163.950 511.050 164.400 ;
        RECT 730.950 163.950 733.050 164.400 ;
        RECT 736.950 165.600 739.050 166.050 ;
        RECT 778.950 165.600 781.050 166.050 ;
        RECT 736.950 164.400 781.050 165.600 ;
        RECT 736.950 163.950 739.050 164.400 ;
        RECT 778.950 163.950 781.050 164.400 ;
        RECT 808.950 165.600 811.050 166.050 ;
        RECT 853.950 165.600 856.050 166.050 ;
        RECT 874.950 165.600 877.050 166.050 ;
        RECT 808.950 164.400 877.050 165.600 ;
        RECT 808.950 163.950 811.050 164.400 ;
        RECT 853.950 163.950 856.050 164.400 ;
        RECT 874.950 163.950 877.050 164.400 ;
        RECT 892.950 165.600 895.050 166.050 ;
        RECT 898.950 165.600 901.050 166.050 ;
        RECT 892.950 164.400 901.050 165.600 ;
        RECT 892.950 163.950 895.050 164.400 ;
        RECT 898.950 163.950 901.050 164.400 ;
        RECT 139.950 162.600 142.050 163.050 ;
        RECT 169.950 162.600 172.050 163.050 ;
        RECT 139.950 161.400 172.050 162.600 ;
        RECT 139.950 160.950 142.050 161.400 ;
        RECT 169.950 160.950 172.050 161.400 ;
        RECT 577.950 162.600 580.050 163.050 ;
        RECT 607.950 162.600 610.050 163.050 ;
        RECT 577.950 161.400 610.050 162.600 ;
        RECT 577.950 160.950 580.050 161.400 ;
        RECT 607.950 160.950 610.050 161.400 ;
        RECT 265.950 159.600 268.050 160.050 ;
        RECT 280.950 159.600 283.050 160.050 ;
        RECT 298.950 159.600 301.050 160.050 ;
        RECT 265.950 158.400 301.050 159.600 ;
        RECT 265.950 157.950 268.050 158.400 ;
        RECT 280.950 157.950 283.050 158.400 ;
        RECT 298.950 157.950 301.050 158.400 ;
        RECT 676.950 159.600 679.050 160.050 ;
        RECT 718.950 159.600 721.050 160.050 ;
        RECT 793.950 159.600 796.050 160.050 ;
        RECT 676.950 158.400 796.050 159.600 ;
        RECT 676.950 157.950 679.050 158.400 ;
        RECT 718.950 157.950 721.050 158.400 ;
        RECT 793.950 157.950 796.050 158.400 ;
        RECT 142.950 156.600 145.050 157.050 ;
        RECT 151.950 156.600 154.050 157.050 ;
        RECT 142.950 155.400 154.050 156.600 ;
        RECT 142.950 154.950 145.050 155.400 ;
        RECT 151.950 154.950 154.050 155.400 ;
        RECT 253.950 156.600 256.050 157.050 ;
        RECT 406.950 156.600 409.050 157.050 ;
        RECT 253.950 155.400 409.050 156.600 ;
        RECT 253.950 154.950 256.050 155.400 ;
        RECT 406.950 154.950 409.050 155.400 ;
        RECT 547.950 156.600 550.050 157.050 ;
        RECT 610.950 156.600 613.050 157.050 ;
        RECT 547.950 155.400 613.050 156.600 ;
        RECT 547.950 154.950 550.050 155.400 ;
        RECT 610.950 154.950 613.050 155.400 ;
        RECT 721.950 156.600 724.050 157.050 ;
        RECT 739.950 156.600 742.050 157.050 ;
        RECT 721.950 155.400 742.050 156.600 ;
        RECT 721.950 154.950 724.050 155.400 ;
        RECT 739.950 154.950 742.050 155.400 ;
        RECT 757.950 156.600 760.050 157.050 ;
        RECT 784.950 156.600 787.050 157.050 ;
        RECT 757.950 155.400 787.050 156.600 ;
        RECT 757.950 154.950 760.050 155.400 ;
        RECT 784.950 154.950 787.050 155.400 ;
        RECT 706.950 153.600 709.050 154.050 ;
        RECT 748.950 153.600 751.050 154.050 ;
        RECT 706.950 152.400 751.050 153.600 ;
        RECT 706.950 151.950 709.050 152.400 ;
        RECT 748.950 151.950 751.050 152.400 ;
        RECT 274.950 150.600 277.050 151.050 ;
        RECT 307.950 150.600 310.050 151.050 ;
        RECT 274.950 149.400 310.050 150.600 ;
        RECT 274.950 148.950 277.050 149.400 ;
        RECT 307.950 148.950 310.050 149.400 ;
        RECT 319.950 150.600 322.050 151.050 ;
        RECT 352.950 150.600 355.050 151.050 ;
        RECT 319.950 149.400 355.050 150.600 ;
        RECT 319.950 148.950 322.050 149.400 ;
        RECT 352.950 148.950 355.050 149.400 ;
        RECT 484.950 150.600 487.050 151.050 ;
        RECT 520.950 150.600 523.050 151.050 ;
        RECT 484.950 149.400 523.050 150.600 ;
        RECT 484.950 148.950 487.050 149.400 ;
        RECT 520.950 148.950 523.050 149.400 ;
        RECT 526.950 150.600 529.050 151.050 ;
        RECT 589.950 150.600 592.050 151.050 ;
        RECT 526.950 149.400 592.050 150.600 ;
        RECT 526.950 148.950 529.050 149.400 ;
        RECT 589.950 148.950 592.050 149.400 ;
        RECT 652.950 150.600 655.050 151.050 ;
        RECT 694.950 150.600 697.050 151.050 ;
        RECT 652.950 149.400 697.050 150.600 ;
        RECT 652.950 148.950 655.050 149.400 ;
        RECT 694.950 148.950 697.050 149.400 ;
        RECT 787.950 150.600 790.050 151.050 ;
        RECT 808.950 150.600 811.050 151.050 ;
        RECT 787.950 149.400 811.050 150.600 ;
        RECT 787.950 148.950 790.050 149.400 ;
        RECT 808.950 148.950 811.050 149.400 ;
        RECT 829.950 150.600 832.050 151.050 ;
        RECT 838.800 150.600 840.900 151.050 ;
        RECT 829.950 149.400 840.900 150.600 ;
        RECT 829.950 148.950 832.050 149.400 ;
        RECT 838.800 148.950 840.900 149.400 ;
        RECT 841.950 150.600 844.050 151.050 ;
        RECT 862.950 150.600 865.050 151.050 ;
        RECT 841.950 149.400 865.050 150.600 ;
        RECT 841.950 148.950 844.050 149.400 ;
        RECT 862.950 148.950 865.050 149.400 ;
        RECT 277.950 147.600 280.050 148.050 ;
        RECT 337.950 147.600 340.050 148.050 ;
        RECT 277.950 146.400 340.050 147.600 ;
        RECT 277.950 145.950 280.050 146.400 ;
        RECT 337.950 145.950 340.050 146.400 ;
        RECT 406.950 147.600 409.050 148.050 ;
        RECT 505.950 147.600 508.050 148.050 ;
        RECT 406.950 146.400 508.050 147.600 ;
        RECT 406.950 145.950 409.050 146.400 ;
        RECT 505.950 145.950 508.050 146.400 ;
        RECT 592.950 147.600 595.050 148.050 ;
        RECT 712.950 147.600 715.050 148.050 ;
        RECT 721.950 147.600 724.050 148.050 ;
        RECT 592.950 146.400 648.600 147.600 ;
        RECT 592.950 145.950 595.050 146.400 ;
        RECT 647.400 145.050 648.600 146.400 ;
        RECT 712.950 146.400 724.050 147.600 ;
        RECT 712.950 145.950 715.050 146.400 ;
        RECT 721.950 145.950 724.050 146.400 ;
        RECT 112.950 144.600 115.050 145.050 ;
        RECT 142.950 144.600 145.050 145.050 ;
        RECT 112.950 143.400 145.050 144.600 ;
        RECT 112.950 142.950 115.050 143.400 ;
        RECT 142.950 142.950 145.050 143.400 ;
        RECT 247.950 144.600 250.050 145.050 ;
        RECT 271.950 144.600 274.050 145.050 ;
        RECT 247.950 143.400 274.050 144.600 ;
        RECT 247.950 142.950 250.050 143.400 ;
        RECT 271.950 142.950 274.050 143.400 ;
        RECT 286.950 144.600 289.050 145.050 ;
        RECT 328.950 144.600 331.050 145.050 ;
        RECT 286.950 143.400 331.050 144.600 ;
        RECT 286.950 142.950 289.050 143.400 ;
        RECT 328.950 142.950 331.050 143.400 ;
        RECT 343.950 144.600 346.050 145.050 ;
        RECT 478.950 144.600 481.050 145.050 ;
        RECT 343.950 143.400 481.050 144.600 ;
        RECT 343.950 142.950 346.050 143.400 ;
        RECT 478.950 142.950 481.050 143.400 ;
        RECT 490.950 144.600 493.050 145.050 ;
        RECT 526.950 144.600 529.050 145.050 ;
        RECT 490.950 143.400 529.050 144.600 ;
        RECT 490.950 142.950 493.050 143.400 ;
        RECT 526.950 142.950 529.050 143.400 ;
        RECT 646.950 144.600 649.050 145.050 ;
        RECT 682.950 144.600 685.050 145.050 ;
        RECT 646.950 143.400 685.050 144.600 ;
        RECT 646.950 142.950 649.050 143.400 ;
        RECT 682.950 142.950 685.050 143.400 ;
        RECT 739.950 144.600 742.050 145.050 ;
        RECT 772.950 144.600 775.050 145.050 ;
        RECT 739.950 143.400 775.050 144.600 ;
        RECT 739.950 142.950 742.050 143.400 ;
        RECT 772.950 142.950 775.050 143.400 ;
        RECT 790.950 144.600 793.050 145.050 ;
        RECT 817.950 144.600 820.050 145.050 ;
        RECT 790.950 143.400 820.050 144.600 ;
        RECT 790.950 142.950 793.050 143.400 ;
        RECT 817.950 142.950 820.050 143.400 ;
        RECT 832.950 144.600 835.050 145.050 ;
        RECT 832.950 143.400 849.600 144.600 ;
        RECT 832.950 142.950 835.050 143.400 ;
        RECT 848.400 142.050 849.600 143.400 ;
        RECT 256.950 141.600 259.050 142.050 ;
        RECT 289.950 141.600 292.050 142.050 ;
        RECT 313.950 141.600 316.050 142.050 ;
        RECT 256.950 140.400 316.050 141.600 ;
        RECT 256.950 139.950 259.050 140.400 ;
        RECT 289.950 139.950 292.050 140.400 ;
        RECT 313.950 139.950 316.050 140.400 ;
        RECT 847.950 141.600 850.050 142.050 ;
        RECT 856.950 141.600 859.050 142.050 ;
        RECT 847.950 140.400 859.050 141.600 ;
        RECT 847.950 139.950 850.050 140.400 ;
        RECT 856.950 139.950 859.050 140.400 ;
        RECT 58.950 138.750 61.050 139.200 ;
        RECT 70.950 138.750 73.050 139.200 ;
        RECT 58.950 137.550 73.050 138.750 ;
        RECT 58.950 137.100 61.050 137.550 ;
        RECT 70.950 137.100 73.050 137.550 ;
        RECT 88.950 138.600 91.050 139.200 ;
        RECT 106.950 138.600 109.050 139.200 ;
        RECT 121.950 138.600 124.050 139.050 ;
        RECT 88.950 137.400 124.050 138.600 ;
        RECT 88.950 137.100 91.050 137.400 ;
        RECT 106.950 137.100 109.050 137.400 ;
        RECT 121.950 136.950 124.050 137.400 ;
        RECT 130.950 138.600 133.050 139.200 ;
        RECT 145.950 138.600 148.050 139.050 ;
        RECT 130.950 137.400 148.050 138.600 ;
        RECT 130.950 137.100 133.050 137.400 ;
        RECT 145.950 136.950 148.050 137.400 ;
        RECT 160.950 138.750 163.050 139.200 ;
        RECT 169.950 138.750 172.050 139.200 ;
        RECT 160.950 137.550 172.050 138.750 ;
        RECT 160.950 137.100 163.050 137.550 ;
        RECT 169.950 137.100 172.050 137.550 ;
        RECT 175.950 138.750 178.050 139.200 ;
        RECT 184.950 138.750 187.050 139.200 ;
        RECT 175.950 137.550 187.050 138.750 ;
        RECT 175.950 137.100 178.050 137.550 ;
        RECT 184.950 137.100 187.050 137.550 ;
        RECT 193.950 136.950 196.050 139.050 ;
        RECT 211.950 138.600 214.050 139.050 ;
        RECT 220.950 138.600 223.050 139.200 ;
        RECT 211.950 137.400 223.050 138.600 ;
        RECT 211.950 136.950 214.050 137.400 ;
        RECT 220.950 137.100 223.050 137.400 ;
        RECT 232.950 138.750 235.050 139.200 ;
        RECT 241.950 138.750 244.050 139.200 ;
        RECT 232.950 137.550 244.050 138.750 ;
        RECT 232.950 137.100 235.050 137.550 ;
        RECT 241.950 137.100 244.050 137.550 ;
        RECT 271.950 138.750 274.050 139.200 ;
        RECT 277.950 138.750 280.050 139.200 ;
        RECT 271.950 137.550 280.050 138.750 ;
        RECT 271.950 137.100 274.050 137.550 ;
        RECT 277.950 137.100 280.050 137.550 ;
        RECT 295.950 138.600 298.050 139.200 ;
        RECT 319.950 138.600 322.050 139.200 ;
        RECT 295.950 137.400 322.050 138.600 ;
        RECT 295.950 137.100 298.050 137.400 ;
        RECT 319.950 137.100 322.050 137.400 ;
        RECT 343.950 137.100 346.050 139.200 ;
        RECT 370.950 138.600 373.050 139.200 ;
        RECT 385.950 138.600 388.050 139.200 ;
        RECT 370.950 137.400 388.050 138.600 ;
        RECT 370.950 137.100 373.050 137.400 ;
        RECT 385.950 137.100 388.050 137.400 ;
        RECT 412.950 138.750 415.050 139.200 ;
        RECT 418.950 138.750 421.050 139.200 ;
        RECT 412.950 137.550 421.050 138.750 ;
        RECT 412.950 137.100 415.050 137.550 ;
        RECT 418.950 137.100 421.050 137.550 ;
        RECT 433.950 138.750 436.050 139.200 ;
        RECT 442.950 138.750 445.050 139.200 ;
        RECT 433.950 137.550 445.050 138.750 ;
        RECT 433.950 137.100 436.050 137.550 ;
        RECT 442.950 137.100 445.050 137.550 ;
        RECT 448.950 137.100 451.050 139.200 ;
        RECT 454.950 138.750 457.050 139.200 ;
        RECT 460.950 138.750 463.050 139.200 ;
        RECT 454.950 137.550 463.050 138.750 ;
        RECT 454.950 137.100 457.050 137.550 ;
        RECT 460.950 137.100 463.050 137.550 ;
        RECT 466.950 138.600 469.050 139.050 ;
        RECT 472.950 138.750 475.050 139.200 ;
        RECT 493.950 138.750 496.050 139.200 ;
        RECT 472.950 138.600 496.050 138.750 ;
        RECT 466.950 137.550 496.050 138.600 ;
        RECT 466.950 137.400 475.050 137.550 ;
        RECT 194.400 135.600 195.600 136.950 ;
        RECT 344.400 135.600 345.600 137.100 ;
        RECT 449.400 135.600 450.600 137.100 ;
        RECT 466.950 136.950 469.050 137.400 ;
        RECT 472.950 137.100 475.050 137.400 ;
        RECT 493.950 137.100 496.050 137.550 ;
        RECT 505.950 138.600 508.050 139.200 ;
        RECT 517.950 138.600 520.050 139.050 ;
        RECT 505.950 137.400 520.050 138.600 ;
        RECT 505.950 137.100 508.050 137.400 ;
        RECT 517.950 136.950 520.050 137.400 ;
        RECT 547.950 136.950 550.050 139.050 ;
        RECT 568.950 137.100 571.050 139.200 ;
        RECT 574.950 138.600 577.050 139.200 ;
        RECT 592.950 138.600 595.050 139.200 ;
        RECT 574.950 137.400 595.050 138.600 ;
        RECT 574.950 137.100 577.050 137.400 ;
        RECT 592.950 137.100 595.050 137.400 ;
        RECT 652.950 138.750 655.050 139.200 ;
        RECT 661.950 138.750 664.050 139.200 ;
        RECT 652.950 137.550 664.050 138.750 ;
        RECT 652.950 137.100 655.050 137.550 ;
        RECT 661.950 137.100 664.050 137.550 ;
        RECT 673.950 138.750 676.050 139.200 ;
        RECT 685.950 138.750 688.050 139.200 ;
        RECT 673.950 137.550 688.050 138.750 ;
        RECT 673.950 137.100 676.050 137.550 ;
        RECT 685.950 137.100 688.050 137.550 ;
        RECT 703.950 138.750 706.050 139.200 ;
        RECT 709.950 138.750 712.050 139.200 ;
        RECT 703.950 137.550 712.050 138.750 ;
        RECT 703.950 137.100 706.050 137.550 ;
        RECT 709.950 137.100 712.050 137.550 ;
        RECT 727.950 137.100 730.050 139.200 ;
        RECT 742.950 138.600 745.050 139.200 ;
        RECT 766.950 138.600 769.050 139.200 ;
        RECT 787.950 138.600 790.050 139.200 ;
        RECT 742.950 137.400 790.050 138.600 ;
        RECT 742.950 137.100 745.050 137.400 ;
        RECT 766.950 137.100 769.050 137.400 ;
        RECT 787.950 137.100 790.050 137.400 ;
        RECT 823.950 137.100 826.050 139.200 ;
        RECT 835.950 138.750 838.050 139.200 ;
        RECT 841.950 138.750 844.050 139.200 ;
        RECT 835.950 137.550 844.050 138.750 ;
        RECT 835.950 137.100 838.050 137.550 ;
        RECT 841.950 137.100 844.050 137.550 ;
        RECT 868.950 138.600 871.050 139.200 ;
        RECT 889.950 138.600 892.050 139.200 ;
        RECT 868.950 137.400 892.050 138.600 ;
        RECT 868.950 137.100 871.050 137.400 ;
        RECT 889.950 137.100 892.050 137.400 ;
        RECT 463.950 135.600 466.050 136.050 ;
        RECT 194.400 134.400 204.600 135.600 ;
        RECT 344.400 134.400 357.600 135.600 ;
        RECT 449.400 134.400 466.050 135.600 ;
        RECT 548.400 135.600 549.600 136.950 ;
        RECT 569.400 135.600 570.600 137.100 ;
        RECT 583.950 135.600 586.050 136.050 ;
        RECT 548.400 134.400 586.050 135.600 ;
        RECT 73.950 132.450 76.050 132.900 ;
        RECT 85.950 132.450 88.050 132.900 ;
        RECT 73.950 131.250 88.050 132.450 ;
        RECT 73.950 130.800 76.050 131.250 ;
        RECT 85.950 130.800 88.050 131.250 ;
        RECT 109.950 132.600 112.050 132.900 ;
        RECT 118.950 132.600 121.050 133.050 ;
        RECT 109.950 131.400 121.050 132.600 ;
        RECT 109.950 130.800 112.050 131.400 ;
        RECT 118.950 130.950 121.050 131.400 ;
        RECT 124.950 132.600 127.050 133.050 ;
        RECT 187.950 132.600 190.050 133.050 ;
        RECT 124.950 131.400 190.050 132.600 ;
        RECT 203.400 132.600 204.600 134.400 ;
        RECT 356.400 133.050 357.600 134.400 ;
        RECT 463.950 133.950 466.050 134.400 ;
        RECT 583.950 133.950 586.050 134.400 ;
        RECT 610.950 135.600 613.050 136.050 ;
        RECT 610.950 134.400 633.600 135.600 ;
        RECT 610.950 133.950 613.050 134.400 ;
        RECT 208.950 132.600 211.050 133.050 ;
        RECT 203.400 131.400 211.050 132.600 ;
        RECT 124.950 130.950 127.050 131.400 ;
        RECT 187.950 130.950 190.050 131.400 ;
        RECT 208.950 130.950 211.050 131.400 ;
        RECT 244.950 132.450 247.050 132.900 ;
        RECT 253.950 132.450 256.050 132.900 ;
        RECT 244.950 131.250 256.050 132.450 ;
        RECT 244.950 130.800 247.050 131.250 ;
        RECT 253.950 130.800 256.050 131.250 ;
        RECT 280.950 132.450 283.050 132.900 ;
        RECT 292.950 132.600 295.050 132.900 ;
        RECT 316.950 132.600 319.050 132.900 ;
        RECT 292.950 132.450 319.050 132.600 ;
        RECT 280.950 131.400 319.050 132.450 ;
        RECT 356.400 131.400 361.050 133.050 ;
        RECT 280.950 131.250 295.050 131.400 ;
        RECT 280.950 130.800 283.050 131.250 ;
        RECT 292.950 130.800 295.050 131.250 ;
        RECT 316.950 130.800 319.050 131.400 ;
        RECT 357.000 130.950 361.050 131.400 ;
        RECT 409.950 132.450 412.050 132.900 ;
        RECT 421.950 132.450 424.050 132.900 ;
        RECT 409.950 131.250 424.050 132.450 ;
        RECT 409.950 130.800 412.050 131.250 ;
        RECT 421.950 130.800 424.050 131.250 ;
        RECT 481.950 132.450 484.050 132.900 ;
        RECT 490.950 132.450 493.050 132.900 ;
        RECT 481.950 131.250 493.050 132.450 ;
        RECT 481.950 130.800 484.050 131.250 ;
        RECT 490.950 130.800 493.050 131.250 ;
        RECT 538.950 132.600 541.050 133.050 ;
        RECT 632.400 132.900 633.600 134.400 ;
        RECT 728.400 133.050 729.600 137.100 ;
        RECT 824.400 135.600 825.600 137.100 ;
        RECT 824.400 134.400 831.600 135.600 ;
        RECT 550.950 132.600 553.050 132.900 ;
        RECT 538.950 131.400 553.050 132.600 ;
        RECT 538.950 130.950 541.050 131.400 ;
        RECT 550.950 130.800 553.050 131.400 ;
        RECT 631.950 130.800 634.050 132.900 ;
        RECT 661.950 132.600 664.050 133.050 ;
        RECT 670.950 132.600 673.050 132.900 ;
        RECT 661.950 131.400 673.050 132.600 ;
        RECT 661.950 130.950 664.050 131.400 ;
        RECT 670.950 130.800 673.050 131.400 ;
        RECT 685.950 132.600 688.050 133.050 ;
        RECT 694.950 132.600 697.050 132.900 ;
        RECT 685.950 131.400 697.050 132.600 ;
        RECT 728.400 131.400 733.050 133.050 ;
        RECT 685.950 130.950 688.050 131.400 ;
        RECT 694.950 130.800 697.050 131.400 ;
        RECT 729.000 130.950 733.050 131.400 ;
        RECT 739.950 132.450 742.050 132.900 ;
        RECT 748.950 132.450 751.050 132.900 ;
        RECT 739.950 131.250 751.050 132.450 ;
        RECT 739.950 130.800 742.050 131.250 ;
        RECT 748.950 130.800 751.050 131.250 ;
        RECT 769.950 132.600 772.050 132.900 ;
        RECT 781.950 132.600 784.050 133.050 ;
        RECT 769.950 131.400 784.050 132.600 ;
        RECT 769.950 130.800 772.050 131.400 ;
        RECT 781.950 130.950 784.050 131.400 ;
        RECT 808.950 132.600 811.050 133.050 ;
        RECT 814.950 132.600 817.050 132.900 ;
        RECT 808.950 131.400 817.050 132.600 ;
        RECT 808.950 130.950 811.050 131.400 ;
        RECT 814.950 130.800 817.050 131.400 ;
        RECT 820.950 132.450 823.050 132.900 ;
        RECT 826.950 132.450 829.050 132.900 ;
        RECT 820.950 131.250 829.050 132.450 ;
        RECT 830.400 132.600 831.600 134.400 ;
        RECT 850.950 132.600 853.050 133.050 ;
        RECT 830.400 131.400 853.050 132.600 ;
        RECT 820.950 130.800 823.050 131.250 ;
        RECT 826.950 130.800 829.050 131.250 ;
        RECT 850.950 130.950 853.050 131.400 ;
        RECT 874.950 132.450 877.050 132.900 ;
        RECT 886.950 132.450 889.050 132.900 ;
        RECT 874.950 131.250 889.050 132.450 ;
        RECT 874.950 130.800 877.050 131.250 ;
        RECT 886.950 130.800 889.050 131.250 ;
        RECT 352.950 129.600 355.050 130.050 ;
        RECT 373.950 129.600 376.050 130.050 ;
        RECT 352.950 128.400 376.050 129.600 ;
        RECT 352.950 127.950 355.050 128.400 ;
        RECT 373.950 127.950 376.050 128.400 ;
        RECT 493.950 129.600 496.050 130.050 ;
        RECT 559.950 129.600 562.050 130.050 ;
        RECT 580.950 129.600 583.050 130.050 ;
        RECT 493.950 128.400 583.050 129.600 ;
        RECT 493.950 127.950 496.050 128.400 ;
        RECT 559.950 127.950 562.050 128.400 ;
        RECT 580.950 127.950 583.050 128.400 ;
        RECT 601.950 129.600 604.050 130.050 ;
        RECT 610.950 129.600 613.050 130.050 ;
        RECT 718.950 129.600 721.050 130.050 ;
        RECT 601.950 128.400 613.050 129.600 ;
        RECT 601.950 127.950 604.050 128.400 ;
        RECT 610.950 127.950 613.050 128.400 ;
        RECT 704.400 128.400 721.050 129.600 ;
        RECT 19.950 126.600 22.050 127.050 ;
        RECT 34.950 126.600 37.050 127.050 ;
        RECT 46.950 126.600 49.050 127.050 ;
        RECT 19.950 125.400 49.050 126.600 ;
        RECT 19.950 124.950 22.050 125.400 ;
        RECT 34.950 124.950 37.050 125.400 ;
        RECT 46.950 124.950 49.050 125.400 ;
        RECT 97.950 126.600 100.050 127.050 ;
        RECT 172.950 126.600 175.050 127.050 ;
        RECT 97.950 125.400 175.050 126.600 ;
        RECT 97.950 124.950 100.050 125.400 ;
        RECT 172.950 124.950 175.050 125.400 ;
        RECT 187.950 126.600 190.050 127.050 ;
        RECT 238.950 126.600 241.050 127.050 ;
        RECT 187.950 125.400 241.050 126.600 ;
        RECT 187.950 124.950 190.050 125.400 ;
        RECT 238.950 124.950 241.050 125.400 ;
        RECT 307.950 126.600 310.050 127.050 ;
        RECT 340.950 126.600 343.050 127.050 ;
        RECT 307.950 125.400 343.050 126.600 ;
        RECT 307.950 124.950 310.050 125.400 ;
        RECT 340.950 124.950 343.050 125.400 ;
        RECT 361.950 126.600 364.050 127.050 ;
        RECT 376.950 126.600 379.050 127.050 ;
        RECT 361.950 125.400 379.050 126.600 ;
        RECT 361.950 124.950 364.050 125.400 ;
        RECT 376.950 124.950 379.050 125.400 ;
        RECT 421.950 126.600 424.050 127.050 ;
        RECT 451.950 126.600 454.050 127.050 ;
        RECT 421.950 125.400 454.050 126.600 ;
        RECT 421.950 124.950 424.050 125.400 ;
        RECT 451.950 124.950 454.050 125.400 ;
        RECT 475.950 126.600 478.050 127.050 ;
        RECT 571.950 126.600 574.050 127.050 ;
        RECT 475.950 125.400 574.050 126.600 ;
        RECT 475.950 124.950 478.050 125.400 ;
        RECT 571.950 124.950 574.050 125.400 ;
        RECT 595.950 126.600 598.050 127.050 ;
        RECT 613.950 126.600 616.050 127.050 ;
        RECT 595.950 125.400 616.050 126.600 ;
        RECT 595.950 124.950 598.050 125.400 ;
        RECT 613.950 124.950 616.050 125.400 ;
        RECT 682.950 126.600 685.050 127.050 ;
        RECT 704.400 126.600 705.600 128.400 ;
        RECT 718.950 127.950 721.050 128.400 ;
        RECT 748.950 129.600 751.050 130.050 ;
        RECT 790.950 129.600 793.050 130.050 ;
        RECT 748.950 128.400 793.050 129.600 ;
        RECT 748.950 127.950 751.050 128.400 ;
        RECT 790.950 127.950 793.050 128.400 ;
        RECT 796.950 129.600 799.050 130.050 ;
        RECT 817.950 129.600 820.050 130.050 ;
        RECT 796.950 128.400 820.050 129.600 ;
        RECT 796.950 127.950 799.050 128.400 ;
        RECT 817.950 127.950 820.050 128.400 ;
        RECT 708.000 126.600 712.050 127.050 ;
        RECT 682.950 125.400 705.600 126.600 ;
        RECT 682.950 124.950 685.050 125.400 ;
        RECT 707.400 124.950 712.050 126.600 ;
        RECT 721.950 126.600 724.050 127.050 ;
        RECT 730.950 126.600 733.050 127.050 ;
        RECT 721.950 125.400 733.050 126.600 ;
        RECT 721.950 124.950 724.050 125.400 ;
        RECT 730.950 124.950 733.050 125.400 ;
        RECT 757.950 126.600 760.050 127.050 ;
        RECT 769.950 126.600 772.050 127.050 ;
        RECT 757.950 125.400 772.050 126.600 ;
        RECT 757.950 124.950 760.050 125.400 ;
        RECT 769.950 124.950 772.050 125.400 ;
        RECT 778.950 126.600 781.050 127.050 ;
        RECT 802.950 126.600 805.050 127.050 ;
        RECT 778.950 125.400 805.050 126.600 ;
        RECT 778.950 124.950 781.050 125.400 ;
        RECT 802.950 124.950 805.050 125.400 ;
        RECT 826.950 126.600 829.050 127.050 ;
        RECT 838.950 126.600 841.050 127.050 ;
        RECT 826.950 125.400 841.050 126.600 ;
        RECT 826.950 124.950 829.050 125.400 ;
        RECT 838.950 124.950 841.050 125.400 ;
        RECT 223.950 123.600 226.050 124.050 ;
        RECT 232.950 123.600 235.050 124.050 ;
        RECT 253.950 123.600 256.050 124.050 ;
        RECT 223.950 122.400 256.050 123.600 ;
        RECT 223.950 121.950 226.050 122.400 ;
        RECT 232.950 121.950 235.050 122.400 ;
        RECT 253.950 121.950 256.050 122.400 ;
        RECT 418.950 123.600 421.050 124.050 ;
        RECT 523.950 123.600 526.050 124.050 ;
        RECT 418.950 122.400 526.050 123.600 ;
        RECT 418.950 121.950 421.050 122.400 ;
        RECT 523.950 121.950 526.050 122.400 ;
        RECT 529.950 123.600 532.050 124.050 ;
        RECT 541.950 123.600 544.050 124.050 ;
        RECT 529.950 122.400 544.050 123.600 ;
        RECT 529.950 121.950 532.050 122.400 ;
        RECT 541.950 121.950 544.050 122.400 ;
        RECT 676.950 123.600 679.050 124.050 ;
        RECT 707.400 123.600 708.600 124.950 ;
        RECT 676.950 122.400 708.600 123.600 ;
        RECT 844.950 123.600 847.050 124.050 ;
        RECT 865.950 123.600 868.050 124.050 ;
        RECT 844.950 122.400 868.050 123.600 ;
        RECT 676.950 121.950 679.050 122.400 ;
        RECT 844.950 121.950 847.050 122.400 ;
        RECT 865.950 121.950 868.050 122.400 ;
        RECT 121.950 120.600 124.050 121.050 ;
        RECT 139.950 120.600 142.050 121.050 ;
        RECT 121.950 119.400 142.050 120.600 ;
        RECT 121.950 118.950 124.050 119.400 ;
        RECT 139.950 118.950 142.050 119.400 ;
        RECT 196.950 120.600 199.050 121.050 ;
        RECT 268.950 120.600 271.050 121.050 ;
        RECT 196.950 119.400 271.050 120.600 ;
        RECT 196.950 118.950 199.050 119.400 ;
        RECT 268.950 118.950 271.050 119.400 ;
        RECT 334.950 120.600 337.050 121.050 ;
        RECT 403.950 120.600 406.050 121.050 ;
        RECT 334.950 119.400 406.050 120.600 ;
        RECT 334.950 118.950 337.050 119.400 ;
        RECT 403.950 118.950 406.050 119.400 ;
        RECT 463.950 120.600 466.050 121.050 ;
        RECT 487.950 120.600 490.050 121.050 ;
        RECT 463.950 119.400 490.050 120.600 ;
        RECT 463.950 118.950 466.050 119.400 ;
        RECT 487.950 118.950 490.050 119.400 ;
        RECT 583.950 120.600 586.050 121.050 ;
        RECT 598.950 120.600 601.050 121.050 ;
        RECT 583.950 119.400 601.050 120.600 ;
        RECT 583.950 118.950 586.050 119.400 ;
        RECT 598.950 118.950 601.050 119.400 ;
        RECT 709.950 120.600 712.050 121.050 ;
        RECT 778.950 120.600 781.050 121.050 ;
        RECT 709.950 119.400 781.050 120.600 ;
        RECT 709.950 118.950 712.050 119.400 ;
        RECT 778.950 118.950 781.050 119.400 ;
        RECT 808.950 120.600 811.050 121.050 ;
        RECT 838.950 120.600 841.050 121.050 ;
        RECT 808.950 119.400 841.050 120.600 ;
        RECT 808.950 118.950 811.050 119.400 ;
        RECT 838.950 118.950 841.050 119.400 ;
        RECT 67.950 117.600 70.050 118.050 ;
        RECT 79.950 117.600 82.050 118.050 ;
        RECT 67.950 116.400 82.050 117.600 ;
        RECT 67.950 115.950 70.050 116.400 ;
        RECT 79.950 115.950 82.050 116.400 ;
        RECT 322.950 117.600 325.050 118.050 ;
        RECT 337.950 117.600 340.050 118.050 ;
        RECT 322.950 116.400 340.050 117.600 ;
        RECT 322.950 115.950 325.050 116.400 ;
        RECT 337.950 115.950 340.050 116.400 ;
        RECT 346.950 117.600 349.050 118.050 ;
        RECT 400.950 117.600 403.050 118.050 ;
        RECT 346.950 116.400 403.050 117.600 ;
        RECT 346.950 115.950 349.050 116.400 ;
        RECT 400.950 115.950 403.050 116.400 ;
        RECT 430.950 117.600 433.050 118.050 ;
        RECT 496.950 117.600 499.050 118.050 ;
        RECT 502.950 117.600 505.050 118.050 ;
        RECT 430.950 116.400 505.050 117.600 ;
        RECT 430.950 115.950 433.050 116.400 ;
        RECT 496.950 115.950 499.050 116.400 ;
        RECT 502.950 115.950 505.050 116.400 ;
        RECT 646.950 117.600 649.050 118.050 ;
        RECT 706.950 117.600 709.050 118.050 ;
        RECT 646.950 116.400 709.050 117.600 ;
        RECT 646.950 115.950 649.050 116.400 ;
        RECT 706.950 115.950 709.050 116.400 ;
        RECT 724.950 117.600 727.050 118.050 ;
        RECT 751.950 117.600 754.050 118.050 ;
        RECT 724.950 116.400 754.050 117.600 ;
        RECT 724.950 115.950 727.050 116.400 ;
        RECT 751.950 115.950 754.050 116.400 ;
        RECT 49.950 114.600 52.050 115.050 ;
        RECT 103.950 114.600 106.050 115.050 ;
        RECT 106.950 114.600 109.050 115.050 ;
        RECT 133.950 114.600 136.050 115.050 ;
        RECT 49.950 113.400 136.050 114.600 ;
        RECT 49.950 112.950 52.050 113.400 ;
        RECT 103.950 112.950 106.050 113.400 ;
        RECT 106.950 112.950 109.050 113.400 ;
        RECT 133.950 112.950 136.050 113.400 ;
        RECT 163.950 114.600 166.050 115.050 ;
        RECT 175.950 114.600 178.050 115.050 ;
        RECT 163.950 113.400 178.050 114.600 ;
        RECT 163.950 112.950 166.050 113.400 ;
        RECT 175.950 112.950 178.050 113.400 ;
        RECT 199.950 114.600 202.050 115.050 ;
        RECT 235.950 114.600 238.050 115.050 ;
        RECT 199.950 113.400 238.050 114.600 ;
        RECT 199.950 112.950 202.050 113.400 ;
        RECT 235.950 112.950 238.050 113.400 ;
        RECT 289.950 114.600 292.050 115.050 ;
        RECT 406.950 114.600 409.050 115.050 ;
        RECT 289.950 113.400 409.050 114.600 ;
        RECT 289.950 112.950 292.050 113.400 ;
        RECT 406.950 112.950 409.050 113.400 ;
        RECT 442.950 114.600 445.050 115.050 ;
        RECT 472.950 114.600 475.050 115.050 ;
        RECT 442.950 113.400 475.050 114.600 ;
        RECT 442.950 112.950 445.050 113.400 ;
        RECT 472.950 112.950 475.050 113.400 ;
        RECT 487.950 114.600 490.050 115.050 ;
        RECT 529.950 114.600 532.050 115.050 ;
        RECT 553.950 114.600 556.050 115.050 ;
        RECT 487.950 113.400 556.050 114.600 ;
        RECT 487.950 112.950 490.050 113.400 ;
        RECT 529.950 112.950 532.050 113.400 ;
        RECT 553.950 112.950 556.050 113.400 ;
        RECT 667.950 114.600 670.050 115.050 ;
        RECT 700.950 114.600 703.050 115.050 ;
        RECT 667.950 113.400 703.050 114.600 ;
        RECT 667.950 112.950 670.050 113.400 ;
        RECT 700.950 112.950 703.050 113.400 ;
        RECT 829.950 114.600 832.050 115.050 ;
        RECT 844.950 114.600 847.050 115.050 ;
        RECT 829.950 113.400 847.050 114.600 ;
        RECT 829.950 112.950 832.050 113.400 ;
        RECT 844.950 112.950 847.050 113.400 ;
        RECT 853.950 114.600 856.050 115.050 ;
        RECT 865.950 114.600 868.050 115.050 ;
        RECT 853.950 113.400 868.050 114.600 ;
        RECT 853.950 112.950 856.050 113.400 ;
        RECT 865.950 112.950 868.050 113.400 ;
        RECT 73.950 111.600 76.050 112.050 ;
        RECT 130.950 111.600 133.050 112.050 ;
        RECT 73.950 110.400 133.050 111.600 ;
        RECT 73.950 109.950 76.050 110.400 ;
        RECT 130.950 109.950 133.050 110.400 ;
        RECT 142.950 111.600 145.050 112.050 ;
        RECT 148.950 111.600 151.050 112.050 ;
        RECT 142.950 110.400 151.050 111.600 ;
        RECT 142.950 109.950 145.050 110.400 ;
        RECT 148.950 109.950 151.050 110.400 ;
        RECT 295.950 111.600 298.050 112.050 ;
        RECT 304.950 111.600 307.050 112.050 ;
        RECT 295.950 110.400 307.050 111.600 ;
        RECT 295.950 109.950 298.050 110.400 ;
        RECT 304.950 109.950 307.050 110.400 ;
        RECT 328.950 111.600 331.050 112.050 ;
        RECT 382.950 111.600 385.050 112.050 ;
        RECT 328.950 110.400 385.050 111.600 ;
        RECT 328.950 109.950 331.050 110.400 ;
        RECT 382.950 109.950 385.050 110.400 ;
        RECT 424.950 111.600 427.050 112.050 ;
        RECT 439.950 111.600 442.050 112.050 ;
        RECT 484.950 111.600 487.050 112.050 ;
        RECT 424.950 110.400 487.050 111.600 ;
        RECT 424.950 109.950 427.050 110.400 ;
        RECT 439.950 109.950 442.050 110.400 ;
        RECT 484.950 109.950 487.050 110.400 ;
        RECT 655.950 111.600 658.050 112.050 ;
        RECT 712.950 111.600 715.050 112.050 ;
        RECT 655.950 110.400 715.050 111.600 ;
        RECT 655.950 109.950 658.050 110.400 ;
        RECT 712.950 109.950 715.050 110.400 ;
        RECT 754.950 111.600 757.050 112.050 ;
        RECT 784.950 111.600 787.050 112.050 ;
        RECT 754.950 110.400 787.050 111.600 ;
        RECT 754.950 109.950 757.050 110.400 ;
        RECT 784.950 109.950 787.050 110.400 ;
        RECT 802.950 111.600 805.050 112.050 ;
        RECT 826.950 111.600 829.050 112.050 ;
        RECT 802.950 110.400 829.050 111.600 ;
        RECT 802.950 109.950 805.050 110.400 ;
        RECT 826.950 109.950 829.050 110.400 ;
        RECT 832.950 111.600 835.050 112.050 ;
        RECT 841.950 111.600 844.050 112.050 ;
        RECT 832.950 110.400 844.050 111.600 ;
        RECT 832.950 109.950 835.050 110.400 ;
        RECT 841.950 109.950 844.050 110.400 ;
        RECT 22.950 108.600 25.050 109.050 ;
        RECT 43.950 108.600 46.050 109.050 ;
        RECT 55.950 108.600 58.050 109.050 ;
        RECT 22.950 107.400 58.050 108.600 ;
        RECT 22.950 106.950 25.050 107.400 ;
        RECT 43.950 106.950 46.050 107.400 ;
        RECT 55.950 106.950 58.050 107.400 ;
        RECT 136.950 108.600 139.050 109.050 ;
        RECT 142.950 108.600 145.050 108.900 ;
        RECT 136.950 107.400 145.050 108.600 ;
        RECT 136.950 106.950 139.050 107.400 ;
        RECT 142.950 106.800 145.050 107.400 ;
        RECT 346.950 108.600 349.050 109.050 ;
        RECT 352.950 108.600 355.050 109.050 ;
        RECT 346.950 107.400 355.050 108.600 ;
        RECT 346.950 106.950 349.050 107.400 ;
        RECT 352.950 106.950 355.050 107.400 ;
        RECT 367.950 108.600 370.050 109.050 ;
        RECT 391.950 108.600 394.050 109.050 ;
        RECT 511.950 108.600 514.050 109.050 ;
        RECT 520.950 108.600 523.050 109.050 ;
        RECT 367.950 107.400 390.600 108.600 ;
        RECT 367.950 106.950 370.050 107.400 ;
        RECT 10.950 105.600 13.050 106.050 ;
        RECT 16.950 105.600 19.050 106.200 ;
        RECT 10.950 104.400 19.050 105.600 ;
        RECT 10.950 103.950 13.050 104.400 ;
        RECT 16.950 104.100 19.050 104.400 ;
        RECT 58.950 105.750 61.050 105.900 ;
        RECT 67.950 105.750 70.050 106.200 ;
        RECT 58.950 105.600 70.050 105.750 ;
        RECT 88.950 105.600 91.050 106.200 ;
        RECT 58.950 104.550 91.050 105.600 ;
        RECT 58.950 103.800 61.050 104.550 ;
        RECT 67.950 104.400 91.050 104.550 ;
        RECT 67.950 104.100 70.050 104.400 ;
        RECT 88.950 104.100 91.050 104.400 ;
        RECT 112.950 105.600 115.050 106.200 ;
        RECT 112.950 104.400 132.600 105.600 ;
        RECT 112.950 104.100 115.050 104.400 ;
        RECT 131.400 99.900 132.600 104.400 ;
        RECT 133.950 104.100 136.050 106.200 ;
        RECT 184.950 105.600 187.050 106.200 ;
        RECT 208.950 105.600 211.050 106.200 ;
        RECT 184.950 104.400 211.050 105.600 ;
        RECT 184.950 104.100 187.050 104.400 ;
        RECT 208.950 104.100 211.050 104.400 ;
        RECT 223.950 105.750 226.050 106.200 ;
        RECT 229.950 105.750 232.050 106.200 ;
        RECT 223.950 104.550 232.050 105.750 ;
        RECT 223.950 104.100 226.050 104.550 ;
        RECT 229.950 104.100 232.050 104.550 ;
        RECT 247.950 105.750 250.050 106.200 ;
        RECT 259.950 105.750 262.050 106.200 ;
        RECT 247.950 104.550 262.050 105.750 ;
        RECT 247.950 104.100 250.050 104.550 ;
        RECT 259.950 104.100 262.050 104.550 ;
        RECT 268.950 105.600 271.050 106.050 ;
        RECT 280.950 105.600 283.050 106.200 ;
        RECT 298.950 105.600 301.050 106.200 ;
        RECT 268.950 104.400 301.050 105.600 ;
        RECT 134.400 102.600 135.600 104.100 ;
        RECT 268.950 103.950 271.050 104.400 ;
        RECT 280.950 104.100 283.050 104.400 ;
        RECT 298.950 104.100 301.050 104.400 ;
        RECT 370.950 105.600 373.050 106.050 ;
        RECT 376.950 105.600 379.050 106.050 ;
        RECT 370.950 104.400 379.050 105.600 ;
        RECT 389.400 105.600 390.600 107.400 ;
        RECT 391.950 107.400 432.600 108.600 ;
        RECT 391.950 106.950 394.050 107.400 ;
        RECT 412.950 105.750 415.050 106.200 ;
        RECT 421.950 105.750 424.050 106.200 ;
        RECT 389.400 104.400 405.600 105.600 ;
        RECT 370.950 103.950 373.050 104.400 ;
        RECT 376.950 103.950 379.050 104.400 ;
        RECT 334.950 102.600 337.050 103.050 ;
        RECT 134.400 101.400 141.600 102.600 ;
        RECT 25.950 99.600 28.050 99.900 ;
        RECT 40.950 99.600 43.050 99.900 ;
        RECT 25.950 98.400 43.050 99.600 ;
        RECT 25.950 97.800 28.050 98.400 ;
        RECT 40.950 97.800 43.050 98.400 ;
        RECT 91.950 99.600 94.050 99.900 ;
        RECT 109.950 99.600 112.050 99.900 ;
        RECT 91.950 98.400 112.050 99.600 ;
        RECT 91.950 97.800 94.050 98.400 ;
        RECT 109.950 97.800 112.050 98.400 ;
        RECT 115.950 99.450 118.050 99.900 ;
        RECT 121.950 99.450 124.050 99.900 ;
        RECT 115.950 98.250 124.050 99.450 ;
        RECT 115.950 97.800 118.050 98.250 ;
        RECT 121.950 97.800 124.050 98.250 ;
        RECT 130.950 97.800 133.050 99.900 ;
        RECT 70.950 96.600 73.050 97.050 ;
        RECT 79.950 96.600 82.050 97.050 ;
        RECT 70.950 95.400 82.050 96.600 ;
        RECT 140.400 96.600 141.600 101.400 ;
        RECT 314.400 101.400 337.050 102.600 ;
        RECT 145.950 99.450 148.050 99.900 ;
        RECT 166.950 99.450 169.050 99.900 ;
        RECT 145.950 98.250 169.050 99.450 ;
        RECT 145.950 97.800 148.050 98.250 ;
        RECT 166.950 97.800 169.050 98.250 ;
        RECT 190.950 99.450 193.050 99.900 ;
        RECT 199.950 99.450 202.050 99.900 ;
        RECT 190.950 98.250 202.050 99.450 ;
        RECT 190.950 97.800 193.050 98.250 ;
        RECT 199.950 97.800 202.050 98.250 ;
        RECT 214.950 99.600 217.050 100.050 ;
        RECT 223.950 99.600 226.050 100.050 ;
        RECT 314.400 99.900 315.600 101.400 ;
        RECT 334.950 100.950 337.050 101.400 ;
        RECT 404.400 100.050 405.600 104.400 ;
        RECT 412.950 104.550 424.050 105.750 ;
        RECT 412.950 104.100 415.050 104.550 ;
        RECT 421.950 104.100 424.050 104.550 ;
        RECT 431.400 105.600 432.600 107.400 ;
        RECT 511.950 107.400 523.050 108.600 ;
        RECT 511.950 106.950 514.050 107.400 ;
        RECT 520.950 106.950 523.050 107.400 ;
        RECT 634.950 108.600 637.050 109.050 ;
        RECT 640.950 108.600 643.050 109.050 ;
        RECT 649.950 108.600 652.050 109.050 ;
        RECT 634.950 107.400 643.050 108.600 ;
        RECT 634.950 106.950 637.050 107.400 ;
        RECT 640.950 106.950 643.050 107.400 ;
        RECT 644.400 107.400 652.050 108.600 ;
        RECT 433.950 105.600 436.050 106.200 ;
        RECT 445.950 105.600 448.050 106.050 ;
        RECT 457.950 105.600 460.050 106.200 ;
        RECT 431.400 104.400 460.050 105.600 ;
        RECT 433.950 104.100 436.050 104.400 ;
        RECT 445.950 103.950 448.050 104.400 ;
        RECT 457.950 104.100 460.050 104.400 ;
        RECT 469.950 105.600 472.050 106.050 ;
        RECT 478.950 105.600 481.050 106.200 ;
        RECT 469.950 104.400 481.050 105.600 ;
        RECT 469.950 103.950 472.050 104.400 ;
        RECT 478.950 104.100 481.050 104.400 ;
        RECT 484.950 105.600 487.050 106.200 ;
        RECT 505.950 105.600 508.050 106.200 ;
        RECT 484.950 104.400 508.050 105.600 ;
        RECT 484.950 104.100 487.050 104.400 ;
        RECT 505.950 104.100 508.050 104.400 ;
        RECT 523.950 105.600 528.000 106.050 ;
        RECT 535.950 105.600 538.050 106.200 ;
        RECT 544.950 105.600 547.050 106.050 ;
        RECT 523.950 103.950 528.600 105.600 ;
        RECT 535.950 104.400 547.050 105.600 ;
        RECT 535.950 104.100 538.050 104.400 ;
        RECT 544.950 103.950 547.050 104.400 ;
        RECT 559.950 105.600 562.050 106.200 ;
        RECT 574.950 105.600 577.050 106.200 ;
        RECT 559.950 104.400 577.050 105.600 ;
        RECT 559.950 104.100 562.050 104.400 ;
        RECT 574.950 104.100 577.050 104.400 ;
        RECT 589.950 105.750 592.050 106.200 ;
        RECT 604.950 105.750 607.050 106.200 ;
        RECT 589.950 104.550 607.050 105.750 ;
        RECT 589.950 104.100 592.050 104.550 ;
        RECT 604.950 104.100 607.050 104.550 ;
        RECT 610.950 105.600 613.050 106.050 ;
        RECT 625.950 105.600 628.050 106.050 ;
        RECT 644.400 105.600 645.600 107.400 ;
        RECT 649.950 106.950 652.050 107.400 ;
        RECT 787.950 108.600 790.050 109.050 ;
        RECT 787.950 107.400 831.600 108.600 ;
        RECT 787.950 106.950 790.050 107.400 ;
        RECT 610.950 104.400 645.600 105.600 ;
        RECT 673.950 105.600 676.050 106.050 ;
        RECT 688.950 105.600 691.050 106.200 ;
        RECT 673.950 104.400 691.050 105.600 ;
        RECT 610.950 103.950 613.050 104.400 ;
        RECT 625.950 103.950 628.050 104.400 ;
        RECT 673.950 103.950 676.050 104.400 ;
        RECT 688.950 104.100 691.050 104.400 ;
        RECT 694.950 105.750 697.050 106.200 ;
        RECT 700.950 105.750 703.050 106.200 ;
        RECT 694.950 104.550 703.050 105.750 ;
        RECT 694.950 104.100 697.050 104.550 ;
        RECT 700.950 104.100 703.050 104.550 ;
        RECT 715.950 105.600 718.050 106.200 ;
        RECT 736.950 105.600 739.050 106.200 ;
        RECT 715.950 104.400 739.050 105.600 ;
        RECT 715.950 104.100 718.050 104.400 ;
        RECT 736.950 104.100 739.050 104.400 ;
        RECT 748.950 105.750 751.050 106.200 ;
        RECT 760.950 105.750 763.050 106.200 ;
        RECT 748.950 105.600 763.050 105.750 ;
        RECT 784.950 105.600 787.050 106.200 ;
        RECT 748.950 104.550 787.050 105.600 ;
        RECT 748.950 104.100 751.050 104.550 ;
        RECT 760.950 104.400 787.050 104.550 ;
        RECT 760.950 104.100 763.050 104.400 ;
        RECT 784.950 104.100 787.050 104.400 ;
        RECT 796.950 105.600 799.050 106.050 ;
        RECT 802.950 105.600 805.050 106.200 ;
        RECT 830.400 105.600 831.600 107.400 ;
        RECT 796.950 104.400 805.050 105.600 ;
        RECT 796.950 103.950 799.050 104.400 ;
        RECT 802.950 104.100 805.050 104.400 ;
        RECT 815.400 104.400 831.600 105.600 ;
        RECT 527.400 102.600 528.600 103.950 ;
        RECT 527.400 101.400 558.600 102.600 ;
        RECT 214.950 98.400 226.050 99.600 ;
        RECT 214.950 97.950 217.050 98.400 ;
        RECT 223.950 97.950 226.050 98.400 ;
        RECT 241.950 99.450 244.050 99.900 ;
        RECT 256.950 99.450 259.050 99.900 ;
        RECT 241.950 98.250 259.050 99.450 ;
        RECT 241.950 97.800 244.050 98.250 ;
        RECT 256.950 97.800 259.050 98.250 ;
        RECT 262.950 99.600 265.050 99.900 ;
        RECT 283.950 99.600 286.050 99.900 ;
        RECT 262.950 99.450 286.050 99.600 ;
        RECT 289.950 99.450 292.050 99.900 ;
        RECT 262.950 98.400 292.050 99.450 ;
        RECT 262.950 97.800 265.050 98.400 ;
        RECT 283.950 98.250 292.050 98.400 ;
        RECT 283.950 97.800 286.050 98.250 ;
        RECT 289.950 97.800 292.050 98.250 ;
        RECT 313.950 97.800 316.050 99.900 ;
        RECT 358.950 99.600 361.050 100.050 ;
        RECT 364.950 99.600 367.050 99.900 ;
        RECT 358.950 98.400 367.050 99.600 ;
        RECT 358.950 97.950 361.050 98.400 ;
        RECT 364.950 97.800 367.050 98.400 ;
        RECT 403.950 97.950 406.050 100.050 ;
        RECT 527.400 99.900 528.600 101.400 ;
        RECT 557.400 99.900 558.600 101.400 ;
        RECT 815.400 100.050 816.600 104.400 ;
        RECT 415.950 99.450 418.050 99.900 ;
        RECT 424.950 99.450 427.050 99.900 ;
        RECT 415.950 98.250 427.050 99.450 ;
        RECT 415.950 97.800 418.050 98.250 ;
        RECT 424.950 97.800 427.050 98.250 ;
        RECT 496.950 99.450 499.050 99.900 ;
        RECT 508.950 99.450 511.050 99.900 ;
        RECT 496.950 98.250 511.050 99.450 ;
        RECT 496.950 97.800 499.050 98.250 ;
        RECT 508.950 97.800 511.050 98.250 ;
        RECT 526.950 97.800 529.050 99.900 ;
        RECT 532.950 99.600 535.050 99.900 ;
        RECT 550.950 99.600 553.050 99.900 ;
        RECT 532.950 98.400 553.050 99.600 ;
        RECT 532.950 97.800 535.050 98.400 ;
        RECT 550.950 97.800 553.050 98.400 ;
        RECT 556.950 97.800 559.050 99.900 ;
        RECT 583.950 99.450 586.050 99.900 ;
        RECT 634.950 99.450 637.050 99.900 ;
        RECT 583.950 98.250 637.050 99.450 ;
        RECT 583.950 97.800 586.050 98.250 ;
        RECT 634.950 97.800 637.050 98.250 ;
        RECT 706.950 99.600 709.050 100.050 ;
        RECT 718.950 99.600 721.050 99.900 ;
        RECT 706.950 98.400 721.050 99.600 ;
        RECT 706.950 97.950 709.050 98.400 ;
        RECT 718.950 97.800 721.050 98.400 ;
        RECT 814.950 97.950 817.050 100.050 ;
        RECT 830.400 99.900 831.600 104.400 ;
        RECT 832.950 105.600 835.050 106.200 ;
        RECT 838.950 105.600 841.050 106.050 ;
        RECT 874.950 105.600 877.050 106.200 ;
        RECT 832.950 104.400 877.050 105.600 ;
        RECT 832.950 104.100 835.050 104.400 ;
        RECT 838.950 103.950 841.050 104.400 ;
        RECT 874.950 104.100 877.050 104.400 ;
        RECT 829.950 97.800 832.050 99.900 ;
        RECT 844.950 99.450 847.050 99.900 ;
        RECT 850.950 99.450 853.050 99.900 ;
        RECT 844.950 98.250 853.050 99.450 ;
        RECT 844.950 97.800 847.050 98.250 ;
        RECT 850.950 97.800 853.050 98.250 ;
        RECT 865.950 99.450 868.050 99.900 ;
        RECT 871.950 99.450 874.050 99.900 ;
        RECT 865.950 98.250 874.050 99.450 ;
        RECT 865.950 97.800 868.050 98.250 ;
        RECT 871.950 97.800 874.050 98.250 ;
        RECT 175.950 96.600 178.050 97.050 ;
        RECT 319.950 96.600 322.050 97.050 ;
        RECT 140.400 95.400 144.600 96.600 ;
        RECT 70.950 94.950 73.050 95.400 ;
        RECT 79.950 94.950 82.050 95.400 ;
        RECT 10.950 93.600 13.050 94.050 ;
        RECT 58.950 93.600 61.050 94.050 ;
        RECT 10.950 92.400 61.050 93.600 ;
        RECT 143.400 93.600 144.600 95.400 ;
        RECT 175.950 95.400 322.050 96.600 ;
        RECT 175.950 94.950 178.050 95.400 ;
        RECT 319.950 94.950 322.050 95.400 ;
        RECT 205.950 93.600 208.050 94.050 ;
        RECT 232.950 93.600 235.050 94.050 ;
        RECT 143.400 92.400 235.050 93.600 ;
        RECT 10.950 91.950 13.050 92.400 ;
        RECT 58.950 91.950 61.050 92.400 ;
        RECT 205.950 91.950 208.050 92.400 ;
        RECT 232.950 91.950 235.050 92.400 ;
        RECT 238.950 93.600 241.050 94.050 ;
        RECT 247.950 93.600 250.050 94.050 ;
        RECT 277.950 93.600 280.050 94.050 ;
        RECT 238.950 92.400 280.050 93.600 ;
        RECT 238.950 91.950 241.050 92.400 ;
        RECT 247.950 91.950 250.050 92.400 ;
        RECT 277.950 91.950 280.050 92.400 ;
        RECT 295.950 93.600 298.050 94.050 ;
        RECT 328.950 93.600 331.050 97.050 ;
        RECT 400.950 96.600 403.050 97.050 ;
        RECT 412.950 96.600 415.050 97.050 ;
        RECT 430.950 96.600 433.050 97.050 ;
        RECT 454.950 96.600 457.050 97.050 ;
        RECT 400.950 95.400 457.050 96.600 ;
        RECT 400.950 94.950 403.050 95.400 ;
        RECT 412.950 94.950 415.050 95.400 ;
        RECT 430.950 94.950 433.050 95.400 ;
        RECT 454.950 94.950 457.050 95.400 ;
        RECT 484.950 96.600 487.050 97.050 ;
        RECT 502.950 96.600 505.050 97.050 ;
        RECT 484.950 95.400 505.050 96.600 ;
        RECT 484.950 94.950 487.050 95.400 ;
        RECT 502.950 94.950 505.050 95.400 ;
        RECT 529.950 96.600 532.050 97.050 ;
        RECT 553.950 96.600 556.050 97.050 ;
        RECT 529.950 95.400 556.050 96.600 ;
        RECT 529.950 94.950 532.050 95.400 ;
        RECT 553.950 94.950 556.050 95.400 ;
        RECT 559.950 96.600 562.050 97.050 ;
        RECT 577.950 96.600 580.050 97.050 ;
        RECT 559.950 95.400 580.050 96.600 ;
        RECT 559.950 94.950 562.050 95.400 ;
        RECT 577.950 94.950 580.050 95.400 ;
        RECT 649.950 96.600 652.050 97.050 ;
        RECT 655.950 96.600 658.050 97.050 ;
        RECT 649.950 95.400 658.050 96.600 ;
        RECT 649.950 94.950 652.050 95.400 ;
        RECT 655.950 94.950 658.050 95.400 ;
        RECT 700.950 96.600 703.050 97.050 ;
        RECT 739.950 96.600 742.050 97.050 ;
        RECT 763.950 96.600 766.050 97.050 ;
        RECT 781.950 96.600 784.050 97.050 ;
        RECT 700.950 95.400 784.050 96.600 ;
        RECT 700.950 94.950 703.050 95.400 ;
        RECT 739.950 94.950 742.050 95.400 ;
        RECT 763.950 94.950 766.050 95.400 ;
        RECT 781.950 94.950 784.050 95.400 ;
        RECT 295.950 93.000 331.050 93.600 ;
        RECT 337.950 93.600 340.050 94.050 ;
        RECT 385.950 93.600 388.050 94.050 ;
        RECT 295.950 92.400 330.600 93.000 ;
        RECT 337.950 92.400 388.050 93.600 ;
        RECT 295.950 91.950 298.050 92.400 ;
        RECT 337.950 91.950 340.050 92.400 ;
        RECT 385.950 91.950 388.050 92.400 ;
        RECT 469.950 93.600 472.050 94.050 ;
        RECT 589.950 93.600 592.050 94.050 ;
        RECT 469.950 92.400 592.050 93.600 ;
        RECT 469.950 91.950 472.050 92.400 ;
        RECT 589.950 91.950 592.050 92.400 ;
        RECT 607.950 93.600 610.050 94.050 ;
        RECT 673.950 93.600 676.050 94.050 ;
        RECT 607.950 92.400 676.050 93.600 ;
        RECT 607.950 91.950 610.050 92.400 ;
        RECT 673.950 91.950 676.050 92.400 ;
        RECT 436.950 90.600 439.050 91.050 ;
        RECT 466.950 90.600 469.050 91.050 ;
        RECT 436.950 89.400 469.050 90.600 ;
        RECT 436.950 88.950 439.050 89.400 ;
        RECT 466.950 88.950 469.050 89.400 ;
        RECT 544.950 90.600 547.050 91.050 ;
        RECT 601.950 90.600 604.050 91.050 ;
        RECT 544.950 89.400 604.050 90.600 ;
        RECT 544.950 88.950 547.050 89.400 ;
        RECT 601.950 88.950 604.050 89.400 ;
        RECT 685.950 90.600 688.050 91.050 ;
        RECT 703.950 90.600 706.050 91.050 ;
        RECT 712.950 90.600 715.050 91.050 ;
        RECT 685.950 89.400 715.050 90.600 ;
        RECT 685.950 88.950 688.050 89.400 ;
        RECT 703.950 88.950 706.050 89.400 ;
        RECT 712.950 88.950 715.050 89.400 ;
        RECT 757.950 90.600 760.050 91.050 ;
        RECT 787.950 90.600 790.050 91.050 ;
        RECT 757.950 89.400 790.050 90.600 ;
        RECT 757.950 88.950 760.050 89.400 ;
        RECT 787.950 88.950 790.050 89.400 ;
        RECT 49.950 87.600 52.050 88.050 ;
        RECT 55.950 87.600 58.050 88.050 ;
        RECT 49.950 86.400 58.050 87.600 ;
        RECT 49.950 85.950 52.050 86.400 ;
        RECT 55.950 85.950 58.050 86.400 ;
        RECT 715.950 87.600 718.050 88.050 ;
        RECT 748.950 87.600 751.050 88.050 ;
        RECT 715.950 86.400 751.050 87.600 ;
        RECT 715.950 85.950 718.050 86.400 ;
        RECT 748.950 85.950 751.050 86.400 ;
        RECT 340.950 84.600 343.050 85.050 ;
        RECT 352.950 84.600 355.050 85.050 ;
        RECT 340.950 83.400 355.050 84.600 ;
        RECT 340.950 82.950 343.050 83.400 ;
        RECT 352.950 82.950 355.050 83.400 ;
        RECT 367.950 84.600 370.050 85.050 ;
        RECT 409.950 84.600 412.050 85.050 ;
        RECT 367.950 83.400 412.050 84.600 ;
        RECT 367.950 82.950 370.050 83.400 ;
        RECT 409.950 82.950 412.050 83.400 ;
        RECT 424.950 84.600 427.050 85.050 ;
        RECT 469.950 84.600 472.050 85.050 ;
        RECT 424.950 83.400 472.050 84.600 ;
        RECT 424.950 82.950 427.050 83.400 ;
        RECT 469.950 82.950 472.050 83.400 ;
        RECT 505.950 84.600 508.050 85.050 ;
        RECT 541.950 84.600 544.050 85.050 ;
        RECT 622.950 84.600 625.050 85.050 ;
        RECT 505.950 83.400 522.600 84.600 ;
        RECT 505.950 82.950 508.050 83.400 ;
        RECT 217.950 81.600 220.050 82.050 ;
        RECT 262.950 81.600 265.050 82.050 ;
        RECT 316.950 81.600 319.050 82.050 ;
        RECT 217.950 80.400 319.050 81.600 ;
        RECT 521.400 81.600 522.600 83.400 ;
        RECT 541.950 83.400 625.050 84.600 ;
        RECT 541.950 82.950 544.050 83.400 ;
        RECT 622.950 82.950 625.050 83.400 ;
        RECT 538.950 81.600 541.050 82.050 ;
        RECT 521.400 80.400 541.050 81.600 ;
        RECT 217.950 79.950 220.050 80.400 ;
        RECT 262.950 79.950 265.050 80.400 ;
        RECT 316.950 79.950 319.050 80.400 ;
        RECT 538.950 79.950 541.050 80.400 ;
        RECT 856.950 81.600 859.050 82.050 ;
        RECT 865.950 81.600 868.050 82.050 ;
        RECT 877.950 81.600 880.050 82.050 ;
        RECT 856.950 80.400 880.050 81.600 ;
        RECT 856.950 79.950 859.050 80.400 ;
        RECT 865.950 79.950 868.050 80.400 ;
        RECT 877.950 79.950 880.050 80.400 ;
        RECT 376.950 78.600 379.050 79.050 ;
        RECT 385.950 78.600 388.050 79.050 ;
        RECT 391.950 78.600 394.050 79.050 ;
        RECT 376.950 77.400 394.050 78.600 ;
        RECT 376.950 76.950 379.050 77.400 ;
        RECT 385.950 76.950 388.050 77.400 ;
        RECT 391.950 76.950 394.050 77.400 ;
        RECT 472.950 78.600 475.050 79.050 ;
        RECT 517.950 78.600 520.050 79.050 ;
        RECT 541.950 78.600 544.050 79.050 ;
        RECT 706.950 78.600 709.050 79.050 ;
        RECT 724.950 78.600 727.050 79.050 ;
        RECT 796.950 78.600 799.050 79.050 ;
        RECT 472.950 77.400 520.050 78.600 ;
        RECT 472.950 76.950 475.050 77.400 ;
        RECT 517.950 76.950 520.050 77.400 ;
        RECT 521.400 77.400 540.600 78.600 ;
        RECT 46.950 75.600 49.050 76.050 ;
        RECT 58.950 75.600 61.050 76.050 ;
        RECT 343.950 75.600 346.050 76.050 ;
        RECT 46.950 74.400 346.050 75.600 ;
        RECT 46.950 73.950 49.050 74.400 ;
        RECT 58.950 73.950 61.050 74.400 ;
        RECT 343.950 73.950 346.050 74.400 ;
        RECT 499.950 75.600 502.050 76.050 ;
        RECT 521.400 75.600 522.600 77.400 ;
        RECT 499.950 74.400 522.600 75.600 ;
        RECT 539.400 75.600 540.600 77.400 ;
        RECT 541.950 77.400 645.600 78.600 ;
        RECT 541.950 76.950 544.050 77.400 ;
        RECT 644.400 76.050 645.600 77.400 ;
        RECT 706.950 77.400 799.050 78.600 ;
        RECT 706.950 76.950 709.050 77.400 ;
        RECT 724.950 76.950 727.050 77.400 ;
        RECT 796.950 76.950 799.050 77.400 ;
        RECT 583.950 75.600 586.050 76.050 ;
        RECT 539.400 74.400 586.050 75.600 ;
        RECT 499.950 73.950 502.050 74.400 ;
        RECT 583.950 73.950 586.050 74.400 ;
        RECT 643.950 75.600 646.050 76.050 ;
        RECT 658.950 75.600 661.050 76.050 ;
        RECT 643.950 74.400 661.050 75.600 ;
        RECT 643.950 73.950 646.050 74.400 ;
        RECT 658.950 73.950 661.050 74.400 ;
        RECT 757.950 75.600 760.050 76.050 ;
        RECT 763.950 75.600 766.050 76.050 ;
        RECT 757.950 74.400 766.050 75.600 ;
        RECT 757.950 73.950 760.050 74.400 ;
        RECT 763.950 73.950 766.050 74.400 ;
        RECT 772.950 75.600 775.050 76.050 ;
        RECT 817.950 75.600 820.050 76.050 ;
        RECT 838.950 75.600 841.050 76.050 ;
        RECT 772.950 74.400 841.050 75.600 ;
        RECT 772.950 73.950 775.050 74.400 ;
        RECT 817.950 73.950 820.050 74.400 ;
        RECT 838.950 73.950 841.050 74.400 ;
        RECT 439.950 72.600 442.050 73.050 ;
        RECT 463.950 72.600 466.050 73.050 ;
        RECT 478.950 72.600 481.050 73.050 ;
        RECT 535.950 72.600 538.050 73.050 ;
        RECT 439.950 71.400 538.050 72.600 ;
        RECT 439.950 70.950 442.050 71.400 ;
        RECT 463.950 70.950 466.050 71.400 ;
        RECT 478.950 70.950 481.050 71.400 ;
        RECT 535.950 70.950 538.050 71.400 ;
        RECT 613.950 72.600 616.050 73.050 ;
        RECT 739.950 72.600 742.050 73.050 ;
        RECT 613.950 71.400 742.050 72.600 ;
        RECT 613.950 70.950 616.050 71.400 ;
        RECT 739.950 70.950 742.050 71.400 ;
        RECT 40.950 69.600 43.050 70.050 ;
        RECT 61.800 69.600 63.900 70.050 ;
        RECT 40.950 68.400 63.900 69.600 ;
        RECT 40.950 67.950 43.050 68.400 ;
        RECT 61.800 67.950 63.900 68.400 ;
        RECT 64.950 69.600 67.050 70.050 ;
        RECT 73.950 69.600 76.050 70.050 ;
        RECT 106.950 69.600 109.050 70.050 ;
        RECT 64.950 68.400 109.050 69.600 ;
        RECT 64.950 67.950 67.050 68.400 ;
        RECT 73.950 67.950 76.050 68.400 ;
        RECT 106.950 67.950 109.050 68.400 ;
        RECT 118.950 69.600 121.050 70.050 ;
        RECT 124.950 69.600 127.050 70.050 ;
        RECT 118.950 68.400 127.050 69.600 ;
        RECT 118.950 67.950 121.050 68.400 ;
        RECT 124.950 67.950 127.050 68.400 ;
        RECT 388.950 69.600 391.050 70.050 ;
        RECT 397.950 69.600 400.050 70.050 ;
        RECT 388.950 68.400 400.050 69.600 ;
        RECT 388.950 67.950 391.050 68.400 ;
        RECT 397.950 67.950 400.050 68.400 ;
        RECT 403.950 69.600 406.050 70.050 ;
        RECT 466.950 69.600 469.050 70.050 ;
        RECT 499.950 69.600 502.050 70.050 ;
        RECT 403.950 68.400 459.600 69.600 ;
        RECT 403.950 67.950 406.050 68.400 ;
        RECT 286.950 66.600 289.050 67.050 ;
        RECT 295.950 66.600 298.050 67.050 ;
        RECT 316.950 66.600 319.050 67.050 ;
        RECT 286.950 65.400 319.050 66.600 ;
        RECT 458.400 66.600 459.600 68.400 ;
        RECT 466.950 68.400 502.050 69.600 ;
        RECT 466.950 67.950 469.050 68.400 ;
        RECT 499.950 67.950 502.050 68.400 ;
        RECT 514.950 69.600 517.050 70.050 ;
        RECT 532.950 69.600 535.050 70.050 ;
        RECT 514.950 68.400 535.050 69.600 ;
        RECT 514.950 67.950 517.050 68.400 ;
        RECT 532.950 67.950 535.050 68.400 ;
        RECT 826.950 69.600 829.050 70.050 ;
        RECT 850.950 69.600 853.050 70.050 ;
        RECT 826.950 68.400 853.050 69.600 ;
        RECT 826.950 67.950 829.050 68.400 ;
        RECT 850.950 67.950 853.050 68.400 ;
        RECT 856.950 69.600 859.050 70.050 ;
        RECT 880.950 69.600 883.050 70.050 ;
        RECT 856.950 68.400 883.050 69.600 ;
        RECT 856.950 67.950 859.050 68.400 ;
        RECT 880.950 67.950 883.050 68.400 ;
        RECT 508.950 66.600 511.050 67.050 ;
        RECT 458.400 65.400 511.050 66.600 ;
        RECT 286.950 64.950 289.050 65.400 ;
        RECT 295.950 64.950 298.050 65.400 ;
        RECT 316.950 64.950 319.050 65.400 ;
        RECT 508.950 64.950 511.050 65.400 ;
        RECT 520.950 66.600 523.050 67.050 ;
        RECT 541.950 66.600 544.050 67.050 ;
        RECT 520.950 65.400 544.050 66.600 ;
        RECT 520.950 64.950 523.050 65.400 ;
        RECT 541.950 64.950 544.050 65.400 ;
        RECT 580.950 66.600 583.050 67.050 ;
        RECT 652.950 66.600 655.050 67.050 ;
        RECT 580.950 65.400 655.050 66.600 ;
        RECT 580.950 64.950 583.050 65.400 ;
        RECT 652.950 64.950 655.050 65.400 ;
        RECT 661.950 66.600 664.050 67.050 ;
        RECT 670.950 66.600 673.050 67.050 ;
        RECT 682.950 66.600 685.050 67.050 ;
        RECT 757.950 66.600 760.050 67.050 ;
        RECT 661.950 65.400 673.050 66.600 ;
        RECT 661.950 64.950 664.050 65.400 ;
        RECT 670.950 64.950 673.050 65.400 ;
        RECT 674.400 65.400 760.050 66.600 ;
        RECT 67.950 63.600 70.050 64.050 ;
        RECT 82.950 63.600 85.050 64.050 ;
        RECT 67.950 62.400 85.050 63.600 ;
        RECT 67.950 61.950 70.050 62.400 ;
        RECT 82.950 61.950 85.050 62.400 ;
        RECT 319.950 63.600 322.050 64.050 ;
        RECT 328.950 63.600 331.050 64.050 ;
        RECT 319.950 62.400 331.050 63.600 ;
        RECT 319.950 61.950 322.050 62.400 ;
        RECT 328.950 61.950 331.050 62.400 ;
        RECT 373.950 63.600 376.050 64.050 ;
        RECT 391.950 63.600 394.050 64.050 ;
        RECT 373.950 62.400 394.050 63.600 ;
        RECT 373.950 61.950 376.050 62.400 ;
        RECT 391.950 61.950 394.050 62.400 ;
        RECT 517.950 63.600 520.050 64.050 ;
        RECT 547.950 63.600 550.050 64.050 ;
        RECT 562.950 63.600 565.050 64.050 ;
        RECT 517.950 62.400 565.050 63.600 ;
        RECT 517.950 61.950 520.050 62.400 ;
        RECT 547.950 61.950 550.050 62.400 ;
        RECT 562.950 61.950 565.050 62.400 ;
        RECT 625.950 63.600 628.050 64.050 ;
        RECT 631.950 63.600 634.050 64.050 ;
        RECT 625.950 62.400 634.050 63.600 ;
        RECT 625.950 61.950 628.050 62.400 ;
        RECT 631.950 61.950 634.050 62.400 ;
        RECT 658.950 63.600 661.050 63.900 ;
        RECT 674.400 63.600 675.600 65.400 ;
        RECT 682.950 64.950 685.050 65.400 ;
        RECT 757.950 64.950 760.050 65.400 ;
        RECT 658.950 62.400 675.600 63.600 ;
        RECT 658.950 61.800 661.050 62.400 ;
        RECT 685.950 61.950 688.050 64.050 ;
        RECT 718.950 63.600 721.050 64.050 ;
        RECT 730.950 63.600 733.050 64.050 ;
        RECT 751.950 63.600 754.050 64.050 ;
        RECT 718.950 62.400 754.050 63.600 ;
        RECT 718.950 61.950 721.050 62.400 ;
        RECT 730.950 61.950 733.050 62.400 ;
        RECT 751.950 61.950 754.050 62.400 ;
        RECT 802.950 63.600 805.050 64.050 ;
        RECT 805.950 63.600 808.050 64.050 ;
        RECT 811.950 63.600 814.050 64.050 ;
        RECT 856.950 63.600 859.050 64.050 ;
        RECT 802.950 62.400 814.050 63.600 ;
        RECT 802.950 61.950 805.050 62.400 ;
        RECT 805.950 61.950 808.050 62.400 ;
        RECT 811.950 61.950 814.050 62.400 ;
        RECT 842.400 62.400 859.050 63.600 ;
        RECT 16.950 60.600 19.050 61.200 ;
        RECT 34.950 60.600 37.050 61.200 ;
        RECT 16.950 59.400 37.050 60.600 ;
        RECT 16.950 59.100 19.050 59.400 ;
        RECT 34.950 59.100 37.050 59.400 ;
        RECT 49.950 60.750 52.050 61.200 ;
        RECT 64.950 60.750 67.050 61.200 ;
        RECT 49.950 59.550 67.050 60.750 ;
        RECT 49.950 59.100 52.050 59.550 ;
        RECT 64.950 59.100 67.050 59.550 ;
        RECT 94.950 60.750 97.050 61.200 ;
        RECT 100.950 60.750 103.050 61.200 ;
        RECT 94.950 59.550 103.050 60.750 ;
        RECT 94.950 59.100 97.050 59.550 ;
        RECT 100.950 59.100 103.050 59.550 ;
        RECT 106.950 60.600 109.050 61.200 ;
        RECT 124.950 60.600 127.050 61.200 ;
        RECT 106.950 59.400 127.050 60.600 ;
        RECT 106.950 59.100 109.050 59.400 ;
        RECT 124.950 59.100 127.050 59.400 ;
        RECT 133.950 60.750 136.050 61.200 ;
        RECT 145.950 60.750 148.050 61.200 ;
        RECT 133.950 59.550 148.050 60.750 ;
        RECT 133.950 59.100 136.050 59.550 ;
        RECT 145.950 59.100 148.050 59.550 ;
        RECT 166.950 59.100 169.050 61.200 ;
        RECT 187.950 60.600 190.050 61.050 ;
        RECT 193.950 60.600 196.050 61.200 ;
        RECT 187.950 59.400 196.050 60.600 ;
        RECT 146.400 57.600 147.600 59.100 ;
        RECT 167.400 57.600 168.600 59.100 ;
        RECT 187.950 58.950 190.050 59.400 ;
        RECT 193.950 59.100 196.050 59.400 ;
        RECT 253.950 60.600 256.050 61.200 ;
        RECT 274.950 60.600 277.050 61.200 ;
        RECT 253.950 59.400 277.050 60.600 ;
        RECT 253.950 59.100 256.050 59.400 ;
        RECT 274.950 59.100 277.050 59.400 ;
        RECT 322.950 59.100 325.050 61.200 ;
        RECT 430.950 60.600 433.050 61.200 ;
        RECT 466.950 60.750 469.050 61.200 ;
        RECT 472.950 60.750 475.050 61.200 ;
        RECT 466.950 60.600 475.050 60.750 ;
        RECT 493.950 60.600 496.050 61.200 ;
        RECT 430.950 59.550 496.050 60.600 ;
        RECT 430.950 59.400 469.050 59.550 ;
        RECT 430.950 59.100 433.050 59.400 ;
        RECT 466.950 59.100 469.050 59.400 ;
        RECT 472.950 59.400 496.050 59.550 ;
        RECT 472.950 59.100 475.050 59.400 ;
        RECT 493.950 59.100 496.050 59.400 ;
        RECT 529.950 60.600 532.050 61.050 ;
        RECT 541.950 60.600 544.050 61.200 ;
        RECT 529.950 59.400 544.050 60.600 ;
        RECT 146.400 56.400 168.600 57.600 ;
        RECT 307.950 57.600 310.050 58.050 ;
        RECT 323.400 57.600 324.600 59.100 ;
        RECT 529.950 58.950 532.050 59.400 ;
        RECT 541.950 59.100 544.050 59.400 ;
        RECT 568.950 60.750 571.050 61.200 ;
        RECT 577.950 60.750 580.050 61.200 ;
        RECT 568.950 59.550 580.050 60.750 ;
        RECT 568.950 59.100 571.050 59.550 ;
        RECT 577.950 59.100 580.050 59.550 ;
        RECT 589.950 59.100 592.050 61.200 ;
        RECT 634.950 60.600 637.050 61.200 ;
        RECT 646.950 60.600 649.050 61.050 ;
        RECT 634.950 59.400 649.050 60.600 ;
        RECT 634.950 59.100 637.050 59.400 ;
        RECT 307.950 56.400 324.600 57.600 ;
        RECT 307.950 55.950 310.050 56.400 ;
        RECT 590.400 55.050 591.600 59.100 ;
        RECT 646.950 58.950 649.050 59.400 ;
        RECT 667.950 60.750 670.050 61.200 ;
        RECT 676.950 60.750 679.050 61.200 ;
        RECT 667.950 59.550 679.050 60.750 ;
        RECT 667.950 59.100 670.050 59.550 ;
        RECT 676.950 59.100 679.050 59.550 ;
        RECT 604.950 57.600 607.050 58.050 ;
        RECT 686.400 57.600 687.600 61.950 ;
        RECT 842.400 61.200 843.600 62.400 ;
        RECT 856.950 61.950 859.050 62.400 ;
        RECT 694.950 60.750 697.050 61.200 ;
        RECT 700.950 60.750 703.050 61.200 ;
        RECT 694.950 59.550 703.050 60.750 ;
        RECT 694.950 59.100 697.050 59.550 ;
        RECT 700.950 59.100 703.050 59.550 ;
        RECT 721.950 58.950 724.050 61.050 ;
        RECT 757.950 59.100 760.050 61.200 ;
        RECT 778.950 60.750 781.050 61.200 ;
        RECT 793.950 60.750 796.050 61.200 ;
        RECT 778.950 59.550 796.050 60.750 ;
        RECT 778.950 59.100 781.050 59.550 ;
        RECT 793.950 59.100 796.050 59.550 ;
        RECT 814.950 60.600 817.050 61.050 ;
        RECT 820.950 60.600 823.050 61.050 ;
        RECT 814.950 59.400 823.050 60.600 ;
        RECT 604.950 56.400 657.600 57.600 ;
        RECT 604.950 55.950 607.050 56.400 ;
        RECT 25.950 54.600 28.050 55.050 ;
        RECT 31.950 54.600 34.050 55.050 ;
        RECT 25.950 53.400 34.050 54.600 ;
        RECT 25.950 52.950 28.050 53.400 ;
        RECT 31.950 52.950 34.050 53.400 ;
        RECT 37.950 54.600 40.050 54.900 ;
        RECT 49.950 54.600 52.050 55.050 ;
        RECT 37.950 53.400 52.050 54.600 ;
        RECT 37.950 52.800 40.050 53.400 ;
        RECT 49.950 52.950 52.050 53.400 ;
        RECT 61.950 54.600 64.050 54.900 ;
        RECT 70.950 54.600 73.050 55.050 ;
        RECT 61.950 53.400 73.050 54.600 ;
        RECT 61.950 52.800 64.050 53.400 ;
        RECT 70.950 52.950 73.050 53.400 ;
        RECT 91.950 54.600 94.050 55.050 ;
        RECT 109.950 54.600 112.050 54.900 ;
        RECT 91.950 54.450 112.050 54.600 ;
        RECT 118.950 54.450 121.050 54.900 ;
        RECT 91.950 53.400 121.050 54.450 ;
        RECT 91.950 52.950 94.050 53.400 ;
        RECT 109.950 53.250 121.050 53.400 ;
        RECT 109.950 52.800 112.050 53.250 ;
        RECT 118.950 52.800 121.050 53.250 ;
        RECT 148.950 54.600 151.050 54.900 ;
        RECT 196.950 54.600 199.050 54.900 ;
        RECT 208.950 54.600 211.050 55.050 ;
        RECT 148.950 53.400 211.050 54.600 ;
        RECT 148.950 52.800 151.050 53.400 ;
        RECT 196.950 52.800 199.050 53.400 ;
        RECT 208.950 52.950 211.050 53.400 ;
        RECT 262.950 54.450 265.050 54.900 ;
        RECT 271.950 54.450 274.050 54.900 ;
        RECT 262.950 53.250 274.050 54.450 ;
        RECT 262.950 52.800 265.050 53.250 ;
        RECT 271.950 52.800 274.050 53.250 ;
        RECT 280.950 54.600 283.050 55.050 ;
        RECT 292.950 54.600 295.050 54.900 ;
        RECT 280.950 53.400 295.050 54.600 ;
        RECT 280.950 52.950 283.050 53.400 ;
        RECT 292.950 52.800 295.050 53.400 ;
        RECT 319.950 54.600 322.050 54.900 ;
        RECT 367.950 54.600 370.050 55.050 ;
        RECT 319.950 53.400 370.050 54.600 ;
        RECT 319.950 52.800 322.050 53.400 ;
        RECT 367.950 52.950 370.050 53.400 ;
        RECT 433.950 54.450 436.050 54.900 ;
        RECT 439.950 54.450 442.050 54.900 ;
        RECT 433.950 53.250 442.050 54.450 ;
        RECT 433.950 52.800 436.050 53.250 ;
        RECT 439.950 52.800 442.050 53.250 ;
        RECT 451.950 54.600 454.050 54.900 ;
        RECT 466.950 54.600 469.050 55.050 ;
        RECT 451.950 53.400 469.050 54.600 ;
        RECT 451.950 52.800 454.050 53.400 ;
        RECT 466.950 52.950 469.050 53.400 ;
        RECT 475.950 54.600 478.050 54.900 ;
        RECT 484.950 54.600 487.050 55.050 ;
        RECT 475.950 53.400 487.050 54.600 ;
        RECT 475.950 52.800 478.050 53.400 ;
        RECT 484.950 52.950 487.050 53.400 ;
        RECT 496.950 54.600 499.050 54.900 ;
        RECT 514.950 54.600 517.050 55.050 ;
        RECT 496.950 53.400 517.050 54.600 ;
        RECT 496.950 52.800 499.050 53.400 ;
        RECT 514.950 52.950 517.050 53.400 ;
        RECT 523.950 54.450 526.050 54.900 ;
        RECT 529.950 54.450 532.050 54.900 ;
        RECT 523.950 53.250 532.050 54.450 ;
        RECT 523.950 52.800 526.050 53.250 ;
        RECT 529.950 52.800 532.050 53.250 ;
        RECT 571.950 54.600 574.050 54.900 ;
        RECT 580.950 54.600 583.050 55.050 ;
        RECT 571.950 53.400 583.050 54.600 ;
        RECT 571.950 52.800 574.050 53.400 ;
        RECT 580.950 52.950 583.050 53.400 ;
        RECT 586.950 54.600 591.600 55.050 ;
        RECT 616.950 54.600 619.050 54.900 ;
        RECT 586.950 53.400 619.050 54.600 ;
        RECT 586.950 52.950 591.000 53.400 ;
        RECT 616.950 52.800 619.050 53.400 ;
        RECT 625.950 54.600 628.050 55.050 ;
        RECT 640.950 54.600 643.050 55.050 ;
        RECT 656.400 54.900 657.600 56.400 ;
        RECT 677.400 56.400 687.600 57.600 ;
        RECT 625.950 53.400 643.050 54.600 ;
        RECT 625.950 52.950 628.050 53.400 ;
        RECT 640.950 52.950 643.050 53.400 ;
        RECT 655.950 52.800 658.050 54.900 ;
        RECT 661.950 54.600 664.050 54.900 ;
        RECT 677.400 54.600 678.600 56.400 ;
        RECT 661.950 53.400 678.600 54.600 ;
        RECT 679.950 54.600 682.050 54.900 ;
        RECT 694.950 54.600 697.050 55.050 ;
        RECT 679.950 53.400 697.050 54.600 ;
        RECT 661.950 52.800 664.050 53.400 ;
        RECT 679.950 52.800 682.050 53.400 ;
        RECT 694.950 52.950 697.050 53.400 ;
        RECT 709.950 54.600 712.050 54.900 ;
        RECT 715.950 54.600 718.050 55.050 ;
        RECT 709.950 53.400 718.050 54.600 ;
        RECT 709.950 52.800 712.050 53.400 ;
        RECT 715.950 52.950 718.050 53.400 ;
        RECT 115.950 51.600 118.050 52.050 ;
        RECT 127.950 51.600 130.050 52.050 ;
        RECT 115.950 50.400 130.050 51.600 ;
        RECT 115.950 49.950 118.050 50.400 ;
        RECT 127.950 49.950 130.050 50.400 ;
        RECT 256.950 51.600 259.050 52.050 ;
        RECT 265.950 51.600 268.050 52.050 ;
        RECT 256.950 50.400 268.050 51.600 ;
        RECT 256.950 49.950 259.050 50.400 ;
        RECT 265.950 49.950 268.050 50.400 ;
        RECT 343.950 51.600 346.050 52.050 ;
        RECT 376.950 51.600 379.050 52.050 ;
        RECT 343.950 50.400 379.050 51.600 ;
        RECT 530.400 51.600 531.600 52.800 ;
        RECT 565.950 51.600 568.050 52.050 ;
        RECT 530.400 50.400 568.050 51.600 ;
        RECT 343.950 49.950 346.050 50.400 ;
        RECT 376.950 49.950 379.050 50.400 ;
        RECT 565.950 49.950 568.050 50.400 ;
        RECT 592.950 51.600 595.050 52.050 ;
        RECT 604.950 51.600 607.050 52.050 ;
        RECT 592.950 50.400 607.050 51.600 ;
        RECT 592.950 49.950 595.050 50.400 ;
        RECT 604.950 49.950 607.050 50.400 ;
        RECT 685.950 51.600 688.050 52.050 ;
        RECT 691.950 51.600 694.050 52.050 ;
        RECT 685.950 50.400 694.050 51.600 ;
        RECT 685.950 49.950 688.050 50.400 ;
        RECT 691.950 49.950 694.050 50.400 ;
        RECT 700.950 51.600 703.050 52.050 ;
        RECT 718.950 51.600 721.050 52.050 ;
        RECT 700.950 50.400 721.050 51.600 ;
        RECT 722.400 51.600 723.600 58.950 ;
        RECT 758.400 57.600 759.600 59.100 ;
        RECT 814.950 58.950 817.050 59.400 ;
        RECT 820.950 58.950 823.050 59.400 ;
        RECT 832.950 60.750 835.050 61.200 ;
        RECT 841.950 60.750 844.050 61.200 ;
        RECT 832.950 59.550 844.050 60.750 ;
        RECT 859.950 60.750 862.050 61.200 ;
        RECT 874.950 60.750 877.050 61.200 ;
        RECT 859.950 60.600 877.050 60.750 ;
        RECT 832.950 59.100 835.050 59.550 ;
        RECT 841.950 59.100 844.050 59.550 ;
        RECT 854.400 59.550 877.050 60.600 ;
        RECT 854.400 59.400 862.050 59.550 ;
        RECT 758.400 56.400 771.600 57.600 ;
        RECT 733.950 54.450 736.050 54.900 ;
        RECT 739.950 54.600 742.050 54.900 ;
        RECT 748.950 54.600 751.050 54.900 ;
        RECT 739.950 54.450 751.050 54.600 ;
        RECT 733.950 53.400 751.050 54.450 ;
        RECT 733.950 53.250 742.050 53.400 ;
        RECT 733.950 52.800 736.050 53.250 ;
        RECT 739.950 52.800 742.050 53.250 ;
        RECT 748.950 52.800 751.050 53.400 ;
        RECT 754.950 54.600 757.050 54.900 ;
        RECT 763.950 54.600 766.050 55.050 ;
        RECT 754.950 53.400 766.050 54.600 ;
        RECT 770.400 54.600 771.600 56.400 ;
        RECT 854.400 54.900 855.600 59.400 ;
        RECT 859.950 59.100 862.050 59.400 ;
        RECT 874.950 59.100 877.050 59.550 ;
        RECT 775.950 54.600 778.050 54.900 ;
        RECT 770.400 53.400 778.050 54.600 ;
        RECT 754.950 52.800 757.050 53.400 ;
        RECT 763.950 52.950 766.050 53.400 ;
        RECT 775.950 52.800 778.050 53.400 ;
        RECT 781.950 54.600 784.050 54.900 ;
        RECT 805.950 54.600 808.050 54.900 ;
        RECT 823.950 54.600 826.050 54.900 ;
        RECT 781.950 53.400 826.050 54.600 ;
        RECT 781.950 52.800 784.050 53.400 ;
        RECT 805.950 52.800 808.050 53.400 ;
        RECT 823.950 52.800 826.050 53.400 ;
        RECT 829.950 54.600 832.050 54.900 ;
        RECT 853.950 54.600 856.050 54.900 ;
        RECT 829.950 53.400 856.050 54.600 ;
        RECT 829.950 52.800 832.050 53.400 ;
        RECT 853.950 52.800 856.050 53.400 ;
        RECT 727.950 51.600 730.050 52.050 ;
        RECT 722.400 50.400 730.050 51.600 ;
        RECT 700.950 49.950 703.050 50.400 ;
        RECT 718.950 49.950 721.050 50.400 ;
        RECT 727.950 49.950 730.050 50.400 ;
        RECT 766.950 51.600 769.050 52.050 ;
        RECT 799.950 51.600 802.050 52.050 ;
        RECT 766.950 50.400 802.050 51.600 ;
        RECT 766.950 49.950 769.050 50.400 ;
        RECT 799.950 49.950 802.050 50.400 ;
        RECT 838.950 51.600 841.050 52.050 ;
        RECT 847.950 51.600 850.050 52.050 ;
        RECT 838.950 50.400 850.050 51.600 ;
        RECT 838.950 49.950 841.050 50.400 ;
        RECT 847.950 49.950 850.050 50.400 ;
        RECT 202.950 48.600 205.050 49.050 ;
        RECT 298.950 48.600 301.050 49.050 ;
        RECT 307.800 48.600 309.900 49.050 ;
        RECT 202.950 47.400 309.900 48.600 ;
        RECT 202.950 46.950 205.050 47.400 ;
        RECT 298.950 46.950 301.050 47.400 ;
        RECT 307.800 46.950 309.900 47.400 ;
        RECT 310.950 48.600 313.050 49.050 ;
        RECT 373.950 48.600 376.050 49.050 ;
        RECT 310.950 47.400 376.050 48.600 ;
        RECT 310.950 46.950 313.050 47.400 ;
        RECT 373.950 46.950 376.050 47.400 ;
        RECT 379.950 48.600 382.050 49.050 ;
        RECT 427.950 48.600 430.050 49.050 ;
        RECT 379.950 47.400 430.050 48.600 ;
        RECT 379.950 46.950 382.050 47.400 ;
        RECT 427.950 46.950 430.050 47.400 ;
        RECT 616.950 48.600 619.050 49.050 ;
        RECT 631.950 48.600 634.050 49.050 ;
        RECT 616.950 47.400 634.050 48.600 ;
        RECT 616.950 46.950 619.050 47.400 ;
        RECT 631.950 46.950 634.050 47.400 ;
        RECT 655.950 48.600 658.050 49.050 ;
        RECT 667.950 48.600 670.050 49.050 ;
        RECT 703.950 48.600 706.050 49.050 ;
        RECT 655.950 47.400 706.050 48.600 ;
        RECT 655.950 46.950 658.050 47.400 ;
        RECT 667.950 46.950 670.050 47.400 ;
        RECT 703.950 46.950 706.050 47.400 ;
        RECT 19.950 45.600 22.050 46.050 ;
        RECT 61.950 45.600 64.050 46.050 ;
        RECT 94.950 45.600 97.050 46.050 ;
        RECT 19.950 44.400 97.050 45.600 ;
        RECT 19.950 43.950 22.050 44.400 ;
        RECT 61.950 43.950 64.050 44.400 ;
        RECT 94.950 43.950 97.050 44.400 ;
        RECT 127.950 45.600 130.050 46.050 ;
        RECT 157.950 45.600 160.050 46.050 ;
        RECT 169.950 45.600 172.050 46.050 ;
        RECT 373.950 45.600 376.050 45.900 ;
        RECT 127.950 44.400 376.050 45.600 ;
        RECT 127.950 43.950 130.050 44.400 ;
        RECT 157.950 43.950 160.050 44.400 ;
        RECT 169.950 43.950 172.050 44.400 ;
        RECT 373.950 43.800 376.050 44.400 ;
        RECT 544.950 45.600 547.050 46.050 ;
        RECT 589.950 45.600 592.050 46.050 ;
        RECT 601.950 45.600 604.050 46.050 ;
        RECT 610.950 45.600 613.050 46.050 ;
        RECT 544.950 44.400 613.050 45.600 ;
        RECT 544.950 43.950 547.050 44.400 ;
        RECT 589.950 43.950 592.050 44.400 ;
        RECT 601.950 43.950 604.050 44.400 ;
        RECT 610.950 43.950 613.050 44.400 ;
        RECT 646.950 45.600 649.050 46.050 ;
        RECT 652.950 45.600 655.050 46.050 ;
        RECT 646.950 44.400 655.050 45.600 ;
        RECT 646.950 43.950 649.050 44.400 ;
        RECT 652.950 43.950 655.050 44.400 ;
        RECT 658.950 45.600 661.050 46.050 ;
        RECT 700.950 45.600 703.050 46.050 ;
        RECT 658.950 44.400 703.050 45.600 ;
        RECT 658.950 43.950 661.050 44.400 ;
        RECT 700.950 43.950 703.050 44.400 ;
        RECT 844.950 45.600 847.050 46.050 ;
        RECT 895.950 45.600 898.050 46.050 ;
        RECT 844.950 44.400 898.050 45.600 ;
        RECT 844.950 43.950 847.050 44.400 ;
        RECT 895.950 43.950 898.050 44.400 ;
        RECT 223.950 42.600 226.050 43.050 ;
        RECT 241.950 42.600 244.050 43.050 ;
        RECT 223.950 41.400 244.050 42.600 ;
        RECT 223.950 40.950 226.050 41.400 ;
        RECT 241.950 40.950 244.050 41.400 ;
        RECT 385.950 42.600 388.050 43.050 ;
        RECT 400.950 42.600 403.050 43.050 ;
        RECT 385.950 41.400 403.050 42.600 ;
        RECT 385.950 40.950 388.050 41.400 ;
        RECT 400.950 40.950 403.050 41.400 ;
        RECT 556.950 42.600 559.050 43.050 ;
        RECT 628.950 42.600 631.050 43.050 ;
        RECT 556.950 41.400 631.050 42.600 ;
        RECT 556.950 40.950 559.050 41.400 ;
        RECT 628.950 40.950 631.050 41.400 ;
        RECT 811.950 42.600 814.050 43.050 ;
        RECT 850.950 42.600 853.050 43.050 ;
        RECT 811.950 41.400 853.050 42.600 ;
        RECT 811.950 40.950 814.050 41.400 ;
        RECT 850.950 40.950 853.050 41.400 ;
        RECT 121.950 39.600 124.050 40.050 ;
        RECT 133.950 39.600 136.050 40.050 ;
        RECT 505.950 39.600 508.050 40.050 ;
        RECT 121.950 38.400 136.050 39.600 ;
        RECT 121.950 37.950 124.050 38.400 ;
        RECT 133.950 37.950 136.050 38.400 ;
        RECT 404.400 38.400 508.050 39.600 ;
        RECT 103.950 36.600 106.050 37.050 ;
        RECT 112.950 36.600 115.050 37.050 ;
        RECT 103.950 35.400 115.050 36.600 ;
        RECT 103.950 34.950 106.050 35.400 ;
        RECT 112.950 34.950 115.050 35.400 ;
        RECT 166.950 36.600 169.050 37.050 ;
        RECT 286.950 36.600 289.050 37.050 ;
        RECT 166.950 35.400 289.050 36.600 ;
        RECT 166.950 34.950 169.050 35.400 ;
        RECT 286.950 34.950 289.050 35.400 ;
        RECT 367.950 36.600 370.050 37.050 ;
        RECT 404.400 36.600 405.600 38.400 ;
        RECT 505.950 37.950 508.050 38.400 ;
        RECT 643.950 39.600 646.050 40.050 ;
        RECT 673.950 39.600 676.050 40.050 ;
        RECT 643.950 38.400 676.050 39.600 ;
        RECT 643.950 37.950 646.050 38.400 ;
        RECT 673.950 37.950 676.050 38.400 ;
        RECT 367.950 35.400 405.600 36.600 ;
        RECT 415.950 36.600 418.050 37.050 ;
        RECT 637.950 36.600 640.050 37.050 ;
        RECT 682.950 36.600 685.050 37.050 ;
        RECT 415.950 35.400 435.600 36.600 ;
        RECT 367.950 34.950 370.050 35.400 ;
        RECT 415.950 34.950 418.050 35.400 ;
        RECT 238.950 33.600 241.050 34.050 ;
        RECT 265.950 33.600 268.050 34.050 ;
        RECT 238.950 32.400 268.050 33.600 ;
        RECT 434.400 33.600 435.600 35.400 ;
        RECT 637.950 35.400 685.050 36.600 ;
        RECT 637.950 34.950 640.050 35.400 ;
        RECT 682.950 34.950 685.050 35.400 ;
        RECT 865.950 36.600 868.050 37.050 ;
        RECT 877.950 36.600 880.050 37.050 ;
        RECT 865.950 35.400 880.050 36.600 ;
        RECT 865.950 34.950 868.050 35.400 ;
        RECT 877.950 34.950 880.050 35.400 ;
        RECT 451.950 33.600 454.050 34.050 ;
        RECT 434.400 32.400 454.050 33.600 ;
        RECT 238.950 31.950 241.050 32.400 ;
        RECT 265.950 31.950 268.050 32.400 ;
        RECT 451.950 31.950 454.050 32.400 ;
        RECT 541.950 33.600 544.050 34.050 ;
        RECT 577.950 33.600 580.050 34.050 ;
        RECT 638.400 33.600 639.600 34.950 ;
        RECT 541.950 32.400 639.600 33.600 ;
        RECT 640.950 33.600 643.050 34.050 ;
        RECT 676.950 33.600 679.050 34.050 ;
        RECT 640.950 32.400 679.050 33.600 ;
        RECT 541.950 31.950 544.050 32.400 ;
        RECT 577.950 31.950 580.050 32.400 ;
        RECT 640.950 31.950 643.050 32.400 ;
        RECT 676.950 31.950 679.050 32.400 ;
        RECT 799.950 33.600 802.050 34.050 ;
        RECT 829.950 33.600 832.050 34.050 ;
        RECT 841.950 33.600 844.050 34.050 ;
        RECT 799.950 32.400 844.050 33.600 ;
        RECT 799.950 31.950 802.050 32.400 ;
        RECT 829.950 31.950 832.050 32.400 ;
        RECT 841.950 31.950 844.050 32.400 ;
        RECT 355.950 30.600 358.050 31.050 ;
        RECT 361.950 30.600 364.050 31.050 ;
        RECT 355.950 29.400 364.050 30.600 ;
        RECT 355.950 28.950 358.050 29.400 ;
        RECT 361.950 28.950 364.050 29.400 ;
        RECT 406.950 30.600 409.050 31.050 ;
        RECT 430.950 30.600 433.050 31.050 ;
        RECT 442.950 30.600 445.050 31.050 ;
        RECT 406.950 29.400 445.050 30.600 ;
        RECT 406.950 28.950 409.050 29.400 ;
        RECT 430.950 28.950 433.050 29.400 ;
        RECT 442.950 28.950 445.050 29.400 ;
        RECT 493.950 30.600 496.050 31.050 ;
        RECT 505.950 30.600 508.050 31.050 ;
        RECT 493.950 29.400 508.050 30.600 ;
        RECT 493.950 28.950 496.050 29.400 ;
        RECT 505.950 28.950 508.050 29.400 ;
        RECT 586.950 28.950 589.050 31.050 ;
        RECT 25.950 27.750 28.050 28.200 ;
        RECT 40.950 27.750 43.050 28.200 ;
        RECT 25.950 27.600 43.050 27.750 ;
        RECT 55.950 27.600 58.050 28.050 ;
        RECT 73.950 27.600 76.050 28.050 ;
        RECT 25.950 26.550 76.050 27.600 ;
        RECT 25.950 26.100 28.050 26.550 ;
        RECT 40.950 26.400 76.050 26.550 ;
        RECT 40.950 26.100 43.050 26.400 ;
        RECT 55.950 25.950 58.050 26.400 ;
        RECT 73.950 25.950 76.050 26.400 ;
        RECT 103.950 27.600 106.050 28.200 ;
        RECT 121.950 27.600 124.050 28.200 ;
        RECT 103.950 26.400 124.050 27.600 ;
        RECT 103.950 26.100 106.050 26.400 ;
        RECT 121.950 26.100 124.050 26.400 ;
        RECT 136.950 27.750 139.050 28.200 ;
        RECT 160.950 27.750 163.050 28.200 ;
        RECT 136.950 27.600 163.050 27.750 ;
        RECT 187.950 27.600 190.050 28.200 ;
        RECT 196.950 27.600 199.050 28.050 ;
        RECT 249.000 27.600 253.050 28.050 ;
        RECT 264.000 27.600 268.050 28.050 ;
        RECT 136.950 26.550 186.600 27.600 ;
        RECT 136.950 26.100 139.050 26.550 ;
        RECT 160.950 26.400 186.600 26.550 ;
        RECT 160.950 26.100 163.050 26.400 ;
        RECT 185.400 24.600 186.600 26.400 ;
        RECT 187.950 26.400 199.050 27.600 ;
        RECT 187.950 26.100 190.050 26.400 ;
        RECT 196.950 25.950 199.050 26.400 ;
        RECT 248.400 25.950 253.050 27.600 ;
        RECT 263.400 25.950 268.050 27.600 ;
        RECT 271.950 27.750 274.050 28.200 ;
        RECT 280.950 27.750 283.050 28.200 ;
        RECT 271.950 26.550 283.050 27.750 ;
        RECT 271.950 26.100 274.050 26.550 ;
        RECT 280.950 26.100 283.050 26.550 ;
        RECT 316.950 27.600 319.050 28.200 ;
        RECT 334.950 27.600 337.050 28.200 ;
        RECT 316.950 26.400 337.050 27.600 ;
        RECT 316.950 26.100 319.050 26.400 ;
        RECT 334.950 26.100 337.050 26.400 ;
        RECT 379.950 27.750 382.050 28.200 ;
        RECT 394.950 27.750 397.050 28.200 ;
        RECT 379.950 26.550 397.050 27.750 ;
        RECT 379.950 26.100 382.050 26.550 ;
        RECT 394.950 26.100 397.050 26.550 ;
        RECT 472.950 27.600 475.050 28.200 ;
        RECT 484.950 27.600 487.050 28.050 ;
        RECT 517.950 27.600 520.050 28.200 ;
        RECT 472.950 26.400 520.050 27.600 ;
        RECT 472.950 26.100 475.050 26.400 ;
        RECT 484.950 25.950 487.050 26.400 ;
        RECT 517.950 26.100 520.050 26.400 ;
        RECT 565.950 27.750 568.050 28.200 ;
        RECT 571.950 27.750 574.050 28.200 ;
        RECT 565.950 26.550 574.050 27.750 ;
        RECT 565.950 26.100 568.050 26.550 ;
        RECT 571.950 26.100 574.050 26.550 ;
        RECT 193.950 24.600 196.050 25.050 ;
        RECT 185.400 23.400 196.050 24.600 ;
        RECT 193.950 22.950 196.050 23.400 ;
        RECT 19.950 21.600 22.050 21.900 ;
        RECT 25.950 21.600 28.050 22.050 ;
        RECT 19.950 20.400 28.050 21.600 ;
        RECT 19.950 19.800 22.050 20.400 ;
        RECT 25.950 19.950 28.050 20.400 ;
        RECT 34.950 21.600 37.050 21.900 ;
        RECT 58.950 21.600 61.050 21.900 ;
        RECT 34.950 20.400 61.050 21.600 ;
        RECT 34.950 19.800 37.050 20.400 ;
        RECT 58.950 19.800 61.050 20.400 ;
        RECT 64.950 21.450 67.050 21.900 ;
        RECT 70.800 21.450 72.900 21.900 ;
        RECT 64.950 20.250 72.900 21.450 ;
        RECT 64.950 19.800 67.050 20.250 ;
        RECT 70.800 19.800 72.900 20.250 ;
        RECT 73.950 21.450 76.050 21.900 ;
        RECT 79.950 21.450 82.050 21.900 ;
        RECT 73.950 20.250 82.050 21.450 ;
        RECT 73.950 19.800 76.050 20.250 ;
        RECT 79.950 19.800 82.050 20.250 ;
        RECT 106.950 21.450 109.050 21.900 ;
        RECT 112.950 21.450 115.050 21.900 ;
        RECT 106.950 20.250 115.050 21.450 ;
        RECT 106.950 19.800 109.050 20.250 ;
        RECT 112.950 19.800 115.050 20.250 ;
        RECT 124.950 21.600 127.050 21.900 ;
        RECT 136.950 21.600 139.050 22.050 ;
        RECT 248.400 21.900 249.600 25.950 ;
        RECT 263.400 21.900 264.600 25.950 ;
        RECT 290.400 23.400 297.600 24.600 ;
        RECT 290.400 21.900 291.600 23.400 ;
        RECT 124.950 20.400 139.050 21.600 ;
        RECT 124.950 19.800 127.050 20.400 ;
        RECT 136.950 19.950 139.050 20.400 ;
        RECT 142.950 21.600 145.050 21.900 ;
        RECT 163.950 21.600 166.050 21.900 ;
        RECT 142.950 20.400 166.050 21.600 ;
        RECT 142.950 19.800 145.050 20.400 ;
        RECT 163.950 19.800 166.050 20.400 ;
        RECT 169.950 21.600 172.050 21.900 ;
        RECT 184.950 21.600 187.050 21.900 ;
        RECT 169.950 20.400 187.050 21.600 ;
        RECT 169.950 19.800 172.050 20.400 ;
        RECT 184.950 19.800 187.050 20.400 ;
        RECT 196.950 21.450 199.050 21.900 ;
        RECT 205.950 21.450 208.050 21.900 ;
        RECT 196.950 20.250 208.050 21.450 ;
        RECT 196.950 19.800 199.050 20.250 ;
        RECT 205.950 19.800 208.050 20.250 ;
        RECT 247.950 19.800 250.050 21.900 ;
        RECT 262.950 19.800 265.050 21.900 ;
        RECT 289.950 19.800 292.050 21.900 ;
        RECT 296.400 21.600 297.600 23.400 ;
        RECT 367.950 21.600 370.050 22.050 ;
        RECT 296.400 20.400 370.050 21.600 ;
        RECT 367.950 19.950 370.050 20.400 ;
        RECT 394.950 21.600 397.050 22.050 ;
        RECT 400.950 21.600 403.050 21.900 ;
        RECT 424.950 21.600 427.050 21.900 ;
        RECT 394.950 20.400 427.050 21.600 ;
        RECT 394.950 19.950 397.050 20.400 ;
        RECT 400.950 19.800 403.050 20.400 ;
        RECT 424.950 19.800 427.050 20.400 ;
        RECT 442.950 21.450 445.050 21.900 ;
        RECT 448.950 21.450 451.050 21.900 ;
        RECT 442.950 20.250 451.050 21.450 ;
        RECT 442.950 19.800 445.050 20.250 ;
        RECT 448.950 19.800 451.050 20.250 ;
        RECT 454.950 21.600 457.050 21.900 ;
        RECT 484.950 21.600 487.050 21.900 ;
        RECT 454.950 21.450 487.050 21.600 ;
        RECT 490.950 21.450 493.050 21.900 ;
        RECT 454.950 20.400 493.050 21.450 ;
        RECT 454.950 19.800 457.050 20.400 ;
        RECT 484.950 20.250 493.050 20.400 ;
        RECT 484.950 19.800 487.050 20.250 ;
        RECT 490.950 19.800 493.050 20.250 ;
        RECT 496.950 21.450 499.050 21.900 ;
        RECT 508.950 21.450 511.050 21.900 ;
        RECT 496.950 20.250 511.050 21.450 ;
        RECT 496.950 19.800 499.050 20.250 ;
        RECT 508.950 19.800 511.050 20.250 ;
        RECT 529.950 21.450 532.050 21.900 ;
        RECT 544.950 21.600 547.050 21.900 ;
        RECT 556.950 21.600 559.050 22.050 ;
        RECT 587.400 21.900 588.600 28.950 ;
        RECT 598.950 27.600 601.050 28.050 ;
        RECT 607.950 27.600 610.050 28.200 ;
        RECT 598.950 26.400 610.050 27.600 ;
        RECT 598.950 25.950 601.050 26.400 ;
        RECT 607.950 26.100 610.050 26.400 ;
        RECT 658.950 27.600 661.050 28.200 ;
        RECT 670.950 27.600 673.050 28.050 ;
        RECT 658.950 26.400 673.050 27.600 ;
        RECT 658.950 26.100 661.050 26.400 ;
        RECT 670.950 25.950 673.050 26.400 ;
        RECT 676.950 27.600 679.050 28.050 ;
        RECT 706.950 27.600 709.050 28.050 ;
        RECT 676.950 26.400 709.050 27.600 ;
        RECT 676.950 25.950 679.050 26.400 ;
        RECT 706.950 25.950 709.050 26.400 ;
        RECT 718.950 26.100 721.050 28.200 ;
        RECT 754.950 27.600 757.050 28.200 ;
        RECT 772.950 27.600 775.050 28.200 ;
        RECT 754.950 26.400 775.050 27.600 ;
        RECT 754.950 26.100 757.050 26.400 ;
        RECT 772.950 26.100 775.050 26.400 ;
        RECT 781.950 27.600 784.050 28.050 ;
        RECT 793.950 27.600 796.050 28.200 ;
        RECT 781.950 26.400 796.050 27.600 ;
        RECT 595.950 24.600 598.050 25.050 ;
        RECT 622.950 24.600 625.050 25.050 ;
        RECT 595.950 23.400 657.600 24.600 ;
        RECT 595.950 22.950 598.050 23.400 ;
        RECT 622.950 22.950 625.050 23.400 ;
        RECT 656.400 21.900 657.600 23.400 ;
        RECT 544.950 21.450 559.050 21.600 ;
        RECT 529.950 20.400 559.050 21.450 ;
        RECT 529.950 20.250 547.050 20.400 ;
        RECT 529.950 19.800 532.050 20.250 ;
        RECT 544.950 19.800 547.050 20.250 ;
        RECT 556.950 19.950 559.050 20.400 ;
        RECT 586.950 19.800 589.050 21.900 ;
        RECT 655.950 19.800 658.050 21.900 ;
        RECT 670.950 21.450 673.050 21.900 ;
        RECT 679.950 21.450 682.050 21.900 ;
        RECT 670.950 20.250 682.050 21.450 ;
        RECT 670.950 19.800 673.050 20.250 ;
        RECT 679.950 19.800 682.050 20.250 ;
        RECT 700.950 21.450 703.050 21.900 ;
        RECT 706.950 21.450 709.050 21.900 ;
        RECT 700.950 20.250 709.050 21.450 ;
        RECT 719.400 21.600 720.600 26.100 ;
        RECT 781.950 25.950 784.050 26.400 ;
        RECT 793.950 26.100 796.050 26.400 ;
        RECT 808.950 27.600 811.050 28.050 ;
        RECT 820.950 27.600 823.050 28.200 ;
        RECT 808.950 26.400 823.050 27.600 ;
        RECT 808.950 25.950 811.050 26.400 ;
        RECT 820.950 26.100 823.050 26.400 ;
        RECT 736.950 21.600 739.050 21.900 ;
        RECT 719.400 20.400 739.050 21.600 ;
        RECT 700.950 19.800 703.050 20.250 ;
        RECT 706.950 19.800 709.050 20.250 ;
        RECT 736.950 19.800 739.050 20.400 ;
        RECT 802.950 21.450 805.050 21.900 ;
        RECT 811.950 21.450 814.050 21.900 ;
        RECT 802.950 20.250 814.050 21.450 ;
        RECT 802.950 19.800 805.050 20.250 ;
        RECT 811.950 19.800 814.050 20.250 ;
        RECT 850.950 21.600 853.050 22.050 ;
        RECT 862.950 21.600 865.050 21.900 ;
        RECT 850.950 20.400 865.050 21.600 ;
        RECT 850.950 19.950 853.050 20.400 ;
        RECT 862.950 19.800 865.050 20.400 ;
        RECT 49.950 18.600 52.050 19.050 ;
        RECT 100.950 18.600 103.050 19.050 ;
        RECT 49.950 17.400 103.050 18.600 ;
        RECT 49.950 16.950 52.050 17.400 ;
        RECT 100.950 16.950 103.050 17.400 ;
        RECT 253.950 18.600 256.050 19.050 ;
        RECT 289.950 18.600 292.050 19.050 ;
        RECT 253.950 17.400 292.050 18.600 ;
        RECT 253.950 16.950 256.050 17.400 ;
        RECT 289.950 16.950 292.050 17.400 ;
        RECT 385.950 18.600 388.050 19.050 ;
        RECT 412.950 18.600 415.050 19.050 ;
        RECT 385.950 17.400 415.050 18.600 ;
        RECT 385.950 16.950 388.050 17.400 ;
        RECT 412.950 16.950 415.050 17.400 ;
        RECT 433.950 18.600 436.050 19.050 ;
        RECT 454.950 18.600 457.050 19.050 ;
        RECT 433.950 17.400 457.050 18.600 ;
        RECT 433.950 16.950 436.050 17.400 ;
        RECT 454.950 16.950 457.050 17.400 ;
        RECT 538.950 18.600 541.050 19.050 ;
        RECT 562.950 18.600 565.050 19.050 ;
        RECT 538.950 17.400 565.050 18.600 ;
        RECT 538.950 16.950 541.050 17.400 ;
        RECT 562.950 16.950 565.050 17.400 ;
        RECT 610.950 18.600 613.050 19.050 ;
        RECT 643.950 18.600 646.050 19.050 ;
        RECT 661.950 18.600 664.050 19.050 ;
        RECT 610.950 17.400 664.050 18.600 ;
        RECT 610.950 16.950 613.050 17.400 ;
        RECT 643.950 16.950 646.050 17.400 ;
        RECT 661.950 16.950 664.050 17.400 ;
        RECT 817.950 18.600 820.050 19.050 ;
        RECT 829.950 18.600 832.050 19.050 ;
        RECT 817.950 17.400 832.050 18.600 ;
        RECT 817.950 16.950 820.050 17.400 ;
        RECT 829.950 16.950 832.050 17.400 ;
        RECT 844.950 18.600 847.050 19.050 ;
        RECT 880.950 18.600 883.050 19.050 ;
        RECT 898.950 18.600 901.050 19.050 ;
        RECT 844.950 17.400 901.050 18.600 ;
        RECT 844.950 16.950 847.050 17.400 ;
        RECT 880.950 16.950 883.050 17.400 ;
        RECT 898.950 16.950 901.050 17.400 ;
        RECT 46.950 15.600 49.050 16.050 ;
        RECT 85.950 15.600 88.050 16.050 ;
        RECT 46.950 14.400 88.050 15.600 ;
        RECT 46.950 13.950 49.050 14.400 ;
        RECT 85.950 13.950 88.050 14.400 ;
        RECT 505.950 15.600 508.050 16.050 ;
        RECT 595.950 15.600 598.050 16.050 ;
        RECT 505.950 14.400 598.050 15.600 ;
        RECT 505.950 13.950 508.050 14.400 ;
        RECT 595.950 13.950 598.050 14.400 ;
        RECT 673.950 15.600 676.050 16.050 ;
        RECT 691.950 15.600 694.050 16.050 ;
        RECT 727.950 15.600 730.050 16.050 ;
        RECT 673.950 14.400 730.050 15.600 ;
        RECT 673.950 13.950 676.050 14.400 ;
        RECT 691.950 13.950 694.050 14.400 ;
        RECT 727.950 13.950 730.050 14.400 ;
        RECT 271.950 12.600 274.050 13.050 ;
        RECT 301.950 12.600 304.050 13.050 ;
        RECT 271.950 11.400 304.050 12.600 ;
        RECT 271.950 10.950 274.050 11.400 ;
        RECT 301.950 10.950 304.050 11.400 ;
        RECT 388.950 12.600 391.050 13.050 ;
        RECT 469.950 12.600 472.050 13.050 ;
        RECT 388.950 11.400 472.050 12.600 ;
        RECT 388.950 10.950 391.050 11.400 ;
        RECT 469.950 10.950 472.050 11.400 ;
        RECT 661.950 12.600 664.050 13.050 ;
        RECT 808.950 12.600 811.050 13.050 ;
        RECT 661.950 11.400 811.050 12.600 ;
        RECT 661.950 10.950 664.050 11.400 ;
        RECT 808.950 10.950 811.050 11.400 ;
        RECT 520.950 9.600 523.050 10.050 ;
        RECT 592.950 9.600 595.050 10.050 ;
        RECT 520.950 8.400 595.050 9.600 ;
        RECT 520.950 7.950 523.050 8.400 ;
        RECT 592.950 7.950 595.050 8.400 ;
        RECT 604.950 9.600 607.050 10.050 ;
        RECT 658.950 9.600 661.050 10.050 ;
        RECT 604.950 8.400 661.050 9.600 ;
        RECT 604.950 7.950 607.050 8.400 ;
        RECT 658.950 7.950 661.050 8.400 ;
        RECT 664.950 9.600 667.050 10.050 ;
        RECT 796.950 9.600 799.050 10.050 ;
        RECT 664.950 8.400 799.050 9.600 ;
        RECT 664.950 7.950 667.050 8.400 ;
        RECT 796.950 7.950 799.050 8.400 ;
        RECT 571.950 6.600 574.050 7.050 ;
        RECT 580.950 6.600 583.050 7.050 ;
        RECT 598.950 6.600 601.050 7.050 ;
        RECT 571.950 5.400 601.050 6.600 ;
        RECT 571.950 4.950 574.050 5.400 ;
        RECT 580.950 4.950 583.050 5.400 ;
        RECT 598.950 4.950 601.050 5.400 ;
        RECT 685.950 6.600 688.050 7.050 ;
        RECT 781.950 6.600 784.050 7.050 ;
        RECT 685.950 5.400 784.050 6.600 ;
        RECT 685.950 4.950 688.050 5.400 ;
        RECT 781.950 4.950 784.050 5.400 ;
  END
END fir_pe
END LIBRARY


/* Verilog module written by vlog2Verilog (qflow) */
/* With explicit power connections */

module fir_pe(
    inout vdd,
    inout gnd,
    input [7:0] Cin,
    input [7:0] Xin,
    output [7:0] Xout,
    input [15:0] Yin,
    output [15:0] Yout,
    input clk
);

wire [15:0] y ;
wire _588_ ;
wire _168_ ;
wire _60_ ;
wire _397_ ;
wire _703_ ;
wire _19_ ;
wire _512_ ;
wire _741_ ;
wire _321_ ;
wire _57_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _415_ ;
wire _95_ ;
wire _644_ ;
wire _224_ ;
wire _453_ ;
wire _509_ ;
wire _682_ ;
wire _262_ ;
wire _738_ ;
wire _318_ ;
wire _491_ ;
wire _547_ ;
wire _127_ ;
wire _356_ ;
wire _585_ ;
wire _165_ ;
wire _394_ ;
wire _679_ ;
wire _259_ ;
wire _488_ ;
wire _700_ ;
wire _297_ ;
wire _16_ ;
wire _54_ ;
wire _603_ ;
wire _412_ ;
wire _92_ ;
wire _641_ ;
wire _221_ ;
wire _450_ ;
wire _506_ ;
wire _735_ ;
wire _315_ ;
wire _544_ ;
wire _124_ ;
wire _353_ ;
wire _409_ ;
wire _89_ ;
wire _582_ ;
wire _162_ ;
wire _638_ ;
wire _218_ ;
wire _391_ ;
wire _447_ ;
wire _676_ ;
wire _256_ ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire _388_ ;
wire _600_ ;
wire _197_ ;
wire _7_ ;
wire _503_ ;
wire _732_ ;
wire _312_ ;
wire _48_ ;
wire _541_ ;
wire _121_ ;
wire _350_ ;
wire _406_ ;
wire _86_ ;
wire _635_ ;
wire _215_ ;
wire _444_ ;
wire _673_ ;
wire _253_ ;
wire _729_ ;
wire _309_ ;
wire _482_ ;
wire _538_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _347_ ;
wire _576_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire _479_ ;
wire _288_ ;
wire _4_ ;
wire _500_ ;
wire _45_ ;
wire _403_ ;
wire _83_ ;
wire _632_ ;
wire _212_ ;
wire _441_ ;
wire _670_ ;
wire _250_ ;
wire _726_ ;
wire _306_ ;
wire _535_ ;
wire _115_ ;
wire _344_ ;
wire _573_ ;
wire _153_ ;
wire _629_ ;
wire _209_ ;
wire Xin_5_bF$buf0 ;
wire Xin_5_bF$buf1 ;
wire Xin_5_bF$buf2 ;
wire Xin_5_bF$buf3 ;
wire _382_ ;
wire _438_ ;
wire _191_ ;
wire _667_ ;
wire _247_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire _285_ ;
wire _1_ ;
wire _42_ ;
wire _379_ ;
wire _188_ ;
wire _400_ ;
wire _80_ ;
wire _723_ ;
wire _303_ ;
wire _39_ ;
wire _532_ ;
wire _112_ ;
wire _341_ ;
wire clk ;
wire _77_ ;
wire _570_ ;
wire _150_ ;
wire _626_ ;
wire _206_ ;
wire _435_ ;
wire _664_ ;
wire _244_ ;
wire _473_ ;
wire _529_ ;
wire _109_ ;
wire _282_ ;
wire _338_ ;
wire _567_ ;
wire _147_ ;
wire _376_ ;
wire _185_ ;
wire _699_ ;
wire _279_ ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire _74_ ;
wire _623_ ;
wire _203_ ;
wire _432_ ;
wire _661_ ;
wire _241_ ;
wire _717_ ;
wire _470_ ;
wire _526_ ;
wire _106_ ;
wire [15:0] _755_ ;
wire _335_ ;
wire _564_ ;
wire _144_ ;
wire _373_ ;
wire _429_ ;
wire _182_ ;
wire _658_ ;
wire _238_ ;
wire _467_ ;
wire _696_ ;
wire _276_ ;
wire _33_ ;
wire _599_ ;
wire _179_ ;
wire _71_ ;
wire _620_ ;
wire _200_ ;
wire _714_ ;
wire _523_ ;
wire _103_ ;
wire [4:4] _752_ ;
wire _332_ ;
wire _68_ ;
wire _561_ ;
wire _141_ ;
wire _617_ ;
wire _370_ ;
wire _426_ ;
wire _655_ ;
wire _235_ ;
wire _464_ ;
wire _693_ ;
wire _273_ ;
wire [1:1] _749_ ;
wire _329_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _367_ ;
wire _596_ ;
wire _176_ ;
wire _499_ ;
wire _711_ ;
wire _27_ ;
wire _520_ ;
wire _100_ ;
wire _65_ ;
wire _614_ ;
wire _423_ ;
wire _652_ ;
wire _232_ ;
wire _708_ ;
wire _461_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _746_ ;
wire _326_ ;
wire _555_ ;
wire _135_ ;
wire _364_ ;
wire _593_ ;
wire _173_ ;
wire _649_ ;
wire _229_ ;
wire _458_ ;
wire _687_ ;
wire _267_ ;
wire _496_ ;
wire _24_ ;
wire _62_ ;
wire _399_ ;
wire _611_ ;
wire _420_ ;
wire _705_ ;
wire _514_ ;
wire _743_ ;
wire _323_ ;
wire _59_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _361_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _646_ ;
wire _226_ ;
wire _455_ ;
wire _684_ ;
wire _264_ ;
wire _493_ ;
wire _549_ ;
wire _129_ ;
wire _21_ ;
wire _358_ ;
wire _587_ ;
wire _167_ ;
wire _396_ ;
wire _702_ ;
wire _299_ ;
wire _18_ ;
wire _511_ ;
wire _740_ ;
wire _320_ ;
wire _56_ ;
wire _605_ ;
wire _414_ ;
wire _94_ ;
wire _643_ ;
wire _223_ ;
wire _452_ ;
wire _508_ ;
wire _681_ ;
wire _261_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _546_ ;
wire _126_ ;
wire _355_ ;
wire _584_ ;
wire _164_ ;
wire _393_ ;
wire _449_ ;
wire _678_ ;
wire _258_ ;
wire _487_ ;
wire _296_ ;
wire _15_ ;
wire _53_ ;
wire _602_ ;
wire _199_ ;
wire _411_ ;
wire _91_ ;
wire _640_ ;
wire _220_ ;
wire _9_ ;
wire _505_ ;
wire _734_ ;
wire _314_ ;
wire _543_ ;
wire _123_ ;
wire _352_ ;
wire _408_ ;
wire _88_ ;
wire _581_ ;
wire _161_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _446_ ;
wire [15:0] Yin ;
wire _675_ ;
wire _255_ ;
wire _484_ ;
wire _293_ ;
wire _12_ ;
wire _349_ ;
wire _578_ ;
wire _158_ ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire _6_ ;
wire _502_ ;
wire _731_ ;
wire _311_ ;
wire _47_ ;
wire _540_ ;
wire _120_ ;
wire _405_ ;
wire _85_ ;
wire _634_ ;
wire _214_ ;
wire _443_ ;
wire _672_ ;
wire _252_ ;
wire _728_ ;
wire _308_ ;
wire _481_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _346_ ;
wire _575_ ;
wire _155_ ;
wire _384_ ;
wire _193_ ;
wire _669_ ;
wire _249_ ;
wire _478_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _402_ ;
wire _82_ ;
wire _631_ ;
wire _211_ ;
wire _440_ ;
wire _725_ ;
wire _305_ ;
wire _534_ ;
wire _114_ ;
wire _343_ ;
wire _79_ ;
wire _572_ ;
wire _152_ ;
wire _628_ ;
wire _208_ ;
wire _381_ ;
wire _437_ ;
wire _190_ ;
wire _666_ ;
wire _246_ ;
wire _475_ ;
wire _284_ ;
wire _0_ ;
wire _569_ ;
wire _149_ ;
wire _41_ ;
wire _378_ ;
wire _187_ ;
wire [15:0] Yout ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _531_ ;
wire _111_ ;
wire _340_ ;
wire _76_ ;
wire _625_ ;
wire _205_ ;
wire _434_ ;
wire _663_ ;
wire _243_ ;
wire _719_ ;
wire _472_ ;
wire _528_ ;
wire _108_ ;
wire _281_ ;
wire _337_ ;
wire _566_ ;
wire _146_ ;
wire _375_ ;
wire _184_ ;
wire _469_ ;
wire _698_ ;
wire _278_ ;
wire _35_ ;
wire [7:0] Xout ;
wire _73_ ;
wire _622_ ;
wire _202_ ;
wire _431_ ;
wire _660_ ;
wire _240_ ;
wire _716_ ;
wire _525_ ;
wire _105_ ;
wire [7:0] _754_ ;
wire _334_ ;
wire _563_ ;
wire _143_ ;
wire _619_ ;
wire _372_ ;
wire _428_ ;
wire _181_ ;
wire _657_ ;
wire _237_ ;
wire _466_ ;
wire _695_ ;
wire _275_ ;
wire _32_ ;
wire _369_ ;
wire _598_ ;
wire _178_ ;
wire _70_ ;
wire _713_ ;
wire _29_ ;
wire _522_ ;
wire _102_ ;
wire [3:3] _751_ ;
wire _331_ ;
wire _67_ ;
wire _560_ ;
wire _140_ ;
wire _616_ ;
wire _425_ ;
wire _654_ ;
wire _234_ ;
wire _463_ ;
wire _519_ ;
wire _692_ ;
wire _272_ ;
wire [0:0] _748_ ;
wire _328_ ;
wire _557_ ;
wire _137_ ;
wire _366_ ;
wire _595_ ;
wire _175_ ;
wire _689_ ;
wire _269_ ;
wire _498_ ;
wire _710_ ;
wire _26_ ;
wire Cin_0_bF$buf0 ;
wire Cin_0_bF$buf1 ;
wire Cin_0_bF$buf2 ;
wire Cin_0_bF$buf3 ;
wire _64_ ;
wire _613_ ;
wire _422_ ;
wire _651_ ;
wire _231_ ;
wire _707_ ;
wire _460_ ;
wire _516_ ;
wire _745_ ;
wire _325_ ;
wire _554_ ;
wire _134_ ;
wire _363_ ;
wire _419_ ;
wire _99_ ;
wire _592_ ;
wire _172_ ;
wire _648_ ;
wire _228_ ;
wire _457_ ;
wire _686_ ;
wire _266_ ;
wire _495_ ;
wire _23_ ;
wire _589_ ;
wire _169_ ;
wire _61_ ;
wire _398_ ;
wire _610_ ;
wire _704_ ;
wire _513_ ;
wire _742_ ;
wire _322_ ;
wire _58_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _360_ ;
wire _416_ ;
wire _96_ ;
wire [7:0] Cin ;
wire _645_ ;
wire _225_ ;
wire _454_ ;
wire _683_ ;
wire _263_ ;
wire _739_ ;
wire _319_ ;
wire _492_ ;
wire _548_ ;
wire _128_ ;
wire _20_ ;
wire _357_ ;
wire _586_ ;
wire _166_ ;
wire _395_ ;
wire _489_ ;
wire _701_ ;
wire _298_ ;
wire _17_ ;
wire _510_ ;
wire _55_ ;
wire _604_ ;
wire _413_ ;
wire _93_ ;
wire _642_ ;
wire _222_ ;
wire _451_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _736_ ;
wire _316_ ;
wire _545_ ;
wire _125_ ;
wire _354_ ;
wire _583_ ;
wire _163_ ;
wire _639_ ;
wire _219_ ;
wire _392_ ;
wire _448_ ;
wire _677_ ;
wire _257_ ;
wire _486_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _601_ ;
wire _198_ ;
wire _410_ ;
wire _90_ ;
wire _8_ ;
wire _504_ ;
wire _733_ ;
wire _313_ ;
wire _49_ ;
wire _542_ ;
wire _122_ ;
wire _351_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _636_ ;
wire _216_ ;
wire _445_ ;
wire _674_ ;
wire _254_ ;
wire _483_ ;
wire _539_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _348_ ;
wire _577_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire _289_ ;
wire _5_ ;
wire _501_ ;
wire _730_ ;
wire _310_ ;
wire _46_ ;
wire _404_ ;
wire _84_ ;
wire _633_ ;
wire _213_ ;
wire _442_ ;
wire _671_ ;
wire _251_ ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire _536_ ;
wire _116_ ;
wire _345_ ;
wire _574_ ;
wire _154_ ;
wire _383_ ;
wire _439_ ;
wire _192_ ;
wire _668_ ;
wire _248_ ;
wire _477_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire _189_ ;
wire _401_ ;
wire _81_ ;
wire _630_ ;
wire _210_ ;
wire _724_ ;
wire _304_ ;
wire _533_ ;
wire _113_ ;
wire _342_ ;
wire _78_ ;
wire _571_ ;
wire _151_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _436_ ;
wire [7:0] Xin ;
wire _665_ ;
wire _245_ ;
wire _474_ ;
wire _283_ ;
wire _339_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire _377_ ;
wire _186_ ;
wire _721_ ;
wire _301_ ;
wire _37_ ;
wire _530_ ;
wire _110_ ;
wire _75_ ;
wire _624_ ;
wire _204_ ;
wire _433_ ;
wire _662_ ;
wire _242_ ;
wire _718_ ;
wire _471_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _336_ ;
wire _565_ ;
wire _145_ ;
wire _374_ ;
wire _183_ ;
wire _659_ ;
wire _239_ ;
wire _468_ ;
wire _697_ ;
wire _277_ ;
wire _34_ ;
wire _72_ ;
wire _621_ ;
wire _201_ ;
wire _430_ ;
wire _715_ ;
wire _524_ ;
wire _104_ ;
wire [15:5] _753_ ;
wire _333_ ;
wire _69_ ;
wire _562_ ;
wire _142_ ;
wire _618_ ;
wire _371_ ;
wire _427_ ;
wire _180_ ;
wire _656_ ;
wire _236_ ;
wire _465_ ;
wire _694_ ;
wire _274_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _368_ ;
wire _597_ ;
wire _177_ ;
wire _712_ ;
wire _28_ ;
wire _521_ ;
wire _101_ ;
wire [2:2] _750_ ;
wire _330_ ;
wire _66_ ;
wire _615_ ;
wire _424_ ;
wire _653_ ;
wire _233_ ;
wire _709_ ;
wire _462_ ;
wire _518_ ;
wire _691_ ;
wire _271_ ;
wire _747_ ;
wire _327_ ;
wire _556_ ;
wire _136_ ;
wire _365_ ;
wire _594_ ;
wire _174_ ;
wire _459_ ;
wire _688_ ;
wire _268_ ;
wire _497_ ;
wire Xin_3_bF$buf0 ;
wire Xin_3_bF$buf1 ;
wire Xin_3_bF$buf2 ;
wire Xin_3_bF$buf3 ;
wire _25_ ;
wire _63_ ;
wire _612_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire _706_ ;
wire _515_ ;
wire _744_ ;
wire _324_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _362_ ;
wire _418_ ;
wire _98_ ;
wire _591_ ;
wire _171_ ;
wire _647_ ;
wire _227_ ;
wire _456_ ;
wire _685_ ;
wire _265_ ;
wire _494_ ;
wire _22_ ;
wire _359_ ;

FILL FILL_0__1241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1259_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1328_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_740_),
    .B(_352_),
    .C(_445_),
    .Y(_451_)
);

FILL FILL_3__1081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__941_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[1]),
    .B(Cin[2]),
    .Y(_741_)
);

FILL FILL_1__1211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1137_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_668_),
    .B(_670_),
    .C(_694_),
    .Y(_696_)
);

OAI21X1 _1066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_740_),
    .B(_151_),
    .C(_250_),
    .Y(_256_)
);

FILL FILL_1__848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1366_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_489_),
    .Y(_491_)
);

FILL FILL_0__1335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1114_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_574_),
    .B(_587_),
    .C(_592_),
    .Y(_593_)
);

FILL FILL_0__1429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1182_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_119_),
    .B(_118_),
    .C(_82_),
    .Y(_124_)
);

FILL FILL_1__1343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1269_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_281_),
    .Y(_388_)
);

FILL FILL_2__1412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89250x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_611_),
    .B(_608_),
    .Y(_616_)
);

FILL FILL_3__882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88950x19650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1208_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[1]),
    .B(Xin_5_bF$buf0),
    .Y(_161_)
);

FILL FILL_1__1381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1085_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_686_),
    .B(_701_),
    .C(_712_),
    .Y(_715_)
);

FILL FILL_0__832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__976_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_18_),
    .B(_16_),
    .C(_9_),
    .Y(_27_)
);

FILL FILL_1__1246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1315_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_506_),
    .Y(_511_)
);

FILL FILL_3__785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__899_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1542_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(y[14]),
    .CLK(clk_bF$buf2),
    .Q(_755_[14])
);

OAI22X1 _1122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_309_),
    .B(_310_),
    .C(_308_),
    .D(_208_),
    .Y(_311_)
);

FILL FILL_0__870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__904_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_57_),
    .B(_58_),
    .C(_55_),
    .Y(_65_)
);

FILL FILL_1__1284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1002_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_81_),
    .B(_116_),
    .C(_120_),
    .Y(_121_)
);

NAND3X1 _1351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_551_),
    .B(_552_),
    .C(_550_),
    .Y(_553_)
);

FILL FILL89550x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1162_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_604_),
    .B(_607_),
    .C(_611_),
    .Y(_613_)
);

FILL FILL_3__879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1149_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_755_[6]),
    .Y(Yout[6])
);

INVX1 _1160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_348_),
    .Y(_349_)
);

FILL FILL_1__942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1391_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_404_),
    .B(_405_),
    .C(_403_),
    .Y(_406_)
);

FILL FILL_0__964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1040_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_154_),
    .B(_157_),
    .Y(_158_)
);

FILL FILL_1__1378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1516_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_650_),
    .B(_651_),
    .Y(_653_)
);

INVX1 _1025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_214_),
    .Y(_215_)
);

FILL FILL_0__773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__807_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_397_),
    .B(_590_),
    .Y(_601_)
);

FILL FILL_1__1187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1325_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _1254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_590_),
    .B(_447_),
    .C(_740_),
    .D(_352_),
    .Y(_448_)
);

FILL FILL_2__823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1134_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_693_),
    .B(_674_),
    .Y(_694_)
);

OAI21X1 _1063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_740_),
    .B(_151_),
    .C(_252_),
    .Y(_253_)
);

FILL FILL_1__845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1294_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1539_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(y[11]),
    .CLK(clk_bF$buf5),
    .Q(_755_[11])
);

XNOR2X1 _1119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_211_),
    .B(_308_),
    .Y(_753_[7])
);

FILL FILL_0__867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1363_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_),
    .B(_488_),
    .C(_486_),
    .Y(_489_)
);

FILL FILL_0__1332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1419_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_439_),
    .B(_463_),
    .C(_466_),
    .Y(_550_)
);

FILL FILL_3__1172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89250x39150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1228_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_755_[3]),
    .Y(Yout[3])
);

AOI21X1 _1157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_270_),
    .B(_267_),
    .C(_260_),
    .Y(_346_)
);

FILL FILL_1__939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1037_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_585_),
    .B(_579_),
    .C(_583_),
    .Y(_589_)
);

FILL FILL_4__1106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1266_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_368_),
    .B(_373_),
    .C(_376_),
    .Y(_384_)
);

FILL FILL_1__977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89550x78150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1014_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_314_),
    .B(_395_),
    .C(_485_),
    .Y(_486_)
);

FILL FILL_2__1503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1082_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _1501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_702_),
    .B(_712_),
    .Y(_713_)
);

FILL FILL_3__973_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_22_),
    .B(_21_),
    .C(_735_),
    .Y(_25_)
);

FILL FILL_1__1243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__760_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_240_),
    .B(_243_),
    .Y(_288_)
);

FILL FILL_2__1312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1138_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_502_),
    .Y(_508_)
);

FILL FILL_3__782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__901_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_57_),
    .B(_58_),
    .C(_61_),
    .Y(_62_)
);

FILL FILL_1__1281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89250x27450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__923_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_113_),
    .B(_114_),
    .C(_112_),
    .Y(_118_)
);

FILL FILL_1__1337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1406_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_573_),
    .B(_608_),
    .Y(_609_)
);

FILL FILL_3__876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1215_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_403_),
    .B(_398_),
    .Y(_404_)
);

FILL FILL_0__961_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_590_),
    .B(_151_),
    .C(_85_),
    .Y(_155_)
);

FILL FILL_1__1375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89550x66450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1513_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[12]),
    .Y(_650_)
);

AOI21X1 _1022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_195_),
    .B(_196_),
    .C(_139_),
    .Y(_212_)
);

FILL FILL_0__770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__804_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_515_),
    .B(_537_),
    .C(_429_),
    .Y(_569_)
);

FILL FILL_1__1184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1322_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_19_),
    .B(_14_),
    .C(_738_),
    .Y(_22_)
);

AND2X2 _1251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[2]),
    .B(Xin[7]),
    .Y(_445_)
);

FILL FILL_2__1309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1062_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_417_),
    .B(_503_),
    .Y(_505_)
);

FILL FILL_3__779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1049_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_689_),
    .B(_690_),
    .Y(_691_)
);

AND2X2 _1060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[2]),
    .B(Xin_5_bF$buf1),
    .Y(_250_)
);

FILL FILL_1__842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1291_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1536_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(y[8]),
    .CLK(clk_bF$buf1),
    .Q(_755_[8])
);

AOI21X1 _1116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297_),
    .B(_292_),
    .C(_215_),
    .Y(_306_)
);

FILL FILL_0__864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1360_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_48_),
    .B(_50_),
    .C(_46_),
    .Y(_59_)
);

FILL FILL_1__1278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1416_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_543_),
    .B(_545_),
    .Y(_546_)
);

FILL FILL_1__1087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1225_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_755_[14]),
    .Y(Yout[14])
);

OAI21X1 _1154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_335_),
    .B(_334_),
    .C(_332_),
    .Y(_343_)
);

FILL FILL_1__936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89250x15750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1034_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_583_),
    .B(_579_),
    .C(_585_),
    .Y(_586_)
);

FILL FILL_4__889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1194_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_646_),
    .Y(_647_)
);

AOI21X1 _1019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_203_),
    .B(_207_),
    .C(_136_),
    .Y(_210_)
);

FILL FILL_0__767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88950x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_380_),
    .B(_374_),
    .C(_345_),
    .Y(_381_)
);

FILL FILL_1__974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1319_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_359_),
    .B(_441_),
    .C(_369_),
    .Y(_442_)
);

FILL FILL_0__996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1072_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_176_),
    .B(_179_),
    .C(_182_),
    .Y(_190_)
);

FILL FILL_1__783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89550x54750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1128_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_686_),
    .B(_685_),
    .C(_646_),
    .Y(_688_)
);

NAND2X1 _1057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin_3_bF$buf1),
    .B(Cin[4]),
    .Y(_247_)
);

FILL FILL_1__839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1357_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_479_),
    .B(_480_),
    .C(_481_),
    .Y(_482_)
);

FILL FILL_2__1500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1166_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254_),
    .B(_257_),
    .C(_275_),
    .D(_271_),
    .Y(_285_)
);

FILL FILL_1__877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__920_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_112_),
    .B(_114_),
    .C(_113_),
    .Y(_115_)
);

FILL FILL_1__1334_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_369_),
    .B(_372_),
    .C(_377_),
    .Y(_378_)
);

FILL FILL_2__1403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__758_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_592_),
    .B(_587_),
    .C(_574_),
    .Y(_606_)
);

FILL FILL_3__873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__929_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_314_),
    .B(_394_),
    .C(_395_),
    .Y(_401_)
);

NAND2X1 _961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin_3_bF$buf2),
    .B(Cin[3]),
    .Y(_152_)
);

FILL FILL_1__1372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__801_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_493_),
    .B(_526_),
    .C(_461_),
    .Y(_537_)
);

FILL FILL_1__1181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_18_),
    .B(_17_),
    .C(_16_),
    .Y(_19_)
);

FILL FILL_1__1237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1306_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_415_),
    .B(_416_),
    .C(_424_),
    .Y(_501_)
);

FILL FILL_3__776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1115_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1533_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(y[5]),
    .CLK(clk_bF$buf3),
    .Q(_755_[5])
);

INVX1 _1113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_200_),
    .Y(_303_)
);

FILL FILL_0__861_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_38_),
    .B(_55_),
    .C(_43_),
    .Y(_56_)
);

FILL FILL_1__1275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1413_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_539_),
    .B(_530_),
    .Y(_543_)
);

FILL FILL_4__848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_755_[11]),
    .Y(Yout[11])
);

NAND3X1 _1151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_318_),
    .B(_333_),
    .C(_339_),
    .Y(_340_)
);

FILL FILL_1__933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89550x19650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1382_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_396_),
    .B(_393_),
    .C(_313_),
    .Y(_398_)
);

FILL FILL_0__955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1031_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[2]),
    .B(Xin[4]),
    .Y(_149_)
);

FILL FILL_1__1369_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_582_),
    .Y(_583_)
);

FILL FILL_2__1438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1507_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin_5_bF$buf3),
    .B(Cin[7]),
    .Y(_643_)
);

NAND3X1 _1016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_204_),
    .B(_205_),
    .C(_206_),
    .Y(_207_)
);

FILL FILL_0__764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1260_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_493_),
    .Y(_504_)
);

FILL FILL_1__1178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1316_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_435_),
    .B(_436_),
    .C(_437_),
    .Y(_438_)
);

FILL FILL_0__993_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_186_),
    .B(_180_),
    .C(_144_),
    .Y(_187_)
);

FILL FILL_1__780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1125_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_652_),
    .B(_657_),
    .C(_683_),
    .Y(_684_)
);

AND2X2 _1054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_240_),
    .B(_243_),
    .Y(_244_)
);

FILL FILL_1__836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1354_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_410_),
    .Y(_479_)
);

FILL FILL_0__1323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1094_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_530_),
    .B(_539_),
    .Y(_540_)
);

FILL FILL_3__1583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1163_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_177_),
    .Y(_282_)
);

FILL FILL_1__874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1219_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_755_[0]),
    .Y(Yout[0])
);

INVX1 _1148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_336_),
    .Y(_337_)
);

FILL FILL_0__896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1392_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[2]),
    .B(Xin_3_bF$buf2),
    .Y(_91_)
);

FILL FILL_4__1041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1028_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_503_),
    .B(_576_),
    .C(_579_),
    .Y(_580_)
);

FILL FILL_0__1417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1188_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_89_),
    .Y(_112_)
);

FILL FILL_1__1331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1257_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_271_),
    .Y(_375_)
);

FILL FILL_1__968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__964_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_15_),
    .B(_732_),
    .C(_742_),
    .Y(_16_)
);

FILL FILL_1__1234_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_267_),
    .B(_270_),
    .C(_272_),
    .Y(_279_)
);

FILL FILL_2__1303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1129_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_428_),
    .B(_434_),
    .Y(_498_)
);

FILL FILL_3__773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1519_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1530_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(y[2]),
    .CLK(clk_bF$buf1),
    .Q(_755_[2])
);

NAND3X1 _1110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_287_),
    .B(_291_),
    .C(_294_),
    .Y(_300_)
);

OAI21X1 _861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_47_),
    .B(_590_),
    .C(_743_),
    .Y(_53_)
);

FILL FILL_1__1272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1410_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_101_),
    .B(_98_),
    .C(_97_),
    .Y(_109_)
);

FILL FILL_1__1328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1206_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_391_),
    .B(_317_),
    .C(_390_),
    .Y(_394_)
);

FILL FILL_0__952_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_112_),
    .B(_145_),
    .C(_106_),
    .Y(_146_)
);

FILL FILL_1__1366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1504_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_77_),
    .B(_447_),
    .C(_576_),
    .Y(_640_)
);

INVX1 _1013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_127_),
    .Y(_204_)
);

FILL FILL_0__761_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_461_),
    .Y(_472_)
);

FILL FILL_1__1175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1313_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_327_),
    .B(_323_),
    .Y(_435_)
);

FILL FILL_0__990_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_177_),
    .B(_178_),
    .C(_183_),
    .Y(_184_)
);

FILL FILL_2__811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1122_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_679_),
    .B(_680_),
    .Y(_681_)
);

NAND3X1 _1051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_226_),
    .B(_230_),
    .C(_238_),
    .Y(_241_)
);

FILL FILL_1__833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1282_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1527_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(Xin[7]),
    .CLK(clk_bF$buf2),
    .Q(_754_[7])
);

OAI21X1 _1107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_295_),
    .B(_296_),
    .C(_294_),
    .Y(_297_)
);

FILL FILL_0__855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1351_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_44_),
    .Y(_50_)
);

FILL FILL_1__1269_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_434_),
    .B(_438_),
    .C(_463_),
    .D(_458_),
    .Y(_476_)
);

FILL FILL_4__1000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1407_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_350_),
    .B(_532_),
    .Y(_536_)
);

FILL FILL_3__1580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88050x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_754_[5]),
    .Y(Xout[5])
);

AOI21X1 _1145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_328_),
    .B(_329_),
    .C(_319_),
    .Y(_334_)
);

FILL FILL_0__893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__927_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_590_),
    .B(_87_),
    .C(_79_),
    .Y(_88_)
);

FILL FILL_2__1376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1025_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin_5_bF$buf3),
    .Y(_577_)
);

FILL FILL_0__1414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1254_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_263_),
    .B(_267_),
    .C(_371_),
    .Y(_372_)
);

FILL FILL_1__965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1223_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_250_),
    .B(_350_),
    .C(_353_),
    .D(_349_),
    .Y(_432_)
);

FILL FILL88350x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1119_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_447_),
    .B(_575_),
    .Y(_678_)
);

AOI21X1 _1048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148_),
    .B(_153_),
    .C(_237_),
    .Y(_238_)
);

FILL FILL_0__796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1292_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[3]),
    .Y(_740_)
);

FILL FILL_0__1508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1348_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_442_),
    .B(_462_),
    .Y(_473_)
);

FILL FILL_0__1317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__961_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_12_),
    .B(_11_),
    .C(_10_),
    .Y(_13_)
);

FILL FILL_1__1231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1157_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_271_),
    .B(_275_),
    .C(_258_),
    .Y(_276_)
);

FILL FILL_1__868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__911_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_95_),
    .B(_102_),
    .C(_105_),
    .Y(_106_)
);

FILL FILL_1__1325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88950x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__978_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_345_),
    .B(_374_),
    .C(_380_),
    .Y(_391_)
);

OAI21X1 _952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_79_),
    .B(_91_),
    .C(_89_),
    .Y(_143_)
);

FILL FILL_1__1363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88350x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1419_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_604_),
    .B(_600_),
    .Y(_637_)
);

OAI21X1 _1010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_187_),
    .B(_191_),
    .C(_194_),
    .Y(_201_)
);

NOR2X1 _761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[0]),
    .B(_407_),
    .Y(_440_)
);

FILL FILL_1__1172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1310_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_746_),
    .Y(_10_)
);

FILL FILL_1__1228_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_106_),
    .Y(_181_)
);

FILL FILL_2__1470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1106_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1524_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(Xin[4]),
    .CLK(clk_bF$buf1),
    .Q(_754_[4])
);

AOI21X1 _1104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_188_),
    .B(_190_),
    .C(_293_),
    .Y(_294_)
);

FILL FILL_0__852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__996_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[2]),
    .Y(_47_)
);

FILL FILL_1__1266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1404_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_350_),
    .B(_532_),
    .C(_531_),
    .Y(_533_)
);

FILL FILL_1__1495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1213_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_754_[2]),
    .Y(Xout[2])
);

AOI22X1 _1142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[2]),
    .B(Xin_5_bF$buf2),
    .C(Cin[3]),
    .D(Xin[4]),
    .Y(_331_)
);

FILL FILL_0__890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__924_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin_3_bF$buf1),
    .B(Cin[3]),
    .Y(_85_)
);

FILL FILL_2__1373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1022_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[1]),
    .B(Cin[6]),
    .Y(_140_)
);

OAI21X1 _1371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_502_),
    .B(_506_),
    .C(_510_),
    .Y(_574_)
);

FILL FILL_4__1511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1182_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_630_),
    .B(_632_),
    .C(_628_),
    .Y(_634_)
);

AOI21X1 _1007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_197_),
    .B(_192_),
    .C(_137_),
    .Y(_198_)
);

FILL FILL_3__899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1251_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_386_),
    .B(_397_),
    .Y(_407_)
);

FILL FILL_1__1169_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_361_),
    .B(_366_),
    .Y(_369_)
);

FILL FILL_1__962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88650x78150 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_425_),
    .B(_420_),
    .C(_427_),
    .Y(_428_)
);

FILL FILL_0__984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1060_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_170_),
    .B(_166_),
    .C(_172_),
    .Y(_178_)
);

FILL FILL_1__1398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_635_),
    .B(_660_),
    .C(_662_),
    .Y(_674_)
);

AOI21X1 _1045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_228_),
    .B(_229_),
    .C(_220_),
    .Y(_235_)
);

FILL FILL_0__793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__827_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_737_),
    .B(_736_),
    .Y(_750_[2])
);

FILL FILL_0__1505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1345_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_412_),
    .B(_464_),
    .C(_468_),
    .Y(_469_)
);

FILL FILL_4__1414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1154_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_269_),
    .B(_268_),
    .C(_261_),
    .Y(_273_)
);

FILL FILL_1__865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88950x31350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__801_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1559_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_753_[15]),
    .CLK(clk_bF$buf2),
    .Q(y[15])
);

OAI21X1 _1139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_87_),
    .B(_77_),
    .C(_321_),
    .Y(_328_)
);

FILL FILL_0__887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1019_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_570_),
    .Y(_571_)
);

FILL FILL_3__1192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1161_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[5]),
    .B(_100_),
    .Y(_103_)
);

FILL FILL_1__1322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1248_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_364_),
    .B(_363_),
    .Y(_366_)
);

FILL FILL_1__959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__955_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf1),
    .B(Xin_3_bF$buf0),
    .C(_2_),
    .Y(_7_)
);

FILL FILL_1__1225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__878_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1521_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(Xin[1]),
    .CLK(clk_bF$buf1),
    .Q(_754_[1])
);

NAND3X1 _1101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_288_),
    .B(_289_),
    .C(_290_),
    .Y(_291_)
);

FILL FILL_3__993_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[0]),
    .B(Cin[4]),
    .Y(_44_)
);

FILL FILL_1__1263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1401_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf3),
    .B(Xin_5_bF$buf0),
    .Y(_100_)
);

FILL FILL_1__1319_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_529_),
    .B(_454_),
    .Y(_530_)
);

FILL FILL_1__1492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__921_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_61_),
    .B(_58_),
    .C(_38_),
    .Y(_82_)
);

FILL FILL_2__1370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88350x15750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__943_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_78_),
    .B(_80_),
    .Y(_137_)
);

FILL FILL_1__1357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1006_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_626_),
    .B(_629_),
    .C(_492_),
    .Y(_630_)
);

NAND3X1 _1004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_188_),
    .B(_189_),
    .C(_190_),
    .Y(_195_)
);

FILL FILL_3__896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1304_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_421_),
    .B(_422_),
    .C(_424_),
    .Y(_425_)
);

FILL FILL_0__981_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_173_),
    .B(_174_),
    .C(_172_),
    .Y(_175_)
);

FILL FILL_1__1395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88650x54750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1113_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _1462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_634_),
    .B(_671_),
    .Y(_753_[12])
);

AND2X2 _1042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_152_),
    .B(_231_),
    .Y(_232_)
);

FILL FILL_0__790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__824_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_559_),
    .B(_734_),
    .C(_731_),
    .Y(_735_)
);

FILL FILL_0__1502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1099_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_739_),
    .B(_20_),
    .C(_24_),
    .Y(_730_)
);

FILL FILL_0__846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1342_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_31_),
    .B(_36_),
    .C(_34_),
    .Y(_41_)
);

NOR2X1 _1271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_460_),
    .B(_462_),
    .Y(_466_)
);

FILL FILL_0__1311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1082_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_523_),
    .B(_524_),
    .C(_525_),
    .Y(_527_)
);

FILL FILL_3__799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1069_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_261_),
    .B(_268_),
    .C(_269_),
    .Y(_270_)
);

FILL FILL_1__862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1207_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1556_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_753_[12]),
    .CLK(clk_bF$buf2),
    .Q(y[12])
);

NAND2X1 _1136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin_3_bF$buf3),
    .B(Cin[5]),
    .Y(_325_)
);

FILL FILL_0__884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1380_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[2]),
    .B(Cin[3]),
    .Y(_79_)
);

FILL FILL_1__1298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1016_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_555_),
    .Y(_567_)
);

FILL FILL_0__1405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1245_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_362_),
    .Y(_363_)
);

FILL FILL_1__956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__914_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_611_),
    .B(_608_),
    .C(_621_),
    .Y(_669_)
);

NAND2X1 _1039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_224_),
    .B(_222_),
    .Y(_229_)
);

FILL FILL_0__787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__930_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_460_),
    .B(_462_),
    .Y(_463_)
);

FILL FILL_3__1092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__952_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_),
    .B(_3_),
    .Y(_4_)
);

FILL FILL_1__1222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1148_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_675_),
    .B(_681_),
    .Y(_709_)
);

NAND3X1 _1077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_263_),
    .B(_262_),
    .C(_266_),
    .Y(_267_)
);

FILL FILL_1__859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__902_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_96_),
    .Y(_97_)
);

FILL FILL_1__1316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88650x19650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__940_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_132_),
    .B(_134_),
    .Y(_135_)
);

FILL FILL_1__1354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__778_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_625_),
    .B(_565_),
    .Y(_627_)
);

OAI21X1 _1001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_191_),
    .B(_187_),
    .C(_139_),
    .Y(_192_)
);

FILL FILL_3__893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1301_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf2),
    .B(Xin_3_bF$buf0),
    .C(Yin[3]),
    .Y(_1_)
);

FILL FILL_1__1219_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_416_),
    .Y(_422_)
);

INVX1 _981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_160_),
    .Y(_172_)
);

FILL FILL_1__1392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88950x58650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__821_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_601_),
    .Y(_732_)
);

FILL FILL_2__1517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1096_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_721_),
    .Y(_727_)
);

FILL FILL_0__843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__987_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_29_),
    .B(_35_),
    .C(_37_),
    .Y(_38_)
);

FILL FILL_1__1257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1326_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_501_),
    .Y(_523_)
);

FILL FILL_3__796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1204_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1553_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_753_[9]),
    .CLK(clk_bF$buf5),
    .Q(y[9])
);

AND2X2 _1133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin_3_bF$buf3),
    .B(Cin[5]),
    .Y(_322_)
);

FILL FILL_0__881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__915_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_744_),
    .B(_70_),
    .C(_63_),
    .Y(_76_)
);

FILL FILL_1__1295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1013_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_564_),
    .B(_558_),
    .Y(_565_)
);

FILL FILL_4__1502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1173_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_624_),
    .B(_618_),
    .Y(_625_)
);

FILL FILL_3__1242_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf0),
    .B(Xin[7]),
    .C(Yin[7]),
    .Y(_360_)
);

FILL FILL_1__953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88350x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_325_),
    .B(_417_),
    .Y(_419_)
);

FILL FILL_0__975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1051_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_164_),
    .B(_162_),
    .Y(_169_)
);

FILL FILL_1__1389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1107_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_635_),
    .B(_660_),
    .C(_664_),
    .Y(_665_)
);

NAND3X1 _1036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_225_),
    .B(_221_),
    .C(_223_),
    .Y(_226_)
);

FILL FILL_0__784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89550x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1280_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_697_),
    .B(_676_),
    .C(_612_),
    .Y(_718_)
);

FILL FILL_1__1198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1336_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_263_),
    .B(_267_),
    .C(_371_),
    .Y(_459_)
);

FILL FILL_4__1405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1145_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_678_),
    .Y(_705_)
);

INVX1 _1074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[7]),
    .Y(_264_)
);

FILL FILL_1__856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1374_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[0]),
    .Y(Cin_0_bF$buf3)
);

BUFX2 BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[0]),
    .Y(Cin_0_bF$buf2)
);

BUFX2 BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[0]),
    .Y(Cin_0_bF$buf1)
);

BUFX2 BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[0]),
    .Y(Cin_0_bF$buf0)
);

FILL FILL_4__1023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1504_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_555_),
    .B(_498_),
    .C(_556_),
    .Y(_562_)
);

FILL FILL_3__1183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1152_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_89_),
    .B(_93_),
    .Y(_94_)
);

FILL FILL_1__1313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1239_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[2]),
    .B(Xin[6]),
    .C(_336_),
    .Y(_357_)
);

FILL FILL_0__1208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89250x78150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1048_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_599_),
    .B(_600_),
    .Y(_602_)
);

FILL FILL_1__759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1190_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_127_),
    .B(_131_),
    .C(_75_),
    .Y(_132_)
);

FILL FILL_1__1351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__946_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_623_),
    .B(_655_),
    .C(_644_),
    .Y(_746_)
);

FILL FILL_1__1216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89550x31350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1093_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_723_),
    .B(_628_),
    .C(_696_),
    .Y(_724_)
);

FILL FILL_0__840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__984_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_30_),
    .B(_34_),
    .C(_32_),
    .Y(_35_)
);

FILL FILL_1__1254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1149_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_444_),
    .B(_448_),
    .C(_519_),
    .Y(_520_)
);

FILL FILL_3__793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1119_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1550_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_753_[6]),
    .CLK(clk_bF$buf0),
    .Q(y[6])
);

NAND2X1 _1130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[1]),
    .B(Cin[7]),
    .Y(_319_)
);

FILL FILL_1__912_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_72_),
    .B(_23_),
    .Y(_73_)
);

FILL FILL_1__1292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1010_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_124_),
    .B(_125_),
    .C(_123_),
    .Y(_129_)
);

FILL FILL_1__1348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1170_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_570_),
    .B(_615_),
    .C(_616_),
    .Y(_621_)
);

FILL FILL_3__887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1226_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[2]),
    .B(Cin[7]),
    .Y(_415_)
);

FILL FILL_0__972_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_165_),
    .B(_163_),
    .C(_161_),
    .Y(_166_)
);

FILL FILL_1__1386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1104_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_637_),
    .B(_659_),
    .Y(_662_)
);

NAND2X1 _1033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_140_),
    .B(_222_),
    .Y(_223_)
);

FILL FILL_0__781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__815_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_644_),
    .Y(_687_)
);

FILL FILL_1__1195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1264_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_717_),
    .B(_720_),
    .Y(_721_)
);

FILL FILL_0__837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1333_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_453_),
    .Y(_456_)
);

FILL FILL_0__1302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1073_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_510_),
    .B(_511_),
    .C(_508_),
    .Y(_517_)
);

FILL FILL_3__1562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1142_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_686_),
    .B(_701_),
    .Y(_702_)
);

NAND2X1 _1071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[1]),
    .B(Xin[6]),
    .Y(_261_)
);

FILL FILL_1__853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1129_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1547_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_751_[3]),
    .CLK(clk_bF$buf3),
    .Q(y[3])
);

AOI21X1 _1127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_276_),
    .B(_280_),
    .C(_246_),
    .Y(_316_)
);

FILL FILL_0__875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1371_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_62_),
    .B(_56_),
    .C(_27_),
    .Y(_70_)
);

FILL FILL_1__1289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1007_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_554_),
    .B(_557_),
    .C(_497_),
    .Y(_558_)
);

FILL FILL_3__1180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1236_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_353_),
    .B(_349_),
    .C(_351_),
    .Y(_354_)
);

FILL FILL_1__947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1045_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _1394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_532_),
    .B(Yin[11]),
    .Y(_598_)
);

FILL FILL_1__756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89250x54750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__921_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _1259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_362_),
    .B(Yin[9]),
    .Y(_453_)
);

FILL FILL_3__1083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__943_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[1]),
    .B(Cin[3]),
    .Y(_743_)
);

FILL FILL_1__1213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1139_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_674_),
    .B(_693_),
    .C(_670_),
    .Y(_699_)
);

AND2X2 _1068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_257_),
    .B(_254_),
    .Y(_258_)
);

FILL FILL_0__1108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1368_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_404_),
    .B(_490_),
    .Y(_494_)
);

FILL FILL_2__1511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__981_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_31_),
    .Y(_32_)
);

FILL FILL_1__1251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__931_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_123_),
    .B(_125_),
    .C(_124_),
    .Y(_126_)
);

FILL FILL_1__1345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__769_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_614_),
    .B(_617_),
    .C(_568_),
    .Y(_618_)
);

FILL FILL_3__884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89250x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__998_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_345_),
    .B(_411_),
    .C(_383_),
    .Y(_412_)
);

NAND2X1 _972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[6]),
    .B(_162_),
    .Y(_163_)
);

FILL FILL_1__1383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1019_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_658_),
    .B(_657_),
    .Y(_659_)
);

NAND2X1 _1030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[0]),
    .B(Cin[7]),
    .Y(_220_)
);

FILL FILL_1__812_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf1),
    .B(Xin[2]),
    .C(Yin[2]),
    .Y(_655_)
);

FILL FILL_1__1192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1087_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_703_),
    .B(_706_),
    .C(_711_),
    .Y(_717_)
);

FILL FILL_0__834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1330_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_747_),
    .B(_28_),
    .C(_1_),
    .Y(_29_)
);

FILL FILL_1__1248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1070_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_350_),
    .B(_445_),
    .Y(_513_)
);

FILL FILL_3__787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1126_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1544_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_748_[0]),
    .CLK(clk_bF$buf4),
    .Q(y[0])
);

AOI21X1 _1124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_215_),
    .B(_297_),
    .C(_312_),
    .Y(_313_)
);

FILL FILL_0__872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__906_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_65_),
    .B(_66_),
    .C(_64_),
    .Y(_67_)
);

FILL FILL_1__1286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89250x19650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1004_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_551_),
    .B(_552_),
    .C(_500_),
    .Y(_555_)
);

FILL FILL_1__1095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1164_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_604_),
    .B(_607_),
    .C(_573_),
    .Y(_615_)
);

FILL FILL_3__1233_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_755_[8]),
    .Y(Yout[8])
);

NAND2X1 _1162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_250_),
    .B(_350_),
    .Y(_351_)
);

FILL FILL_1__944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1393_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_315_),
    .B(_408_),
    .C(_394_),
    .Y(_409_)
);

FILL FILL_0__966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1042_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_96_),
    .B(_159_),
    .C(_98_),
    .Y(_160_)
);

NAND3X1 _1391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_588_),
    .B(_581_),
    .C(_586_),
    .Y(_595_)
);

FILL FILL_0__1431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89550x58650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1518_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_654_),
    .Y(_656_)
);

OAI21X1 _1027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_144_),
    .B(_216_),
    .C(_189_),
    .Y(_217_)
);

FILL FILL_0__775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1271_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[1]),
    .B(Cin[1]),
    .Y(_623_)
);

FILL FILL_1__1189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1327_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_590_),
    .B(_447_),
    .C(_350_),
    .Y(_450_)
);

FILL FILL_3__1080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1136_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_674_),
    .B(_693_),
    .Y(_695_)
);

NAND2X1 _1065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_252_),
    .B(_249_),
    .Y(_255_)
);

FILL FILL_1__847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1365_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _1294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_406_),
    .B(_490_),
    .Y(_753_[9])
);

FILL FILL_4__1014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_755_[5]),
    .Y(Yout[5])
);

FILL FILL_0_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[4]),
    .B(Cin[4]),
    .Y(_348_)
);

FILL FILL_0_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1039_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_591_),
    .B(_589_),
    .C(_588_),
    .Y(_592_)
);

FILL FILL_0__1428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1199_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_80_),
    .B(_122_),
    .Y(_123_)
);

FILL FILL_1__1342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1268_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_381_),
    .B(_385_),
    .C(_317_),
    .Y(_387_)
);

FILL FILL_1__979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89550x46950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1084_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_700_),
    .B(_714_),
    .Y(_753_[14])
);

FILL FILL_0__831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__975_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_744_),
    .Y(_26_)
);

FILL FILL_1__1245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1314_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_423_),
    .B(_509_),
    .Y(_510_)
);

FILL FILL_3__784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__898_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1541_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(y[13]),
    .CLK(clk_bF$buf5),
    .Q(_755_[13])
);

AND2X2 _1121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_302_),
    .B(_207_),
    .Y(_310_)
);

FILL FILL_1__903_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_745_),
    .B(_13_),
    .C(_17_),
    .Y(_64_)
);

FILL FILL_1__1283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1001_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_119_),
    .B(_118_),
    .C(_117_),
    .Y(_120_)
);

FILL FILL_1__1339_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_528_),
    .B(_540_),
    .Y(_552_)
);

FILL FILL_1__1092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1087_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_542_),
    .B(_546_),
    .C(_610_),
    .Y(_611_)
);

FILL FILL_3__878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1390_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_311_),
    .Y(_405_)
);

FILL FILL_0__963_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_147_),
    .B(_155_),
    .C(_156_),
    .Y(_157_)
);

FILL FILL_1__1377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1515_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_651_),
    .B(_650_),
    .Y(_652_)
);

NAND2X1 _1024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_142_),
    .B(_143_),
    .Y(_214_)
);

FILL FILL_0__772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__806_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[2]),
    .Y(_590_)
);

FILL FILL_1__1186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1324_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[7]),
    .Y(_447_)
);

FILL FILL_2__822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1064_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_506_),
    .B(_505_),
    .C(_502_),
    .Y(_507_)
);

FILL FILL_3__1133_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_692_),
    .B(_688_),
    .Y(_693_)
);

NAND2X1 _1062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[2]),
    .B(Xin_5_bF$buf2),
    .Y(_252_)
);

FILL FILL_1__844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1293_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1538_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(y[10]),
    .CLK(clk_bF$buf5),
    .Q(_755_[10])
);

NAND2X1 _1118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_302_),
    .B(_307_),
    .Y(_308_)
);

FILL FILL_0__866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1362_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_59_),
    .B(_60_),
    .Y(_61_)
);

AOI21X1 _1291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_477_),
    .B(_469_),
    .C(_410_),
    .Y(_488_)
);

FILL FILL_4__797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1418_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_541_),
    .B(_547_),
    .C(_500_),
    .Y(_549_)
);

FILL FILL_3__1171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1227_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_755_[2]),
    .Y(Yout[2])
);

NAND2X1 _1156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_340_),
    .B(_344_),
    .Y(_345_)
);

FILL FILL_1__938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88050x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1036_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_536_),
    .Y(_588_)
);

FILL FILL_0__1425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1265_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_379_),
    .B(_347_),
    .C(_378_),
    .Y(_383_)
);

FILL FILL_1__976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1204_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_683_),
    .Y(_690_)
);

AND2X2 _1059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[3]),
    .B(Xin[4]),
    .Y(_249_)
);

FILL FILL_0__1519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1359_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_394_),
    .Y(_485_)
);

FILL FILL_2__1502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1081_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _1500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_711_),
    .B(_707_),
    .Y(_712_)
);

FILL FILL_3__972_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_23_),
    .Y(_24_)
);

FILL FILL_1__1242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1168_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_281_),
    .B(_286_),
    .C(_244_),
    .Y(_287_)
);

FILL FILL_1__879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__922_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_43_),
    .B(_55_),
    .C(_57_),
    .Y(_117_)
);

FILL FILL_1__1336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1405_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_604_),
    .B(_607_),
    .Y(_608_)
);

FILL FILL_3__875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__989_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_400_),
    .B(_401_),
    .C(_402_),
    .Y(_403_)
);

FILL FILL_0__960_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_153_),
    .B(_148_),
    .C(_150_),
    .Y(_154_)
);

FILL FILL_1__1374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1512_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_648_),
    .B(_647_),
    .Y(_649_)
);

NAND2X1 _1021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_207_),
    .B(_208_),
    .Y(_211_)
);

FILL FILL_1__803_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_548_),
    .Y(_559_)
);

FILL FILL_1__1183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1321_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_739_),
    .B(_20_),
    .Y(_21_)
);

FILL FILL_1__1239_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_443_),
    .Y(_444_)
);

FILL FILL_2__1308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1061_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin_5_bF$buf3),
    .B(Cin[5]),
    .Y(_503_)
);

FILL FILL_3__778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1290_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1535_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(y[7]),
    .CLK(clk_bF$buf0),
    .Q(_755_[7])
);

AOI21X1 _1115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_300_),
    .B(_299_),
    .C(_214_),
    .Y(_305_)
);

FILL FILL_0__863_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_37_),
    .B(_35_),
    .C(_29_),
    .Y(_58_)
);

FILL FILL_1__1277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1415_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_529_),
    .B(_454_),
    .C(_544_),
    .Y(_545_)
);

FILL FILL_1__1086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1224_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_755_[13]),
    .Y(Yout[13])
);

NAND3X1 _1153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_327_),
    .B(_338_),
    .C(_330_),
    .Y(_342_)
);

FILL FILL_1__935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1384_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_214_),
    .B(_399_),
    .C(_292_),
    .Y(_400_)
);

FILL FILL88350x78150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1033_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_584_),
    .Y(_585_)
);

FILL FILL_0__1422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89250x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1509_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_638_),
    .B(_642_),
    .C(_645_),
    .Y(_646_)
);

INVX1 _1018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_208_),
    .Y(_209_)
);

FILL FILL_0__766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1262_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_483_),
    .Y(_526_)
);

NAND3X1 _1191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_378_),
    .B(_379_),
    .C(_376_),
    .Y(_380_)
);

FILL FILL_1__973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1318_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_361_),
    .B(_366_),
    .Y(_441_)
);

FILL FILL_0__995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1071_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_146_),
    .B(_185_),
    .C(_184_),
    .Y(_189_)
);

FILL FILL_1__782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1127_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_652_),
    .B(_657_),
    .C(_683_),
    .Y(_686_)
);

OAI21X1 _1056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_245_),
    .B(_158_),
    .C(_177_),
    .Y(_246_)
);

FILL FILL_1__838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1356_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_464_),
    .B(_468_),
    .C(_471_),
    .Y(_481_)
);

FILL FILL_4__1005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1165_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_278_),
    .B(_279_),
    .C(_277_),
    .Y(_284_)
);

FILL FILL_1__876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1104_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[4]),
    .B(Cin[7]),
    .Y(_582_)
);

FILL FILL_0__1419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1172_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_102_),
    .B(_105_),
    .C(_107_),
    .Y(_114_)
);

FILL FILL_1__1333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1259_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_354_),
    .B(_358_),
    .Y(_377_)
);

FILL FILL_2__1402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__757_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_596_),
    .B(_595_),
    .C(_594_),
    .Y(_605_)
);

FILL FILL_3__872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__928_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[4]),
    .Y(_151_)
);

FILL FILL_1__1371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__966_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8_),
    .B(_5_),
    .C(_746_),
    .Y(_18_)
);

FILL FILL_1__1236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1305_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_467_),
    .B(_465_),
    .C(_458_),
    .Y(_500_)
);

FILL FILL_3__775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__889_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1532_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(y[4]),
    .CLK(clk_bF$buf3),
    .Q(_755_[4])
);

NAND3X1 _1112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_213_),
    .B(_298_),
    .C(_301_),
    .Y(_302_)
);

FILL FILL_0__860_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_49_),
    .B(_54_),
    .Y(_55_)
);

FILL FILL_1__1274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1412_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_106_),
    .B(_110_),
    .C(_94_),
    .Y(_111_)
);

AND2X2 _1341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_522_),
    .B(_527_),
    .Y(_542_)
);

FILL FILL_1__1083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1139_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_755_[10]),
    .Y(Yout[10])
);

OAI21X1 _1150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_335_),
    .B(_334_),
    .C(_338_),
    .Y(_339_)
);

FILL FILL_1__932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1381_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_395_),
    .B(_394_),
    .C(_314_),
    .Y(_396_)
);

FILL FILL_0__954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1030_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_147_),
    .Y(_148_)
);

FILL FILL_1__1368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88350x54750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1506_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_577_),
    .B(_575_),
    .C(_641_),
    .Y(_642_)
);

NAND3X1 _1015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_137_),
    .B(_192_),
    .C(_197_),
    .Y(_206_)
);

FILL FILL_0__763_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf1),
    .B(Xin[1]),
    .C(Yin[1]),
    .Y(_493_)
);

FILL FILL_1__1177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1315_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_430_),
    .B(_431_),
    .C(_427_),
    .Y(_437_)
);

FILL FILL_0__992_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_184_),
    .B(_185_),
    .C(_182_),
    .Y(_186_)
);

FILL FILL_2__813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1124_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _1473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_682_),
    .B(Yin[13]),
    .Y(_683_)
);

NAND3X1 _1053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_218_),
    .B(_241_),
    .C(_242_),
    .Y(_243_)
);

FILL FILL_1__835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88950x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1284_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1529_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(y[1]),
    .CLK(clk_bF$buf4),
    .Q(_755_[1])
);

OAI21X1 _1109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_295_),
    .B(_296_),
    .C(_217_),
    .Y(_299_)
);

FILL FILL_0__857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1353_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_410_),
    .B(_469_),
    .C(_477_),
    .Y(_478_)
);

FILL FILL_4__788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1409_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_534_),
    .B(_538_),
    .Y(_539_)
);

FILL FILL_3__1582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1162_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_280_),
    .B(_246_),
    .C(_276_),
    .Y(_281_)
);

FILL FILL_1__873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1218_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_754_[7]),
    .Y(Xout[7])
);

NAND2X1 _1147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[3]),
    .B(Xin_5_bF$buf1),
    .Y(_336_)
);

FILL FILL_0__895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1391_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[2]),
    .B(Xin_3_bF$buf2),
    .C(_79_),
    .Y(_90_)
);

FILL FILL_4__1460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1027_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_577_),
    .B(_324_),
    .C(_578_),
    .Y(_579_)
);

FILL FILL_4__1516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1256_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_373_),
    .B(_368_),
    .C(_347_),
    .Y(_374_)
);

FILL FILL_1__967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1004_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_473_),
    .B(_474_),
    .C(_465_),
    .Y(_475_)
);

FILL FILL_4__1419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__963_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[1]),
    .B(Cin[3]),
    .Y(_15_)
);

FILL FILL_1__1233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88950x23550 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_274_),
    .B(_273_),
    .C(_260_),
    .Y(_278_)
);

FILL FILL_2__1302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1128_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_410_),
    .B(_477_),
    .C(_496_),
    .Y(_497_)
);

FILL FILL_3__772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1518_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_51_),
    .B(_740_),
    .C(_45_),
    .Y(_52_)
);

FILL FILL_1__1271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88350x19650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__913_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_104_),
    .B(_103_),
    .C(_96_),
    .Y(_108_)
);

FILL FILL_1__1327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1205_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_392_),
    .B(_387_),
    .C(_315_),
    .Y(_393_)
);

FILL FILL_0__951_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_105_),
    .B(_102_),
    .C(_95_),
    .Y(_145_)
);

FILL FILL_1__1365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88650x58650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1503_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[6]),
    .B(Xin[7]),
    .Y(_639_)
);

OAI21X1 _1012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_202_),
    .B(_198_),
    .C(_127_),
    .Y(_203_)
);

FILL FILL_0__760_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[0]),
    .B(Cin[1]),
    .Y(_461_)
);

FILL FILL_1__1174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1312_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4_),
    .B(_1_),
    .C(_0_),
    .Y(_12_)
);

NAND3X1 _1241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_414_),
    .B(_428_),
    .C(_433_),
    .Y(_434_)
);

AND2X2 _992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_157_),
    .B(_154_),
    .Y(_183_)
);

FILL FILL_2__810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1039_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_352_),
    .B(_575_),
    .C(_639_),
    .Y(_680_)
);

NAND3X1 _1050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_219_),
    .B(_234_),
    .C(_239_),
    .Y(_240_)
);

FILL FILL_1__832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1281_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1526_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(Xin[6]),
    .CLK(clk_bF$buf3),
    .Q(_754_[6])
);

AOI21X1 _1106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_281_),
    .B(_286_),
    .C(_244_),
    .Y(_296_)
);

FILL FILL_0__854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1350_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_44_),
    .B(_48_),
    .C(_46_),
    .Y(_49_)
);

FILL FILL_1__1268_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1406_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[10]),
    .Y(_535_)
);

FILL FILL_1__1497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1215_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_754_[4]),
    .Y(Xout[4])
);

NAND3X1 _1144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_332_),
    .B(_327_),
    .C(_330_),
    .Y(_333_)
);

FILL FILL_0__892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__926_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin_3_bF$buf1),
    .Y(_87_)
);

FILL FILL_2__1375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[6]),
    .B(Cin[6]),
    .Y(_576_)
);

FILL FILL_0__1413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1184_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_635_),
    .Y(_636_)
);

NAND3X1 _1009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_195_),
    .B(_196_),
    .C(_139_),
    .Y(_200_)
);

FILL FILL_0__757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1253_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_362_),
    .B(_370_),
    .Y(_371_)
);

FILL FILL_1__964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1309_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _1238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_415_),
    .B(_416_),
    .C(_419_),
    .Y(_431_)
);

FILL FILL_0__986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1062_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_179_),
    .B(_176_),
    .C(_146_),
    .Y(_180_)
);

FILL FILL_1__773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1118_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_576_),
    .Y(_677_)
);

NOR2X1 _1047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_152_),
    .B(_231_),
    .Y(_237_)
);

FILL FILL_0__795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1291_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_738_),
    .Y(_739_)
);

FILL FILL_0__1507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1347_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_382_),
    .B(_384_),
    .C(_470_),
    .Y(_471_)
);

FILL FILL_0__1316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1156_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_274_),
    .B(_273_),
    .C(_272_),
    .Y(_275_)
);

FILL FILL_1__867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88950x85950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__910_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_96_),
    .B(_103_),
    .C(_104_),
    .Y(_105_)
);

FILL FILL_1__1324_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_367_),
    .B(_365_),
    .C(_359_),
    .Y(_368_)
);

FILL FILL_0__1219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__919_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_383_),
    .B(_384_),
    .C(_382_),
    .Y(_390_)
);

FILL FILL89250x31350 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_78_),
    .B(_140_),
    .C(_141_),
    .Y(_142_)
);

FILL FILL_1__1362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__935_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_418_),
    .Y(_429_)
);

FILL FILL_1__1171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__957_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_746_),
    .B(_5_),
    .C(_8_),
    .Y(_9_)
);

FILL FILL_1__1227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1105_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1523_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(Xin_3_bF$buf1),
    .CLK(clk_bF$buf4),
    .Q(_754_[3])
);

INVX1 _1103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_189_),
    .Y(_293_)
);

FILL FILL_0__851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__995_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_743_),
    .B(_45_),
    .Y(_46_)
);

FILL FILL_1__1265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1403_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[4]),
    .B(Xin[7]),
    .Y(_532_)
);

FILL FILL_4__838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1212_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_754_[1]),
    .Y(Xout[1])
);

NAND3X1 _1141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_319_),
    .B(_328_),
    .C(_329_),
    .Y(_330_)
);

FILL FILL_1__923_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_83_),
    .Y(_84_)
);

FILL FILL_2__1372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1021_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_123_),
    .B(_138_),
    .C(_116_),
    .Y(_139_)
);

FILL FILL_1__1359_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_528_),
    .B(_540_),
    .C(_572_),
    .Y(_573_)
);

FILL FILL_2__1428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1181_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_618_),
    .B(_631_),
    .Y(_632_)
);

NAND3X1 _1006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_195_),
    .B(_196_),
    .C(_194_),
    .Y(_197_)
);

FILL FILL_3__898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1250_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[0]),
    .Y(_397_)
);

FILL FILL_1__1168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1306_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_348_),
    .B(_426_),
    .C(_351_),
    .Y(_427_)
);

FILL FILL_0__983_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_160_),
    .B(_173_),
    .C(_174_),
    .Y(_177_)
);

FILL FILL_1__1397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1115_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_671_),
    .B(_672_),
    .C(_670_),
    .Y(_673_)
);

NAND3X1 _1044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_226_),
    .B(_230_),
    .C(_233_),
    .Y(_234_)
);

FILL FILL_0__792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__826_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_731_),
    .B(_734_),
    .C(_559_),
    .Y(_737_)
);

FILL FILL_0__1504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1344_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_467_),
    .B(_466_),
    .C(_465_),
    .Y(_468_)
);

FILL FILL_0__1313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1084_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[9]),
    .B(_363_),
    .Y(_529_)
);

FILL FILL_3__1573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1153_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_260_),
    .Y(_272_)
);

FILL FILL_1__864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1209_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1558_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_753_[14]),
    .CLK(clk_bF$buf2),
    .Q(y[14])
);

NAND3X1 _1138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_326_),
    .B(_320_),
    .C(_323_),
    .Y(_327_)
);

FILL FILL_0__886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1382_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_80_),
    .B(_78_),
    .Y(_81_)
);

FILL FILL_4__1451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1018_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_516_),
    .B(_522_),
    .Y(_570_)
);

FILL FILL_3__1191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1160_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_98_),
    .B(_97_),
    .C(_101_),
    .Y(_102_)
);

FILL FILL_1__1321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1247_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_363_),
    .B(_364_),
    .C(_361_),
    .Y(_365_)
);

FILL FILL_1__958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89550x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__954_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[3]),
    .B(_3_),
    .Y(_6_)
);

FILL FILL_1__1224_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_709_),
    .B(_710_),
    .Y(_711_)
);

NAND3X1 _1079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf0),
    .B(Xin[7]),
    .C(_264_),
    .Y(_269_)
);

FILL FILL_0__1119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1509_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1520_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(Xin[0]),
    .CLK(clk_bF$buf1),
    .Q(_754_[0])
);

NAND3X1 _1100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_276_),
    .B(_280_),
    .C(_283_),
    .Y(_290_)
);

FILL FILL_3__992_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_42_),
    .B(_41_),
    .C(_40_),
    .Y(_43_)
);

FILL FILL_1__1262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1400_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[5]),
    .Y(_99_)
);

FILL FILL_1__1318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__942_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_73_),
    .B(_133_),
    .C(_132_),
    .Y(_136_)
);

FILL FILL_1__1356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1005_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_565_),
    .Y(_629_)
);

AOI21X1 _1003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_81_),
    .B(_120_),
    .C(_193_),
    .Y(_194_)
);

FILL FILL_3__895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89550x23550 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_322_),
    .B(_423_),
    .Y(_424_)
);

FILL FILL_0__980_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_161_),
    .B(_163_),
    .C(_165_),
    .Y(_174_)
);

FILL FILL_1__1394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1112_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_670_),
    .B(_668_),
    .Y(_671_)
);

NAND2X1 _1041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[2]),
    .B(Xin[4]),
    .Y(_231_)
);

FILL FILL_1__823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__967_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_718_),
    .B(_733_),
    .C(_732_),
    .Y(_734_)
);

FILL FILL_2__1519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1098_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_728_),
    .B(_722_),
    .Y(_753_[15])
);

FILL FILL_0__845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1341_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_),
    .B(_4_),
    .C(_39_),
    .Y(_40_)
);

FILL FILL_1__1259_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_434_),
    .B(_438_),
    .Y(_465_)
);

FILL FILL_4__1410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1081_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_517_),
    .B(_518_),
    .C(_514_),
    .Y(_525_)
);

FILL FILL_3__798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1206_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1555_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_753_[11]),
    .CLK(clk_bF$buf5),
    .Q(y[11])
);

INVX1 _1135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[6]),
    .Y(_324_)
);

FILL FILL_0__883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__917_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_397_),
    .B(_77_),
    .Y(_78_)
);

FILL FILL_1__1297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1015_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_565_),
    .B(_495_),
    .C(_564_),
    .Y(_566_)
);

FILL FILL_0__1404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89250x58650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1244_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[1]),
    .B(Xin[7]),
    .C(Yin[8]),
    .Y(_362_)
);

FILL FILL_1__955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1213_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_415_),
    .Y(_421_)
);

FILL FILL_0__977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1109_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_615_),
    .B(_621_),
    .C(_667_),
    .Y(_668_)
);

NAND2X1 _1038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_227_),
    .B(_140_),
    .Y(_228_)
);

FILL FILL_0__786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1282_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_601_),
    .B(_708_),
    .C(_729_),
    .Y(_731_)
);

FILL FILL_1__993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89550x11850 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1338_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_454_),
    .B(_457_),
    .Y(_462_)
);

FILL FILL_3__1091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__951_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf2),
    .B(Xin_3_bF$buf0),
    .Y(_3_)
);

FILL FILL_1__1221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1147_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_703_),
    .B(_706_),
    .Y(_707_)
);

NAND2X1 _1076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_264_),
    .B(_265_),
    .Y(_266_)
);

FILL FILL_1__858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__901_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[1]),
    .B(Xin[4]),
    .Y(_96_)
);

FILL FILL_1__1315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1124_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_593_),
    .B(_597_),
    .C(_603_),
    .Y(_604_)
);

FILL FILL_0__1439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1192_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_133_),
    .Y(_134_)
);

FILL FILL_1__1353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1409_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_566_),
    .B(_626_),
    .Y(_753_[11])
);

AOI21X1 _1000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_190_),
    .B(_189_),
    .C(_188_),
    .Y(_191_)
);

FILL FILL_3__892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1300_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_747_),
    .Y(_0_)
);

FILL FILL_1__1218_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_170_),
    .B(_166_),
    .C(_160_),
    .Y(_171_)
);

FILL FILL_1__1391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89550x85950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1095_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_725_),
    .B(_724_),
    .C(_713_),
    .Y(_726_)
);

FILL FILL_0__842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__986_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_31_),
    .B(_36_),
    .C(_33_),
    .Y(_37_)
);

FILL FILL_1__1256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1325_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_501_),
    .B(_516_),
    .C(_521_),
    .Y(_522_)
);

FILL FILL_3__795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1203_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1552_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_753_[8]),
    .CLK(clk_bF$buf1),
    .Q(y[8])
);

AND2X2 _1132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[2]),
    .B(Cin[6]),
    .Y(_321_)
);

FILL FILL_0__880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__914_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_74_),
    .Y(_75_)
);

FILL FILL_1__1294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1012_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .B(_130_),
    .C(_128_),
    .Y(_131_)
);

NAND3X1 _1361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_562_),
    .B(_563_),
    .C(_561_),
    .Y(_564_)
);

FILL FILL_2__1419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1172_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_620_),
    .B(_621_),
    .C(_622_),
    .Y(_624_)
);

FILL FILL_3__889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1159_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_358_),
    .B(_354_),
    .Y(_359_)
);

FILL FILL_1__952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1228_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[4]),
    .B(Cin[6]),
    .Y(_417_)
);

FILL FILL_0__974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1050_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf3),
    .B(Xin[6]),
    .C(Yin[6]),
    .Y(_168_)
);

FILL FILL_1__1388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1106_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_659_),
    .B(_637_),
    .Y(_664_)
);

OAI21X1 _1035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_47_),
    .B(_77_),
    .C(_224_),
    .Y(_225_)
);

FILL FILL_0__783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__817_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_612_),
    .B(_676_),
    .C(_697_),
    .Y(_708_)
);

FILL FILL_1__1197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1335_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_454_),
    .B(_457_),
    .C(_442_),
    .Y(_458_)
);

FILL FILL_0__1304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1144_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[14]),
    .Y(_704_)
);

NAND3X1 _1073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf0),
    .B(Xin[7]),
    .C(Yin[7]),
    .Y(_263_)
);

FILL FILL_1__855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1113_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1549_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_753_[5]),
    .CLK(clk_bF$buf3),
    .Q(y[5])
);

OAI21X1 _1129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_224_),
    .B(_227_),
    .C(_226_),
    .Y(_318_)
);

FILL FILL_0__877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1009_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_479_),
    .B(_560_),
    .C(_469_),
    .Y(_561_)
);

FILL FILL_3__1182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1169_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_83_),
    .B(_90_),
    .C(_92_),
    .Y(_93_)
);

FILL FILL_1__1312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1238_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[3]),
    .B(Xin_5_bF$buf1),
    .C(_355_),
    .Y(_356_)
);

FILL FILL_1__949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1047_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_534_),
    .B(_598_),
    .Y(_600_)
);

FILL FILL_1__758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__945_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_744_),
    .B(_742_),
    .Y(_745_)
);

FILL FILL_1__1215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1024_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _1299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_475_),
    .B(_476_),
    .C(_471_),
    .Y(_496_)
);

FILL FILL_2__1513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1092_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_618_),
    .B(_631_),
    .C(_627_),
    .D(_492_),
    .Y(_723_)
);

FILL FILL_3__983_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_33_),
    .Y(_34_)
);

FILL FILL_1__1253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1309_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_350_),
    .B(_445_),
    .Y(_519_)
);

FILL FILL_3__792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__911_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_71_),
    .B(_68_),
    .Y(_72_)
);

FILL FILL_1__1291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__933_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_67_),
    .B(_26_),
    .C(_69_),
    .Y(_128_)
);

FILL FILL_1__1347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1416_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_499_),
    .B(_619_),
    .C(_555_),
    .Y(_620_)
);

FILL FILL_3__886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1225_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_227_),
    .B(_413_),
    .C(_327_),
    .Y(_414_)
);

FILL FILL_0__971_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf3),
    .B(Xin[6]),
    .C(_164_),
    .Y(_165_)
);

FILL FILL_1__1385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1103_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_660_),
    .Y(_661_)
);

AND2X2 _1032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[2]),
    .B(Cin[5]),
    .Y(_222_)
);

FILL FILL_0__780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_633_),
    .B(_644_),
    .C(_666_),
    .Y(_676_)
);

FILL FILL_1__1194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1089_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _1508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_719_),
    .B(Yin[15]),
    .Y(_720_)
);

FILL FILL_0__836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1332_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf2),
    .B(Xin[4]),
    .C(Yin[4]),
    .Y(_31_)
);

NAND2X1 _1261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_449_),
    .B(_452_),
    .Y(_455_)
);

FILL FILL_4__1401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1072_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_507_),
    .B(_512_),
    .C(_514_),
    .Y(_516_)
);

FILL FILL_3__789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1059_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_692_),
    .Y(_701_)
);

OAI21X1 _1070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_161_),
    .B(_259_),
    .C(_168_),
    .Y(_260_)
);

FILL FILL_1__852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1128_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1546_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_750_[2]),
    .CLK(clk_bF$buf4),
    .Q(y[2])
);

INVX1 _1126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_314_),
    .Y(_315_)
);

FILL FILL_0__874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1370_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9_),
    .B(_14_),
    .C(_65_),
    .D(_66_),
    .Y(_69_)
);

FILL FILL_1__1288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88050x78150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1006_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_556_),
    .B(_555_),
    .C(_498_),
    .Y(_557_)
);

FILL FILL_1__1097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1235_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_590_),
    .B(_352_),
    .C(_336_),
    .Y(_353_)
);

FILL FILL_1__946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1044_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_594_),
    .B(_595_),
    .C(_596_),
    .Y(_597_)
);

FILL FILL_0__1433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__904_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_648_),
    .B(_647_),
    .C(_654_),
    .Y(_658_)
);

INVX1 _1029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_218_),
    .Y(_219_)
);

FILL FILL_0__777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1329_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_443_),
    .B(_450_),
    .C(_451_),
    .Y(_452_)
);

FILL FILL_3__1082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__942_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_397_),
    .B(_740_),
    .C(_741_),
    .Y(_742_)
);

FILL FILL_1__1212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1138_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_696_),
    .Y(_698_)
);

NAND3X1 _1067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_247_),
    .B(_255_),
    .C(_256_),
    .Y(_257_)
);

FILL FILL_1__849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1367_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_403_),
    .B(_491_),
    .C(_484_),
    .Y(_492_)
);

FILL FILL_2__1510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__930_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_115_),
    .B(_111_),
    .C(_117_),
    .Y(_125_)
);

FILL FILL_1__1344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__861_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_244_),
    .B(_286_),
    .C(_388_),
    .Y(_389_)
);

FILL FILL_2__1413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1092_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_616_),
    .B(_615_),
    .C(_570_),
    .Y(_617_)
);

FILL FILL_3__883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1209_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_378_),
    .B(_379_),
    .C(_347_),
    .Y(_411_)
);

NAND2X1 _971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf3),
    .B(Xin[6]),
    .Y(_162_)
);

FILL FILL_1__1382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__811_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf1),
    .B(Xin[2]),
    .C(Yin[2]),
    .Y(_644_)
);

FILL FILL_1__1191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1086_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_714_),
    .B(_700_),
    .C(_715_),
    .Y(_716_)
);

FILL FILL_0__833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__977_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf2),
    .B(Xin_3_bF$buf0),
    .C(Yin[3]),
    .Y(_28_)
);

FILL FILL_1__1247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89250x150 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_508_),
    .B(_511_),
    .C(_510_),
    .Y(_512_)
);

FILL FILL_3__786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1125_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1543_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(y[15]),
    .CLK(clk_bF$buf2),
    .Q(_755_[15])
);

INVX1 _1123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_292_),
    .Y(_312_)
);

FILL FILL_0__871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__905_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_38_),
    .B(_61_),
    .C(_43_),
    .Y(_66_)
);

FILL FILL_1__1285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1003_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549_),
    .B(_553_),
    .C(_499_),
    .Y(_554_)
);

FILL FILL_1__1094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88050x54750 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_609_),
    .B(_613_),
    .C(_571_),
    .Y(_614_)
);

FILL FILL_3__1232_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_755_[7]),
    .Y(Yout[7])
);

AND2X2 _1161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[3]),
    .B(Xin[6]),
    .Y(_350_)
);

FILL FILL_1__943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1392_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_390_),
    .B(_391_),
    .C(_317_),
    .Y(_408_)
);

FILL FILL_0__965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1041_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf3),
    .B(Xin_5_bF$buf0),
    .C(Yin[5]),
    .Y(_159_)
);

FILL FILL_1__1379_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_574_),
    .Y(_594_)
);

FILL FILL_4__1110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1517_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_653_),
    .B(_652_),
    .Y(_654_)
);

AOI21X1 _1026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_184_),
    .B(_185_),
    .C(_146_),
    .Y(_216_)
);

FILL FILL_0__774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1270_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_461_),
    .B(_493_),
    .C(_483_),
    .Y(_612_)
);

FILL FILL88650x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1326_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_444_),
    .B(_448_),
    .C(_446_),
    .Y(_449_)
);

FILL FILL_1__790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1135_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_673_),
    .B(_694_),
    .Y(_753_[13])
);

NAND3X1 _1064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_253_),
    .B(_248_),
    .C(_251_),
    .Y(_254_)
);

FILL FILL_1__846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88950x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_484_),
    .B(_489_),
    .Y(_490_)
);

FILL FILL_4__1433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__804_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_522_),
    .B(_527_),
    .C(_546_),
    .Y(_551_)
);

FILL FILL_3__1173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__820_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_755_[4]),
    .Y(Yout[4])
);

OAI21X1 _1158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_346_),
    .B(_277_),
    .C(_271_),
    .Y(_347_)
);

FILL FILL_4__1051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1038_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_582_),
    .B(_580_),
    .Y(_591_)
);

FILL FILL_0__1427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1180_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_78_),
    .Y(_122_)
);

FILL FILL_1__1341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1267_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_383_),
    .B(_384_),
    .C(_382_),
    .Y(_385_)
);

FILL FILL_1__978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1076_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[3]),
    .Y(Xin_3_bF$buf3)
);

BUFX2 BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[3]),
    .Y(Xin_3_bF$buf2)
);

BUFX2 BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[3]),
    .Y(Xin_3_bF$buf1)
);

BUFX2 BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[3]),
    .Y(Xin_3_bF$buf0)
);

BUFX2 BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[5]),
    .Y(Xin_5_bF$buf3)
);

BUFX2 BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[5]),
    .Y(Xin_5_bF$buf2)
);

BUFX2 BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[5]),
    .Y(Xin_5_bF$buf1)
);

BUFX2 BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[5]),
    .Y(Xin_5_bF$buf0)
);

FILL FILL_1__787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88650x23550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1083_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_713_),
    .Y(_714_)
);

FILL FILL_0__830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__974_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24_),
    .B(_25_),
    .Y(_751_[3])
);

FILL FILL_1__1244_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_285_),
    .B(_284_),
    .C(_246_),
    .Y(_289_)
);

FILL FILL_2__1313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88050x19650 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin_5_bF$buf3),
    .B(Cin[5]),
    .Y(_509_)
);

FILL FILL_3__783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1109_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1540_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(y[12]),
    .CLK(clk_bF$buf2),
    .Q(_755_[12])
);

INVX1 _1120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_307_),
    .Y(_309_)
);

FILL FILL_1__902_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_27_),
    .B(_56_),
    .C(_62_),
    .Y(_63_)
);

FILL FILL_1__1282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1000_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_89_),
    .B(_93_),
    .C(_110_),
    .D(_106_),
    .Y(_119_)
);

FILL FILL_1__1338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1160_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_572_),
    .Y(_610_)
);

FILL FILL_3__877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1216_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _1214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_311_),
    .B(_404_),
    .Y(_753_[8])
);

FILL FILL_0__962_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_87_),
    .B(_740_),
    .C(_149_),
    .Y(_156_)
);

FILL FILL_1__1376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1514_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[11]),
    .B(_532_),
    .Y(_651_)
);

OAI21X1 _1023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_137_),
    .B(_212_),
    .C(_200_),
    .Y(_213_)
);

FILL FILL_0__771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88950x39150 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_569_),
    .B(_559_),
    .Y(_749_[1])
);

FILL FILL_1__1185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1323_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_350_),
    .B(_445_),
    .Y(_446_)
);

FILL FILL_2__821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1063_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin_5_bF$buf3),
    .B(Cin[5]),
    .C(Xin[4]),
    .D(Cin[6]),
    .Y(_506_)
);

FILL FILL_3__1132_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_647_),
    .B(_684_),
    .C(_691_),
    .Y(_692_)
);

NAND2X1 _1061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_249_),
    .B(_250_),
    .Y(_251_)
);

FILL FILL_1__843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1292_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1537_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(y[9]),
    .CLK(clk_bF$buf0),
    .Q(_755_[9])
);

OAI21X1 _1117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_306_),
    .B(_305_),
    .C(_304_),
    .Y(_307_)
);

FILL FILL_0__865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1361_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_44_),
    .B(_52_),
    .C(_53_),
    .Y(_60_)
);

FILL FILL_1__1279_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_481_),
    .B(_480_),
    .C(_479_),
    .Y(_487_)
);

FILL FILL_2__1348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1417_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_546_),
    .B(_542_),
    .Y(_547_)
);

FILL FILL_3__1170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1226_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_755_[15]),
    .Y(Yout[15])
);

NAND3X1 _1155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_341_),
    .B(_342_),
    .C(_343_),
    .Y(_344_)
);

FILL FILL_1__937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1035_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_536_),
    .B(_581_),
    .C(_586_),
    .Y(_587_)
);

FILL FILL_0__1424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1264_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_340_),
    .B(_344_),
    .Y(_382_)
);

FILL FILL_1__975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__762_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin_5_bF$buf1),
    .B(Cin[4]),
    .Y(_443_)
);

FILL FILL_0__997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88950x27450 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_650_),
    .B(_651_),
    .C(_657_),
    .Y(_689_)
);

INVX1 _1058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_247_),
    .Y(_248_)
);

FILL FILL_0__1518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88650x85950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1358_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_409_),
    .B(_478_),
    .C(_482_),
    .Y(_484_)
);

FILL FILL_2__1501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__971_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_735_),
    .B(_22_),
    .C(_21_),
    .Y(_23_)
);

FILL FILL_1__1241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1167_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_284_),
    .B(_285_),
    .C(_283_),
    .Y(_286_)
);

FILL FILL_1__878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__921_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_115_),
    .B(_111_),
    .C(_82_),
    .Y(_116_)
);

FILL FILL_1__1335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1083_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_605_),
    .B(_606_),
    .C(_602_),
    .Y(_607_)
);

FILL FILL_3__874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__988_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_315_),
    .B(_387_),
    .C(_392_),
    .Y(_402_)
);

OAI21X1 _962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_590_),
    .B(_151_),
    .C(_152_),
    .Y(_153_)
);

FILL FILL_1__1373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1268_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1009_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_645_),
    .B(_642_),
    .C(_638_),
    .Y(_648_)
);

NOR2X1 _1020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_210_),
    .B(_209_),
    .Y(_753_[6])
);

FILL FILL_1__802_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_515_),
    .B(_537_),
    .C(_429_),
    .Y(_548_)
);

FILL FILL_1__1182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1320_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_14_),
    .B(_19_),
    .Y(_20_)
);

FILL FILL_1__1238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88950x15750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1060_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin_3_bF$buf3),
    .B(Cin[7]),
    .Y(_502_)
);

FILL FILL_3__777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1116_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1534_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(y[6]),
    .CLK(clk_bF$buf0),
    .Q(_755_[6])
);

AOI21X1 _1114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_199_),
    .B(_201_),
    .C(_303_),
    .Y(_304_)
);

FILL FILL_0__862_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_41_),
    .B(_42_),
    .C(_40_),
    .Y(_57_)
);

FILL FILL_1__1276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1414_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_538_),
    .B(_534_),
    .Y(_544_)
);

FILL FILL_1__1085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1223_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_755_[12]),
    .Y(Yout[12])
);

AND2X2 _1152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_226_),
    .B(_223_),
    .Y(_341_)
);

FILL FILL_1__934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1383_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_287_),
    .B(_291_),
    .C(_217_),
    .Y(_399_)
);

FILL FILL_0__956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1032_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_85_),
    .B(_149_),
    .Y(_150_)
);

NOR2X1 _1381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_503_),
    .B(_576_),
    .Y(_584_)
);

FILL FILL_4__1101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1508_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_641_),
    .B(_643_),
    .Y(_645_)
);

NAND3X1 _1017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_136_),
    .B(_207_),
    .C(_203_),
    .Y(_208_)
);

FILL FILL_0__765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1261_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_472_),
    .B(_483_),
    .C(_504_),
    .Y(_515_)
);

FILL FILL_1__1179_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_365_),
    .B(_359_),
    .C(_367_),
    .Y(_379_)
);

FILL FILL_1__972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1317_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_434_),
    .B(_438_),
    .Y(_439_)
);

FILL FILL_0__994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1070_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_143_),
    .B(_142_),
    .Y(_188_)
);

FILL FILL_1__781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1126_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_684_),
    .Y(_685_)
);

AOI21X1 _1055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_174_),
    .B(_173_),
    .C(_160_),
    .Y(_245_)
);

FILL FILL_1__837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1355_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_476_),
    .B(_475_),
    .C(_412_),
    .Y(_480_)
);

FILL FILL_4__1424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1164_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_183_),
    .B(_178_),
    .C(_282_),
    .Y(_283_)
);

FILL FILL_1__875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__811_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_755_[1]),
    .Y(Yout[1])
);

AOI22X1 _1149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_149_),
    .B(_337_),
    .C(_253_),
    .D(_248_),
    .Y(_338_)
);

FILL FILL_0__897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1029_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_151_),
    .B(_575_),
    .C(_580_),
    .Y(_581_)
);

FILL FILL_0__1418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89550x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88650x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89250x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_109_),
    .B(_108_),
    .C(_95_),
    .Y(_113_)
);

FILL FILL_1__1332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1258_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_258_),
    .B(_275_),
    .C(_375_),
    .Y(_376_)
);

FILL FILL_1__969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89550x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__965_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9_),
    .Y(_17_)
);

FILL FILL_1__1235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1304_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_498_),
    .Y(_499_)
);

FILL FILL_3__774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__888_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1531_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(y[3]),
    .CLK(clk_bF$buf3),
    .Q(_755_[3])
);

NAND3X1 _1111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_214_),
    .B(_299_),
    .C(_300_),
    .Y(_301_)
);

NAND3X1 _862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_50_),
    .B(_52_),
    .C(_53_),
    .Y(_54_)
);

FILL FILL_1__1273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1411_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_109_),
    .B(_108_),
    .C(_107_),
    .Y(_110_)
);

FILL FILL_1__1329_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_528_),
    .B(_540_),
    .Y(_541_)
);

FILL FILL_1__1082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89250x23550 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_381_),
    .B(_385_),
    .C(_389_),
    .Y(_395_)
);

FILL FILL_0__953_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[2]),
    .B(Cin[4]),
    .Y(_147_)
);

FILL FILL_1__1367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1505_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_578_),
    .B(_639_),
    .C(_640_),
    .Y(_641_)
);

NAND3X1 _1014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_199_),
    .B(_200_),
    .C(_201_),
    .Y(_205_)
);

FILL FILL_0__762_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf1),
    .B(Xin[1]),
    .C(Yin[1]),
    .Y(_483_)
);

FILL FILL_1__1176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1314_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_425_),
    .B(_432_),
    .C(_420_),
    .Y(_436_)
);

FILL FILL_0__991_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_158_),
    .B(_171_),
    .C(_175_),
    .Y(_185_)
);

FILL FILL_2__812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1123_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_681_),
    .B(_675_),
    .Y(_682_)
);

OAI21X1 _1052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_236_),
    .B(_235_),
    .C(_233_),
    .Y(_242_)
);

FILL FILL_1__834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1283_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1528_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(y[0]),
    .CLK(clk_bF$buf4),
    .Q(_755_[0])
);

NAND3X1 _1108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_215_),
    .B(_292_),
    .C(_297_),
    .Y(_298_)
);

FILL FILL_0__856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1352_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[1]),
    .Y(_51_)
);

OAI21X1 _1281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_475_),
    .B(_476_),
    .C(_471_),
    .Y(_477_)
);

FILL FILL_0__1321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1408_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_531_),
    .B(_536_),
    .C(_535_),
    .Y(_538_)
);

FILL FILL_3__1581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1079_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_277_),
    .B(_279_),
    .C(_278_),
    .Y(_280_)
);

FILL FILL_1__872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1217_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_754_[6]),
    .Y(Xout[6])
);

AOI21X1 _1146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_323_),
    .B(_326_),
    .C(_320_),
    .Y(_335_)
);

FILL FILL_0__894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1390_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_84_),
    .B(_88_),
    .C(_86_),
    .Y(_89_)
);

FILL FILL_2__1377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1026_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[5]),
    .B(Xin[6]),
    .Y(_578_)
);

FILL FILL_0__1415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89550x39150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1255_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_354_),
    .B(_358_),
    .C(_369_),
    .D(_372_),
    .Y(_373_)
);

FILL FILL_1__966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89250x11850 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__924_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_677_),
    .B(_678_),
    .Y(_679_)
);

OAI21X1 _1049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_236_),
    .B(_235_),
    .C(_238_),
    .Y(_239_)
);

FILL FILL_0__797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__940_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_454_),
    .B(_457_),
    .C(_460_),
    .Y(_474_)
);

FILL FILL_0__1318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__962_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9_),
    .B(_13_),
    .C(_745_),
    .Y(_14_)
);

FILL FILL_1__1232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1158_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254_),
    .B(_257_),
    .Y(_277_)
);

FILL FILL_1__869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__912_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_95_),
    .Y(_107_)
);

FILL FILL_1__1326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89550x27450 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_390_),
    .B(_391_),
    .C(_389_),
    .Y(_392_)
);

FILL FILL_0__950_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_143_),
    .B(_142_),
    .Y(_144_)
);

FILL FILL_1__1364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89250x85950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1259_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1502_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_582_),
    .B(_580_),
    .C(_585_),
    .Y(_638_)
);

AOI21X1 _1011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_201_),
    .B(_200_),
    .C(_199_),
    .Y(_202_)
);

NOR2X1 _762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_440_),
    .B(_429_),
    .Y(_748_[0])
);

FILL FILL_1__1173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1311_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7_),
    .B(_6_),
    .C(_747_),
    .Y(_11_)
);

FILL FILL_1__1229_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_430_),
    .B(_431_),
    .C(_432_),
    .Y(_433_)
);

AOI21X1 _991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_94_),
    .B(_110_),
    .C(_181_),
    .Y(_182_)
);

FILL FILL_2__1471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1280_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1525_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(Xin_5_bF$buf2),
    .CLK(clk_bF$buf0),
    .Q(_754_[5])
);

AOI21X1 _1105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_290_),
    .B(_289_),
    .C(_288_),
    .Y(_295_)
);

FILL FILL_0__853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__997_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_47_),
    .B(_590_),
    .C(_15_),
    .Y(_48_)
);

FILL FILL_1__1267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1405_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[10]),
    .B(_533_),
    .Y(_534_)
);

FILL FILL_1__1496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1214_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_754_[3]),
    .Y(Xout[3])
);

OAI21X1 _1143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_247_),
    .B(_331_),
    .C(_251_),
    .Y(_332_)
);

FILL FILL_0__891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__925_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_45_),
    .B(_85_),
    .Y(_86_)
);

FILL FILL_2__1374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1023_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[7]),
    .Y(_575_)
);

FILL FILL_0__1412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1183_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_587_),
    .B(_593_),
    .Y(_635_)
);

INVX1 _1008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_137_),
    .Y(_199_)
);

FILL FILL_0__756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1252_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[0]),
    .B(_407_),
    .Y(_418_)
);

INVX1 _1181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_364_),
    .Y(_370_)
);

FILL FILL_1__963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89550x15750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1308_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_424_),
    .B(_422_),
    .C(_421_),
    .Y(_430_)
);

FILL FILL_0__985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1061_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_154_),
    .B(_157_),
    .C(_178_),
    .D(_177_),
    .Y(_179_)
);

FILL FILL_1__1399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1117_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _1466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_578_),
    .B(_639_),
    .C(_643_),
    .D(_641_),
    .Y(_675_)
);

AOI22X1 _1046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[0]),
    .B(Cin[7]),
    .C(_223_),
    .D(_225_),
    .Y(_236_)
);

FILL FILL_0__794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1290_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_732_),
    .B(_718_),
    .C(_708_),
    .Y(_738_)
);

FILL FILL_0__1506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1346_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_383_),
    .Y(_470_)
);

FILL FILL_0__1315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1155_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_266_),
    .B(_263_),
    .C(_262_),
    .Y(_274_)
);

FILL FILL_1__866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1514_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_544_),
    .B(_530_),
    .Y(_572_)
);

FILL FILL_3__1193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1162_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf2),
    .B(Xin_5_bF$buf2),
    .C(_99_),
    .Y(_104_)
);

FILL FILL_1__1323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1249_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_263_),
    .B(_267_),
    .C(_366_),
    .Y(_367_)
);

FILL FILL_4__1318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__918_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[0]),
    .B(Cin[6]),
    .C(Xin[1]),
    .D(Cin[5]),
    .Y(_141_)
);

FILL FILL_1__1361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__956_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_747_),
    .B(_6_),
    .C(_7_),
    .Y(_8_)
);

FILL FILL_1__1226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__879_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1522_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(Xin[2]),
    .CLK(clk_bF$buf4),
    .Q(_754_[2])
);

NAND3X1 _1102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_291_),
    .B(_287_),
    .C(_217_),
    .Y(_292_)
);

FILL FILL_0__850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__994_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[2]),
    .B(Cin[2]),
    .Y(_45_)
);

FILL FILL_1__1264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1402_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_99_),
    .B(_100_),
    .Y(_101_)
);

AOI22X1 _1331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[3]),
    .B(Xin[7]),
    .C(Cin[4]),
    .D(Xin[6]),
    .Y(_531_)
);

FILL FILL_1__1493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88650x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1129_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_754_[0]),
    .Y(Xout[0])
);

OAI21X1 _1140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_47_),
    .B(_324_),
    .C(_322_),
    .Y(_329_)
);

FILL FILL_1__922_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[1]),
    .B(Cin[4]),
    .Y(_83_)
);

FILL FILL_2__1371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1020_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_111_),
    .B(_115_),
    .C(_82_),
    .Y(_138_)
);

FILL FILL_1__1358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1180_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_624_),
    .B(_564_),
    .Y(_631_)
);

NAND3X1 _1005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_144_),
    .B(_180_),
    .C(_186_),
    .Y(_196_)
);

FILL FILL_3__897_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf1),
    .Y(_386_)
);

FILL FILL_1__1167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1305_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_336_),
    .B(_355_),
    .Y(_426_)
);

FILL FILL_0__982_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_171_),
    .B(_175_),
    .C(_158_),
    .Y(_176_)
);

FILL FILL_1__1396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1114_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_634_),
    .Y(_672_)
);

OAI21X1 _1043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_147_),
    .B(_232_),
    .C(_150_),
    .Y(_233_)
);

FILL FILL_0__791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__825_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_735_),
    .Y(_736_)
);

FILL FILL_0__1503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1274_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_730_),
    .B(_72_),
    .Y(_752_[4])
);

FILL FILL_0__847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1343_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_454_),
    .B(_457_),
    .C(_442_),
    .Y(_467_)
);

FILL FILL_4__778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1083_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_522_),
    .B(_527_),
    .Y(_528_)
);

FILL FILL_3__1572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1152_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_260_),
    .B(_267_),
    .C(_270_),
    .Y(_271_)
);

FILL FILL_1__863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1208_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1557_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_753_[13]),
    .CLK(clk_bF$buf5),
    .Q(y[13])
);

OAI21X1 _1137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_47_),
    .B(_324_),
    .C(_325_),
    .Y(_326_)
);

FILL FILL_0__885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1381_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_741_),
    .B(_79_),
    .C(_59_),
    .Y(_80_)
);

FILL FILL_1__1299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1017_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_498_),
    .B(_556_),
    .C(_567_),
    .Y(_568_)
);

FILL FILL_3__1190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1246_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[1]),
    .B(Xin[7]),
    .C(Yin[8]),
    .Y(_364_)
);

FILL FILL_1__957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1414_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_458_),
    .B(_463_),
    .C(_439_),
    .Y(_464_)
);

FILL FILL_3__1093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__953_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_),
    .B(_0_),
    .C(_4_),
    .Y(_5_)
);

FILL FILL_1__1223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1149_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[13]),
    .B(_682_),
    .Y(_710_)
);

NAND2X1 _1078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[7]),
    .B(_265_),
    .Y(_268_)
);

FILL FILL_0__1118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__991_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_30_),
    .B(_33_),
    .C(_32_),
    .Y(_42_)
);

FILL FILL_1__1261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__903_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf3),
    .B(Xin_5_bF$buf0),
    .C(Yin[5]),
    .Y(_98_)
);

FILL FILL_1__1317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__941_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135_),
    .B(_73_),
    .Y(_753_[5])
);

FILL FILL_1__1355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__779_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_494_),
    .B(_311_),
    .C(_627_),
    .Y(_628_)
);

INVX1 _1002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_116_),
    .Y(_193_)
);

FILL FILL_3__894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1302_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[3]),
    .Y(_2_)
);

AND2X2 _1231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[4]),
    .B(Cin[6]),
    .Y(_423_)
);

NAND3X1 _982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_168_),
    .B(_167_),
    .C(_169_),
    .Y(_173_)
);

FILL FILL_1__1393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1029_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_669_),
    .B(_665_),
    .C(_663_),
    .Y(_670_)
);

NAND3X1 _1040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_220_),
    .B(_228_),
    .C(_229_),
    .Y(_230_)
);

FILL FILL_1__822_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_708_),
    .Y(_733_)
);

FILL FILL_2__1518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1097_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_715_),
    .B(_727_),
    .C(_726_),
    .Y(_728_)
);

FILL FILL_0__844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1340_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_),
    .Y(_39_)
);

FILL FILL_1__1258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88950x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1080_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_512_),
    .B(_507_),
    .C(_520_),
    .Y(_524_)
);

FILL FILL_3__797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1205_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1554_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_753_[10]),
    .CLK(clk_bF$buf5),
    .Q(y[10])
);

NAND2X1 _1134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_321_),
    .B(_322_),
    .Y(_323_)
);

FILL FILL_0__882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__916_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[5]),
    .Y(_77_)
);

FILL FILL_1__1296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1014_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_495_),
    .B(_565_),
    .Y(_753_[10])
);

FILL FILL_0__1403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1174_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_625_),
    .Y(_626_)
);

FILL FILL_3__1243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88350x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_261_),
    .B(_360_),
    .C(_263_),
    .Y(_361_)
);

FILL FILL_1__954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1212_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_416_),
    .B(_419_),
    .C(_415_),
    .Y(_420_)
);

FILL FILL_0__976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1052_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_169_),
    .B(_168_),
    .C(_167_),
    .Y(_170_)
);

FILL FILL_1__763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1108_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_665_),
    .B(_663_),
    .Y(_667_)
);

NAND2X1 _1037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[2]),
    .B(Cin[5]),
    .Y(_227_)
);

FILL FILL_0__785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1281_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_718_),
    .Y(_729_)
);

FILL FILL_1__1199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1268_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88650x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_377_),
    .B(_372_),
    .C(_459_),
    .Y(_460_)
);

FILL FILL_3__1090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1146_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_677_),
    .B(_705_),
    .C(_704_),
    .Y(_706_)
);

NAND2X1 _1075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf0),
    .B(Xin[7]),
    .Y(_265_)
);

FILL FILL_1__857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__900_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_33_),
    .B(_31_),
    .C(_30_),
    .Y(_95_)
);

FILL FILL_1__1314_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_348_),
    .B(_356_),
    .C(_357_),
    .Y(_358_)
);

FILL FILL_4__1309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL89550x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1049_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_602_),
    .Y(_603_)
);

FILL FILL_0__1438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1191_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_127_),
    .B(_131_),
    .C(_72_),
    .D(_21_),
    .Y(_133_)
);

FILL FILL88350x23550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__947_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[1]),
    .B(Xin[2]),
    .Y(_747_)
);

FILL FILL_1__1217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1094_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_699_),
    .B(_695_),
    .Y(_725_)
);

FILL FILL_0__841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__985_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_30_),
    .Y(_36_)
);

FILL FILL_1__1255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1324_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_517_),
    .B(_518_),
    .C(_520_),
    .Y(_521_)
);

FILL FILL_3__794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1202_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1551_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_753_[7]),
    .CLK(clk_bF$buf0),
    .Q(y[7])
);

INVX1 _1131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_319_),
    .Y(_320_)
);

FILL FILL_1__913_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_68_),
    .B(_21_),
    .C(_71_),
    .Y(_74_)
);

FILL FILL_1__1293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1011_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_120_),
    .B(_116_),
    .C(_81_),
    .Y(_130_)
);

FILL FILL_1__1349_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_499_),
    .B(_553_),
    .C(_549_),
    .Y(_563_)
);

FILL FILL_4__866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1097_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_571_),
    .B(_613_),
    .C(_609_),
    .Y(_622_)
);

FILL FILL_3__888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88650x39150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1227_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin_3_bF$buf3),
    .B(Cin[6]),
    .C(Xin[4]),
    .D(Cin[5]),
    .Y(_416_)
);

FILL FILL_0__973_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_161_),
    .Y(_167_)
);

FILL FILL_1__1387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1105_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_662_),
    .B(_661_),
    .C(_636_),
    .Y(_663_)
);

NAND2X1 _1034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[1]),
    .B(Cin[6]),
    .Y(_224_)
);

FILL FILL_0__782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__816_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_655_),
    .B(_687_),
    .C(_623_),
    .Y(_697_)
);

FILL FILL_1__1196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88950x78150 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_456_),
    .B(_455_),
    .Y(_457_)
);

FILL FILL_4__769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1074_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _1319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_502_),
    .B(_506_),
    .C(_505_),
    .Y(_518_)
);

FILL FILL_3__1563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1143_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[14]),
    .B(_576_),
    .C(_678_),
    .Y(_703_)
);

INVX1 _1072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_261_),
    .Y(_262_)
);

FILL FILL_1__854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1112_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1548_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_752_[4]),
    .CLK(clk_bF$buf3),
    .Q(y[4])
);

OAI21X1 _1128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_288_),
    .B(_316_),
    .C(_281_),
    .Y(_317_)
);

FILL FILL_0__876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1372_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_69_),
    .B(_70_),
    .C(_744_),
    .Y(_71_)
);

FILL FILL_2__1359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1008_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_468_),
    .B(_464_),
    .C(_412_),
    .Y(_560_)
);

FILL FILL_3__1181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1168_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[2]),
    .B(Cin[3]),
    .C(_91_),
    .Y(_92_)
);

FILL FILL_1__1311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88050x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[2]),
    .B(Xin[6]),
    .Y(_355_)
);

FILL FILL_1__948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1046_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert5 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf0)
);

NAND2X1 _1395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_598_),
    .B(_534_),
    .Y(_599_)
);

FILL FILL_1__757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88350x85950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__944_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_743_),
    .B(_601_),
    .Y(_744_)
);

FILL FILL_1__1214_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_695_),
    .B(_699_),
    .C(_634_),
    .D(_698_),
    .Y(_700_)
);

AOI21X1 _1069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf0),
    .B(Xin[6]),
    .C(Yin[6]),
    .Y(_259_)
);

FILL FILL_0__1109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1369_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_311_),
    .B(_494_),
    .C(_492_),
    .Y(_495_)
);

FILL FILL_2__1512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1091_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_721_),
    .B(_716_),
    .Y(_722_)
);

FILL FILL_3__982_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[1]),
    .B(Xin_3_bF$buf2),
    .Y(_33_)
);

FILL FILL_1__1252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__932_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_121_),
    .B(_126_),
    .C(_76_),
    .Y(_127_)
);

FILL FILL_1__1346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1415_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_552_),
    .B(_551_),
    .C(_500_),
    .Y(_619_)
);

FILL FILL_3__885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88650x15750 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin_3_bF$buf3),
    .B(Cin[6]),
    .Y(_413_)
);

FILL FILL_0__970_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[6]),
    .Y(_164_)
);

FILL FILL_1__1384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1102_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_637_),
    .B(_659_),
    .Y(_660_)
);

INVX1 _1031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_220_),
    .Y(_221_)
);

FILL FILL_1__813_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_655_),
    .Y(_666_)
);

FILL FILL_1__1193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1088_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[14]),
    .B(_677_),
    .C(_678_),
    .Y(_719_)
);

FILL FILL_0__835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1331_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf2),
    .B(Xin[4]),
    .C(Yin[4]),
    .Y(_30_)
);

FILL FILL_1__1249_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_453_),
    .B(_449_),
    .C(_452_),
    .Y(_454_)
);

FILL FILL_2__1318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL88950x54750 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_443_),
    .B(_513_),
    .C(_446_),
    .Y(_514_)
);

FILL FILL_3__788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1127_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1545_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_749_[1]),
    .CLK(clk_bF$buf4),
    .Q(y[1])
);

NAND2X1 _1125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_234_),
    .B(_240_),
    .Y(_314_)
);

FILL FILL_0__873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__907_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_26_),
    .B(_63_),
    .C(_67_),
    .Y(_68_)
);

FILL FILL_1__1287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1005_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_541_),
    .B(_547_),
    .C(_550_),
    .Y(_556_)
);

FILL FILL_1__1096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1234_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_755_[9]),
    .Y(Yout[9])
);

INVX1 _1163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[6]),
    .Y(_352_)
);

FILL FILL_1__945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1394_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_333_),
    .B(_340_),
    .Y(_410_)
);

FILL FILL_0__967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1043_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_591_),
    .B(_589_),
    .C(_536_),
    .Y(_596_)
);

FILL FILL_4__898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1519_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_656_),
    .B(_649_),
    .Y(_657_)
);

NAND2X1 _1028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_140_),
    .B(_78_),
    .Y(_218_)
);

FILL FILL_0__776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1272_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_623_),
    .Y(_633_)
);

FILL FILL_1__983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1341_ (
    .gnd(gnd),
    .vdd(vdd)
);

endmodule

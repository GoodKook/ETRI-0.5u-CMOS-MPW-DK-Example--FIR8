* NGSPICE file created from fir_pe.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL vdd gnd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 D CLK Q vdd gnd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A Y vdd gnd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D Y vdd gnd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A Y vdd gnd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D Y vdd gnd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B Y vdd gnd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B Y vdd gnd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A Y vdd gnd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A Y vdd gnd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C Y vdd gnd
.ends

.subckt fir_pe gnd vdd Cin[7] Cin[6] Cin[5] Cin[4] Cin[3] Cin[2] Cin[1] Cin[0] Xin[7]
+ Xin[6] Xin[5] Xin[4] Xin[3] Xin[2] Xin[1] Xin[0] Xout[7] Xout[6] Xout[5] Xout[4]
+ Xout[3] Xout[2] Xout[1] Xout[0] Yin[15] Yin[14] Yin[13] Yin[12] Yin[11] Yin[10]
+ Yin[9] Yin[8] Yin[7] Yin[6] Yin[5] Yin[4] Yin[3] Yin[2] Yin[1] Yin[0] Yout[15] Yout[14]
+ Yout[13] Yout[12] Yout[11] Yout[10] Yout[9] Yout[8] Yout[7] Yout[6] Yout[5] Yout[4]
+ Yout[3] Yout[2] Yout[1] Yout[0] clk
XFILL_3__1468_ vdd gnd FILL
XFILL_1__1104_ vdd gnd FILL
XFILL_2__992_ vdd gnd FILL
XFILL_3__1399_ vdd gnd FILL
XFILL_1__1035_ vdd gnd FILL
XFILL_2__1213_ vdd gnd FILL
XFILL_0__815_ vdd gnd FILL
XFILL_2__1144_ vdd gnd FILL
XFILL_2__1075_ vdd gnd FILL
XFILL_3__888_ vdd gnd FILL
XFILL_3__957_ vdd gnd FILL
X_1270_ _1301_/B _1280_/B _1303_/B vdd gnd NAND2X1
XFILL_3__1322_ vdd gnd FILL
XFILL_0__1475_ vdd gnd FILL
XFILL_3__1253_ vdd gnd FILL
XFILL_3__1184_ vdd gnd FILL
X_1537_ _1553_/Q _1551_/CLK _1583_/A vdd gnd DFFPOSX1
X_1399_ _1428_/B _1399_/B _1399_/C _1430_/A vdd gnd NAND3X1
X_1468_ _1468_/A _1470_/B _1507_/C vdd gnd NOR2X1
XFILL_2__975_ vdd gnd FILL
XFILL_3__811_ vdd gnd FILL
X_981_ _986_/A _987_/C vdd gnd INVX1
XFILL_1__1018_ vdd gnd FILL
XFILL88350x54750 vdd gnd FILL
XFILL_0__1260_ vdd gnd FILL
XFILL_2__1127_ vdd gnd FILL
XFILL_2__1058_ vdd gnd FILL
XFILL_0__1191_ vdd gnd FILL
XFILL_1__993_ vdd gnd FILL
X_1322_ _1326_/A _1326_/B _1325_/C _1323_/C vdd gnd OAI21X1
X_1253_ Xin[7] _1468_/A vdd gnd INVX1
XFILL_3__1236_ vdd gnd FILL
XFILL_3__1305_ vdd gnd FILL
X_1184_ _1188_/A _1188_/B _1248_/C _1266_/B _1195_/B vdd gnd AOI22X1
XFILL_2__760_ vdd gnd FILL
XFILL_3__1098_ vdd gnd FILL
XFILL_0__1458_ vdd gnd FILL
XFILL_0__1389_ vdd gnd FILL
XFILL_3__1167_ vdd gnd FILL
XFILL_4__1345_ vdd gnd FILL
XFILL_4__1414_ vdd gnd FILL
XFILL_1__1567_ vdd gnd FILL
XFILL_4__1276_ vdd gnd FILL
XFILL_1__1498_ vdd gnd FILL
XFILL_2__889_ vdd gnd FILL
XFILL_2__958_ vdd gnd FILL
X_964_ _964_/A _964_/B _964_/C _966_/B vdd gnd OAI21X1
X_895_ _895_/A _965_/A vdd gnd INVX1
XFILL_3__1021_ vdd gnd FILL
XFILL_0__1174_ vdd gnd FILL
XFILL_0__1312_ vdd gnd FILL
XFILL_0__1243_ vdd gnd FILL
XFILL_1__976_ vdd gnd FILL
X_1236_ _1243_/A _1243_/C _1244_/C _1301_/A vdd gnd NAND3X1
X_1305_ _1305_/A Cin[7] _1371_/A vdd gnd NAND2X1
X_1098_ _1125_/B _1098_/B _1128_/A vdd gnd NAND2X1
XFILL_3__1219_ vdd gnd FILL
XFILL_1__1352_ vdd gnd FILL
XFILL_1__1421_ vdd gnd FILL
XFILL_1__1283_ vdd gnd FILL
X_1167_ Cin[3] _1249_/A _1234_/B _1169_/B vdd gnd NAND3X1
XFILL_2__812_ vdd gnd FILL
XFILL_2__1461_ vdd gnd FILL
XFILL_2__1392_ vdd gnd FILL
XFILL_0__994_ vdd gnd FILL
XFILL88350x78150 vdd gnd FILL
X_947_ _947_/A _947_/B _947_/C _948_/B vdd gnd AOI21X1
XFILL_1__830_ vdd gnd FILL
X_878_ _878_/A _878_/B _878_/C _884_/B vdd gnd AOI21X1
XFILL_1__761_ vdd gnd FILL
XFILL_3__1570_ vdd gnd FILL
XFILL_4__972_ vdd gnd FILL
X_1021_ _1121_/B _1122_/D _1119_/A vdd gnd NAND2X1
XFILL_3__1004_ vdd gnd FILL
XFILL_0__1157_ vdd gnd FILL
XFILL_0__1226_ vdd gnd FILL
XFILL_0__1088_ vdd gnd FILL
XFILL_1__959_ vdd gnd FILL
X_1219_ _1219_/A _1219_/B _1300_/A vdd gnd NAND2X1
XFILL_1__1404_ vdd gnd FILL
XFILL_1__1335_ vdd gnd FILL
XFILL_1__1266_ vdd gnd FILL
XFILL_3__990_ vdd gnd FILL
XFILL_1__1197_ vdd gnd FILL
X_801_ _886_/A _965_/B _888_/A _823_/C vdd gnd OAI21X1
XFILL_2__1513_ vdd gnd FILL
XFILL_2__1375_ vdd gnd FILL
XFILL_2__1444_ vdd gnd FILL
XFILL_0__977_ vdd gnd FILL
XFILL_0__1011_ vdd gnd FILL
X_1570_ _1570_/A Yout[10] vdd gnd BUFX2
XFILL_1__813_ vdd gnd FILL
XFILL_3__1484_ vdd gnd FILL
X_1004_ _997_/Y _998_/Y _999_/Y _1022_/A vdd gnd NAND3X1
XFILL_1__1120_ vdd gnd FILL
XFILL_0__1209_ vdd gnd FILL
XFILL_1__1051_ vdd gnd FILL
XFILL_2__1160_ vdd gnd FILL
XFILL_0__831_ vdd gnd FILL
XFILL_0__900_ vdd gnd FILL
XFILL_0__762_ vdd gnd FILL
XFILL_2__1091_ vdd gnd FILL
XFILL_1__1249_ vdd gnd FILL
XFILL_1__1318_ vdd gnd FILL
XFILL_3__973_ vdd gnd FILL
XFILL_0__1560_ vdd gnd FILL
XFILL_2__1289_ vdd gnd FILL
XFILL_0__1491_ vdd gnd FILL
XFILL_2__1427_ vdd gnd FILL
XFILL_2__1358_ vdd gnd FILL
XFILL_1_CLKBUF1_insert0 vdd gnd FILL
X_1553_ _1553_/D _1557_/CLK _1553_/Q vdd gnd DFFPOSX1
XFILL_2_BUFX2_insert14 vdd gnd FILL
X_1484_ _1484_/A _1486_/C _1557_/D vdd gnd XOR2X1
XFILL_3__1467_ vdd gnd FILL
XFILL_3__1398_ vdd gnd FILL
XFILL_1__1103_ vdd gnd FILL
XFILL_2__991_ vdd gnd FILL
XFILL_1__1034_ vdd gnd FILL
XFILL_2__1143_ vdd gnd FILL
XFILL_2__1212_ vdd gnd FILL
XFILL_0__814_ vdd gnd FILL
XFILL_2__1074_ vdd gnd FILL
XFILL_3__956_ vdd gnd FILL
XFILL_3__887_ vdd gnd FILL
XFILL_3__1252_ vdd gnd FILL
XFILL_3__1321_ vdd gnd FILL
XFILL_0__1474_ vdd gnd FILL
XFILL_3__1183_ vdd gnd FILL
X_1536_ _1552_/Q _1552_/CLK _1582_/A vdd gnd DFFPOSX1
XFILL_1__1583_ vdd gnd FILL
X_1467_ _1492_/B _1507_/B vdd gnd INVX1
X_1398_ _1402_/C _1399_/C vdd gnd INVX1
XFILL_3__1519_ vdd gnd FILL
XFILL_2__974_ vdd gnd FILL
XFILL_1__1017_ vdd gnd FILL
XFILL_3__810_ vdd gnd FILL
X_980_ _987_/A _987_/B _986_/A _994_/B vdd gnd OAI21X1
XFILL_2__1126_ vdd gnd FILL
XFILL_0__1190_ vdd gnd FILL
XFILL_2__1057_ vdd gnd FILL
XFILL_3__939_ vdd gnd FILL
XFILL_1__992_ vdd gnd FILL
X_1252_ _1336_/A _1320_/B _1316_/C vdd gnd NAND2X1
X_1321_ _1321_/A _1321_/B _1321_/C _1325_/C vdd gnd AOI21X1
XFILL_3__1235_ vdd gnd FILL
XFILL_0__1457_ vdd gnd FILL
X_1183_ _1265_/A _1265_/B _1265_/C _1266_/B vdd gnd NAND3X1
XFILL_3__1304_ vdd gnd FILL
XFILL_3__1097_ vdd gnd FILL
XFILL_0__1388_ vdd gnd FILL
XFILL_3__1166_ vdd gnd FILL
X_1519_ _1519_/A _941_/C _1548_/D vdd gnd XOR2X1
XFILL_1__1566_ vdd gnd FILL
XFILL_2__957_ vdd gnd FILL
XFILL_1__1497_ vdd gnd FILL
XFILL_2__888_ vdd gnd FILL
XFILL88950x15750 vdd gnd FILL
X_963_ _963_/A _963_/B _963_/C _992_/B vdd gnd NAND3X1
X_894_ _894_/A _964_/C _897_/C vdd gnd NAND2X1
XFILL_3__1020_ vdd gnd FILL
XFILL_0__1311_ vdd gnd FILL
XFILL_2__1109_ vdd gnd FILL
XFILL_0__1242_ vdd gnd FILL
XFILL_0__1173_ vdd gnd FILL
XFILL_1__975_ vdd gnd FILL
X_1235_ _1235_/A _1235_/B _1235_/C _1244_/C vdd gnd OAI21X1
XFILL_1__1420_ vdd gnd FILL
X_1304_ _1304_/A _1304_/B _1304_/C _1324_/A vdd gnd OAI21X1
X_1166_ Cin[2] Xin[6] _1234_/B vdd gnd NAND2X1
XFILL_2__811_ vdd gnd FILL
X_1097_ _1198_/A _1199_/B _1199_/A _1208_/A vdd gnd NAND3X1
XFILL_3__1149_ vdd gnd FILL
XFILL_3__1218_ vdd gnd FILL
XFILL_4__1060_ vdd gnd FILL
XFILL_1__1351_ vdd gnd FILL
XFILL_0__1509_ vdd gnd FILL
XFILL_1__1282_ vdd gnd FILL
XFILL_2__1460_ vdd gnd FILL
XFILL_2__1391_ vdd gnd FILL
XFILL_4__1327_ vdd gnd FILL
XFILL_4__1258_ vdd gnd FILL
XFILL_0__993_ vdd gnd FILL
XFILL_4__1189_ vdd gnd FILL
XFILL88950x27450 vdd gnd FILL
X_1020_ _1020_/A _1020_/B _1550_/D vdd gnd NOR2X1
X_877_ _877_/A _877_/B _877_/C _877_/D _936_/C vdd gnd AOI22X1
X_946_ _951_/A _946_/B _946_/Y vdd gnd NAND2X1
XFILL_1__760_ vdd gnd FILL
XFILL_3__1003_ vdd gnd FILL
XFILL_0__1087_ vdd gnd FILL
XFILL_0__1156_ vdd gnd FILL
XFILL_0__1225_ vdd gnd FILL
XFILL_1__889_ vdd gnd FILL
X_1149_ _965_/C _1149_/B _1149_/C _1149_/D _1153_/B vdd gnd AOI22X1
XFILL_1__958_ vdd gnd FILL
X_1218_ _1218_/A _1218_/B _1288_/A _1287_/A vdd gnd OAI21X1
XFILL_1__1403_ vdd gnd FILL
XFILL_1__1196_ vdd gnd FILL
XFILL_1__1334_ vdd gnd FILL
XFILL_1__1265_ vdd gnd FILL
X_800_ Xin[1] Cin[2] _888_/A vdd gnd NAND2X1
XFILL88950x39150 vdd gnd FILL
XFILL_2__1512_ vdd gnd FILL
XFILL_2__1374_ vdd gnd FILL
XFILL_2__1443_ vdd gnd FILL
XFILL_0__976_ vdd gnd FILL
XFILL_0__1010_ vdd gnd FILL
XFILL_1__812_ vdd gnd FILL
X_1003_ _938_/C _938_/A _1003_/C _1010_/C vdd gnd AOI21X1
X_929_ _938_/C _948_/C _938_/A _935_/A vdd gnd NAND3X1
XFILL_3__1483_ vdd gnd FILL
XFILL_1__1050_ vdd gnd FILL
XFILL_0__1208_ vdd gnd FILL
XFILL_0__1139_ vdd gnd FILL
XFILL_1__1317_ vdd gnd FILL
XFILL_0__830_ vdd gnd FILL
XFILL_0__761_ vdd gnd FILL
XFILL_2__1090_ vdd gnd FILL
XFILL_1__1248_ vdd gnd FILL
XFILL_1__1179_ vdd gnd FILL
XFILL_3__972_ vdd gnd FILL
XFILL_0__1490_ vdd gnd FILL
XFILL_2__1426_ vdd gnd FILL
XFILL_1_CLKBUF1_insert1 vdd gnd FILL
XFILL_2__1288_ vdd gnd FILL
XFILL_2__1357_ vdd gnd FILL
XFILL_2_BUFX2_insert15 vdd gnd FILL
XFILL_0__959_ vdd gnd FILL
X_1552_ _1552_/D _1552_/CLK _1552_/Q vdd gnd DFFPOSX1
X_1483_ _1488_/B _1488_/A _1486_/C vdd gnd XOR2X1
XFILL_2__990_ vdd gnd FILL
XFILL_3__1466_ vdd gnd FILL
XFILL_3__1397_ vdd gnd FILL
XFILL_1__1102_ vdd gnd FILL
XFILL_1__1033_ vdd gnd FILL
XFILL_4__1009_ vdd gnd FILL
XFILL_2__1142_ vdd gnd FILL
XFILL_2__1211_ vdd gnd FILL
XFILL_2__1073_ vdd gnd FILL
XFILL_0__813_ vdd gnd FILL
XFILL_3__955_ vdd gnd FILL
XFILL_3__886_ vdd gnd FILL
XFILL_2__1409_ vdd gnd FILL
XFILL_0__1473_ vdd gnd FILL
XFILL_3__1320_ vdd gnd FILL
XFILL_3__1251_ vdd gnd FILL
XFILL_3__1182_ vdd gnd FILL
X_1535_ _1551_/Q _1551_/CLK _1581_/A vdd gnd DFFPOSX1
XFILL_3__1518_ vdd gnd FILL
X_1466_ _1466_/A _1470_/C _1466_/C _1466_/D _1497_/A vdd gnd OAI22X1
XFILL_1__1582_ vdd gnd FILL
X_1397_ _1397_/A _1430_/B _1402_/C vdd gnd NAND2X1
XFILL_2__973_ vdd gnd FILL
XFILL_3__1449_ vdd gnd FILL
XFILL_1__1016_ vdd gnd FILL
XFILL_2__1056_ vdd gnd FILL
XFILL_2__1125_ vdd gnd FILL
X_1320_ _1336_/A _1320_/B _1321_/C vdd gnd AND2X2
XFILL_1__991_ vdd gnd FILL
XFILL_3__938_ vdd gnd FILL
XFILL_3__869_ vdd gnd FILL
X_1251_ Cin[2] Xin[7] _1320_/B vdd gnd AND2X2
X_1182_ _1259_/A _1182_/B _1265_/C vdd gnd NAND2X1
XFILL_3__1303_ vdd gnd FILL
XFILL_0__1456_ vdd gnd FILL
XFILL_3__1165_ vdd gnd FILL
XFILL_3__1234_ vdd gnd FILL
XFILL_3__1096_ vdd gnd FILL
XFILL_0__1387_ vdd gnd FILL
X_1518_ _828_/A _828_/B _833_/A _1519_/A vdd gnd OAI21X1
X_1449_ _1449_/A _1481_/A _1449_/C _1450_/A vdd gnd OAI21X1
XFILL_1__1565_ vdd gnd FILL
XFILL_1__1496_ vdd gnd FILL
XFILL_2__956_ vdd gnd FILL
XFILL_2__887_ vdd gnd FILL
X_962_ _964_/A _964_/B _962_/C _963_/A vdd gnd OAI21X1
X_893_ _895_/A Cin[3] _964_/C vdd gnd AND2X2
XFILL_0__1310_ vdd gnd FILL
XFILL_0__1241_ vdd gnd FILL
XFILL_2__1108_ vdd gnd FILL
XFILL_2__1039_ vdd gnd FILL
XFILL_0__1172_ vdd gnd FILL
XFILL_1__974_ vdd gnd FILL
X_1303_ _1303_/A _1303_/B _1303_/C _1413_/C vdd gnd OAI21X1
X_1096_ _1099_/B _1099_/A _1100_/C _1199_/B vdd gnd OAI21X1
XFILL_1__1350_ vdd gnd FILL
X_1165_ _1239_/C _1239_/D _1235_/C _1188_/A vdd gnd NAND3X1
X_1234_ _1234_/A _1234_/B _1235_/B vdd gnd AND2X2
XFILL_2__810_ vdd gnd FILL
XFILL_3__1148_ vdd gnd FILL
XFILL_3__1217_ vdd gnd FILL
XFILL_0__1439_ vdd gnd FILL
XFILL_0__1508_ vdd gnd FILL
XFILL_1__1281_ vdd gnd FILL
XFILL_3__1079_ vdd gnd FILL
XFILL89250x74250 vdd gnd FILL
XFILL_1__1479_ vdd gnd FILL
XFILL_2__1390_ vdd gnd FILL
XFILL_2__939_ vdd gnd FILL
XFILL_0__992_ vdd gnd FILL
X_945_ _945_/A _945_/B _945_/C _945_/Y vdd gnd OAI21X1
X_876_ _936_/B _884_/C _936_/A _882_/A vdd gnd NAND3X1
XFILL_3__1002_ vdd gnd FILL
XFILL_0__1224_ vdd gnd FILL
XFILL_0__1086_ vdd gnd FILL
XFILL_0__1155_ vdd gnd FILL
XFILL_1__957_ vdd gnd FILL
XFILL_1__888_ vdd gnd FILL
X_1148_ _1234_/A _1149_/B vdd gnd INVX1
X_1079_ _1171_/A Xin[7] _1079_/C _1083_/A vdd gnd NAND3X1
X_1217_ _1217_/A _1217_/B _1217_/C _1218_/B vdd gnd AOI21X1
XFILL_1__1402_ vdd gnd FILL
XFILL_1__1333_ vdd gnd FILL
XFILL_1__1195_ vdd gnd FILL
XFILL_1__1264_ vdd gnd FILL
XFILL_2__1442_ vdd gnd FILL
XFILL_2__1511_ vdd gnd FILL
XFILL_2__1373_ vdd gnd FILL
XFILL_4__1309_ vdd gnd FILL
XFILL_0__975_ vdd gnd FILL
XFILL_1__811_ vdd gnd FILL
X_928_ _932_/A _932_/B _933_/C _938_/A vdd gnd OAI21X1
X_1002_ _948_/C _1003_/C vdd gnd INVX1
XFILL_4__953_ vdd gnd FILL
X_859_ Xin[1] _860_/A vdd gnd INVX1
XFILL_3__1482_ vdd gnd FILL
XFILL_4__884_ vdd gnd FILL
XFILL_0__1207_ vdd gnd FILL
XFILL88950x150 vdd gnd FILL
XFILL_0__1069_ vdd gnd FILL
XFILL_0__1138_ vdd gnd FILL
XFILL_1__1316_ vdd gnd FILL
XFILL_0__760_ vdd gnd FILL
XFILL_1__1247_ vdd gnd FILL
XFILL_1__1178_ vdd gnd FILL
XFILL_3__971_ vdd gnd FILL
XFILL_2__1425_ vdd gnd FILL
XFILL_2__1356_ vdd gnd FILL
XFILL_1_CLKBUF1_insert2 vdd gnd FILL
XFILL_0__958_ vdd gnd FILL
XFILL_2__1287_ vdd gnd FILL
X_1551_ _1551_/D _1551_/CLK _1551_/Q vdd gnd DFFPOSX1
XFILL_0__889_ vdd gnd FILL
XFILL_2_BUFX2_insert16 vdd gnd FILL
X_1482_ _1490_/A _1482_/B _1488_/B vdd gnd NAND2X1
XFILL_3__1465_ vdd gnd FILL
XFILL_1__1101_ vdd gnd FILL
XFILL_3__1396_ vdd gnd FILL
XFILL_1__1032_ vdd gnd FILL
XFILL_4__1574_ vdd gnd FILL
XFILL_2__1210_ vdd gnd FILL
XFILL_0__812_ vdd gnd FILL
XFILL_2__1141_ vdd gnd FILL
XFILL_2__1072_ vdd gnd FILL
XFILL_3__954_ vdd gnd FILL
XFILL_3__885_ vdd gnd FILL
XFILL_3__1181_ vdd gnd FILL
XFILL_2__1339_ vdd gnd FILL
XFILL_2__1408_ vdd gnd FILL
XFILL_3__1250_ vdd gnd FILL
XFILL_0__1472_ vdd gnd FILL
X_1534_ _1550_/Q _1551_/CLK _1580_/A vdd gnd DFFPOSX1
X_1465_ _1465_/A _1465_/B _1465_/C _1488_/A vdd gnd AOI21X1
XFILL_1__1581_ vdd gnd FILL
X_1396_ _1396_/A _1396_/B _1430_/B vdd gnd OR2X2
XFILL_3__1448_ vdd gnd FILL
XFILL_3__1517_ vdd gnd FILL
XFILL_4__1290_ vdd gnd FILL
XFILL_2__972_ vdd gnd FILL
XFILL_3__1379_ vdd gnd FILL
XFILL_1__1015_ vdd gnd FILL
XFILL_4__1488_ vdd gnd FILL
XFILL_2__1055_ vdd gnd FILL
XFILL_2__1124_ vdd gnd FILL
XFILL_1__990_ vdd gnd FILL
X_1181_ _1181_/A _1182_/B vdd gnd INVX1
XFILL_3__937_ vdd gnd FILL
XFILL_3__868_ vdd gnd FILL
XFILL_3__1302_ vdd gnd FILL
X_1250_ _1316_/A _1321_/A vdd gnd INVX1
XFILL_3__799_ vdd gnd FILL
XFILL_3__1095_ vdd gnd FILL
XFILL_3__1233_ vdd gnd FILL
XFILL_0__1455_ vdd gnd FILL
XFILL_0__1386_ vdd gnd FILL
XFILL_3__1164_ vdd gnd FILL
X_1448_ _1448_/A _1448_/B _1478_/C vdd gnd NAND2X1
X_1517_ _1517_/A _1517_/B _1559_/D vdd gnd NAND2X1
XFILL89550x46950 vdd gnd FILL
XFILL_1__1564_ vdd gnd FILL
XFILL_1__1495_ vdd gnd FILL
X_1379_ Xin[4] Cin[7] _1431_/A vdd gnd NAND2X1
XFILL_2__955_ vdd gnd FILL
XFILL_2__886_ vdd gnd FILL
X_961_ _961_/A Cin[3] _962_/C vdd gnd NAND2X1
X_892_ _901_/A _897_/A vdd gnd INVX1
XFILL_0__1240_ vdd gnd FILL
XFILL_2__1107_ vdd gnd FILL
XFILL_2__1038_ vdd gnd FILL
XFILL_0__1171_ vdd gnd FILL
XFILL_1__973_ vdd gnd FILL
X_1233_ _1237_/C _1237_/B _1304_/C _1243_/A vdd gnd NAND3X1
X_1302_ _1366_/A _1414_/A vdd gnd INVX1
X_1095_ _1095_/A _1095_/B _1187_/B _1186_/A _1099_/A vdd gnd AOI22X1
XFILL_1__1280_ vdd gnd FILL
XFILL_0__1507_ vdd gnd FILL
X_1164_ _964_/A _1470_/A _1234_/A _1239_/C vdd gnd OAI21X1
XFILL_3__1078_ vdd gnd FILL
XFILL_3__1216_ vdd gnd FILL
XFILL_3__1147_ vdd gnd FILL
XFILL_0__1369_ vdd gnd FILL
XFILL_0__1438_ vdd gnd FILL
XFILL89550x58650 vdd gnd FILL
XFILL_0__991_ vdd gnd FILL
XFILL_1__1478_ vdd gnd FILL
XFILL_2__938_ vdd gnd FILL
XFILL_2__869_ vdd gnd FILL
X_944_ _944_/A _945_/A _944_/Y vdd gnd XOR2X1
X_875_ _877_/C _877_/D _875_/C _936_/A vdd gnd NAND3X1
XFILL_3__1001_ vdd gnd FILL
XFILL_0__1154_ vdd gnd FILL
XFILL_0__1223_ vdd gnd FILL
XFILL_0__1085_ vdd gnd FILL
XFILL_1__956_ vdd gnd FILL
XFILL_1__887_ vdd gnd FILL
X_1216_ _1297_/A _1216_/B _1296_/A _1294_/A vdd gnd OAI21X1
XFILL_4__1110_ vdd gnd FILL
XFILL_4__1041_ vdd gnd FILL
X_1078_ Yin[7] _1078_/B _1083_/B vdd gnd NAND2X1
X_1147_ Cin[3] _1249_/A _1234_/A vdd gnd NAND2X1
XFILL_1__1401_ vdd gnd FILL
XFILL_1__1263_ vdd gnd FILL
XFILL_1__1332_ vdd gnd FILL
XFILL_1__1194_ vdd gnd FILL
XFILL_2__1441_ vdd gnd FILL
XFILL_2__1510_ vdd gnd FILL
XFILL_2__1372_ vdd gnd FILL
XFILL_0__974_ vdd gnd FILL
XFILL_4__1239_ vdd gnd FILL
XFILL_1__810_ vdd gnd FILL
X_927_ _952_/C _927_/B _991_/B _990_/A _932_/A vdd gnd AOI22X1
X_858_ _868_/A _867_/B vdd gnd INVX1
XFILL_3__1481_ vdd gnd FILL
X_1001_ _1010_/B _996_/Y _948_/Y _1015_/B vdd gnd OAI21X1
X_789_ _803_/B _797_/C _789_/C _795_/A vdd gnd NAND3X1
XFILL_0__1206_ vdd gnd FILL
XFILL_0__1137_ vdd gnd FILL
XFILL_0__1068_ vdd gnd FILL
XFILL_1__939_ vdd gnd FILL
XFILL_1__1246_ vdd gnd FILL
XFILL_1__1315_ vdd gnd FILL
XFILL_1__1177_ vdd gnd FILL
XFILL_3__970_ vdd gnd FILL
XFILL_2__1424_ vdd gnd FILL
XFILL_2__1355_ vdd gnd FILL
XFILL_0__957_ vdd gnd FILL
XFILL_1_CLKBUF1_insert3 vdd gnd FILL
XFILL_2__1286_ vdd gnd FILL
XFILL_2_BUFX2_insert17 vdd gnd FILL
X_1550_ _1550_/D _1551_/CLK _1550_/Q vdd gnd DFFPOSX1
XFILL_0__888_ vdd gnd FILL
X_1481_ _1481_/A _1481_/B _1481_/C _1490_/A vdd gnd NAND3X1
XFILL_3__1464_ vdd gnd FILL
XFILL_4__866_ vdd gnd FILL
XFILL_4__935_ vdd gnd FILL
XFILL_1__1100_ vdd gnd FILL
XFILL_3__1395_ vdd gnd FILL
XFILL_4__797_ vdd gnd FILL
XFILL_1__1031_ vdd gnd FILL
XFILL_2__1140_ vdd gnd FILL
XFILL_0__811_ vdd gnd FILL
XFILL_2__1071_ vdd gnd FILL
XFILL_1__1229_ vdd gnd FILL
XFILL_3__953_ vdd gnd FILL
XFILL88350x74250 vdd gnd FILL
XFILL_3__884_ vdd gnd FILL
XFILL_2__1338_ vdd gnd FILL
XFILL_2__1407_ vdd gnd FILL
XFILL_2__1269_ vdd gnd FILL
XFILL_3__1180_ vdd gnd FILL
XFILL_0__1471_ vdd gnd FILL
X_1533_ _1549_/Q _1549_/CLK _1579_/A vdd gnd DFFPOSX1
X_1395_ _1396_/B _1396_/A _1397_/A vdd gnd NAND2X1
X_1464_ _1464_/A _1464_/B _1488_/C _1484_/A vdd gnd OAI21X1
XFILL_1__1580_ vdd gnd FILL
XFILL_3__1447_ vdd gnd FILL
XFILL_3__1516_ vdd gnd FILL
XFILL_3__1378_ vdd gnd FILL
XFILL_2__971_ vdd gnd FILL
XFILL_1__1014_ vdd gnd FILL
XFILL_2__1123_ vdd gnd FILL
XFILL_2__1054_ vdd gnd FILL
XFILL_3__936_ vdd gnd FILL
XFILL_3__798_ vdd gnd FILL
XFILL_3__867_ vdd gnd FILL
XFILL_3__1232_ vdd gnd FILL
X_1180_ _1247_/A _1247_/B _1248_/C vdd gnd NAND2X1
XFILL_3__1301_ vdd gnd FILL
XFILL_3__1094_ vdd gnd FILL
XFILL_0__1454_ vdd gnd FILL
XFILL_0__1385_ vdd gnd FILL
XFILL_3__1163_ vdd gnd FILL
X_1516_ _1516_/A _1516_/B _1516_/C _1517_/A vdd gnd NAND3X1
XFILL_4__1341_ vdd gnd FILL
XFILL_4__1410_ vdd gnd FILL
X_1447_ _1449_/C _1448_/A vdd gnd INVX1
X_1378_ _964_/B _1470_/B _1431_/B _1391_/B vdd gnd OAI21X1
XFILL_1__1563_ vdd gnd FILL
XFILL_4__1272_ vdd gnd FILL
XFILL_1__1494_ vdd gnd FILL
XFILL_2__954_ vdd gnd FILL
XFILL_2__885_ vdd gnd FILL
X_891_ Xin[1] Cin[4] _901_/A vdd gnd NAND2X1
X_960_ Xin[4] _964_/B vdd gnd INVX2
XFILL_2__1106_ vdd gnd FILL
XFILL_0__1170_ vdd gnd FILL
XFILL_2__1037_ vdd gnd FILL
XFILL88350x4050 vdd gnd FILL
XFILL_1__972_ vdd gnd FILL
XFILL_3__919_ vdd gnd FILL
X_1232_ _1232_/A _1312_/A _1304_/C vdd gnd NAND2X1
X_1301_ _1301_/A _1301_/B _1366_/A vdd gnd NAND2X1
X_1094_ _1094_/A _1094_/B _1158_/B _1099_/B vdd gnd AOI21X1
XFILL_3__1215_ vdd gnd FILL
XFILL_0__1437_ vdd gnd FILL
XFILL_0__1506_ vdd gnd FILL
X_1163_ Xin[6] _1470_/A vdd gnd INVX1
XFILL_3__1077_ vdd gnd FILL
XFILL_3__1146_ vdd gnd FILL
XFILL_0__1368_ vdd gnd FILL
XFILL_0__1299_ vdd gnd FILL
XFILL_0__990_ vdd gnd FILL
XFILL_2__937_ vdd gnd FILL
XFILL_1__1477_ vdd gnd FILL
XFILL_2__868_ vdd gnd FILL
XFILL_2__799_ vdd gnd FILL
X_943_ _945_/C _943_/B _944_/A vdd gnd NAND2X1
X_874_ _890_/C _890_/A _925_/A _877_/D vdd gnd NAND3X1
XFILL_3__1000_ vdd gnd FILL
XFILL_0__1153_ vdd gnd FILL
XFILL_0__1084_ vdd gnd FILL
XFILL_0__1222_ vdd gnd FILL
XFILL_1__955_ vdd gnd FILL
XFILL_1__886_ vdd gnd FILL
X_1146_ _1242_/B _1146_/B _1146_/C _1154_/A vdd gnd AOI21X1
X_1215_ _1422_/B _1216_/B vdd gnd INVX1
XFILL_1__1400_ vdd gnd FILL
XFILL_3__1129_ vdd gnd FILL
X_1077_ _1265_/A _1084_/C _1084_/A _1265_/B vdd gnd NAND3X1
XFILL_1__1193_ vdd gnd FILL
XFILL_1__1262_ vdd gnd FILL
XFILL_1__1331_ vdd gnd FILL
XFILL_2__1440_ vdd gnd FILL
XFILL_2__1371_ vdd gnd FILL
XFILL_0__973_ vdd gnd FILL
X_926_ _926_/A _926_/B _955_/A _932_/B vdd gnd AOI21X1
X_1000_ _999_/Y _998_/Y _997_/Y _1010_/B vdd gnd AOI21X1
X_788_ _797_/B _789_/C vdd gnd INVX1
X_857_ _868_/A _867_/A _867_/C _863_/A vdd gnd NAND3X1
XFILL_3__1480_ vdd gnd FILL
XFILL_2__1569_ vdd gnd FILL
XFILL_0__1067_ vdd gnd FILL
XFILL_0__1136_ vdd gnd FILL
XFILL_0__1205_ vdd gnd FILL
XFILL_1__938_ vdd gnd FILL
XFILL_1__869_ vdd gnd FILL
X_1129_ _1129_/A _1223_/A _1152_/A _1151_/A vdd gnd OAI21X1
XFILL_4__1023_ vdd gnd FILL
XFILL_1__1245_ vdd gnd FILL
XFILL_1__1314_ vdd gnd FILL
XFILL_1__1176_ vdd gnd FILL
XFILL_2__1354_ vdd gnd FILL
XFILL_2__1423_ vdd gnd FILL
XFILL_2__1285_ vdd gnd FILL
XFILL_0__956_ vdd gnd FILL
XFILL_0__887_ vdd gnd FILL
XFILL_1_CLKBUF1_insert4 vdd gnd FILL
X_1480_ _1480_/A _1480_/B _1481_/C vdd gnd NAND2X1
X_909_ _912_/C _911_/B _917_/A vdd gnd NAND2X1
XFILL_3__1394_ vdd gnd FILL
XFILL_3__1463_ vdd gnd FILL
XFILL_1__1030_ vdd gnd FILL
XFILL_0__1119_ vdd gnd FILL
XFILL_0__810_ vdd gnd FILL
XFILL_2__1070_ vdd gnd FILL
XFILL_1__1159_ vdd gnd FILL
XFILL_1__1228_ vdd gnd FILL
XFILL88950x23550 vdd gnd FILL
XFILL_3__883_ vdd gnd FILL
XFILL_3__952_ vdd gnd FILL
XFILL88650x58650 vdd gnd FILL
XFILL_2__1406_ vdd gnd FILL
XFILL_0__1470_ vdd gnd FILL
XFILL_4_BUFX2_insert8 vdd gnd FILL
XFILL_2__1268_ vdd gnd FILL
XFILL_2__1337_ vdd gnd FILL
X_1532_ _1548_/Q _1549_/CLK _1578_/A vdd gnd DFFPOSX1
XFILL_0__939_ vdd gnd FILL
XFILL_2__1199_ vdd gnd FILL
X_1394_ _1443_/B Yin[11] _1396_/B vdd gnd XNOR2X1
X_1463_ _1489_/C _1464_/B vdd gnd INVX1
XFILL_3__1515_ vdd gnd FILL
XFILL_2__970_ vdd gnd FILL
XFILL_3__1446_ vdd gnd FILL
XFILL_3__1377_ vdd gnd FILL
XFILL_4__917_ vdd gnd FILL
XFILL_4__848_ vdd gnd FILL
XFILL_1__1013_ vdd gnd FILL
XFILL_2__1122_ vdd gnd FILL
XFILL_2__1053_ vdd gnd FILL
XFILL88950x35250 vdd gnd FILL
XFILL_3__866_ vdd gnd FILL
XFILL_3__935_ vdd gnd FILL
XFILL_3__797_ vdd gnd FILL
XFILL_3__1231_ vdd gnd FILL
XFILL_0__1453_ vdd gnd FILL
XFILL_3__1300_ vdd gnd FILL
XFILL_3__1162_ vdd gnd FILL
XFILL_3__1093_ vdd gnd FILL
XFILL_0__1384_ vdd gnd FILL
X_1515_ _1515_/A _1516_/B vdd gnd INVX1
XFILL_1__1562_ vdd gnd FILL
X_1446_ _1446_/A _1476_/A _1449_/C vdd gnd NAND2X1
X_1377_ _1381_/A _1492_/B _1386_/B _1431_/B vdd gnd OAI21X1
XFILL_2__953_ vdd gnd FILL
XFILL_3__1429_ vdd gnd FILL
XFILL_1__1493_ vdd gnd FILL
XFILL_2__884_ vdd gnd FILL
X_890_ _890_/A _890_/B _890_/C _947_/C vdd gnd OAI21X1
XFILL_2__1105_ vdd gnd FILL
XFILL_2__1036_ vdd gnd FILL
XFILL_1__971_ vdd gnd FILL
XFILL_3__918_ vdd gnd FILL
XFILL_3__849_ vdd gnd FILL
X_1231_ Xin[4] Cin[6] _1312_/A vdd gnd AND2X2
X_1300_ _1300_/A _1300_/B _1300_/C _1356_/C vdd gnd AOI21X1
X_1162_ _1239_/A _1336_/A _1235_/C vdd gnd NAND2X1
X_1093_ _993_/C _993_/B _1093_/C _1100_/C vdd gnd AOI21X1
XFILL_3__1145_ vdd gnd FILL
XFILL_3__1214_ vdd gnd FILL
XFILL_0__1436_ vdd gnd FILL
XFILL_0__1505_ vdd gnd FILL
XFILL_3__1076_ vdd gnd FILL
XFILL_0__1367_ vdd gnd FILL
XFILL_0__1298_ vdd gnd FILL
X_1429_ _1465_/A _1454_/C vdd gnd INVX1
XFILL_1__1476_ vdd gnd FILL
XFILL_2__936_ vdd gnd FILL
XFILL_2__798_ vdd gnd FILL
XFILL_2__867_ vdd gnd FILL
X_942_ _945_/B _943_/B vdd gnd INVX1
X_873_ _925_/C _890_/B _925_/B _877_/C vdd gnd OAI21X1
XFILL_0__1221_ vdd gnd FILL
XFILL_2__1019_ vdd gnd FILL
XFILL_0__1152_ vdd gnd FILL
XFILL_0__1083_ vdd gnd FILL
XFILL_1__954_ vdd gnd FILL
X_1145_ _1145_/A _1145_/B _1145_/C _1154_/B vdd gnd AOI21X1
XFILL_1__885_ vdd gnd FILL
X_1214_ _1422_/B _1297_/A _1552_/D vdd gnd XNOR2X1
XFILL_1__1330_ vdd gnd FILL
XFILL_3__1128_ vdd gnd FILL
XFILL_1__1192_ vdd gnd FILL
X_1076_ _1079_/C _1078_/B _1084_/A vdd gnd NAND2X1
XFILL_0__1419_ vdd gnd FILL
XFILL_1__1261_ vdd gnd FILL
XFILL_3__1059_ vdd gnd FILL
XFILL_2__1370_ vdd gnd FILL
XFILL_1__1459_ vdd gnd FILL
XFILL_0__972_ vdd gnd FILL
XFILL_2__919_ vdd gnd FILL
X_925_ _925_/A _925_/B _925_/C _933_/C vdd gnd AOI21X1
X_787_ _787_/A _787_/B _787_/C _797_/B vdd gnd AOI21X1
X_856_ _861_/A _964_/A _856_/C _867_/A vdd gnd OAI21X1
XFILL_2__1568_ vdd gnd FILL
XFILL_0__1204_ vdd gnd FILL
XFILL_2__1499_ vdd gnd FILL
XFILL_0__1066_ vdd gnd FILL
XFILL_0__1135_ vdd gnd FILL
XFILL_1__937_ vdd gnd FILL
XFILL_1__868_ vdd gnd FILL
X_1128_ _1128_/A _1128_/B _1198_/A _1217_/C vdd gnd OAI21X1
X_1059_ Cin[3] Xin[4] _1065_/B vdd gnd AND2X2
XFILL_1__799_ vdd gnd FILL
XFILL_1__1313_ vdd gnd FILL
XFILL_1__1244_ vdd gnd FILL
XFILL_1__1175_ vdd gnd FILL
XFILL_2__1422_ vdd gnd FILL
XFILL_2__1353_ vdd gnd FILL
XFILL_2__1284_ vdd gnd FILL
XFILL_1_CLKBUF1_insert5 vdd gnd FILL
XFILL_0__955_ vdd gnd FILL
XFILL_0__886_ vdd gnd FILL
X_908_ _977_/A _970_/B _911_/B vdd gnd NAND2X1
X_839_ _912_/A Xin[4] Yin[4] _903_/B vdd gnd AOI21X1
XFILL_3__1462_ vdd gnd FILL
XFILL_3__1393_ vdd gnd FILL
XFILL_0__1118_ vdd gnd FILL
XFILL_0__1049_ vdd gnd FILL
XFILL_4__1005_ vdd gnd FILL
XFILL_1__1089_ vdd gnd FILL
XFILL_1__1158_ vdd gnd FILL
XFILL_1__1227_ vdd gnd FILL
XFILL_3__882_ vdd gnd FILL
XFILL_3__951_ vdd gnd FILL
XFILL_2__1405_ vdd gnd FILL
XFILL_0__938_ vdd gnd FILL
XFILL_2__1198_ vdd gnd FILL
XFILL_2__1267_ vdd gnd FILL
XFILL_2__1336_ vdd gnd FILL
X_1531_ _1547_/Q _1549_/CLK _1577_/A vdd gnd DFFPOSX1
XFILL_0__869_ vdd gnd FILL
X_1462_ _1489_/C _1464_/A _1556_/D vdd gnd XNOR2X1
XFILL_3__1445_ vdd gnd FILL
XFILL_3__1514_ vdd gnd FILL
X_1393_ _1400_/C _1400_/B _1400_/A _1399_/B vdd gnd NAND3X1
XFILL_3__1376_ vdd gnd FILL
XFILL_1__1012_ vdd gnd FILL
XFILL_4__778_ vdd gnd FILL
XFILL_2__1121_ vdd gnd FILL
XFILL_2__1052_ vdd gnd FILL
XFILL_3__865_ vdd gnd FILL
XFILL_3__934_ vdd gnd FILL
XFILL_3__796_ vdd gnd FILL
XFILL_3__1092_ vdd gnd FILL
XFILL_3__1230_ vdd gnd FILL
XFILL_0__1452_ vdd gnd FILL
XFILL_0__1383_ vdd gnd FILL
XFILL_2__1319_ vdd gnd FILL
XFILL_3__1161_ vdd gnd FILL
X_1445_ _1478_/A _1478_/B _1446_/A vdd gnd NAND2X1
X_1514_ _1514_/A _1514_/B _1514_/C _1516_/C vdd gnd OAI21X1
XFILL_1__1561_ vdd gnd FILL
X_1376_ _1435_/A _1376_/B _1466_/A _1386_/B vdd gnd OAI21X1
XFILL_3__1428_ vdd gnd FILL
XFILL_1__1492_ vdd gnd FILL
XFILL_2__883_ vdd gnd FILL
XFILL_2__952_ vdd gnd FILL
XFILL_3__1359_ vdd gnd FILL
XFILL_2__1104_ vdd gnd FILL
XFILL_2__1035_ vdd gnd FILL
XFILL_1__970_ vdd gnd FILL
XBUFX2_insert6 Cin[0] _977_/A vdd gnd BUFX2
XFILL_3__917_ vdd gnd FILL
XFILL_3__848_ vdd gnd FILL
X_1092_ _993_/A _1093_/C vdd gnd INVX1
XFILL_3__779_ vdd gnd FILL
X_1230_ _1304_/B _1237_/B vdd gnd INVX1
X_1161_ Cin[3] Xin[6] _1336_/A vdd gnd AND2X2
XFILL_3__1144_ vdd gnd FILL
XFILL_3__1213_ vdd gnd FILL
XFILL_3__1075_ vdd gnd FILL
XFILL_0__1366_ vdd gnd FILL
XFILL_0__1504_ vdd gnd FILL
XFILL_0__1435_ vdd gnd FILL
XFILL_0__1297_ vdd gnd FILL
XFILL_1_BUFX2_insert10 vdd gnd FILL
X_1428_ _1428_/A _1428_/B _1465_/A vdd gnd NAND2X1
XFILL_1__1475_ vdd gnd FILL
X_1359_ _1414_/C _1366_/A _1366_/B _1361_/A vdd gnd NAND3X1
XFILL_4__1322_ vdd gnd FILL
XFILL_4__1253_ vdd gnd FILL
XFILL_4__1184_ vdd gnd FILL
XFILL_2__866_ vdd gnd FILL
XFILL_2__935_ vdd gnd FILL
X_941_ _941_/A _941_/B _941_/C _941_/D _945_/B vdd gnd AOI22X1
XFILL_2__797_ vdd gnd FILL
X_872_ _872_/A _872_/B _872_/C _875_/C vdd gnd AOI21X1
XFILL_0__1220_ vdd gnd FILL
XFILL_2__1018_ vdd gnd FILL
XFILL_0__1082_ vdd gnd FILL
XFILL_0__1151_ vdd gnd FILL
XFILL_1__953_ vdd gnd FILL
X_1213_ _1296_/A _1213_/B _1297_/A vdd gnd NAND2X1
XFILL_1__884_ vdd gnd FILL
X_1144_ _1154_/C _1242_/A _1153_/C _1219_/A vdd gnd NAND3X1
X_1075_ _1171_/A Xin[7] _1078_/B vdd gnd NAND2X1
XFILL_1__1260_ vdd gnd FILL
XFILL_3__1127_ vdd gnd FILL
XFILL_3__1058_ vdd gnd FILL
XFILL_1__1191_ vdd gnd FILL
XFILL_0__1349_ vdd gnd FILL
XFILL_0__1418_ vdd gnd FILL
XFILL_0__971_ vdd gnd FILL
XFILL_1__1458_ vdd gnd FILL
XFILL_1__1389_ vdd gnd FILL
XFILL_2__918_ vdd gnd FILL
XFILL_2__849_ vdd gnd FILL
X_924_ _947_/B _947_/A _947_/C _948_/C vdd gnd NAND3X1
X_786_ _787_/C _787_/B _787_/A _797_/C vdd gnd NAND3X1
X_855_ Xin[2] _861_/A vdd gnd INVX2
XFILL_2__1567_ vdd gnd FILL
XFILL_2__1498_ vdd gnd FILL
XFILL_4__880_ vdd gnd FILL
XFILL_0__1203_ vdd gnd FILL
XFILL_0__1134_ vdd gnd FILL
XFILL_0__1065_ vdd gnd FILL
XFILL_1__936_ vdd gnd FILL
XFILL_1__867_ vdd gnd FILL
XFILL_1__798_ vdd gnd FILL
X_1127_ _1127_/A _1127_/B _1127_/C _1128_/B vdd gnd AOI21X1
X_1058_ _1143_/A _1149_/D vdd gnd INVX1
XFILL_1__1312_ vdd gnd FILL
XFILL_1__1243_ vdd gnd FILL
XFILL_1__1174_ vdd gnd FILL
XFILL_2__1352_ vdd gnd FILL
XFILL_2__1421_ vdd gnd FILL
XFILL_0__954_ vdd gnd FILL
XFILL_2__1283_ vdd gnd FILL
XFILL_0__885_ vdd gnd FILL
X_907_ Yin[5] _912_/C vdd gnd INVX1
X_838_ _912_/A Xin[4] Yin[4] _903_/C vdd gnd NAND3X1
XFILL_3__1461_ vdd gnd FILL
X_769_ _777_/C _770_/B vdd gnd INVX1
XFILL88950x4050 vdd gnd FILL
XFILL_3__1392_ vdd gnd FILL
XFILL_0__1117_ vdd gnd FILL
XFILL_0__1048_ vdd gnd FILL
XFILL_4__1570_ vdd gnd FILL
XFILL_1_BUFX2_insert6 vdd gnd FILL
XFILL_1__919_ vdd gnd FILL
XFILL89550x54750 vdd gnd FILL
XFILL_1__1226_ vdd gnd FILL
XFILL_1__1088_ vdd gnd FILL
XFILL_1__1157_ vdd gnd FILL
XFILL_3__950_ vdd gnd FILL
XFILL_3__881_ vdd gnd FILL
XFILL_2__1404_ vdd gnd FILL
XFILL_2__1335_ vdd gnd FILL
XFILL_0__937_ vdd gnd FILL
XFILL_2__1197_ vdd gnd FILL
XFILL_2__1266_ vdd gnd FILL
XFILL_0__868_ vdd gnd FILL
X_1530_ _1546_/Q _1552_/CLK _1576_/A vdd gnd DFFPOSX1
X_1461_ _1488_/C _1486_/A _1464_/A vdd gnd NAND2X1
X_1392_ _1392_/A _1392_/B _1392_/C _1400_/A vdd gnd OAI21X1
XFILL_0__799_ vdd gnd FILL
XFILL_3__1444_ vdd gnd FILL
XFILL_3__1513_ vdd gnd FILL
XFILL_3__1375_ vdd gnd FILL
XFILL_1__1011_ vdd gnd FILL
XFILL_4__1484_ vdd gnd FILL
XFILL89550x66450 vdd gnd FILL
XFILL_2__1120_ vdd gnd FILL
XFILL_1__1209_ vdd gnd FILL
XFILL_2__1051_ vdd gnd FILL
XFILL_3__933_ vdd gnd FILL
XFILL_3__864_ vdd gnd FILL
XFILL_3__795_ vdd gnd FILL
XFILL_3__1091_ vdd gnd FILL
XFILL_0__1451_ vdd gnd FILL
XFILL_0__1382_ vdd gnd FILL
XFILL_2__1249_ vdd gnd FILL
XFILL_2__1318_ vdd gnd FILL
XFILL_3__1160_ vdd gnd FILL
X_1375_ Cin[5] Xin[6] _1466_/A vdd gnd NAND2X1
X_1444_ _1478_/B _1478_/A _1476_/A vdd gnd OR2X2
X_1513_ _1513_/A _1513_/B _1514_/A vdd gnd AND2X2
XFILL_1__1560_ vdd gnd FILL
XFILL_1__1491_ vdd gnd FILL
XFILL_3__1427_ vdd gnd FILL
XFILL_3__1358_ vdd gnd FILL
XFILL_2__882_ vdd gnd FILL
XFILL_4__829_ vdd gnd FILL
XFILL_2__951_ vdd gnd FILL
XFILL_3__1289_ vdd gnd FILL
XFILL89550x78150 vdd gnd FILL
XFILL_2__1103_ vdd gnd FILL
XFILL_2__1034_ vdd gnd FILL
XFILL_3__916_ vdd gnd FILL
XBUFX2_insert7 Cin[0] _912_/A vdd gnd BUFX2
XFILL_3__847_ vdd gnd FILL
XFILL_3__778_ vdd gnd FILL
X_1091_ _1127_/B _1127_/C _1127_/A _1198_/A vdd gnd NAND3X1
XFILL_3__1212_ vdd gnd FILL
XFILL_0__1503_ vdd gnd FILL
X_1160_ _1235_/A _1239_/D vdd gnd INVX1
XFILL_3__1143_ vdd gnd FILL
XFILL_3__1074_ vdd gnd FILL
XFILL_0__1434_ vdd gnd FILL
XFILL_0__1365_ vdd gnd FILL
XFILL_0__1296_ vdd gnd FILL
XFILL_1_BUFX2_insert11 vdd gnd FILL
X_1427_ _1427_/A _1427_/B _1512_/B _1489_/C vdd gnd NAND3X1
X_1358_ _1358_/A _1358_/B _1358_/C _1361_/C vdd gnd OAI21X1
X_1289_ _1289_/A _1289_/B _1289_/C _1292_/C vdd gnd AOI21X1
XFILL_1__1474_ vdd gnd FILL
XFILL_2__865_ vdd gnd FILL
XFILL_2__934_ vdd gnd FILL
XFILL_2__796_ vdd gnd FILL
X_940_ _941_/A _941_/B _940_/C _945_/C vdd gnd NAND3X1
X_871_ _878_/C _878_/B _878_/A _884_/C vdd gnd NAND3X1
XFILL_2__1583_ vdd gnd FILL
XFILL_0__1150_ vdd gnd FILL
XFILL_2__1017_ vdd gnd FILL
XFILL_0__1081_ vdd gnd FILL
XFILL_1__883_ vdd gnd FILL
XFILL_1__952_ vdd gnd FILL
X_1212_ _1212_/A _1212_/B _1212_/C _1296_/A vdd gnd NAND3X1
X_1143_ _1143_/A _1143_/B _1143_/C _1154_/C vdd gnd OAI21X1
X_1074_ Yin[7] _1079_/C vdd gnd INVX1
XFILL_0__1417_ vdd gnd FILL
XFILL_3__1057_ vdd gnd FILL
XFILL_3__1126_ vdd gnd FILL
XFILL_0__1348_ vdd gnd FILL
XFILL_0__1279_ vdd gnd FILL
XFILL_1__1190_ vdd gnd FILL
XFILL_4__1304_ vdd gnd FILL
XFILL_2__917_ vdd gnd FILL
XFILL_0__970_ vdd gnd FILL
XFILL_4__1097_ vdd gnd FILL
XFILL_4__1235_ vdd gnd FILL
XFILL_1__1457_ vdd gnd FILL
XFILL_1__1388_ vdd gnd FILL
XFILL_4__1166_ vdd gnd FILL
XFILL_2__848_ vdd gnd FILL
XFILL_2__779_ vdd gnd FILL
X_923_ _955_/A _926_/B _926_/A _947_/B vdd gnd NAND3X1
X_854_ _861_/C _894_/A _867_/C vdd gnd NAND2X1
XFILL_2__1566_ vdd gnd FILL
X_785_ _805_/B _785_/B _805_/A _787_/A vdd gnd OAI21X1
XFILL_2_CLKBUF1_insert0 vdd gnd FILL
XFILL_2__1497_ vdd gnd FILL
XFILL_0__1202_ vdd gnd FILL
XFILL_0__1133_ vdd gnd FILL
XFILL_0__1064_ vdd gnd FILL
XFILL_1__866_ vdd gnd FILL
XFILL_1__935_ vdd gnd FILL
XFILL_1__797_ vdd gnd FILL
X_1126_ _1289_/A _1218_/A vdd gnd INVX1
XFILL_3__1109_ vdd gnd FILL
X_1057_ _895_/A Cin[4] _1143_/A vdd gnd NAND2X1
XFILL_1__1242_ vdd gnd FILL
XFILL_1__1311_ vdd gnd FILL
XFILL_1__1173_ vdd gnd FILL
XFILL_2__1351_ vdd gnd FILL
XFILL_2__1420_ vdd gnd FILL
XFILL_1__1509_ vdd gnd FILL
XFILL_2__1282_ vdd gnd FILL
XFILL_0__953_ vdd gnd FILL
XFILL_0__884_ vdd gnd FILL
X_906_ _977_/A _970_/B Yin[5] _969_/C vdd gnd NAND3X1
X_837_ _837_/A _837_/B _847_/A _866_/C vdd gnd OAI21X1
X_768_ _768_/A _777_/C _768_/C _773_/A vdd gnd NAND3X1
XFILL_3__1460_ vdd gnd FILL
XFILL_3__1391_ vdd gnd FILL
XFILL_0__1116_ vdd gnd FILL
XFILL_0__1047_ vdd gnd FILL
XFILL_1_BUFX2_insert7 vdd gnd FILL
XFILL_1__918_ vdd gnd FILL
XFILL_1__849_ vdd gnd FILL
X_1109_ _1109_/A _1109_/B _1208_/C _1115_/B vdd gnd OAI21X1
XFILL_1__1156_ vdd gnd FILL
XFILL_1__1225_ vdd gnd FILL
XFILL_1__1087_ vdd gnd FILL
XFILL89550x4050 vdd gnd FILL
XFILL_3__880_ vdd gnd FILL
XFILL_2__1334_ vdd gnd FILL
XFILL_2__1403_ vdd gnd FILL
XFILL_2__1265_ vdd gnd FILL
XFILL_0__936_ vdd gnd FILL
XFILL_0__867_ vdd gnd FILL
XFILL_2__1196_ vdd gnd FILL
XFILL_0__798_ vdd gnd FILL
X_1460_ _1460_/A _1460_/B _1460_/C _1488_/C vdd gnd NAND3X1
X_1391_ _1391_/A _1391_/B _1391_/C _1400_/B vdd gnd NAND3X1
XFILL_3__1374_ vdd gnd FILL
XFILL_3__1443_ vdd gnd FILL
XFILL_3__1512_ vdd gnd FILL
XFILL_1__1010_ vdd gnd FILL
XFILL_1__1208_ vdd gnd FILL
XFILL_2__1050_ vdd gnd FILL
XFILL_1__1139_ vdd gnd FILL
XFILL_3__932_ vdd gnd FILL
XFILL_3__863_ vdd gnd FILL
XFILL_3__794_ vdd gnd FILL
XFILL_0__1450_ vdd gnd FILL
XFILL_3__1090_ vdd gnd FILL
XFILL_2__1317_ vdd gnd FILL
XFILL_2__1248_ vdd gnd FILL
XFILL_0__1381_ vdd gnd FILL
XFILL_0__919_ vdd gnd FILL
X_1512_ _1512_/A _1512_/B _1512_/C _1514_/B vdd gnd AOI21X1
XFILL_2__1179_ vdd gnd FILL
X_1374_ _1436_/A _1435_/A vdd gnd INVX1
X_1443_ Yin[11] _1443_/B _1478_/B vdd gnd NAND2X1
XFILL_0__1579_ vdd gnd FILL
XFILL_2__950_ vdd gnd FILL
XFILL_3__1288_ vdd gnd FILL
XFILL_1__1490_ vdd gnd FILL
XFILL_3__1426_ vdd gnd FILL
XFILL_3__1357_ vdd gnd FILL
XFILL_2__881_ vdd gnd FILL
XFILL_2__1102_ vdd gnd FILL
XFILL_2__1033_ vdd gnd FILL
XFILL_3__915_ vdd gnd FILL
XFILL_3__846_ vdd gnd FILL
XBUFX2_insert8 Cin[0] _814_/A vdd gnd BUFX2
XFILL_3__1142_ vdd gnd FILL
X_1090_ _1158_/B _1094_/B _1094_/A _1127_/B vdd gnd NAND3X1
XFILL_3__1211_ vdd gnd FILL
XFILL_3__777_ vdd gnd FILL
XFILL_0__1433_ vdd gnd FILL
XFILL_0__1502_ vdd gnd FILL
XFILL_3__1073_ vdd gnd FILL
XFILL_0__1364_ vdd gnd FILL
XFILL_0__1295_ vdd gnd FILL
XFILL_1_BUFX2_insert12 vdd gnd FILL
X_1288_ _1288_/A _1289_/C vdd gnd INVX1
X_1426_ _1511_/A _1511_/B _1427_/B vdd gnd NAND2X1
X_1357_ _1357_/A _1357_/B _1357_/C _1358_/B vdd gnd AOI21X1
XFILL_2__933_ vdd gnd FILL
XFILL_3__1409_ vdd gnd FILL
XFILL_1__1473_ vdd gnd FILL
XFILL_2__864_ vdd gnd FILL
XFILL_2__795_ vdd gnd FILL
X_870_ _925_/C _890_/B _890_/A _878_/A vdd gnd OAI21X1
XFILL_2__1582_ vdd gnd FILL
XFILL_2__1016_ vdd gnd FILL
XFILL88650x54750 vdd gnd FILL
XFILL_0__1080_ vdd gnd FILL
XFILL_1__882_ vdd gnd FILL
X_999_ _999_/A _999_/B _999_/C _999_/Y vdd gnd OAI21X1
XFILL_3__829_ vdd gnd FILL
X_1142_ Cin[2] _912_/B Cin[3] Xin[4] _1143_/B vdd gnd AOI22X1
XFILL_1__951_ vdd gnd FILL
X_1211_ _1218_/A _1211_/B _1211_/C _1212_/C vdd gnd NAND3X1
XFILL_3__1125_ vdd gnd FILL
X_1073_ _1171_/A Xin[7] Yin[7] _1265_/A vdd gnd NAND3X1
XFILL_0__1416_ vdd gnd FILL
XFILL_3__1056_ vdd gnd FILL
XFILL_0__1347_ vdd gnd FILL
XFILL_0__1278_ vdd gnd FILL
X_1409_ _1430_/A _1409_/B _1409_/C _1458_/A vdd gnd NAND3X1
XFILL_2__916_ vdd gnd FILL
XFILL_1__1456_ vdd gnd FILL
XFILL_1__1387_ vdd gnd FILL
XFILL_2__847_ vdd gnd FILL
XFILL_2__778_ vdd gnd FILL
XFILL88950x31350 vdd gnd FILL
XFILL88050x19650 vdd gnd FILL
XFILL_2__1565_ vdd gnd FILL
X_922_ _954_/B _954_/A _922_/C _926_/B vdd gnd NAND3X1
X_784_ _805_/C _785_/B vdd gnd INVX1
X_853_ Xin[2] Cin[2] _894_/A vdd gnd AND2X2
XFILL_2_CLKBUF1_insert1 vdd gnd FILL
XFILL_0__1201_ vdd gnd FILL
XFILL88350x7950 vdd gnd FILL
XFILL_2__1496_ vdd gnd FILL
XFILL_0__1063_ vdd gnd FILL
XFILL_0__1132_ vdd gnd FILL
XCLKBUF1_insert0 clk _1557_/CLK vdd gnd CLKBUF1
XFILL_1__934_ vdd gnd FILL
XFILL_1__865_ vdd gnd FILL
XFILL_1__796_ vdd gnd FILL
X_1125_ _1125_/A _1125_/B _1289_/A vdd gnd NAND2X1
XFILL_1__1310_ vdd gnd FILL
X_1056_ _1056_/A _994_/A _993_/A _1127_/C vdd gnd OAI21X1
XFILL_3__1108_ vdd gnd FILL
XFILL_1__1172_ vdd gnd FILL
XFILL_1__1241_ vdd gnd FILL
XFILL_3__1039_ vdd gnd FILL
XFILL_2__1350_ vdd gnd FILL
XFILL_1__1439_ vdd gnd FILL
XFILL_1__1508_ vdd gnd FILL
XFILL_2__1281_ vdd gnd FILL
XFILL_0__883_ vdd gnd FILL
XFILL_0__952_ vdd gnd FILL
XFILL88650x78150 vdd gnd FILL
X_905_ _969_/A _917_/C vdd gnd INVX1
X_836_ _912_/A _836_/B Yin[3] _837_/B vdd gnd AOI21X1
X_767_ _777_/B _768_/C vdd gnd INVX1
XFILL_3__1390_ vdd gnd FILL
XFILL_4__930_ vdd gnd FILL
XFILL_4__792_ vdd gnd FILL
XFILL_4__861_ vdd gnd FILL
XFILL_2__1479_ vdd gnd FILL
XFILL_0__1115_ vdd gnd FILL
XFILL_0__1046_ vdd gnd FILL
XFILL_1__917_ vdd gnd FILL
XFILL_1_BUFX2_insert8 vdd gnd FILL
XFILL_1__848_ vdd gnd FILL
XFILL_1__779_ vdd gnd FILL
X_1108_ _1124_/A _1209_/C _1124_/B _1112_/B vdd gnd NAND3X1
X_1039_ _1129_/A _1039_/B _1045_/B vdd gnd NAND2X1
XFILL_1__1086_ vdd gnd FILL
XFILL_1__1155_ vdd gnd FILL
XFILL_1__1224_ vdd gnd FILL
XFILL_2__1402_ vdd gnd FILL
XFILL_2__1195_ vdd gnd FILL
XFILL_2__1264_ vdd gnd FILL
XFILL_2__1333_ vdd gnd FILL
XFILL_0__866_ vdd gnd FILL
XFILL_0__935_ vdd gnd FILL
XFILL_0__797_ vdd gnd FILL
XFILL_3__1511_ vdd gnd FILL
X_1390_ _1401_/C _1400_/C vdd gnd INVX1
X_819_ _848_/B _847_/A _848_/A _820_/A vdd gnd AOI21X1
XFILL_3__1373_ vdd gnd FILL
XFILL_3__1442_ vdd gnd FILL
XFILL_0__1029_ vdd gnd FILL
XFILL_1__1069_ vdd gnd FILL
XFILL_1__1207_ vdd gnd FILL
XFILL_1__1138_ vdd gnd FILL
XFILL_3__931_ vdd gnd FILL
XFILL_3__862_ vdd gnd FILL
XFILL_3__793_ vdd gnd FILL
XFILL_0__1380_ vdd gnd FILL
XFILL_2__1316_ vdd gnd FILL
XFILL_2__1247_ vdd gnd FILL
XFILL_2__1178_ vdd gnd FILL
XFILL_0__918_ vdd gnd FILL
XFILL_0__849_ vdd gnd FILL
X_1442_ Yin[12] _1478_/A vdd gnd INVX1
X_1511_ _1511_/A _1511_/B _1511_/C _1511_/D _1512_/A vdd gnd AOI22X1
X_1373_ Xin[6] Cin[6] _1492_/B vdd gnd NAND2X1
XFILL_3__1425_ vdd gnd FILL
XFILL_0__1578_ vdd gnd FILL
XFILL_2__880_ vdd gnd FILL
XFILL_3__1356_ vdd gnd FILL
XFILL_3__1287_ vdd gnd FILL
XFILL_4__1396_ vdd gnd FILL
XFILL_4__1465_ vdd gnd FILL
XFILL_2__1101_ vdd gnd FILL
XFILL_2__1032_ vdd gnd FILL
XFILL_3__914_ vdd gnd FILL
XFILL_3__845_ vdd gnd FILL
XFILL_3__776_ vdd gnd FILL
XFILL_3__1141_ vdd gnd FILL
XFILL_3__1210_ vdd gnd FILL
XFILL_0__1432_ vdd gnd FILL
XBUFX2_insert9 Cin[0] _1171_/A vdd gnd BUFX2
XFILL_0__1501_ vdd gnd FILL
XFILL_0__1363_ vdd gnd FILL
XFILL_3__1072_ vdd gnd FILL
XFILL_0__1294_ vdd gnd FILL
XFILL_1_BUFX2_insert13 vdd gnd FILL
X_1425_ _1425_/A _1425_/B _1511_/B vdd gnd NAND2X1
XFILL_3__1408_ vdd gnd FILL
X_1356_ _1356_/A _1356_/B _1356_/C _1362_/B vdd gnd OAI21X1
X_1287_ _1287_/A _1287_/B _1287_/C _1296_/C vdd gnd NAND3X1
XFILL_1__1472_ vdd gnd FILL
XFILL_2__932_ vdd gnd FILL
XFILL_2__863_ vdd gnd FILL
XFILL_3__1339_ vdd gnd FILL
XFILL_2__794_ vdd gnd FILL
XFILL_2__1581_ vdd gnd FILL
XFILL_2__1015_ vdd gnd FILL
XFILL_1__950_ vdd gnd FILL
XFILL_1__881_ vdd gnd FILL
X_998_ _998_/A _998_/B _998_/C _998_/Y vdd gnd NAND3X1
XFILL_3__828_ vdd gnd FILL
XFILL_3__759_ vdd gnd FILL
X_1141_ _1145_/C _1145_/A _1145_/B _1153_/C vdd gnd NAND3X1
X_1072_ _1172_/A _1084_/C vdd gnd INVX1
X_1210_ _1289_/A _1288_/A _1289_/B _1212_/B vdd gnd NAND3X1
XFILL_3__1055_ vdd gnd FILL
XFILL_3__1124_ vdd gnd FILL
XFILL_0__1346_ vdd gnd FILL
XFILL_0__1415_ vdd gnd FILL
XFILL_0__1277_ vdd gnd FILL
X_1408_ _1416_/C _1416_/B _1416_/A _1412_/A vdd gnd AOI21X1
X_1339_ _1369_/B _1342_/A _1370_/B vdd gnd XOR2X1
XFILL_1__1455_ vdd gnd FILL
XFILL_2__915_ vdd gnd FILL
XFILL_2__846_ vdd gnd FILL
XFILL_1__1386_ vdd gnd FILL
X_921_ _921_/A _921_/B _954_/C _926_/A vdd gnd OAI21X1
XFILL_2__777_ vdd gnd FILL
X_783_ _783_/A _805_/C _783_/C _787_/B vdd gnd NAND3X1
X_852_ Xin[0] Cin[4] _868_/A vdd gnd NAND2X1
XFILL_2__1564_ vdd gnd FILL
XFILL_2_CLKBUF1_insert2 vdd gnd FILL
XFILL_0__1200_ vdd gnd FILL
XFILL_2__1495_ vdd gnd FILL
XFILL_0__1062_ vdd gnd FILL
XCLKBUF1_insert1 clk _1546_/CLK vdd gnd CLKBUF1
XFILL_0__1131_ vdd gnd FILL
XFILL_1__933_ vdd gnd FILL
XFILL_1__864_ vdd gnd FILL
X_1055_ _986_/C _986_/B _986_/A _1056_/A vdd gnd AOI21X1
XFILL_1__795_ vdd gnd FILL
X_1124_ _1124_/A _1124_/B _1124_/C _1207_/C vdd gnd AOI21X1
XFILL_3__1107_ vdd gnd FILL
XFILL_3__1038_ vdd gnd FILL
XFILL_1__1171_ vdd gnd FILL
XFILL_1__1240_ vdd gnd FILL
XFILL_0__1329_ vdd gnd FILL
XFILL_0__951_ vdd gnd FILL
XFILL_4__1216_ vdd gnd FILL
XFILL_4__1147_ vdd gnd FILL
XFILL_1__1369_ vdd gnd FILL
XFILL_2__1280_ vdd gnd FILL
XFILL_1__1438_ vdd gnd FILL
XFILL_1__1507_ vdd gnd FILL
XFILL_0__882_ vdd gnd FILL
XFILL_2__829_ vdd gnd FILL
XFILL_4__1078_ vdd gnd FILL
X_904_ Cin[1] Xin[4] _969_/A vdd gnd NAND2X1
X_835_ _835_/A _835_/B _877_/A _878_/C vdd gnd OAI21X1
X_766_ _814_/A Xin[1] Yin[1] _777_/B vdd gnd AOI21X1
XFILL_2__1478_ vdd gnd FILL
XFILL_0__1114_ vdd gnd FILL
XFILL_0__1045_ vdd gnd FILL
XFILL_1__916_ vdd gnd FILL
XFILL_1__847_ vdd gnd FILL
XFILL_1_BUFX2_insert9 vdd gnd FILL
XFILL_1__778_ vdd gnd FILL
X_1107_ _1109_/A _1109_/B _1110_/C _1124_/B vdd gnd OAI21X1
X_1038_ _1223_/A _951_/B _1045_/A vdd gnd NAND2X1
XFILL_1__1223_ vdd gnd FILL
XFILL_1__1085_ vdd gnd FILL
XFILL_1__1154_ vdd gnd FILL
XFILL_2__1401_ vdd gnd FILL
XFILL_2__1332_ vdd gnd FILL
XFILL_0__934_ vdd gnd FILL
XFILL_2__1194_ vdd gnd FILL
XFILL_2__1263_ vdd gnd FILL
XFILL_0__865_ vdd gnd FILL
XFILL_0__796_ vdd gnd FILL
X_818_ _818_/A _818_/B _837_/A _820_/B vdd gnd AOI21X1
XFILL_3__1441_ vdd gnd FILL
XFILL_3__1510_ vdd gnd FILL
XFILL_4__912_ vdd gnd FILL
XFILL_3__1372_ vdd gnd FILL
XFILL_4__843_ vdd gnd FILL
XFILL_4__774_ vdd gnd FILL
XFILL_0__1028_ vdd gnd FILL
XFILL_1__1206_ vdd gnd FILL
XFILL_1__1068_ vdd gnd FILL
XFILL_1__1137_ vdd gnd FILL
XFILL_3__930_ vdd gnd FILL
XFILL_3__792_ vdd gnd FILL
XFILL_3__861_ vdd gnd FILL
XFILL_2__1315_ vdd gnd FILL
XFILL_2__1177_ vdd gnd FILL
XFILL_0__917_ vdd gnd FILL
XFILL_2__1246_ vdd gnd FILL
XFILL_0__848_ vdd gnd FILL
XFILL_0__779_ vdd gnd FILL
X_1441_ _1449_/A _1481_/A _1448_/B vdd gnd NOR2X1
X_1510_ _1515_/A _1510_/B _1517_/B vdd gnd NAND2X1
XFILL_3__1424_ vdd gnd FILL
X_1372_ Cin[7] _1470_/B vdd gnd INVX1
XFILL_0__1577_ vdd gnd FILL
XFILL_3__1355_ vdd gnd FILL
XFILL_3__1286_ vdd gnd FILL
XFILL_2__1100_ vdd gnd FILL
XFILL_2__1031_ vdd gnd FILL
XFILL_3__913_ vdd gnd FILL
XFILL_3__844_ vdd gnd FILL
XFILL_3__775_ vdd gnd FILL
XFILL_0__1500_ vdd gnd FILL
XFILL_3__1140_ vdd gnd FILL
XFILL_3__1071_ vdd gnd FILL
XFILL_0__1362_ vdd gnd FILL
XFILL_0__1431_ vdd gnd FILL
XFILL_0__1293_ vdd gnd FILL
XFILL_2__1229_ vdd gnd FILL
XFILL_1_BUFX2_insert14 vdd gnd FILL
X_1424_ _1424_/A _1424_/B _1511_/D _1427_/A vdd gnd NAND3X1
X_1355_ _1366_/B _1414_/C _1366_/A _1356_/B vdd gnd AOI21X1
XFILL_3__1338_ vdd gnd FILL
XFILL_3__1407_ vdd gnd FILL
X_1286_ _1358_/A _1290_/B _1290_/A _1287_/C vdd gnd NAND3X1
XFILL_4__1180_ vdd gnd FILL
XFILL_1__1471_ vdd gnd FILL
XFILL_2__931_ vdd gnd FILL
XFILL_2__862_ vdd gnd FILL
XFILL_2__793_ vdd gnd FILL
XFILL_3__1269_ vdd gnd FILL
XFILL89250x85950 vdd gnd FILL
XFILL_2__1580_ vdd gnd FILL
XFILL_4__1447_ vdd gnd FILL
XFILL_4__1516_ vdd gnd FILL
XFILL_4__1378_ vdd gnd FILL
XFILL_2__1014_ vdd gnd FILL
XFILL_1__880_ vdd gnd FILL
X_997_ _997_/A _997_/B _997_/Y vdd gnd XOR2X1
XFILL_3__827_ vdd gnd FILL
XFILL_3__758_ vdd gnd FILL
X_1140_ _861_/A _1376_/B _1232_/A _1145_/B vdd gnd OAI21X1
X_1071_ Cin[1] Xin[6] _1172_/A vdd gnd NAND2X1
XFILL_3__1123_ vdd gnd FILL
XFILL_3__1054_ vdd gnd FILL
XFILL_0__1276_ vdd gnd FILL
XFILL_0__1345_ vdd gnd FILL
XFILL_0__1414_ vdd gnd FILL
X_1338_ _1396_/A _1343_/A _1342_/A vdd gnd NAND2X1
X_1407_ _1430_/A _1409_/B _1459_/A _1416_/B vdd gnd NAND3X1
XFILL_1__1454_ vdd gnd FILL
X_1269_ _1303_/C _1348_/B _1348_/A _1357_/B vdd gnd NAND3X1
XFILL_1__1385_ vdd gnd FILL
XFILL_2__914_ vdd gnd FILL
XFILL_2__845_ vdd gnd FILL
XFILL_2__776_ vdd gnd FILL
X_851_ _865_/B _865_/A _865_/C _925_/A vdd gnd NAND3X1
X_920_ _927_/B _952_/C _955_/A vdd gnd NAND2X1
X_782_ _805_/B _783_/C vdd gnd INVX1
XFILL_2__1563_ vdd gnd FILL
XFILL_2__1494_ vdd gnd FILL
XFILL_0__1130_ vdd gnd FILL
XFILL_2_CLKBUF1_insert3 vdd gnd FILL
XCLKBUF1_insert2 clk _1549_/CLK vdd gnd CLKBUF1
XFILL_0__1061_ vdd gnd FILL
XFILL_1__932_ vdd gnd FILL
XFILL_1__863_ vdd gnd FILL
X_1123_ _1209_/C _1124_/C vdd gnd INVX1
XFILL_1__794_ vdd gnd FILL
X_1054_ _1125_/B _1098_/B _1199_/A vdd gnd AND2X2
XFILL_3__1106_ vdd gnd FILL
XFILL_3__1037_ vdd gnd FILL
XFILL_0__1328_ vdd gnd FILL
XFILL_0__1259_ vdd gnd FILL
XFILL_1__1170_ vdd gnd FILL
XFILL_1__1506_ vdd gnd FILL
XFILL89550x74250 vdd gnd FILL
XFILL_0__950_ vdd gnd FILL
XFILL_1__1437_ vdd gnd FILL
XFILL_1__1368_ vdd gnd FILL
XFILL_0__881_ vdd gnd FILL
XFILL_2__828_ vdd gnd FILL
XFILL_2__759_ vdd gnd FILL
XFILL_1__1299_ vdd gnd FILL
X_903_ _903_/A _903_/B _903_/C _954_/C vdd gnd OAI21X1
X_834_ _884_/A _936_/B vdd gnd INVX1
X_765_ _814_/A Xin[1] Yin[1] _777_/C vdd gnd NAND3X1
XFILL_2__1477_ vdd gnd FILL
XFILL_0__1113_ vdd gnd FILL
XFILL_0__1044_ vdd gnd FILL
XFILL_1__915_ vdd gnd FILL
XFILL_1__846_ vdd gnd FILL
X_1106_ _1198_/A _1199_/B _1199_/A _1109_/B vdd gnd AOI21X1
XFILL_1__777_ vdd gnd FILL
XFILL_4__1000_ vdd gnd FILL
XFILL_1__1153_ vdd gnd FILL
X_1037_ Xin[2] Cin[5] _1223_/A vdd gnd NAND2X1
XFILL_1__1222_ vdd gnd FILL
XFILL_1__1084_ vdd gnd FILL
XFILL_2__1262_ vdd gnd FILL
XFILL_2__1400_ vdd gnd FILL
XFILL_2__1331_ vdd gnd FILL
XFILL_0__933_ vdd gnd FILL
XFILL_0__864_ vdd gnd FILL
XFILL_4__1129_ vdd gnd FILL
XFILL_2__1193_ vdd gnd FILL
XFILL_0__795_ vdd gnd FILL
X_817_ _825_/C _820_/C vdd gnd INVX1
XFILL_3__1440_ vdd gnd FILL
XFILL_3__1371_ vdd gnd FILL
XFILL_0__1027_ vdd gnd FILL
XFILL_1__829_ vdd gnd FILL
XFILL_3__1569_ vdd gnd FILL
XFILL_1__1136_ vdd gnd FILL
XFILL_1__1205_ vdd gnd FILL
XFILL_1__1067_ vdd gnd FILL
XFILL_3__791_ vdd gnd FILL
XFILL_3__860_ vdd gnd FILL
XFILL_2__1245_ vdd gnd FILL
XFILL_2__1314_ vdd gnd FILL
XFILL_0__916_ vdd gnd FILL
XFILL_0__847_ vdd gnd FILL
XFILL_2__1176_ vdd gnd FILL
XFILL_0__778_ vdd gnd FILL
XFILL88950x7950 vdd gnd FILL
X_1440_ _1440_/A _1440_/B _1440_/C _1449_/A vdd gnd AOI21X1
X_1371_ _1371_/A _1371_/B _1371_/C _1401_/C vdd gnd OAI21X1
XFILL_3__989_ vdd gnd FILL
XFILL_3__1354_ vdd gnd FILL
XFILL_3__1423_ vdd gnd FILL
XFILL_0__1576_ vdd gnd FILL
XFILL_3__1285_ vdd gnd FILL
X_1569_ _1569_/A Yout[1] vdd gnd BUFX2
XFILL_1__1119_ vdd gnd FILL
XFILL_2__1030_ vdd gnd FILL
XFILL_3__912_ vdd gnd FILL
XFILL_3__843_ vdd gnd FILL
XFILL_3__774_ vdd gnd FILL
XFILL_0__1430_ vdd gnd FILL
XFILL_3__1070_ vdd gnd FILL
XFILL_2__1228_ vdd gnd FILL
XFILL_0__1361_ vdd gnd FILL
XFILL_0__1292_ vdd gnd FILL
XFILL_2__1159_ vdd gnd FILL
XFILL_1_BUFX2_insert15 vdd gnd FILL
X_1354_ _1354_/A _1354_/B _1354_/C _1366_/B vdd gnd OAI21X1
X_1423_ _1423_/A _1424_/B vdd gnd INVX1
X_1285_ _1357_/B _1357_/A _1299_/C _1290_/A vdd gnd NAND3X1
XFILL_2__930_ vdd gnd FILL
XFILL_3__1406_ vdd gnd FILL
XFILL_3__1337_ vdd gnd FILL
XFILL_1__1470_ vdd gnd FILL
XFILL_2__792_ vdd gnd FILL
XFILL_2__861_ vdd gnd FILL
XFILL_3__1199_ vdd gnd FILL
XFILL_3__1268_ vdd gnd FILL
XFILL_2__1013_ vdd gnd FILL
X_996_ _996_/A _996_/B _996_/C _996_/Y vdd gnd AOI21X1
XFILL_3__826_ vdd gnd FILL
X_1070_ _983_/A _1070_/B _982_/A _1157_/C vdd gnd OAI21X1
XFILL_3__1122_ vdd gnd FILL
XFILL_3__757_ vdd gnd FILL
XFILL_0__1413_ vdd gnd FILL
XFILL_3__1053_ vdd gnd FILL
XFILL_0__1275_ vdd gnd FILL
XFILL_0__1344_ vdd gnd FILL
X_1406_ _1406_/A _1406_/B _1406_/C _1459_/A vdd gnd AOI21X1
X_1268_ _1278_/C _1277_/B _1348_/B vdd gnd NAND2X1
X_1337_ _1337_/A _1392_/C _1337_/C _1343_/A vdd gnd OAI21X1
XFILL_2__913_ vdd gnd FILL
X_1199_ _1199_/A _1199_/B _1199_/C _1205_/C vdd gnd AOI21X1
XFILL_1__1453_ vdd gnd FILL
XFILL_1__1384_ vdd gnd FILL
XFILL_2__844_ vdd gnd FILL
XFILL_2__775_ vdd gnd FILL
X_850_ _903_/C _903_/A _850_/C _865_/B vdd gnd NAND3X1
X_781_ _814_/A Xin[2] Yin[2] _805_/B vdd gnd AOI21X1
XFILL_2__1562_ vdd gnd FILL
XFILL_2__1493_ vdd gnd FILL
XFILL_2_CLKBUF1_insert4 vdd gnd FILL
XFILL_0__1060_ vdd gnd FILL
XCLKBUF1_insert3 clk _1559_/CLK vdd gnd CLKBUF1
XFILL_3__809_ vdd gnd FILL
X_979_ _982_/C _982_/A _982_/B _987_/A vdd gnd AOI21X1
X_1122_ _1122_/A _1122_/B _1122_/C _1122_/D _1422_/B vdd gnd OAI22X1
XFILL_1__931_ vdd gnd FILL
XFILL_1__862_ vdd gnd FILL
XFILL_1__793_ vdd gnd FILL
XFILL_3__1105_ vdd gnd FILL
X_1053_ _1053_/A _1053_/B _1053_/C _1098_/B vdd gnd NAND3X1
XFILL_3__1036_ vdd gnd FILL
XFILL_0__1327_ vdd gnd FILL
XFILL_0__1258_ vdd gnd FILL
XFILL_0__1189_ vdd gnd FILL
XFILL_1__1505_ vdd gnd FILL
XFILL_0__880_ vdd gnd FILL
XFILL_1__1436_ vdd gnd FILL
XFILL_1__1367_ vdd gnd FILL
XFILL_1__1298_ vdd gnd FILL
XFILL_2__827_ vdd gnd FILL
XFILL_2__758_ vdd gnd FILL
X_833_ _833_/A _833_/B _833_/Y vdd gnd AND2X2
X_902_ _952_/C _927_/B _991_/A vdd gnd AND2X2
X_764_ _777_/A _768_/A vdd gnd INVX1
XFILL_2__1476_ vdd gnd FILL
XFILL_0__1112_ vdd gnd FILL
XFILL_0__1043_ vdd gnd FILL
XFILL_1__914_ vdd gnd FILL
XFILL_1__845_ vdd gnd FILL
X_1105_ _1105_/A _1105_/B _1128_/A _1109_/A vdd gnd AOI21X1
XFILL_1__776_ vdd gnd FILL
XFILL_1__1152_ vdd gnd FILL
X_1036_ _1046_/D _1036_/B _1152_/B _1152_/A vdd gnd NAND3X1
XFILL_1__1221_ vdd gnd FILL
XFILL_3__1019_ vdd gnd FILL
XFILL_1__1083_ vdd gnd FILL
XFILL_2__1330_ vdd gnd FILL
XFILL_1__1419_ vdd gnd FILL
XFILL_2__1261_ vdd gnd FILL
XFILL_0__932_ vdd gnd FILL
XFILL_0__863_ vdd gnd FILL
XFILL_2__1192_ vdd gnd FILL
XFILL_0__794_ vdd gnd FILL
XFILL88350x85950 vdd gnd FILL
X_816_ _825_/C _825_/B _825_/A _877_/A vdd gnd NAND3X1
XFILL_3__1370_ vdd gnd FILL
XFILL_2__1459_ vdd gnd FILL
XFILL_0__1026_ vdd gnd FILL
X_1019_ _1019_/A _1121_/B _945_/Y _1020_/A vdd gnd AOI21X1
XFILL_1__828_ vdd gnd FILL
XFILL_1__759_ vdd gnd FILL
XFILL_3__1568_ vdd gnd FILL
XFILL_3__1499_ vdd gnd FILL
XFILL_1__1204_ vdd gnd FILL
XFILL_1__1066_ vdd gnd FILL
XFILL_1__1135_ vdd gnd FILL
XFILL_3__790_ vdd gnd FILL
XFILL_2__1244_ vdd gnd FILL
XFILL_2__1313_ vdd gnd FILL
XFILL_2__1175_ vdd gnd FILL
XFILL_0__915_ vdd gnd FILL
XFILL_0__846_ vdd gnd FILL
XFILL_0__777_ vdd gnd FILL
XFILL_3__988_ vdd gnd FILL
X_1370_ _1370_/A _1370_/B _1405_/A _1409_/C vdd gnd OAI21X1
XFILL_0__1575_ vdd gnd FILL
XFILL_3__1353_ vdd gnd FILL
XFILL_3__1422_ vdd gnd FILL
XFILL_3__1284_ vdd gnd FILL
XFILL_4__824_ vdd gnd FILL
XFILL_0__1009_ vdd gnd FILL
X_1568_ _1568_/A Yout[0] vdd gnd BUFX2
X_1499_ _1499_/A _1499_/B _1506_/C vdd gnd NAND2X1
XFILL_1__1118_ vdd gnd FILL
XFILL_1__1049_ vdd gnd FILL
XFILL89550x7950 vdd gnd FILL
XFILL_3__911_ vdd gnd FILL
XFILL_3__842_ vdd gnd FILL
XFILL88650x74250 vdd gnd FILL
XFILL_3__773_ vdd gnd FILL
XFILL_2__1158_ vdd gnd FILL
XFILL_2__1227_ vdd gnd FILL
XFILL_0__1360_ vdd gnd FILL
XFILL_0__1291_ vdd gnd FILL
XFILL_0__829_ vdd gnd FILL
XFILL_2__1089_ vdd gnd FILL
X_1422_ _1422_/A _1422_/B _1511_/C _1512_/B vdd gnd NAND3X1
XFILL_1_BUFX2_insert16 vdd gnd FILL
X_1353_ _1413_/B _1413_/A _1413_/C _1414_/C vdd gnd NAND3X1
XFILL_3__1405_ vdd gnd FILL
X_1284_ _1299_/B _1299_/A _1357_/C _1290_/B vdd gnd OAI21X1
XFILL_2__860_ vdd gnd FILL
XFILL_3__1267_ vdd gnd FILL
XFILL_0__1489_ vdd gnd FILL
XFILL_3__1336_ vdd gnd FILL
XFILL_2__791_ vdd gnd FILL
XFILL_3__1198_ vdd gnd FILL
XFILL_2__1012_ vdd gnd FILL
XFILL_2__989_ vdd gnd FILL
X_995_ _998_/C _998_/B _999_/C _996_/A vdd gnd NAND3X1
XFILL_3__825_ vdd gnd FILL
XFILL_3__756_ vdd gnd FILL
XFILL_3__1121_ vdd gnd FILL
XFILL_0__1343_ vdd gnd FILL
XFILL_0__1412_ vdd gnd FILL
XFILL_3__1052_ vdd gnd FILL
XFILL_0__1274_ vdd gnd FILL
X_1405_ _1405_/A _1406_/C vdd gnd INVX1
X_1198_ _1198_/A _1199_/C vdd gnd INVX1
XFILL_4__1230_ vdd gnd FILL
X_1267_ _1344_/B _1278_/B _1277_/B vdd gnd NAND2X1
XFILL_1__1452_ vdd gnd FILL
X_1336_ _1336_/A _1443_/B _1392_/C vdd gnd AND2X2
XFILL_4__1161_ vdd gnd FILL
XFILL_2__912_ vdd gnd FILL
XFILL_2__843_ vdd gnd FILL
XFILL_4__1092_ vdd gnd FILL
XFILL_1__1383_ vdd gnd FILL
XFILL_3__1319_ vdd gnd FILL
XFILL_2__774_ vdd gnd FILL
X_780_ _814_/A Xin[2] Yin[2] _805_/C vdd gnd NAND3X1
XFILL_2__1561_ vdd gnd FILL
XFILL_2_CLKBUF1_insert5 vdd gnd FILL
XFILL_4__1359_ vdd gnd FILL
XFILL_4__1428_ vdd gnd FILL
XFILL_2__1492_ vdd gnd FILL
XFILL_1__930_ vdd gnd FILL
XCLKBUF1_insert4 clk _1552_/CLK vdd gnd CLKBUF1
X_978_ _978_/A _978_/B _982_/C vdd gnd NAND2X1
XFILL_3__808_ vdd gnd FILL
X_1121_ _1121_/A _1121_/B _1122_/B vdd gnd AND2X2
XFILL_1__792_ vdd gnd FILL
XFILL_1__861_ vdd gnd FILL
X_1052_ _1052_/A _1052_/B _1052_/C _1053_/C vdd gnd OAI21X1
XFILL_3__1104_ vdd gnd FILL
XFILL_3__1035_ vdd gnd FILL
XFILL_0__1326_ vdd gnd FILL
XFILL_0__1257_ vdd gnd FILL
XFILL_0__1188_ vdd gnd FILL
XFILL_1__1504_ vdd gnd FILL
X_1319_ _1371_/A _1371_/B _1319_/C _1326_/B vdd gnd NOR3X1
XFILL_1__1435_ vdd gnd FILL
XFILL_2__826_ vdd gnd FILL
XFILL_1__1366_ vdd gnd FILL
XFILL_1__1297_ vdd gnd FILL
X_901_ _901_/A _901_/B _901_/C _927_/B vdd gnd NAND3X1
XFILL_2__757_ vdd gnd FILL
X_832_ _832_/A _941_/D _832_/C _833_/B vdd gnd OAI21X1
X_763_ Xin[0] Cin[1] _777_/A vdd gnd NAND2X1
XFILL_2__1475_ vdd gnd FILL
XFILL_0__1111_ vdd gnd FILL
XFILL_0__1042_ vdd gnd FILL
XFILL_1__913_ vdd gnd FILL
XFILL_1__844_ vdd gnd FILL
X_1104_ _997_/Y _999_/Y _1104_/C _1110_/C vdd gnd AOI21X1
XFILL_1__775_ vdd gnd FILL
X_1035_ _861_/A _886_/B _1129_/A _1046_/D vdd gnd OAI21X1
XFILL_4__986_ vdd gnd FILL
XFILL_3__1018_ vdd gnd FILL
XFILL_1__1082_ vdd gnd FILL
XFILL_1__1151_ vdd gnd FILL
XFILL_1__1220_ vdd gnd FILL
XFILL_0__1309_ vdd gnd FILL
XFILL_0__931_ vdd gnd FILL
XFILL_2__1191_ vdd gnd FILL
XFILL_1__1349_ vdd gnd FILL
XFILL_1__1418_ vdd gnd FILL
XFILL_2__1260_ vdd gnd FILL
XFILL_2__809_ vdd gnd FILL
XFILL_0__862_ vdd gnd FILL
XFILL_0__793_ vdd gnd FILL
X_815_ _837_/A _818_/B _818_/A _825_/A vdd gnd NAND3X1
XFILL_2__1458_ vdd gnd FILL
XFILL_2__1389_ vdd gnd FILL
XFILL_0__1025_ vdd gnd FILL
XFILL_1__827_ vdd gnd FILL
XFILL_3__1567_ vdd gnd FILL
X_1018_ _1122_/D _1020_/B vdd gnd INVX1
XFILL_1__758_ vdd gnd FILL
XFILL_1__1203_ vdd gnd FILL
XFILL_3__1498_ vdd gnd FILL
XFILL_1__1065_ vdd gnd FILL
XFILL_1__1134_ vdd gnd FILL
XFILL_2__1312_ vdd gnd FILL
XFILL_0__914_ vdd gnd FILL
XFILL_2__1174_ vdd gnd FILL
XFILL_2__1243_ vdd gnd FILL
XFILL_0__845_ vdd gnd FILL
XFILL_0__776_ vdd gnd FILL
XFILL_3__987_ vdd gnd FILL
XFILL_3__1421_ vdd gnd FILL
XFILL_0__1574_ vdd gnd FILL
XFILL_3__1352_ vdd gnd FILL
XFILL_3__1283_ vdd gnd FILL
XFILL_0__1008_ vdd gnd FILL
X_1567_ _1567_/A Xout[7] vdd gnd BUFX2
X_1498_ Yin[13] _1498_/B _1499_/B vdd gnd NAND2X1
XFILL_1__1117_ vdd gnd FILL
XFILL_1__1048_ vdd gnd FILL
XFILL_3__910_ vdd gnd FILL
XFILL_3__841_ vdd gnd FILL
XFILL_3__772_ vdd gnd FILL
XFILL88950x58650 vdd gnd FILL
XFILL_2__1088_ vdd gnd FILL
XFILL_2__1157_ vdd gnd FILL
XFILL_2__1226_ vdd gnd FILL
XFILL_0__1290_ vdd gnd FILL
XFILL_0__828_ vdd gnd FILL
XFILL_0__759_ vdd gnd FILL
X_1421_ _1421_/A _1423_/A _1511_/C vdd gnd NOR2X1
XFILL_1_BUFX2_insert17 vdd gnd FILL
XFILL_3__1404_ vdd gnd FILL
X_1352_ _1360_/C _1360_/B _1414_/A _1356_/A vdd gnd AOI21X1
X_1283_ _1300_/A _1358_/A vdd gnd INVX1
XFILL_4__806_ vdd gnd FILL
XFILL_3__1197_ vdd gnd FILL
XFILL_0__1488_ vdd gnd FILL
XFILL_3__1335_ vdd gnd FILL
XFILL_3__1266_ vdd gnd FILL
XFILL_2__790_ vdd gnd FILL
XFILL_2__1011_ vdd gnd FILL
XFILL_2__988_ vdd gnd FILL
X_994_ _994_/A _994_/B _994_/C _998_/B vdd gnd NAND3X1
XFILL_3__824_ vdd gnd FILL
XFILL_3__1120_ vdd gnd FILL
XFILL_3__1051_ vdd gnd FILL
XFILL_0__1273_ vdd gnd FILL
XFILL_0__1342_ vdd gnd FILL
XFILL_0__1411_ vdd gnd FILL
XFILL_2__1209_ vdd gnd FILL
X_1404_ _1409_/C _1459_/B _1416_/C vdd gnd NAND2X1
X_1335_ Yin[10] _1337_/C vdd gnd INVX1
X_1197_ _1205_/A _1205_/B _1217_/C _1211_/B vdd gnd OAI21X1
XFILL_1__1451_ vdd gnd FILL
XFILL_1__1382_ vdd gnd FILL
X_1266_ _1266_/A _1266_/B _1266_/C _1278_/C vdd gnd AOI21X1
XFILL_3__1318_ vdd gnd FILL
XFILL_2__911_ vdd gnd FILL
XFILL_2__842_ vdd gnd FILL
XFILL_2__773_ vdd gnd FILL
XFILL_3__1249_ vdd gnd FILL
XFILL_2__1560_ vdd gnd FILL
XFILL_2__1491_ vdd gnd FILL
XCLKBUF1_insert5 clk _1551_/CLK vdd gnd CLKBUF1
X_977_ _977_/A Xin[6] Yin[6] _982_/A vdd gnd NAND3X1
XFILL_1__860_ vdd gnd FILL
XFILL_3__807_ vdd gnd FILL
X_1120_ _1120_/A _1122_/A vdd gnd INVX1
XFILL_1__791_ vdd gnd FILL
X_1051_ _1152_/A _1051_/B _1051_/C _1053_/B vdd gnd NAND3X1
XFILL_3__1103_ vdd gnd FILL
XFILL_3__1034_ vdd gnd FILL
XFILL_0__1325_ vdd gnd FILL
XFILL_0__1256_ vdd gnd FILL
XFILL_0__1187_ vdd gnd FILL
XFILL_1__989_ vdd gnd FILL
X_1318_ _1371_/C _1318_/B _1318_/C _1326_/A vdd gnd AOI21X1
XFILL_4__1143_ vdd gnd FILL
XFILL_4__1212_ vdd gnd FILL
XFILL_4__1074_ vdd gnd FILL
XFILL_1__1434_ vdd gnd FILL
XFILL_1__1365_ vdd gnd FILL
XFILL_1__1503_ vdd gnd FILL
X_1249_ _1249_/A Cin[4] _1316_/A vdd gnd NAND2X1
XFILL_2__825_ vdd gnd FILL
XFILL_2__756_ vdd gnd FILL
XFILL_1__1296_ vdd gnd FILL
X_831_ _881_/B _833_/A vdd gnd INVX1
X_900_ Xin[2] Cin[3] _952_/B _901_/C vdd gnd NAND3X1
X_762_ _762_/A _773_/C _762_/Y vdd gnd NOR2X1
XFILL_2__1474_ vdd gnd FILL
XFILL_0__1110_ vdd gnd FILL
XFILL_0__1041_ vdd gnd FILL
XFILL_1__912_ vdd gnd FILL
XFILL_3__1583_ vdd gnd FILL
XFILL_1__843_ vdd gnd FILL
X_1103_ _998_/Y _1104_/C vdd gnd INVX1
XFILL_1__774_ vdd gnd FILL
X_1034_ Xin[1] Cin[6] _1129_/A vdd gnd NAND2X1
XFILL_3__1017_ vdd gnd FILL
XFILL_1__1081_ vdd gnd FILL
XFILL_1__1150_ vdd gnd FILL
XFILL_0__1308_ vdd gnd FILL
XFILL_0__1239_ vdd gnd FILL
XFILL_0__930_ vdd gnd FILL
XFILL_1__1417_ vdd gnd FILL
XFILL_1__1348_ vdd gnd FILL
XFILL_2__1190_ vdd gnd FILL
XFILL_2__808_ vdd gnd FILL
XFILL_0__792_ vdd gnd FILL
XFILL_0__861_ vdd gnd FILL
XFILL_1__1279_ vdd gnd FILL
X_814_ _814_/A _836_/B _814_/C _818_/A vdd gnd NAND3X1
XFILL_2__1457_ vdd gnd FILL
XFILL_2__1388_ vdd gnd FILL
X_1583_ _1583_/A Yout[9] vdd gnd BUFX2
XFILL_0__1024_ vdd gnd FILL
XFILL_3__1566_ vdd gnd FILL
XFILL_1__826_ vdd gnd FILL
XFILL_3__1497_ vdd gnd FILL
X_1017_ _945_/Y _1121_/B _1019_/A _1122_/D vdd gnd NAND3X1
XFILL_1__757_ vdd gnd FILL
XFILL_1__1202_ vdd gnd FILL
XFILL_1__1064_ vdd gnd FILL
XFILL_1__1133_ vdd gnd FILL
XFILL_2__1242_ vdd gnd FILL
XFILL_2__1311_ vdd gnd FILL
XFILL_0__844_ vdd gnd FILL
XFILL_0__913_ vdd gnd FILL
XFILL_2__1173_ vdd gnd FILL
XFILL_0__775_ vdd gnd FILL
XFILL_3__986_ vdd gnd FILL
XFILL_3__1351_ vdd gnd FILL
XFILL_3__1420_ vdd gnd FILL
XFILL_0__1573_ vdd gnd FILL
XFILL_2__1509_ vdd gnd FILL
XFILL_3__1282_ vdd gnd FILL
XFILL_0__1007_ vdd gnd FILL
XFILL89550x150 vdd gnd FILL
X_1566_ _1566_/A Xout[6] vdd gnd BUFX2
XFILL_4__1460_ vdd gnd FILL
X_1497_ _1497_/A _1497_/B _1499_/A vdd gnd NAND2X1
XFILL_1__809_ vdd gnd FILL
XFILL_4__1391_ vdd gnd FILL
XFILL_1__1116_ vdd gnd FILL
XFILL_1__1047_ vdd gnd FILL
XFILL_3__840_ vdd gnd FILL
XFILL_3__771_ vdd gnd FILL
XFILL_2__1225_ vdd gnd FILL
XFILL_0__827_ vdd gnd FILL
XFILL_2__1087_ vdd gnd FILL
XFILL_2__1156_ vdd gnd FILL
XFILL_0__758_ vdd gnd FILL
X_1351_ _1413_/B _1413_/A _1354_/C _1360_/B vdd gnd NAND3X1
X_1420_ _1420_/A _1424_/A _1555_/D vdd gnd XOR2X1
XFILL_3__969_ vdd gnd FILL
XFILL_3__1334_ vdd gnd FILL
XFILL_3__1403_ vdd gnd FILL
X_1282_ _1300_/A _1358_/C _1300_/B _1287_/B vdd gnd NAND3X1
XFILL_3__1196_ vdd gnd FILL
XFILL_0__1487_ vdd gnd FILL
XFILL_3__1265_ vdd gnd FILL
X_1549_ _944_/Y _1549_/CLK _1549_/Q vdd gnd DFFPOSX1
XFILL_2__987_ vdd gnd FILL
XFILL_2__1010_ vdd gnd FILL
XBUFX2_insert10 Xin[3] _1305_/A vdd gnd BUFX2
X_993_ _993_/A _993_/B _993_/C _998_/C vdd gnd NAND3X1
XFILL_3__823_ vdd gnd FILL
XFILL_3_CLKBUF1_insert0 vdd gnd FILL
XFILL_0__1410_ vdd gnd FILL
XFILL_2__1208_ vdd gnd FILL
XFILL_3__1050_ vdd gnd FILL
XFILL_0__1272_ vdd gnd FILL
XFILL_0__1341_ vdd gnd FILL
XFILL_2__1139_ vdd gnd FILL
X_1334_ Yin[10] _1334_/B _1396_/A vdd gnd NAND2X1
X_1403_ _1430_/A _1409_/B _1459_/B vdd gnd NAND2X1
X_1265_ _1265_/A _1265_/B _1265_/C _1266_/C vdd gnd AOI21X1
XFILL_2__910_ vdd gnd FILL
X_1196_ _1275_/A _1276_/B _1276_/A _1205_/B vdd gnd AOI21X1
XFILL_1__1450_ vdd gnd FILL
XFILL_3__1317_ vdd gnd FILL
XFILL_1__1381_ vdd gnd FILL
XFILL_2__841_ vdd gnd FILL
XFILL_2__772_ vdd gnd FILL
XFILL_3__1248_ vdd gnd FILL
XFILL_3__1179_ vdd gnd FILL
XFILL_2__1490_ vdd gnd FILL
XFILL_1__1579_ vdd gnd FILL
X_976_ _983_/A _982_/B vdd gnd INVX1
XFILL_3__806_ vdd gnd FILL
XFILL_1__790_ vdd gnd FILL
XFILL_3__1102_ vdd gnd FILL
X_1050_ _1050_/A _1125_/A _1050_/C _1125_/B vdd gnd NAND3X1
XFILL_3__1033_ vdd gnd FILL
XFILL_0__1186_ vdd gnd FILL
XFILL_0__1255_ vdd gnd FILL
XFILL_0__1324_ vdd gnd FILL
XFILL_1__988_ vdd gnd FILL
XFILL_1__1502_ vdd gnd FILL
X_1317_ _1325_/B _1325_/A _1326_/C _1367_/A vdd gnd NAND3X1
X_1248_ _1248_/A _1248_/B _1248_/C _1277_/A vdd gnd OAI21X1
XFILL_1__1433_ vdd gnd FILL
XFILL_1__1364_ vdd gnd FILL
XFILL_1__1295_ vdd gnd FILL
X_1179_ _1190_/C _1190_/A _1248_/A _1195_/A vdd gnd AOI21X1
XFILL_2__824_ vdd gnd FILL
X_830_ _832_/C _832_/A _941_/D _881_/B vdd gnd NOR3X1
X_761_ Yin[0] _761_/B _762_/A vdd gnd NOR2X1
XFILL_2__1473_ vdd gnd FILL
XFILL_0__1040_ vdd gnd FILL
XFILL_1__911_ vdd gnd FILL
XFILL_1__842_ vdd gnd FILL
X_1102_ _1208_/B _1208_/A _1208_/C _1209_/C vdd gnd NAND3X1
X_959_ _964_/C _965_/C _963_/C vdd gnd NAND2X1
XFILL_1__773_ vdd gnd FILL
XFILL_3__1582_ vdd gnd FILL
X_1033_ _951_/B _1039_/B _1152_/B vdd gnd NAND2X1
XFILL_3__1016_ vdd gnd FILL
XFILL_1__1080_ vdd gnd FILL
XFILL_0__1238_ vdd gnd FILL
XFILL_0__1307_ vdd gnd FILL
XFILL_0__1169_ vdd gnd FILL
XFILL_0__860_ vdd gnd FILL
XFILL_1__1347_ vdd gnd FILL
XFILL_1__1416_ vdd gnd FILL
XFILL_1__1278_ vdd gnd FILL
XFILL_2__807_ vdd gnd FILL
XFILL_0__791_ vdd gnd FILL
X_813_ Yin[3] _813_/B _818_/B vdd gnd NAND2X1
XFILL_2__1456_ vdd gnd FILL
XFILL_2__1387_ vdd gnd FILL
XFILL_0__989_ vdd gnd FILL
XFILL_0__1023_ vdd gnd FILL
X_1582_ _1582_/A Yout[8] vdd gnd BUFX2
XFILL_3__1565_ vdd gnd FILL
XFILL_1__825_ vdd gnd FILL
XFILL_1__756_ vdd gnd FILL
XFILL_3__1496_ vdd gnd FILL
X_1016_ _1016_/A _1016_/B _1016_/C _1121_/B vdd gnd NAND3X1
XFILL_4__967_ vdd gnd FILL
XFILL_4__898_ vdd gnd FILL
XFILL_1__1201_ vdd gnd FILL
XFILL_1__1132_ vdd gnd FILL
XFILL_1__1063_ vdd gnd FILL
XFILL_2__1310_ vdd gnd FILL
XFILL_2__1241_ vdd gnd FILL
XFILL_0__912_ vdd gnd FILL
XFILL_0__843_ vdd gnd FILL
XFILL_2__1172_ vdd gnd FILL
XFILL_3__985_ vdd gnd FILL
XFILL_0__774_ vdd gnd FILL
XFILL_3__1350_ vdd gnd FILL
XFILL_0__1572_ vdd gnd FILL
XFILL_2__1508_ vdd gnd FILL
XFILL_3__1281_ vdd gnd FILL
XFILL_2__1439_ vdd gnd FILL
XFILL_0__1006_ vdd gnd FILL
X_1565_ _1565_/A Xout[5] vdd gnd BUFX2
X_1496_ _1506_/A _1506_/B _1500_/B vdd gnd NAND2X1
XFILL_1__808_ vdd gnd FILL
XFILL_3__1479_ vdd gnd FILL
XFILL_1__1115_ vdd gnd FILL
XFILL_1__1046_ vdd gnd FILL
XFILL_3__770_ vdd gnd FILL
XFILL_2__1155_ vdd gnd FILL
XFILL_2__1224_ vdd gnd FILL
XFILL_0__826_ vdd gnd FILL
XFILL_0__757_ vdd gnd FILL
XFILL_2__1086_ vdd gnd FILL
XFILL_3__968_ vdd gnd FILL
X_1350_ _1370_/A _1370_/B _1413_/A vdd gnd NAND2X1
X_1281_ _1299_/A _1299_/B _1299_/C _1300_/B vdd gnd OAI21X1
XFILL_3__899_ vdd gnd FILL
XFILL_3__1264_ vdd gnd FILL
XFILL_3__1402_ vdd gnd FILL
XFILL_3__1333_ vdd gnd FILL
XFILL_3__1195_ vdd gnd FILL
XFILL_0__1486_ vdd gnd FILL
X_1548_ _1548_/D _1549_/CLK _1548_/Q vdd gnd DFFPOSX1
XFILL_4__1373_ vdd gnd FILL
XFILL_4__1442_ vdd gnd FILL
X_1479_ _1479_/A _1480_/B vdd gnd INVX1
XFILL_4__1511_ vdd gnd FILL
XFILL89250x19650 vdd gnd FILL
XFILL_2__986_ vdd gnd FILL
XBUFX2_insert11 Xin[3] _961_/A vdd gnd BUFX2
XFILL_1__1029_ vdd gnd FILL
XFILL_3__822_ vdd gnd FILL
X_992_ _992_/A _992_/B _993_/C vdd gnd AND2X2
XFILL_3_CLKBUF1_insert1 vdd gnd FILL
XFILL_2__1207_ vdd gnd FILL
XFILL_2__1138_ vdd gnd FILL
XFILL_0__1271_ vdd gnd FILL
XFILL_0__1340_ vdd gnd FILL
XFILL_0__809_ vdd gnd FILL
XFILL_2__1069_ vdd gnd FILL
X_1402_ _1402_/A _1402_/B _1402_/C _1409_/B vdd gnd OAI21X1
X_1264_ _1344_/B _1278_/B _1277_/A _1303_/C vdd gnd NAND3X1
X_1333_ _1336_/A _1443_/B _1337_/A _1334_/B vdd gnd AOI21X1
X_1195_ _1195_/A _1195_/B _1195_/C _1276_/B vdd gnd OAI21X1
XFILL_1__1380_ vdd gnd FILL
XFILL_3__1316_ vdd gnd FILL
XFILL_3__1247_ vdd gnd FILL
XFILL_0__1469_ vdd gnd FILL
XFILL_2__840_ vdd gnd FILL
XFILL_2__771_ vdd gnd FILL
XFILL_3__1178_ vdd gnd FILL
XFILL_1__1578_ vdd gnd FILL
XFILL_2__969_ vdd gnd FILL
X_975_ _983_/C _983_/B _983_/A _987_/B vdd gnd AOI21X1
XFILL_3__805_ vdd gnd FILL
XFILL_3__1101_ vdd gnd FILL
XFILL_0__1323_ vdd gnd FILL
XFILL_3__1032_ vdd gnd FILL
XFILL_0__1185_ vdd gnd FILL
XFILL_0__1254_ vdd gnd FILL
XFILL_1__987_ vdd gnd FILL
XFILL_1__1432_ vdd gnd FILL
XFILL_1__1501_ vdd gnd FILL
X_1316_ _1316_/A _1316_/B _1316_/C _1326_/C vdd gnd OAI21X1
X_1247_ _1247_/A _1247_/B _1248_/B vdd gnd NOR2X1
X_1178_ _1265_/A _1265_/B _1247_/B _1190_/C vdd gnd NAND3X1
XFILL_2__823_ vdd gnd FILL
XFILL_1__1294_ vdd gnd FILL
XFILL_1__1363_ vdd gnd FILL
X_760_ _760_/A _773_/C vdd gnd INVX1
XFILL_2__1472_ vdd gnd FILL
XFILL_1__910_ vdd gnd FILL
XFILL_1__841_ vdd gnd FILL
XFILL_3__1581_ vdd gnd FILL
X_889_ _946_/B _951_/A _938_/C vdd gnd XOR2X1
X_1101_ _1128_/A _1105_/B _1105_/A _1208_/B vdd gnd NAND3X1
XFILL_1__772_ vdd gnd FILL
X_958_ Cin[2] Xin[4] _965_/C vdd gnd AND2X2
X_1032_ Xin[2] Cin[5] _1039_/B vdd gnd AND2X2
XFILL_3__1015_ vdd gnd FILL
XFILL_0__1306_ vdd gnd FILL
XFILL_0__1099_ vdd gnd FILL
XFILL_0__1237_ vdd gnd FILL
XFILL_0__1168_ vdd gnd FILL
XFILL_4__1124_ vdd gnd FILL
XFILL_0_BUFX2_insert10 vdd gnd FILL
XFILL_1__1415_ vdd gnd FILL
XFILL_2__806_ vdd gnd FILL
XFILL_4__1055_ vdd gnd FILL
XFILL_0__790_ vdd gnd FILL
XFILL_1__1346_ vdd gnd FILL
XFILL_1__1277_ vdd gnd FILL
X_812_ _847_/A _848_/A _848_/B _825_/B vdd gnd NAND3X1
XFILL88050x35250 vdd gnd FILL
XFILL_2__1455_ vdd gnd FILL
XFILL_2__1386_ vdd gnd FILL
XFILL_0__988_ vdd gnd FILL
XFILL_0__1022_ vdd gnd FILL
X_1581_ _1581_/A Yout[7] vdd gnd BUFX2
X_1015_ _946_/Y _1015_/B _1015_/C _1016_/C vdd gnd NAND3X1
XFILL_1__824_ vdd gnd FILL
XFILL_3__1564_ vdd gnd FILL
XFILL_3__1495_ vdd gnd FILL
XFILL_1__1062_ vdd gnd FILL
XFILL_1__1131_ vdd gnd FILL
XFILL_1__1200_ vdd gnd FILL
XFILL_2__1171_ vdd gnd FILL
XFILL_2__1240_ vdd gnd FILL
XFILL_0__911_ vdd gnd FILL
XFILL_0__842_ vdd gnd FILL
XFILL_0__773_ vdd gnd FILL
XFILL_1__1329_ vdd gnd FILL
XFILL_3__984_ vdd gnd FILL
XFILL_0__1571_ vdd gnd FILL
XFILL_3__1280_ vdd gnd FILL
XFILL_2__1438_ vdd gnd FILL
XFILL_2__1507_ vdd gnd FILL
XFILL_4__820_ vdd gnd FILL
XFILL_2__1369_ vdd gnd FILL
XFILL_0__1005_ vdd gnd FILL
X_1564_ _1564_/A Xout[4] vdd gnd BUFX2
XFILL_1__807_ vdd gnd FILL
X_1495_ _1507_/B _1495_/B _1495_/C _1506_/B vdd gnd OAI21X1
XFILL_3__1478_ vdd gnd FILL
XFILL_3_BUFX2_insert6 vdd gnd FILL
XFILL_1__1114_ vdd gnd FILL
XFILL_1__1045_ vdd gnd FILL
XFILL_4__949_ vdd gnd FILL
XFILL_2__1154_ vdd gnd FILL
XFILL_2__1223_ vdd gnd FILL
XFILL_0__825_ vdd gnd FILL
XFILL_0__756_ vdd gnd FILL
XFILL_2__1085_ vdd gnd FILL
XFILL_3__967_ vdd gnd FILL
XFILL_3__898_ vdd gnd FILL
XFILL_3__1401_ vdd gnd FILL
X_1280_ _1301_/B _1280_/B _1348_/B _1303_/C _1299_/B vdd gnd AOI22X1
XFILL_3__1194_ vdd gnd FILL
XFILL_0__1485_ vdd gnd FILL
XFILL_3__1263_ vdd gnd FILL
XFILL_3__1332_ vdd gnd FILL
X_1547_ _833_/Y _1549_/CLK _1547_/Q vdd gnd DFFPOSX1
X_1478_ _1478_/A _1478_/B _1478_/C _1480_/A vdd gnd OAI21X1
XFILL_2__985_ vdd gnd FILL
XFILL_1__1028_ vdd gnd FILL
XBUFX2_insert12 Xin[3] _895_/A vdd gnd BUFX2
X_991_ _991_/A _991_/B _991_/C _999_/C vdd gnd AOI21X1
XFILL_3__821_ vdd gnd FILL
XFILL_3_CLKBUF1_insert2 vdd gnd FILL
XFILL_2__1068_ vdd gnd FILL
XFILL_2__1206_ vdd gnd FILL
XFILL_2__1137_ vdd gnd FILL
XFILL_0__1270_ vdd gnd FILL
XFILL_0__808_ vdd gnd FILL
X_1401_ _1401_/A _1428_/A _1401_/C _1402_/B vdd gnd AOI21X1
X_1194_ _1220_/B _1220_/C _1220_/A _1275_/A vdd gnd NAND3X1
X_1263_ _1263_/A _1263_/B _1278_/B vdd gnd NAND2X1
X_1332_ Cin[4] Xin[7] _1443_/B vdd gnd AND2X2
XFILL_3__1177_ vdd gnd FILL
XFILL_3__1246_ vdd gnd FILL
XFILL_3__1315_ vdd gnd FILL
XFILL_0__1468_ vdd gnd FILL
XFILL_2__770_ vdd gnd FILL
XFILL_0__1399_ vdd gnd FILL
XFILL_1__1577_ vdd gnd FILL
XFILL_4__1424_ vdd gnd FILL
XFILL_4__1355_ vdd gnd FILL
XFILL_2__968_ vdd gnd FILL
XFILL_2__899_ vdd gnd FILL
X_974_ _977_/A Xin[6] _978_/A _983_/C vdd gnd NAND3X1
XFILL_3__804_ vdd gnd FILL
XFILL_3__1100_ vdd gnd FILL
XFILL_3__1031_ vdd gnd FILL
XFILL_0__1322_ vdd gnd FILL
XFILL_4_BUFX2_insert13 vdd gnd FILL
XFILL_0__1253_ vdd gnd FILL
XFILL_0__1184_ vdd gnd FILL
XFILL_1__986_ vdd gnd FILL
X_1315_ _1336_/A _1320_/B _1316_/B vdd gnd NOR2X1
X_1177_ _1181_/A _1329_/B _1247_/B vdd gnd NOR2X1
XFILL_1__1362_ vdd gnd FILL
X_1246_ _1301_/B _1280_/B _1348_/A vdd gnd AND2X2
XFILL_1__1500_ vdd gnd FILL
XFILL_1__1431_ vdd gnd FILL
XFILL_2__822_ vdd gnd FILL
XFILL_1__1293_ vdd gnd FILL
XFILL_3__1229_ vdd gnd FILL
XFILL_2__1471_ vdd gnd FILL
XFILL88950x54750 vdd gnd FILL
XFILL_3__1580_ vdd gnd FILL
XFILL_1__840_ vdd gnd FILL
X_957_ _966_/A _963_/B vdd gnd INVX1
X_888_ _888_/A _952_/A _888_/C _946_/B vdd gnd OAI21X1
X_1100_ _1127_/A _1127_/B _1100_/C _1105_/A vdd gnd NAND3X1
XFILL_1__771_ vdd gnd FILL
X_1031_ _1045_/C _1036_/B vdd gnd INVX1
XFILL_3__1014_ vdd gnd FILL
XFILL_0__1236_ vdd gnd FILL
XFILL_0__1305_ vdd gnd FILL
XFILL_0__1098_ vdd gnd FILL
XFILL_0__1167_ vdd gnd FILL
XFILL_1__969_ vdd gnd FILL
XFILL_0_BUFX2_insert11 vdd gnd FILL
XFILL_1__1345_ vdd gnd FILL
XFILL_1__1414_ vdd gnd FILL
X_1229_ _1304_/A _1237_/C vdd gnd INVX1
XFILL_2__805_ vdd gnd FILL
XFILL_1__1276_ vdd gnd FILL
X_811_ _814_/C _813_/B _848_/B vdd gnd NAND2X1
XFILL_2__1454_ vdd gnd FILL
XFILL88350x19650 vdd gnd FILL
XFILL_2__1385_ vdd gnd FILL
X_1580_ _1580_/A Yout[6] vdd gnd BUFX2
XFILL_0__987_ vdd gnd FILL
XFILL_0__1021_ vdd gnd FILL
XFILL_1__823_ vdd gnd FILL
XFILL_3__1563_ vdd gnd FILL
X_1014_ _1114_/A _1113_/A _1114_/B _1016_/B vdd gnd NAND3X1
XFILL_3__1494_ vdd gnd FILL
XFILL_1__1061_ vdd gnd FILL
XFILL_1__1130_ vdd gnd FILL
XFILL_0__1219_ vdd gnd FILL
XFILL_0__910_ vdd gnd FILL
XFILL_4__1106_ vdd gnd FILL
XFILL_4__1037_ vdd gnd FILL
XFILL_1__1328_ vdd gnd FILL
XFILL_2__1170_ vdd gnd FILL
XFILL_0__841_ vdd gnd FILL
XFILL_0__772_ vdd gnd FILL
XFILL_1__1259_ vdd gnd FILL
XFILL88950x78150 vdd gnd FILL
XFILL_3__983_ vdd gnd FILL
XFILL_2__1437_ vdd gnd FILL
XFILL_2__1506_ vdd gnd FILL
XFILL_0__1570_ vdd gnd FILL
XFILL_2__1368_ vdd gnd FILL
XFILL_2__1299_ vdd gnd FILL
XFILL_0__1004_ vdd gnd FILL
X_1563_ _1563_/A Xout[3] vdd gnd BUFX2
X_1494_ _1507_/C _1495_/B vdd gnd INVX1
XFILL_1__806_ vdd gnd FILL
XFILL_3__1477_ vdd gnd FILL
XFILL_3_BUFX2_insert7 vdd gnd FILL
XFILL_1__1113_ vdd gnd FILL
XFILL_1__1044_ vdd gnd FILL
XFILL_2__1222_ vdd gnd FILL
XFILL_0__824_ vdd gnd FILL
XFILL_2__1153_ vdd gnd FILL
XFILL_2__1084_ vdd gnd FILL
XFILL_3__897_ vdd gnd FILL
XFILL_3__966_ vdd gnd FILL
XFILL_3__1400_ vdd gnd FILL
XFILL_3__1331_ vdd gnd FILL
XFILL_3__1193_ vdd gnd FILL
XFILL_0__1484_ vdd gnd FILL
XFILL_3__1262_ vdd gnd FILL
X_1546_ _796_/Y _1546_/CLK _1546_/Q vdd gnd DFFPOSX1
X_1477_ _1504_/A _1477_/B _1477_/C _1482_/B vdd gnd OAI21X1
XBUFX2_insert13 Xin[3] _836_/B vdd gnd BUFX2
XFILL_2__984_ vdd gnd FILL
X_990_ _990_/A _991_/C vdd gnd INVX1
XFILL_1__1027_ vdd gnd FILL
XFILL_3__820_ vdd gnd FILL
XFILL_2__1205_ vdd gnd FILL
XFILL_3_CLKBUF1_insert3 vdd gnd FILL
XFILL_0__807_ vdd gnd FILL
XFILL_2__1067_ vdd gnd FILL
XFILL_2__1136_ vdd gnd FILL
X_1400_ _1400_/A _1400_/B _1400_/C _1402_/A vdd gnd AOI21X1
X_1331_ Cin[3] Xin[7] Cin[4] Xin[6] _1337_/A vdd gnd AOI22X1
XFILL_3__949_ vdd gnd FILL
X_1193_ _1219_/B _1193_/B _1276_/A vdd gnd AND2X2
X_1262_ _1262_/A _1263_/A vdd gnd INVX1
XFILL_3__1314_ vdd gnd FILL
XFILL_3__1245_ vdd gnd FILL
XFILL_0__1467_ vdd gnd FILL
XFILL_0__1398_ vdd gnd FILL
XFILL_3__1176_ vdd gnd FILL
X_1529_ _1545_/Q _1546_/CLK _1569_/A vdd gnd DFFPOSX1
XFILL_1__1576_ vdd gnd FILL
XFILL_4__1285_ vdd gnd FILL
XFILL_2__967_ vdd gnd FILL
XFILL_2__898_ vdd gnd FILL
X_973_ Yin[6] _978_/A vdd gnd INVX1
XFILL_3__803_ vdd gnd FILL
XFILL_3__1030_ vdd gnd FILL
XFILL_0__1252_ vdd gnd FILL
XFILL_0__1321_ vdd gnd FILL
XFILL_2__1119_ vdd gnd FILL
XFILL_0__1183_ vdd gnd FILL
XFILL_1__985_ vdd gnd FILL
X_1314_ _1318_/C _1318_/B _1371_/C _1325_/A vdd gnd NAND3X1
XFILL_0__1519_ vdd gnd FILL
X_1245_ _1245_/A _1245_/B _1245_/C _1280_/B vdd gnd NAND3X1
XFILL_1__1430_ vdd gnd FILL
XFILL_1__1361_ vdd gnd FILL
X_1176_ _1329_/B _1181_/A _1247_/A _1190_/A vdd gnd OAI21X1
XFILL_2__821_ vdd gnd FILL
XFILL_3__1159_ vdd gnd FILL
XFILL_3__1228_ vdd gnd FILL
XFILL_1__1292_ vdd gnd FILL
XFILL_2__1470_ vdd gnd FILL
X_956_ Xin[2] Cin[4] _966_/A vdd gnd NAND2X1
XFILL_1__770_ vdd gnd FILL
XFILL_4__981_ vdd gnd FILL
X_887_ Xin[2] Cin[3] _952_/A vdd gnd NAND2X1
X_1030_ Xin[0] Cin[7] _1045_/C vdd gnd NAND2X1
XFILL_3__1013_ vdd gnd FILL
XFILL_0__1235_ vdd gnd FILL
XFILL_0__1304_ vdd gnd FILL
XFILL_0__1166_ vdd gnd FILL
XFILL_0__1097_ vdd gnd FILL
XFILL_1__968_ vdd gnd FILL
XFILL_1__899_ vdd gnd FILL
XFILL_0_BUFX2_insert12 vdd gnd FILL
X_1228_ _1304_/B _1238_/C _1304_/A _1243_/C vdd gnd OAI21X1
XFILL_1__1275_ vdd gnd FILL
X_1159_ Xin[4] Cin[4] _1235_/A vdd gnd NAND2X1
XFILL_1__1344_ vdd gnd FILL
XFILL_1__1413_ vdd gnd FILL
XFILL_2__804_ vdd gnd FILL
X_810_ _912_/A _836_/B _813_/B vdd gnd NAND2X1
XFILL_2__1453_ vdd gnd FILL
XFILL_2__1384_ vdd gnd FILL
XFILL_0__1020_ vdd gnd FILL
XFILL_0__986_ vdd gnd FILL
X_939_ _939_/A _939_/B _939_/C _941_/B vdd gnd OAI21X1
XFILL_3__1562_ vdd gnd FILL
XFILL_1__822_ vdd gnd FILL
XFILL_3__1493_ vdd gnd FILL
X_1013_ _941_/A _1016_/A vdd gnd INVX1
XFILL89250x150 vdd gnd FILL
XFILL_0__1149_ vdd gnd FILL
XFILL_0__1218_ vdd gnd FILL
XFILL_1__1060_ vdd gnd FILL
XFILL_0__840_ vdd gnd FILL
XFILL_1__1327_ vdd gnd FILL
XFILL_1__1258_ vdd gnd FILL
XFILL_0__771_ vdd gnd FILL
XFILL_1__1189_ vdd gnd FILL
XFILL_3__982_ vdd gnd FILL
XFILL_2__1436_ vdd gnd FILL
XFILL_2__1367_ vdd gnd FILL
XFILL_2__1505_ vdd gnd FILL
XFILL_0__969_ vdd gnd FILL
XFILL_0__1003_ vdd gnd FILL
XFILL_2__1298_ vdd gnd FILL
X_1562_ _1562_/A Xout[2] vdd gnd BUFX2
X_1493_ Yin[14] _1495_/C vdd gnd INVX1
XFILL_1__805_ vdd gnd FILL
XFILL_3__1476_ vdd gnd FILL
XFILL_1__1112_ vdd gnd FILL
XFILL_3_BUFX2_insert8 vdd gnd FILL
XFILL_1__1043_ vdd gnd FILL
XFILL_2__1221_ vdd gnd FILL
XFILL_0__823_ vdd gnd FILL
XFILL_2__1152_ vdd gnd FILL
XFILL_2__1083_ vdd gnd FILL
XFILL_3__965_ vdd gnd FILL
XFILL_3__896_ vdd gnd FILL
XFILL_3__1330_ vdd gnd FILL
XFILL_4__801_ vdd gnd FILL
XFILL_3__1192_ vdd gnd FILL
XFILL_0__1483_ vdd gnd FILL
XFILL_2__1419_ vdd gnd FILL
XFILL_3__1261_ vdd gnd FILL
X_1545_ _774_/Y _1546_/CLK _1545_/Q vdd gnd DFFPOSX1
X_1476_ _1476_/A _1478_/C _1479_/A _1504_/A vdd gnd AOI21X1
XFILL_3__1459_ vdd gnd FILL
XFILL_2__983_ vdd gnd FILL
XBUFX2_insert14 Xin[5] _1436_/A vdd gnd BUFX2
XFILL_1__1026_ vdd gnd FILL
XFILL_3_CLKBUF1_insert4 vdd gnd FILL
XFILL_2__1204_ vdd gnd FILL
XFILL_2__1135_ vdd gnd FILL
XFILL_0__806_ vdd gnd FILL
XFILL_2__1066_ vdd gnd FILL
XFILL_3__948_ vdd gnd FILL
X_1330_ _1344_/A _1344_/B _1369_/B vdd gnd NAND2X1
X_1261_ _1261_/A _1261_/B _1263_/B vdd gnd NAND2X1
XFILL_3__879_ vdd gnd FILL
X_1192_ _1201_/C _1201_/B _1221_/A _1205_/A vdd gnd AOI21X1
XFILL_3__1244_ vdd gnd FILL
XFILL_3__1313_ vdd gnd FILL
XFILL_0__1466_ vdd gnd FILL
XFILL_0__1397_ vdd gnd FILL
XFILL_3__1175_ vdd gnd FILL
X_1528_ _1544_/Q _1546_/CLK _1568_/A vdd gnd DFFPOSX1
X_1459_ _1459_/A _1459_/B _1459_/C _1460_/A vdd gnd OAI21X1
XFILL_1__1575_ vdd gnd FILL
XFILL_1__1009_ vdd gnd FILL
XFILL_2__897_ vdd gnd FILL
XFILL_2__966_ vdd gnd FILL
X_972_ Yin[6] _978_/B _983_/B vdd gnd NAND2X1
XFILL_3__802_ vdd gnd FILL
XFILL_2__1118_ vdd gnd FILL
XFILL_0__1320_ vdd gnd FILL
XFILL_0__1251_ vdd gnd FILL
XFILL_0__1182_ vdd gnd FILL
XFILL_2__1049_ vdd gnd FILL
XFILL_1__984_ vdd gnd FILL
X_1244_ _1244_/A _1244_/B _1244_/C _1245_/C vdd gnd OAI21X1
X_1313_ _1371_/B _1318_/B vdd gnd INVX1
XFILL_0__1518_ vdd gnd FILL
XFILL_3__1227_ vdd gnd FILL
XFILL_1__1360_ vdd gnd FILL
XFILL_1__1291_ vdd gnd FILL
X_1175_ Cin[1] Xin[7] Yin[8] _1181_/A vdd gnd AOI21X1
XFILL_2__820_ vdd gnd FILL
XFILL_3__1089_ vdd gnd FILL
XFILL_3__1158_ vdd gnd FILL
XFILL_0__1449_ vdd gnd FILL
XFILL89550x85950 vdd gnd FILL
XFILL_4__1405_ vdd gnd FILL
XFILL_4__1336_ vdd gnd FILL
XFILL_4__1198_ vdd gnd FILL
XFILL_2__949_ vdd gnd FILL
XFILL_4__1267_ vdd gnd FILL
XFILL_1__1489_ vdd gnd FILL
X_955_ _955_/A _955_/B _990_/A _998_/A vdd gnd OAI21X1
X_886_ _886_/A _886_/B _951_/A vdd gnd NOR2X1
XFILL_0__1303_ vdd gnd FILL
XFILL_3__1012_ vdd gnd FILL
XFILL_0__1165_ vdd gnd FILL
XFILL_0__1234_ vdd gnd FILL
XFILL_0__1096_ vdd gnd FILL
XFILL_0_BUFX2_insert13 vdd gnd FILL
XFILL_1__967_ vdd gnd FILL
XFILL_1__898_ vdd gnd FILL
X_1158_ _1158_/A _1158_/B _1186_/A _1220_/C vdd gnd OAI21X1
X_1227_ _1227_/A _1307_/A _1238_/C vdd gnd NOR2X1
XFILL_1__1412_ vdd gnd FILL
XFILL_2__803_ vdd gnd FILL
X_1089_ _1265_/B _1157_/A _1089_/C _1094_/B vdd gnd NAND3X1
XFILL_1__1343_ vdd gnd FILL
XFILL_1__1274_ vdd gnd FILL
XFILL89250x15750 vdd gnd FILL
XFILL_2__1452_ vdd gnd FILL
XFILL_2__1383_ vdd gnd FILL
XFILL_0__985_ vdd gnd FILL
X_1012_ _1012_/A _1012_/B _941_/A _1019_/A vdd gnd OAI21X1
X_938_ _938_/A _948_/C _938_/C _939_/B vdd gnd AOI21X1
XFILL_1__821_ vdd gnd FILL
X_869_ _888_/C _869_/B _890_/A vdd gnd NAND2X1
XFILL_3__1561_ vdd gnd FILL
XFILL_3__1492_ vdd gnd FILL
XFILL_4__963_ vdd gnd FILL
XFILL_4__894_ vdd gnd FILL
XFILL_0__1148_ vdd gnd FILL
XFILL_0__1079_ vdd gnd FILL
XFILL_0__1217_ vdd gnd FILL
XFILL89250x27450 vdd gnd FILL
XFILL_0__770_ vdd gnd FILL
XFILL_1__1326_ vdd gnd FILL
XFILL_1__1257_ vdd gnd FILL
XFILL_1__1188_ vdd gnd FILL
XFILL_3__981_ vdd gnd FILL
XFILL_2__1504_ vdd gnd FILL
XFILL_2__1366_ vdd gnd FILL
XFILL_2__1297_ vdd gnd FILL
XFILL_2__1435_ vdd gnd FILL
XFILL_0__968_ vdd gnd FILL
XFILL_0__1002_ vdd gnd FILL
XFILL_0__899_ vdd gnd FILL
X_1561_ _1561_/A Xout[1] vdd gnd BUFX2
X_1492_ Yin[14] _1492_/B _1507_/C _1506_/A vdd gnd NAND3X1
XFILL_1__804_ vdd gnd FILL
XFILL_3__1475_ vdd gnd FILL
XFILL_1__1111_ vdd gnd FILL
XFILL_1__1042_ vdd gnd FILL
XFILL89250x39150 vdd gnd FILL
XFILL_3_BUFX2_insert9 vdd gnd FILL
XFILL_2__1151_ vdd gnd FILL
XFILL_2__1220_ vdd gnd FILL
XFILL_4__1018_ vdd gnd FILL
XFILL_0__822_ vdd gnd FILL
XFILL_2__1082_ vdd gnd FILL
XFILL_1__1309_ vdd gnd FILL
XFILL_3__964_ vdd gnd FILL
XFILL_3__895_ vdd gnd FILL
XFILL_0__1482_ vdd gnd FILL
XFILL_2__1418_ vdd gnd FILL
XFILL_3__1260_ vdd gnd FILL
XFILL_3__1191_ vdd gnd FILL
XFILL_2__1349_ vdd gnd FILL
X_1544_ _762_/Y _1546_/CLK _1544_/Q vdd gnd DFFPOSX1
X_1475_ _1481_/B _1477_/B vdd gnd INVX1
XFILL_2__982_ vdd gnd FILL
XFILL_3__1458_ vdd gnd FILL
XFILL_3__1389_ vdd gnd FILL
XBUFX2_insert15 Xin[5] _912_/B vdd gnd BUFX2
XFILL_1__1025_ vdd gnd FILL
XFILL_3_CLKBUF1_insert5 vdd gnd FILL
XFILL_2__1203_ vdd gnd FILL
XFILL_2__1134_ vdd gnd FILL
XFILL_0__805_ vdd gnd FILL
XFILL_2__1065_ vdd gnd FILL
XFILL_3__947_ vdd gnd FILL
XFILL_3__878_ vdd gnd FILL
X_1191_ _1220_/A _1220_/B _1195_/C _1201_/C vdd gnd NAND3X1
X_1260_ _1262_/A _1261_/A _1261_/B _1344_/B vdd gnd NAND3X1
XFILL_3__1174_ vdd gnd FILL
XFILL_3__1312_ vdd gnd FILL
XFILL_3__1243_ vdd gnd FILL
XFILL_0__1465_ vdd gnd FILL
XFILL_0__1396_ vdd gnd FILL
X_1527_ Xin[7] _1559_/CLK _1567_/A vdd gnd DFFPOSX1
XFILL_1__1574_ vdd gnd FILL
X_1458_ _1458_/A _1459_/C _1458_/C _1486_/A vdd gnd NAND3X1
X_1389_ _1401_/C _1428_/A _1401_/A _1428_/B vdd gnd NAND3X1
XFILL_2__965_ vdd gnd FILL
XFILL_1__1008_ vdd gnd FILL
XFILL_2__896_ vdd gnd FILL
X_971_ _977_/A Xin[6] _978_/B vdd gnd NAND2X1
XFILL_3__801_ vdd gnd FILL
XFILL_0__1181_ vdd gnd FILL
XFILL_2__1117_ vdd gnd FILL
XFILL_2__1048_ vdd gnd FILL
XFILL_0__1250_ vdd gnd FILL
XFILL_1__983_ vdd gnd FILL
X_1174_ _1259_/A _1329_/B vdd gnd INVX1
X_1312_ _1312_/A _1312_/B _1371_/C vdd gnd NAND2X1
X_1243_ _1243_/A _1243_/B _1243_/C _1245_/B vdd gnd NAND3X1
XFILL_3__1157_ vdd gnd FILL
XFILL_3__1226_ vdd gnd FILL
XFILL_0__1448_ vdd gnd FILL
XFILL_0__1517_ vdd gnd FILL
XFILL_1__1290_ vdd gnd FILL
XFILL_3__1088_ vdd gnd FILL
XFILL_0__1379_ vdd gnd FILL
XFILL_2__948_ vdd gnd FILL
XFILL_1__1488_ vdd gnd FILL
XFILL_2__879_ vdd gnd FILL
X_954_ _954_/A _954_/B _954_/C _955_/B vdd gnd AOI21X1
X_885_ Cin[5] _886_/B vdd gnd INVX1
XFILL_3__1011_ vdd gnd FILL
XFILL_0__1302_ vdd gnd FILL
XFILL_0__1095_ vdd gnd FILL
XFILL_0__1233_ vdd gnd FILL
XFILL_0__1164_ vdd gnd FILL
XFILL_1__966_ vdd gnd FILL
XFILL_4__1120_ vdd gnd FILL
XFILL_1__897_ vdd gnd FILL
X_1157_ _1157_/A _1265_/B _1157_/C _1158_/A vdd gnd AOI21X1
XFILL_0_BUFX2_insert14 vdd gnd FILL
X_1226_ Xin[4] Cin[6] _1307_/A vdd gnd NAND2X1
XFILL_1__1342_ vdd gnd FILL
XFILL_1__1411_ vdd gnd FILL
XFILL_3__1209_ vdd gnd FILL
XFILL_2__802_ vdd gnd FILL
X_1088_ _1088_/A _1088_/B _1157_/C _1094_/A vdd gnd OAI21X1
XFILL_4__1051_ vdd gnd FILL
XFILL_1__1273_ vdd gnd FILL
XFILL_2__1451_ vdd gnd FILL
XFILL_2__1382_ vdd gnd FILL
XFILL_4__1249_ vdd gnd FILL
XFILL_4__1318_ vdd gnd FILL
XFILL_0__984_ vdd gnd FILL
XFILL_1__820_ vdd gnd FILL
XFILL_3__1560_ vdd gnd FILL
X_937_ _937_/A _937_/B _948_/A _939_/A vdd gnd AOI21X1
X_1011_ _1114_/B _1113_/A _1114_/A _1012_/A vdd gnd AOI21X1
X_868_ _868_/A _868_/B _868_/C _869_/B vdd gnd NAND3X1
XFILL_3__1491_ vdd gnd FILL
X_799_ Cin[3] _965_/B vdd gnd INVX2
XFILL_0__1216_ vdd gnd FILL
XFILL_0__1078_ vdd gnd FILL
XFILL_0__1147_ vdd gnd FILL
XFILL_1__949_ vdd gnd FILL
X_1209_ _1209_/A _1209_/B _1209_/C _1212_/A vdd gnd OAI21X1
XFILL_1__1325_ vdd gnd FILL
XFILL_1__1187_ vdd gnd FILL
XFILL_1__1256_ vdd gnd FILL
XFILL_3__980_ vdd gnd FILL
XFILL_2__1434_ vdd gnd FILL
XFILL_2__1503_ vdd gnd FILL
XFILL_0_BUFX2_insert6 vdd gnd FILL
XFILL_2__1365_ vdd gnd FILL
XFILL_2__1296_ vdd gnd FILL
XFILL_0__1001_ vdd gnd FILL
XFILL_0__967_ vdd gnd FILL
XFILL_0__898_ vdd gnd FILL
X_1560_ _1560_/A Xout[0] vdd gnd BUFX2
XFILL_1__803_ vdd gnd FILL
X_1491_ _1504_/A _1504_/B _1501_/A vdd gnd NOR2X1
XFILL_3__1474_ vdd gnd FILL
XFILL_1__1110_ vdd gnd FILL
XFILL_1__1041_ vdd gnd FILL
XFILL_4__1583_ vdd gnd FILL
XFILL_2__1081_ vdd gnd FILL
XFILL_2__1150_ vdd gnd FILL
XFILL_1__1308_ vdd gnd FILL
XFILL_0__821_ vdd gnd FILL
XFILL_1__1239_ vdd gnd FILL
XFILL_3__963_ vdd gnd FILL
XFILL_3__894_ vdd gnd FILL
XFILL88650x85950 vdd gnd FILL
XFILL_0__1481_ vdd gnd FILL
XFILL_2__1417_ vdd gnd FILL
XFILL_3__1190_ vdd gnd FILL
XFILL_2__1348_ vdd gnd FILL
XFILL_2__1279_ vdd gnd FILL
X_1543_ _1559_/Q _1559_/CLK _1575_/A vdd gnd DFFPOSX1
X_1474_ _1476_/A _1478_/C _1479_/A _1481_/B vdd gnd NAND3X1
XFILL_2__981_ vdd gnd FILL
XFILL_3__1457_ vdd gnd FILL
XFILL_3__1388_ vdd gnd FILL
XFILL_1__1024_ vdd gnd FILL
XBUFX2_insert16 Xin[5] _1249_/A vdd gnd BUFX2
XFILL88350x15750 vdd gnd FILL
XFILL_4__1497_ vdd gnd FILL
XFILL_0__804_ vdd gnd FILL
XFILL_2__1064_ vdd gnd FILL
XFILL_2__1202_ vdd gnd FILL
XFILL_2__1133_ vdd gnd FILL
XFILL_3__877_ vdd gnd FILL
XFILL_3__946_ vdd gnd FILL
XFILL_3__1311_ vdd gnd FILL
X_1190_ _1190_/A _1248_/A _1190_/C _1220_/B vdd gnd NAND3X1
XFILL_3__1242_ vdd gnd FILL
XFILL_0__1395_ vdd gnd FILL
XFILL_0__1464_ vdd gnd FILL
XFILL_3__1173_ vdd gnd FILL
X_1526_ Xin[6] _1549_/CLK _1566_/A vdd gnd DFFPOSX1
X_1457_ _1460_/B _1460_/C _1458_/C vdd gnd NAND2X1
XFILL_1__1573_ vdd gnd FILL
X_1388_ _1392_/A _1392_/B _1391_/A _1401_/A vdd gnd OAI21X1
XFILL_3__1509_ vdd gnd FILL
XFILL_2__964_ vdd gnd FILL
XFILL_2__895_ vdd gnd FILL
X_970_ Cin[1] _970_/B _983_/A vdd gnd NAND2X1
XFILL_1__1007_ vdd gnd FILL
XFILL_3__800_ vdd gnd FILL
XFILL88950x74250 vdd gnd FILL
XFILL_4_BUFX2_insert17 vdd gnd FILL
XFILL_2__1116_ vdd gnd FILL
XFILL_2__1047_ vdd gnd FILL
XFILL_0__1180_ vdd gnd FILL
XFILL_1__982_ vdd gnd FILL
X_1311_ _1436_/A Cin[5] _1312_/B vdd gnd AND2X2
XFILL_3__929_ vdd gnd FILL
X_1242_ _1242_/A _1242_/B _1245_/A vdd gnd AND2X2
X_1173_ Cin[1] Xin[7] Yin[8] _1259_/A vdd gnd NAND3X1
XFILL_3__1087_ vdd gnd FILL
XFILL_3__1156_ vdd gnd FILL
XFILL_3__1225_ vdd gnd FILL
XFILL_0__1447_ vdd gnd FILL
XFILL_0__1516_ vdd gnd FILL
XFILL_0__1378_ vdd gnd FILL
X_1509_ _1509_/A _1509_/B _1515_/A vdd gnd XOR2X1
XFILL_1__1487_ vdd gnd FILL
XFILL_2__947_ vdd gnd FILL
XFILL_2__878_ vdd gnd FILL
X_953_ _997_/A _997_/B _996_/C vdd gnd XNOR2X1
X_884_ _884_/A _884_/B _884_/C _935_/C vdd gnd OAI21X1
XFILL_3__1010_ vdd gnd FILL
XFILL_0__1232_ vdd gnd FILL
XFILL_0__1301_ vdd gnd FILL
XFILL_0__1094_ vdd gnd FILL
XFILL_0__1163_ vdd gnd FILL
XFILL_0_BUFX2_insert15 vdd gnd FILL
XFILL_1__965_ vdd gnd FILL
XFILL_1__896_ vdd gnd FILL
X_1087_ _1095_/A _1095_/B _1158_/B vdd gnd NAND2X1
X_1156_ _1219_/B _1193_/B _1221_/A vdd gnd NAND2X1
X_1225_ _1305_/A Cin[6] Xin[4] Cin[5] _1304_/B vdd gnd AOI22X1
XFILL_1__1341_ vdd gnd FILL
XFILL_1__1410_ vdd gnd FILL
XFILL_2__801_ vdd gnd FILL
XFILL_3__1208_ vdd gnd FILL
XFILL_3__1139_ vdd gnd FILL
XFILL_1__1272_ vdd gnd FILL
XFILL_2__1450_ vdd gnd FILL
XFILL_0__983_ vdd gnd FILL
XFILL_2__1381_ vdd gnd FILL
X_936_ _936_/A _936_/B _936_/C _939_/C vdd gnd AOI21X1
XFILL_3__1490_ vdd gnd FILL
XFILL_2__1579_ vdd gnd FILL
X_798_ _829_/C _828_/A vdd gnd INVX1
X_1010_ _996_/Y _1010_/B _1010_/C _1114_/B vdd gnd OAI21X1
X_867_ _867_/A _867_/B _867_/C _888_/C vdd gnd NAND3X1
XFILL_0__1215_ vdd gnd FILL
XFILL_0__1077_ vdd gnd FILL
XFILL_0__1146_ vdd gnd FILL
XFILL_1__948_ vdd gnd FILL
XFILL_1__879_ vdd gnd FILL
X_1208_ _1208_/A _1208_/B _1208_/C _1209_/B vdd gnd AOI21X1
X_1139_ _965_/A _886_/B _1139_/C _1145_/A vdd gnd OAI21X1
XFILL_1__1255_ vdd gnd FILL
XFILL_1__1324_ vdd gnd FILL
XFILL_1__1186_ vdd gnd FILL
XFILL_0_BUFX2_insert7 vdd gnd FILL
XFILL_2__1433_ vdd gnd FILL
XFILL_2__1502_ vdd gnd FILL
XFILL_2__1364_ vdd gnd FILL
XFILL_0__1000_ vdd gnd FILL
XFILL_0__966_ vdd gnd FILL
XFILL_2__1295_ vdd gnd FILL
XFILL_0__897_ vdd gnd FILL
X_1490_ _1490_/A _1504_/B vdd gnd INVX1
X_919_ _990_/A _991_/B _991_/A _947_/A vdd gnd NAND3X1
XFILL_1__802_ vdd gnd FILL
XFILL_3__1473_ vdd gnd FILL
XFILL_4__944_ vdd gnd FILL
XFILL_4__875_ vdd gnd FILL
XFILL_1__1040_ vdd gnd FILL
XFILL_0__1129_ vdd gnd FILL
XFILL_0__820_ vdd gnd FILL
XFILL_2__1080_ vdd gnd FILL
XFILL_1__1238_ vdd gnd FILL
XFILL_1__1307_ vdd gnd FILL
XFILL_1__1169_ vdd gnd FILL
XFILL_3__962_ vdd gnd FILL
XFILL_3__893_ vdd gnd FILL
XFILL_2__1347_ vdd gnd FILL
XFILL_2__1416_ vdd gnd FILL
XFILL_0__1480_ vdd gnd FILL
XFILL_0__949_ vdd gnd FILL
XFILL_2__1278_ vdd gnd FILL
X_1542_ _1558_/Q _1559_/CLK _1574_/A vdd gnd DFFPOSX1
X_1473_ _1498_/B Yin[13] _1479_/A vdd gnd XNOR2X1
XFILL_3__1456_ vdd gnd FILL
XFILL_2__980_ vdd gnd FILL
XFILL_3__1387_ vdd gnd FILL
XBUFX2_insert17 Xin[5] _970_/B vdd gnd BUFX2
XFILL_1__1023_ vdd gnd FILL
XFILL_4__1565_ vdd gnd FILL
XFILL_2__1201_ vdd gnd FILL
XFILL_0__803_ vdd gnd FILL
XFILL_2__1063_ vdd gnd FILL
XFILL_2__1132_ vdd gnd FILL
XFILL_3__945_ vdd gnd FILL
XFILL_3__876_ vdd gnd FILL
XFILL_3__1310_ vdd gnd FILL
XFILL_3__1172_ vdd gnd FILL
XFILL_0__1394_ vdd gnd FILL
XFILL_0__1463_ vdd gnd FILL
XFILL_3__1241_ vdd gnd FILL
X_1525_ _912_/B _1551_/CLK _1565_/A vdd gnd DFFPOSX1
XFILL_4__1350_ vdd gnd FILL
X_1456_ _1465_/A _1465_/B _1456_/C _1460_/B vdd gnd NAND3X1
X_1387_ _1431_/A _1431_/B _1392_/A vdd gnd NOR2X1
XFILL_1__1572_ vdd gnd FILL
XFILL_3__1439_ vdd gnd FILL
XFILL_3__1508_ vdd gnd FILL
XFILL_4__1281_ vdd gnd FILL
XFILL_2__963_ vdd gnd FILL
XFILL_2__894_ vdd gnd FILL
XFILL_1__1006_ vdd gnd FILL
XFILL_4__1479_ vdd gnd FILL
XFILL_2__1115_ vdd gnd FILL
XFILL_2__1046_ vdd gnd FILL
XFILL_3__928_ vdd gnd FILL
XFILL_1__981_ vdd gnd FILL
X_1310_ _1371_/A _1318_/C vdd gnd INVX1
X_1241_ _1241_/A _1301_/A _1241_/C _1301_/B vdd gnd NAND3X1
XFILL_3__859_ vdd gnd FILL
XFILL_3__1224_ vdd gnd FILL
X_1172_ _1172_/A _1172_/B _1265_/A _1247_/A vdd gnd OAI21X1
XFILL_0__1515_ vdd gnd FILL
XFILL_3__1086_ vdd gnd FILL
XFILL_3__1155_ vdd gnd FILL
XFILL_0__1446_ vdd gnd FILL
XFILL_0__1377_ vdd gnd FILL
X_1439_ _1477_/C _1481_/A vdd gnd INVX1
X_1508_ _1508_/A Yin[15] _1509_/B vdd gnd XNOR2X1
XFILL_1__1486_ vdd gnd FILL
XFILL_2__877_ vdd gnd FILL
XFILL_2__946_ vdd gnd FILL
X_883_ _883_/A _940_/C vdd gnd INVX1
X_952_ _952_/A _952_/B _952_/C _997_/A vdd gnd OAI21X1
XFILL_0__1231_ vdd gnd FILL
XFILL_0__1300_ vdd gnd FILL
XFILL_0__1162_ vdd gnd FILL
XFILL_0__1093_ vdd gnd FILL
XFILL_2__1029_ vdd gnd FILL
XFILL_1__964_ vdd gnd FILL
XFILL_1__895_ vdd gnd FILL
X_1224_ Xin[2] Cin[7] _1304_/A vdd gnd NAND2X1
XFILL_0_BUFX2_insert16 vdd gnd FILL
X_1086_ _1186_/A _1187_/B _1187_/A _1127_/A vdd gnd NAND3X1
XFILL_3__1207_ vdd gnd FILL
X_1155_ _1155_/A _1155_/B _1155_/C _1193_/B vdd gnd NAND3X1
XFILL_1__1271_ vdd gnd FILL
XFILL_1__1340_ vdd gnd FILL
XFILL_3__1069_ vdd gnd FILL
XFILL_2__800_ vdd gnd FILL
XFILL_3__1138_ vdd gnd FILL
XFILL_0__1429_ vdd gnd FILL
XFILL_2__1380_ vdd gnd FILL
XFILL_0__982_ vdd gnd FILL
XFILL_1__1469_ vdd gnd FILL
XFILL_2__929_ vdd gnd FILL
X_866_ _866_/A _866_/B _866_/C _890_/B vdd gnd AOI21X1
X_935_ _935_/A _935_/B _935_/C _941_/A vdd gnd NAND3X1
XFILL_2__1578_ vdd gnd FILL
X_797_ _823_/B _797_/B _797_/C _829_/C vdd gnd OAI21X1
XFILL_0__1145_ vdd gnd FILL
XFILL_0__1214_ vdd gnd FILL
XFILL_0__1076_ vdd gnd FILL
XFILL_1__947_ vdd gnd FILL
XFILL_1__878_ vdd gnd FILL
X_1207_ _1207_/A _1207_/B _1207_/C _1213_/B vdd gnd OAI21X1
X_1069_ _1171_/A Xin[6] Yin[6] _1070_/B vdd gnd AOI21X1
XFILL_4__1101_ vdd gnd FILL
XFILL_4__1032_ vdd gnd FILL
X_1138_ _1146_/B _1146_/C _1242_/B _1242_/A vdd gnd NAND3X1
XFILL_1__1323_ vdd gnd FILL
XFILL_1__1254_ vdd gnd FILL
XFILL_1__1185_ vdd gnd FILL
XFILL_2__1501_ vdd gnd FILL
XFILL_0_BUFX2_insert8 vdd gnd FILL
XFILL_2__1294_ vdd gnd FILL
XFILL_2__1432_ vdd gnd FILL
XFILL_2__1363_ vdd gnd FILL
XFILL_0__896_ vdd gnd FILL
XFILL_0__965_ vdd gnd FILL
X_918_ _921_/A _921_/B _922_/C _991_/B vdd gnd OAI21X1
X_849_ _903_/B _849_/B _849_/C _865_/A vdd gnd OAI21X1
XFILL_1__801_ vdd gnd FILL
XFILL_3__1472_ vdd gnd FILL
XFILL_0__1128_ vdd gnd FILL
XFILL_0__1059_ vdd gnd FILL
XFILL_1__1306_ vdd gnd FILL
XFILL_1__1237_ vdd gnd FILL
XFILL_1__1168_ vdd gnd FILL
XFILL_3__961_ vdd gnd FILL
XFILL_1__1099_ vdd gnd FILL
XFILL_3__892_ vdd gnd FILL
XFILL_2__1346_ vdd gnd FILL
XFILL_2__1415_ vdd gnd FILL
XFILL_2__1277_ vdd gnd FILL
XFILL_0__948_ vdd gnd FILL
XFILL_0__879_ vdd gnd FILL
X_1541_ _1557_/Q _1557_/CLK _1573_/A vdd gnd DFFPOSX1
X_1472_ _1497_/B _1497_/A _1498_/B vdd gnd XOR2X1
XFILL_3__1455_ vdd gnd FILL
XFILL_3__1386_ vdd gnd FILL
XFILL_4__926_ vdd gnd FILL
XFILL_1__1022_ vdd gnd FILL
XFILL_4__857_ vdd gnd FILL
XFILL_4__788_ vdd gnd FILL
XFILL89250x11850 vdd gnd FILL
XFILL_2__1131_ vdd gnd FILL
XFILL_2__1200_ vdd gnd FILL
XFILL_0__802_ vdd gnd FILL
XFILL_2__1062_ vdd gnd FILL
XFILL_3__944_ vdd gnd FILL
XFILL_3__875_ vdd gnd FILL
XFILL_3__1240_ vdd gnd FILL
XFILL_0__1462_ vdd gnd FILL
XFILL_3__1171_ vdd gnd FILL
XFILL_0__1393_ vdd gnd FILL
XFILL_2__1329_ vdd gnd FILL
X_1524_ Xin[4] _1552_/CLK _1564_/A vdd gnd DFFPOSX1
XFILL_1__1571_ vdd gnd FILL
X_1455_ _1455_/A _1455_/B _1456_/C vdd gnd OR2X2
X_1386_ _1431_/C _1386_/B _1386_/C _1392_/B vdd gnd AOI21X1
XFILL_3__1507_ vdd gnd FILL
XFILL_2__962_ vdd gnd FILL
XFILL_3__1369_ vdd gnd FILL
XFILL_3__1438_ vdd gnd FILL
XFILL_1__1005_ vdd gnd FILL
XFILL_2__893_ vdd gnd FILL
XFILL89250x23550 vdd gnd FILL
XFILL_2__1114_ vdd gnd FILL
XFILL_2__1045_ vdd gnd FILL
XFILL_3__927_ vdd gnd FILL
XFILL_1__980_ vdd gnd FILL
XFILL_3__858_ vdd gnd FILL
X_1171_ _1171_/A Xin[7] Yin[7] _1172_/B vdd gnd AOI21X1
X_1240_ _1244_/A _1244_/B _1243_/B _1241_/C vdd gnd OAI21X1
XFILL_3__789_ vdd gnd FILL
XFILL_3__1154_ vdd gnd FILL
XFILL_3__1223_ vdd gnd FILL
XFILL_0__1445_ vdd gnd FILL
XFILL_0__1514_ vdd gnd FILL
XFILL_3__1085_ vdd gnd FILL
XFILL_0__1376_ vdd gnd FILL
X_1507_ Yin[14] _1507_/B _1507_/C _1508_/A vdd gnd OAI21X1
XFILL89250x35250 vdd gnd FILL
X_1369_ _1369_/A _1369_/B _1405_/A vdd gnd NAND2X1
XFILL_4__1401_ vdd gnd FILL
XFILL_4__1332_ vdd gnd FILL
X_1438_ _1440_/C _1440_/B _1440_/A _1477_/C vdd gnd NAND3X1
XFILL_2__945_ vdd gnd FILL
XFILL_1__1485_ vdd gnd FILL
XFILL_2__876_ vdd gnd FILL
X_882_ _882_/A _941_/D _882_/C _883_/A vdd gnd NAND3X1
X_951_ _951_/A _951_/B _951_/C _997_/B vdd gnd AOI21X1
XFILL_0__1092_ vdd gnd FILL
XFILL_2__1028_ vdd gnd FILL
XFILL_0__1230_ vdd gnd FILL
XFILL_0__1161_ vdd gnd FILL
XFILL_0_BUFX2_insert17 vdd gnd FILL
XFILL_1__963_ vdd gnd FILL
XFILL_1__894_ vdd gnd FILL
X_1154_ _1154_/A _1154_/B _1154_/C _1155_/C vdd gnd OAI21X1
X_1223_ _1223_/A _1223_/B _1242_/A _1241_/A vdd gnd OAI21X1
X_1085_ _1088_/A _1088_/B _1089_/C _1187_/B vdd gnd OAI21X1
XFILL_3__1206_ vdd gnd FILL
XFILL_3__1137_ vdd gnd FILL
XFILL_0__1428_ vdd gnd FILL
XFILL_1__1270_ vdd gnd FILL
XFILL_3__1068_ vdd gnd FILL
XFILL_0__1359_ vdd gnd FILL
XFILL_2__928_ vdd gnd FILL
XFILL_0__981_ vdd gnd FILL
XFILL_1__1399_ vdd gnd FILL
XFILL_1__1468_ vdd gnd FILL
XFILL_2__859_ vdd gnd FILL
X_865_ _865_/A _865_/B _865_/C _925_/C vdd gnd AOI21X1
X_934_ _948_/A _937_/B _937_/A _935_/B vdd gnd NAND3X1
X_796_ _796_/A _796_/B _796_/Y vdd gnd NOR2X1
XFILL_2__1577_ vdd gnd FILL
XFILL_0__1144_ vdd gnd FILL
XFILL_0__1213_ vdd gnd FILL
XFILL_0__1075_ vdd gnd FILL
XFILL_1__877_ vdd gnd FILL
XFILL_1__946_ vdd gnd FILL
X_1206_ _1289_/B _1288_/A _1289_/A _1207_/A vdd gnd AOI21X1
X_1137_ _861_/A _1376_/B _1227_/A _1146_/B vdd gnd OAI21X1
X_1068_ _1095_/B _1095_/A _1187_/A vdd gnd AND2X2
XFILL_1__1322_ vdd gnd FILL
XFILL_1__1253_ vdd gnd FILL
XFILL_1__1184_ vdd gnd FILL
XFILL_2__1500_ vdd gnd FILL
XFILL_2__1431_ vdd gnd FILL
XFILL_0_BUFX2_insert9 vdd gnd FILL
XFILL_2__1362_ vdd gnd FILL
XFILL_2__1293_ vdd gnd FILL
XFILL_0__964_ vdd gnd FILL
XFILL_0__895_ vdd gnd FILL
XFILL_1__800_ vdd gnd FILL
X_917_ _917_/A _969_/C _917_/C _921_/A vdd gnd AOI21X1
X_848_ _848_/A _848_/B _848_/C _865_/C vdd gnd AOI21X1
X_779_ _805_/A _783_/A vdd gnd INVX1
XFILL_3__1471_ vdd gnd FILL
XFILL_0__1127_ vdd gnd FILL
XFILL_0__1058_ vdd gnd FILL
XFILL_3_BUFX2_insert10 vdd gnd FILL
XFILL_1__929_ vdd gnd FILL
XFILL_1__1305_ vdd gnd FILL
XFILL_4__1014_ vdd gnd FILL
XFILL_1__1098_ vdd gnd FILL
XFILL_1__1236_ vdd gnd FILL
XFILL_1__1167_ vdd gnd FILL
XFILL_3__891_ vdd gnd FILL
XFILL_3__960_ vdd gnd FILL
XFILL_2__1414_ vdd gnd FILL
XFILL_2__1276_ vdd gnd FILL
XFILL_2__1345_ vdd gnd FILL
XFILL_0__947_ vdd gnd FILL
XFILL_0__878_ vdd gnd FILL
X_1540_ _1556_/Q _1559_/CLK _1572_/A vdd gnd DFFPOSX1
X_1471_ _1471_/A _1471_/B _1497_/B vdd gnd AND2X2
XFILL_3__1454_ vdd gnd FILL
XFILL_3__1385_ vdd gnd FILL
XFILL_1__1021_ vdd gnd FILL
XFILL_2__1061_ vdd gnd FILL
XFILL_2__1130_ vdd gnd FILL
XFILL_0__801_ vdd gnd FILL
XFILL_1__1219_ vdd gnd FILL
XFILL_3__943_ vdd gnd FILL
XFILL_3__874_ vdd gnd FILL
XFILL_0__1461_ vdd gnd FILL
XFILL_3__1170_ vdd gnd FILL
XFILL88650x4050 vdd gnd FILL
XFILL_2__1328_ vdd gnd FILL
XFILL_0__1392_ vdd gnd FILL
XFILL_2__1259_ vdd gnd FILL
X_1523_ _895_/A _1546_/CLK _1563_/A vdd gnd DFFPOSX1
X_1454_ _1465_/C _1454_/B _1454_/C _1460_/C vdd gnd OAI21X1
X_1385_ _1392_/C _1391_/A vdd gnd INVX1
XFILL_3__1506_ vdd gnd FILL
XFILL_1__1570_ vdd gnd FILL
XFILL_2__961_ vdd gnd FILL
XFILL_3__1437_ vdd gnd FILL
XFILL_3__1368_ vdd gnd FILL
XFILL_3__1299_ vdd gnd FILL
XFILL_1__1004_ vdd gnd FILL
XFILL_2__892_ vdd gnd FILL
XFILL_2__1113_ vdd gnd FILL
XFILL_2__1044_ vdd gnd FILL
XFILL_3__926_ vdd gnd FILL
XFILL_3__788_ vdd gnd FILL
XFILL_3__857_ vdd gnd FILL
X_1170_ _1188_/B _1188_/A _1248_/A vdd gnd NAND2X1
XFILL_3__1153_ vdd gnd FILL
XFILL_3__1222_ vdd gnd FILL
XFILL_0__1375_ vdd gnd FILL
XFILL_0__1444_ vdd gnd FILL
XFILL_0__1513_ vdd gnd FILL
XFILL_3__1084_ vdd gnd FILL
X_1437_ _1466_/D _1466_/C _1440_/A vdd gnd OR2X2
X_1506_ _1506_/A _1506_/B _1506_/C _1509_/A vdd gnd NAND3X1
XFILL_1__1484_ vdd gnd FILL
X_1368_ _1415_/A _1416_/A vdd gnd INVX1
XFILL_4__1262_ vdd gnd FILL
X_1299_ _1299_/A _1299_/B _1299_/C _1300_/C vdd gnd NOR3X1
XFILL89550x19650 vdd gnd FILL
XFILL_2__944_ vdd gnd FILL
XFILL_2__875_ vdd gnd FILL
XFILL_4__1193_ vdd gnd FILL
X_950_ Xin[0] Cin[6] Xin[1] Cin[5] _951_/C vdd gnd AOI22X1
X_881_ _941_/C _881_/B _945_/A vdd gnd NAND2X1
XFILL_2__1027_ vdd gnd FILL
XFILL_0__1091_ vdd gnd FILL
XFILL_0__1160_ vdd gnd FILL
XFILL_1__962_ vdd gnd FILL
XFILL_3__909_ vdd gnd FILL
XFILL_1__893_ vdd gnd FILL
X_1153_ _1242_/A _1153_/B _1153_/C _1155_/B vdd gnd NAND3X1
X_1084_ _1084_/A _1265_/A _1084_/C _1088_/A vdd gnd AOI21X1
X_1222_ _1305_/A Cin[6] _1223_/B vdd gnd NAND2X1
XFILL_3__1067_ vdd gnd FILL
XFILL_3__1136_ vdd gnd FILL
XFILL_3__1205_ vdd gnd FILL
XFILL_0__1427_ vdd gnd FILL
XFILL_0__1358_ vdd gnd FILL
XFILL_0__1289_ vdd gnd FILL
XFILL_1__1467_ vdd gnd FILL
XFILL_2__927_ vdd gnd FILL
XFILL_0__980_ vdd gnd FILL
XFILL_2__858_ vdd gnd FILL
XFILL_1__1398_ vdd gnd FILL
X_933_ _947_/B _947_/A _933_/C _937_/B vdd gnd NAND3X1
XFILL_2__789_ vdd gnd FILL
X_864_ _890_/C _925_/B _925_/A _878_/B vdd gnd NAND3X1
X_795_ _795_/A _795_/B _795_/C _796_/A vdd gnd AOI21X1
XFILL_2__1576_ vdd gnd FILL
XFILL_0__1212_ vdd gnd FILL
XFILL_0__1143_ vdd gnd FILL
XFILL_0__1074_ vdd gnd FILL
XFILL_1__945_ vdd gnd FILL
XFILL_1__876_ vdd gnd FILL
X_1067_ _1143_/A _1067_/B _1067_/C _1095_/B vdd gnd NAND3X1
X_1136_ _1305_/A Cin[5] _1227_/A vdd gnd NAND2X1
X_1205_ _1205_/A _1205_/B _1205_/C _1289_/B vdd gnd OAI21X1
XFILL_1__1321_ vdd gnd FILL
XFILL_3__1119_ vdd gnd FILL
XFILL_1__1252_ vdd gnd FILL
XFILL_1__1183_ vdd gnd FILL
XFILL_2__1430_ vdd gnd FILL
XFILL_1__1519_ vdd gnd FILL
XFILL_2__1361_ vdd gnd FILL
XFILL_2__1292_ vdd gnd FILL
XFILL88350x23550 vdd gnd FILL
XFILL_0__963_ vdd gnd FILL
XFILL_0__894_ vdd gnd FILL
X_916_ _916_/A _916_/B _969_/A _921_/B vdd gnd AOI21X1
XFILL_3__1470_ vdd gnd FILL
X_847_ _847_/A _848_/C vdd gnd INVX1
X_778_ Xin[1] Cin[1] _805_/A vdd gnd NAND2X1
XFILL_3_BUFX2_insert11 vdd gnd FILL
XFILL_0__1057_ vdd gnd FILL
XFILL_0__1126_ vdd gnd FILL
XFILL_1__928_ vdd gnd FILL
XFILL_1__859_ vdd gnd FILL
X_1119_ _1119_/A _1122_/C _1551_/D vdd gnd XNOR2X1
XFILL_1__1235_ vdd gnd FILL
XFILL_1__1304_ vdd gnd FILL
XFILL_1__1097_ vdd gnd FILL
XFILL_1__1166_ vdd gnd FILL
XFILL_3__890_ vdd gnd FILL
XFILL88350x35250 vdd gnd FILL
XFILL_2__1344_ vdd gnd FILL
XFILL_2__1413_ vdd gnd FILL
XFILL_0__946_ vdd gnd FILL
XFILL_2__1275_ vdd gnd FILL
XFILL_0__877_ vdd gnd FILL
X_1470_ _1470_/A _1470_/B _1470_/C _1471_/B vdd gnd OAI21X1
XFILL_3__1453_ vdd gnd FILL
XFILL_3__1384_ vdd gnd FILL
XFILL_1__1020_ vdd gnd FILL
XFILL_0__1109_ vdd gnd FILL
XFILL_4__1493_ vdd gnd FILL
XFILL_0__800_ vdd gnd FILL
XFILL_1__1218_ vdd gnd FILL
XFILL_2__1060_ vdd gnd FILL
XFILL_1__1149_ vdd gnd FILL
XFILL_3__942_ vdd gnd FILL
XFILL_3__873_ vdd gnd FILL
XFILL_0__1460_ vdd gnd FILL
XFILL_0__1391_ vdd gnd FILL
XFILL_2__1327_ vdd gnd FILL
XFILL_0__929_ vdd gnd FILL
XFILL_2__1258_ vdd gnd FILL
XFILL_2__1189_ vdd gnd FILL
X_1522_ Xin[2] _1546_/CLK _1562_/A vdd gnd DFFPOSX1
X_1453_ _1455_/B _1455_/A _1465_/C vdd gnd NOR2X1
XFILL_3__1436_ vdd gnd FILL
XFILL_3__1505_ vdd gnd FILL
X_1384_ _1392_/C _1391_/B _1391_/C _1428_/A vdd gnd NAND3X1
XFILL_4__907_ vdd gnd FILL
XFILL_2__891_ vdd gnd FILL
XFILL_2__960_ vdd gnd FILL
XFILL_3__1367_ vdd gnd FILL
XFILL_3__1298_ vdd gnd FILL
XFILL_4__838_ vdd gnd FILL
XFILL_1__1003_ vdd gnd FILL
XFILL_4__769_ vdd gnd FILL
XFILL89250x4050 vdd gnd FILL
XFILL_2__1112_ vdd gnd FILL
XFILL_2__1043_ vdd gnd FILL
XFILL_3__925_ vdd gnd FILL
XFILL_3__787_ vdd gnd FILL
XFILL_3__856_ vdd gnd FILL
XFILL_0__1512_ vdd gnd FILL
XFILL_3__1152_ vdd gnd FILL
XFILL_3__1083_ vdd gnd FILL
XFILL_3__1221_ vdd gnd FILL
XFILL_0__1374_ vdd gnd FILL
XFILL_0__1443_ vdd gnd FILL
X_1436_ _1436_/A Cin[7] _1466_/C vdd gnd NAND2X1
X_1367_ _1367_/A _1367_/B _1415_/A vdd gnd NAND2X1
X_1505_ _1505_/A _1505_/B _1516_/A _1510_/B vdd gnd OAI21X1
XFILL_1__1483_ vdd gnd FILL
XFILL_3__1419_ vdd gnd FILL
X_1298_ _1422_/B _1422_/A _1511_/D _1364_/B vdd gnd AOI21X1
XFILL_2__943_ vdd gnd FILL
XFILL_2__874_ vdd gnd FILL
X_880_ _882_/C _882_/A _941_/C vdd gnd AND2X2
XFILL_2__1026_ vdd gnd FILL
XFILL_0__1090_ vdd gnd FILL
XFILL_3__908_ vdd gnd FILL
XFILL_1__961_ vdd gnd FILL
XFILL_1__892_ vdd gnd FILL
X_1221_ _1221_/A _1221_/B _1275_/A _1357_/C vdd gnd OAI21X1
XFILL_3__839_ vdd gnd FILL
X_1152_ _1152_/A _1152_/B _1155_/A vdd gnd AND2X2
X_1083_ _1083_/A _1083_/B _1172_/A _1088_/B vdd gnd AOI21X1
XFILL_3__1204_ vdd gnd FILL
XFILL_3__1066_ vdd gnd FILL
XFILL_3__1135_ vdd gnd FILL
XFILL_0__1288_ vdd gnd FILL
XFILL_0__1426_ vdd gnd FILL
XFILL_0__1357_ vdd gnd FILL
X_1419_ _1421_/A _1424_/A vdd gnd INVX1
XFILL_4__1313_ vdd gnd FILL
XFILL_1__1466_ vdd gnd FILL
XFILL_4__1244_ vdd gnd FILL
XFILL_1__1397_ vdd gnd FILL
XFILL_4__1175_ vdd gnd FILL
XFILL_2__926_ vdd gnd FILL
XFILL_2__788_ vdd gnd FILL
XFILL_2__857_ vdd gnd FILL
X_932_ _932_/A _932_/B _947_/C _937_/A vdd gnd OAI21X1
X_863_ _863_/A _863_/B _925_/B vdd gnd NAND2X1
X_794_ _832_/C _796_/B vdd gnd INVX1
XFILL_2__1575_ vdd gnd FILL
XFILL_0__1142_ vdd gnd FILL
XFILL_0__1211_ vdd gnd FILL
XFILL_2__1009_ vdd gnd FILL
XFILL_0__1073_ vdd gnd FILL
XFILL_1__944_ vdd gnd FILL
XFILL_1__875_ vdd gnd FILL
X_1204_ _1217_/B _1217_/C _1217_/A _1288_/A vdd gnd NAND3X1
X_1066_ _965_/B _964_/B _1239_/A _1067_/C vdd gnd OAI21X1
X_1135_ Cin[6] _1376_/B vdd gnd INVX1
XFILL_1__1320_ vdd gnd FILL
XFILL_1__1251_ vdd gnd FILL
XFILL_3__1118_ vdd gnd FILL
XFILL_3__1049_ vdd gnd FILL
XFILL_0__1409_ vdd gnd FILL
XFILL_1__1182_ vdd gnd FILL
XFILL_2__1360_ vdd gnd FILL
XFILL_1__1518_ vdd gnd FILL
XFILL_0__962_ vdd gnd FILL
XFILL_1__1449_ vdd gnd FILL
XFILL_2__1291_ vdd gnd FILL
XFILL_2__909_ vdd gnd FILL
XFILL_0__893_ vdd gnd FILL
X_915_ _954_/C _922_/C vdd gnd INVX1
X_846_ _866_/C _866_/B _866_/A _890_/C vdd gnd NAND3X1
XFILL_4__940_ vdd gnd FILL
XFILL_4__871_ vdd gnd FILL
X_777_ _777_/A _777_/B _777_/C _787_/C vdd gnd OAI21X1
XFILL_2__1489_ vdd gnd FILL
XFILL_0__1125_ vdd gnd FILL
XFILL_3_BUFX2_insert12 vdd gnd FILL
XFILL_0__1056_ vdd gnd FILL
XFILL_1__927_ vdd gnd FILL
XFILL_1__858_ vdd gnd FILL
X_1118_ _1121_/A _1120_/A _1122_/C vdd gnd NAND2X1
XFILL_1__789_ vdd gnd FILL
X_1049_ _1052_/A _1052_/B _1051_/C _1050_/C vdd gnd OAI21X1
XFILL_1__1303_ vdd gnd FILL
XFILL_1__1234_ vdd gnd FILL
XFILL_1__1096_ vdd gnd FILL
XFILL_1__1165_ vdd gnd FILL
XFILL_4_CLKBUF1_insert4 vdd gnd FILL
XFILL_2__1343_ vdd gnd FILL
XFILL_2__1412_ vdd gnd FILL
XFILL_2__1274_ vdd gnd FILL
XFILL88650x19650 vdd gnd FILL
XFILL_0__945_ vdd gnd FILL
XFILL_0__876_ vdd gnd FILL
XFILL88050x7950 vdd gnd FILL
X_829_ _829_/A _877_/B _829_/C _832_/A vdd gnd AOI21X1
XFILL_3__1452_ vdd gnd FILL
XFILL_3__1383_ vdd gnd FILL
XFILL_0__1108_ vdd gnd FILL
XFILL_0__1039_ vdd gnd FILL
XFILL_1__1148_ vdd gnd FILL
XFILL_1__1217_ vdd gnd FILL
XFILL_3__941_ vdd gnd FILL
XFILL_1__1079_ vdd gnd FILL
XFILL_3__872_ vdd gnd FILL
XFILL_0__1390_ vdd gnd FILL
XFILL_2__1326_ vdd gnd FILL
XFILL_2__1257_ vdd gnd FILL
XFILL_0__928_ vdd gnd FILL
XFILL_0__859_ vdd gnd FILL
XFILL_2__1188_ vdd gnd FILL
X_1521_ Xin[1] _1552_/CLK _1561_/A vdd gnd DFFPOSX1
X_1452_ _1465_/B _1454_/B vdd gnd INVX1
X_1383_ _1386_/C _1386_/B _1431_/C _1391_/C vdd gnd NAND3X1
XFILL_3__1366_ vdd gnd FILL
XFILL_3__1504_ vdd gnd FILL
XFILL_3__1435_ vdd gnd FILL
XFILL_2__890_ vdd gnd FILL
XFILL_1__1002_ vdd gnd FILL
XFILL_3__1297_ vdd gnd FILL
XFILL_2__1111_ vdd gnd FILL
XFILL_2__1042_ vdd gnd FILL
XFILL_3__924_ vdd gnd FILL
XFILL_3__786_ vdd gnd FILL
XFILL_3__855_ vdd gnd FILL
XFILL_3__1220_ vdd gnd FILL
XFILL_0__1511_ vdd gnd FILL
XFILL_3__1082_ vdd gnd FILL
XFILL_3__1151_ vdd gnd FILL
XFILL_0__1373_ vdd gnd FILL
XFILL_0__1442_ vdd gnd FILL
XFILL_2__1309_ vdd gnd FILL
X_1504_ _1504_/A _1504_/B _1504_/C _1516_/A vdd gnd OAI21X1
X_1366_ _1366_/A _1366_/B _1366_/C _1412_/C vdd gnd AOI21X1
X_1435_ _1435_/A _1470_/B _1466_/D _1440_/B vdd gnd OAI21X1
XFILL_2__942_ vdd gnd FILL
XFILL_3__1349_ vdd gnd FILL
XFILL_1__1482_ vdd gnd FILL
XFILL_3__1418_ vdd gnd FILL
X_1297_ _1297_/A _1297_/B _1422_/A vdd gnd NOR2X1
XFILL_2__873_ vdd gnd FILL
XFILL_2__1025_ vdd gnd FILL
XFILL_3__907_ vdd gnd FILL
XFILL_3__838_ vdd gnd FILL
XFILL_1__891_ vdd gnd FILL
XFILL_1__960_ vdd gnd FILL
X_1151_ _1151_/A _1219_/A _1151_/C _1219_/B vdd gnd NAND3X1
X_1220_ _1220_/A _1220_/B _1220_/C _1221_/B vdd gnd AOI21X1
X_1082_ _1157_/C _1089_/C vdd gnd INVX1
XFILL_3__1203_ vdd gnd FILL
XFILL_3__769_ vdd gnd FILL
XFILL_0__1425_ vdd gnd FILL
XFILL_3__1065_ vdd gnd FILL
XFILL_3__1134_ vdd gnd FILL
XFILL_0__1356_ vdd gnd FILL
XFILL_0__1287_ vdd gnd FILL
X_1349_ _1367_/B _1349_/B _1406_/B _1413_/B vdd gnd NAND3X1
X_1418_ _1425_/A _1511_/A _1421_/A vdd gnd NAND2X1
XFILL_2__925_ vdd gnd FILL
XFILL_1__1396_ vdd gnd FILL
XFILL_1__1465_ vdd gnd FILL
XFILL_2__787_ vdd gnd FILL
XFILL_2__856_ vdd gnd FILL
X_931_ _946_/B _931_/B _948_/A vdd gnd XOR2X1
X_862_ _867_/B _868_/B _868_/C _863_/B vdd gnd NAND3X1
X_793_ _795_/C _795_/B _795_/A _832_/C vdd gnd NAND3X1
XFILL_2__1574_ vdd gnd FILL
XFILL_2__1008_ vdd gnd FILL
XFILL_0__1141_ vdd gnd FILL
XFILL_0__1072_ vdd gnd FILL
XFILL_0__1210_ vdd gnd FILL
XFILL_1__943_ vdd gnd FILL
XFILL_1__874_ vdd gnd FILL
X_1203_ _1211_/C _1211_/B _1218_/A _1207_/B vdd gnd AOI21X1
X_1134_ _1139_/C _1232_/A _1242_/B vdd gnd NAND2X1
XFILL_1__1181_ vdd gnd FILL
XFILL_3__1117_ vdd gnd FILL
X_1065_ _1065_/A _1065_/B _1067_/B vdd gnd NAND2X1
XFILL_0__1408_ vdd gnd FILL
XFILL_1__1250_ vdd gnd FILL
XFILL_3__1048_ vdd gnd FILL
XFILL_0__1339_ vdd gnd FILL
XFILL_4__1226_ vdd gnd FILL
XFILL_1__1517_ vdd gnd FILL
XFILL_2__1290_ vdd gnd FILL
XFILL_2__908_ vdd gnd FILL
XFILL_0__961_ vdd gnd FILL
XFILL_0__892_ vdd gnd FILL
XFILL_4__1157_ vdd gnd FILL
XFILL_1__1448_ vdd gnd FILL
XFILL_1__1379_ vdd gnd FILL
XFILL_2__839_ vdd gnd FILL
X_914_ _954_/C _954_/B _954_/A _990_/A vdd gnd NAND3X1
X_845_ _903_/B _849_/B _903_/A _866_/A vdd gnd OAI21X1
X_776_ _886_/A _964_/A _803_/B vdd gnd NOR2X1
XFILL_2__1488_ vdd gnd FILL
XFILL_3_BUFX2_insert13 vdd gnd FILL
XFILL_0__1055_ vdd gnd FILL
XFILL_0__1124_ vdd gnd FILL
XFILL_1__926_ vdd gnd FILL
X_1117_ _1117_/A _1117_/B _1117_/C _1120_/A vdd gnd OAI21X1
XFILL_1__788_ vdd gnd FILL
XFILL_1__857_ vdd gnd FILL
XFILL_4__999_ vdd gnd FILL
X_1048_ _963_/B _963_/A _1048_/C _1051_/C vdd gnd AOI21X1
XFILL89250x31350 vdd gnd FILL
XFILL_1__1233_ vdd gnd FILL
XFILL_1__1302_ vdd gnd FILL
XFILL_1__1164_ vdd gnd FILL
XFILL_1__1095_ vdd gnd FILL
XFILL_2__1411_ vdd gnd FILL
XFILL_2__1273_ vdd gnd FILL
XFILL_2__1342_ vdd gnd FILL
XFILL_0__944_ vdd gnd FILL
XFILL_0__875_ vdd gnd FILL
X_828_ _828_/A _828_/B _941_/D vdd gnd NOR2X1
X_759_ Yin[0] _761_/B _760_/A vdd gnd NAND2X1
XFILL_3__1451_ vdd gnd FILL
XFILL_3__1382_ vdd gnd FILL
XFILL_0__1107_ vdd gnd FILL
XFILL_0__1038_ vdd gnd FILL
XFILL_1__909_ vdd gnd FILL
XFILL_4__1560_ vdd gnd FILL
XFILL_1__1216_ vdd gnd FILL
XFILL_1__1147_ vdd gnd FILL
XFILL_3__940_ vdd gnd FILL
XFILL_3__871_ vdd gnd FILL
XFILL_1__1078_ vdd gnd FILL
XFILL_2__1187_ vdd gnd FILL
XFILL_2__1325_ vdd gnd FILL
XFILL_2__1256_ vdd gnd FILL
XFILL_0__927_ vdd gnd FILL
XFILL_0__858_ vdd gnd FILL
XFILL_0__789_ vdd gnd FILL
X_1520_ Xin[0] _1552_/CLK _1560_/A vdd gnd DFFPOSX1
X_1451_ _1455_/B _1455_/A _1465_/B vdd gnd NAND2X1
XFILL_3__1503_ vdd gnd FILL
X_1382_ _1382_/A _1431_/C vdd gnd INVX1
XFILL_3__1434_ vdd gnd FILL
XFILL_3__1365_ vdd gnd FILL
XFILL_3__1296_ vdd gnd FILL
XFILL_1__1001_ vdd gnd FILL
XFILL_4__1474_ vdd gnd FILL
XFILL_2__1110_ vdd gnd FILL
XFILL_2__1041_ vdd gnd FILL
XFILL_3__923_ vdd gnd FILL
XFILL_3__854_ vdd gnd FILL
XFILL_3__785_ vdd gnd FILL
XFILL_3__1150_ vdd gnd FILL
XFILL_0__1441_ vdd gnd FILL
XFILL_0__1510_ vdd gnd FILL
XFILL_3__1081_ vdd gnd FILL
XFILL_2__1308_ vdd gnd FILL
XFILL_0__1372_ vdd gnd FILL
XFILL_2__1239_ vdd gnd FILL
X_1503_ _1505_/B _1505_/A _1558_/D vdd gnd XOR2X1
X_1434_ _1466_/A _1470_/C _1434_/C _1466_/D vdd gnd OAI21X1
X_1365_ _1414_/C _1366_/C vdd gnd INVX1
X_1296_ _1296_/A _1296_/B _1296_/C _1511_/D vdd gnd OAI21X1
XFILL_2__941_ vdd gnd FILL
XFILL_1__1481_ vdd gnd FILL
XFILL_3__1417_ vdd gnd FILL
XFILL_3__1348_ vdd gnd FILL
XFILL_3__1279_ vdd gnd FILL
XFILL_2__872_ vdd gnd FILL
XFILL_2__1024_ vdd gnd FILL
XFILL_3__906_ vdd gnd FILL
XFILL_3__837_ vdd gnd FILL
XFILL_1__890_ vdd gnd FILL
X_1150_ _1154_/A _1154_/B _1153_/B _1151_/C vdd gnd OAI21X1
XFILL_3__768_ vdd gnd FILL
X_1081_ _1157_/C _1265_/B _1157_/A _1186_/A vdd gnd NAND3X1
XFILL_3__1202_ vdd gnd FILL
XFILL_3__1133_ vdd gnd FILL
XFILL_0__1424_ vdd gnd FILL
XFILL_0__1355_ vdd gnd FILL
XFILL_3__1064_ vdd gnd FILL
XFILL_0__1286_ vdd gnd FILL
X_1417_ _1417_/A _1459_/C _1417_/C _1425_/A vdd gnd NAND3X1
XFILL_1__1464_ vdd gnd FILL
X_1348_ _1348_/A _1348_/B _1348_/C _1354_/C vdd gnd AOI21X1
X_1279_ _1279_/A _1279_/B _1303_/B _1299_/A vdd gnd AOI21X1
XFILL_2__924_ vdd gnd FILL
XFILL_2__855_ vdd gnd FILL
XFILL_1__1395_ vdd gnd FILL
X_930_ _951_/A _931_/B vdd gnd INVX1
XFILL_2__786_ vdd gnd FILL
X_792_ _797_/B _792_/B _823_/B _795_/B vdd gnd OAI21X1
X_861_ _861_/A _964_/A _861_/C _868_/C vdd gnd OAI21X1
XFILL_2__1573_ vdd gnd FILL
XFILL_2__1007_ vdd gnd FILL
XFILL_0__1140_ vdd gnd FILL
XFILL_0__1071_ vdd gnd FILL
XFILL_1__942_ vdd gnd FILL
XFILL_1__873_ vdd gnd FILL
X_1064_ _1149_/C _1149_/D _1143_/C _1095_/A vdd gnd NAND3X1
X_1202_ _1217_/A _1217_/B _1205_/C _1211_/C vdd gnd NAND3X1
X_1133_ _1305_/A Cin[5] _1232_/A vdd gnd AND2X2
XFILL_3__1116_ vdd gnd FILL
XFILL_3__1047_ vdd gnd FILL
XFILL_0__1338_ vdd gnd FILL
XFILL_0__1407_ vdd gnd FILL
XFILL_1__1180_ vdd gnd FILL
XFILL_0__1269_ vdd gnd FILL
XFILL_1__1447_ vdd gnd FILL
XFILL_1__1516_ vdd gnd FILL
XFILL_2__907_ vdd gnd FILL
XFILL_2__838_ vdd gnd FILL
XFILL_0__891_ vdd gnd FILL
XFILL_4__1087_ vdd gnd FILL
XFILL_0__960_ vdd gnd FILL
XFILL_1__1378_ vdd gnd FILL
X_913_ _969_/A _916_/B _916_/A _954_/A vdd gnd NAND3X1
XFILL_2__769_ vdd gnd FILL
X_844_ _903_/C _849_/B vdd gnd INVX1
X_775_ Cin[2] _964_/A vdd gnd INVX2
XFILL_2__1487_ vdd gnd FILL
XFILL_0__1123_ vdd gnd FILL
XFILL_0__1054_ vdd gnd FILL
XFILL_3_BUFX2_insert14 vdd gnd FILL
XFILL_1__925_ vdd gnd FILL
XFILL_1__787_ vdd gnd FILL
X_1116_ _1124_/B _1209_/C _1124_/A _1117_/A vdd gnd AOI21X1
X_1047_ _962_/C _1047_/B _1048_/C vdd gnd NOR2X1
XFILL_1__856_ vdd gnd FILL
XFILL_1__1301_ vdd gnd FILL
XFILL_1__1094_ vdd gnd FILL
XFILL_1__1232_ vdd gnd FILL
XFILL89550x15750 vdd gnd FILL
XFILL_1__1163_ vdd gnd FILL
XFILL_2__1410_ vdd gnd FILL
XFILL_2__1272_ vdd gnd FILL
XFILL_2__1341_ vdd gnd FILL
XFILL_0__943_ vdd gnd FILL
XFILL_0__874_ vdd gnd FILL
XFILL_3__1450_ vdd gnd FILL
XFILL_4__921_ vdd gnd FILL
X_827_ _877_/B _829_/A _828_/B vdd gnd NAND2X1
X_758_ _758_/A _886_/A _761_/B vdd gnd NOR2X1
XFILL_3__1381_ vdd gnd FILL
XFILL_4__783_ vdd gnd FILL
XFILL_4__852_ vdd gnd FILL
XFILL_0__1106_ vdd gnd FILL
XFILL_0__1037_ vdd gnd FILL
XFILL_1__908_ vdd gnd FILL
XFILL_3__1579_ vdd gnd FILL
XFILL_1__839_ vdd gnd FILL
XFILL_1__1215_ vdd gnd FILL
XFILL89550x27450 vdd gnd FILL
XFILL_1__1077_ vdd gnd FILL
XFILL_1__1146_ vdd gnd FILL
XFILL_3__870_ vdd gnd FILL
XFILL_2__1324_ vdd gnd FILL
XFILL_0__926_ vdd gnd FILL
XFILL_2__1186_ vdd gnd FILL
XFILL_2__1255_ vdd gnd FILL
XFILL_0__788_ vdd gnd FILL
XFILL_0__857_ vdd gnd FILL
X_1450_ _1450_/A _1478_/C _1455_/A vdd gnd NAND2X1
XFILL_3__999_ vdd gnd FILL
XFILL_3__1433_ vdd gnd FILL
XFILL_3__1502_ vdd gnd FILL
X_1381_ _1381_/A _1492_/B _1382_/A vdd gnd NOR2X1
XFILL_3__1364_ vdd gnd FILL
XFILL_3__1295_ vdd gnd FILL
XFILL_1__1000_ vdd gnd FILL
X_1579_ _1579_/A Yout[5] vdd gnd BUFX2
XFILL89550x39150 vdd gnd FILL
XFILL_2__1040_ vdd gnd FILL
XFILL_1__1129_ vdd gnd FILL
XFILL_3__922_ vdd gnd FILL
XFILL_3__784_ vdd gnd FILL
XFILL88050x54750 vdd gnd FILL
XFILL_3__853_ vdd gnd FILL
XFILL_3__1080_ vdd gnd FILL
XFILL_0__1440_ vdd gnd FILL
XFILL_0__1371_ vdd gnd FILL
XFILL_2__1307_ vdd gnd FILL
XFILL_0__909_ vdd gnd FILL
XFILL_2__1238_ vdd gnd FILL
XFILL_2__1169_ vdd gnd FILL
X_1433_ _886_/B _1468_/A _1492_/B _1434_/C vdd gnd OAI21X1
X_1502_ _1514_/C _1505_/A vdd gnd INVX1
XFILL_3__1416_ vdd gnd FILL
XFILL_1__1480_ vdd gnd FILL
X_1364_ _1423_/A _1364_/B _1425_/B _1420_/A vdd gnd OAI21X1
X_1295_ _1295_/A _1296_/B vdd gnd INVX1
XFILL_2__940_ vdd gnd FILL
XFILL_2__871_ vdd gnd FILL
XFILL_0__1569_ vdd gnd FILL
XFILL_3__1347_ vdd gnd FILL
XFILL_3__1278_ vdd gnd FILL
XFILL_4__1456_ vdd gnd FILL
XFILL_4__1387_ vdd gnd FILL
XFILL_2__1023_ vdd gnd FILL
XFILL_3__905_ vdd gnd FILL
XFILL_3__836_ vdd gnd FILL
XFILL_3__767_ vdd gnd FILL
X_1080_ _1172_/A _1083_/B _1083_/A _1157_/A vdd gnd NAND3X1
XFILL88650x7950 vdd gnd FILL
XFILL_3__1063_ vdd gnd FILL
XFILL_3__1201_ vdd gnd FILL
XFILL_3__1132_ vdd gnd FILL
XFILL_0__1354_ vdd gnd FILL
XFILL_0__1423_ vdd gnd FILL
XFILL_0__1285_ vdd gnd FILL
X_1347_ _1354_/A _1354_/B _1413_/C _1360_/C vdd gnd OAI21X1
X_1416_ _1416_/A _1416_/B _1416_/C _1417_/C vdd gnd NAND3X1
XFILL_1__1394_ vdd gnd FILL
XFILL_1__1463_ vdd gnd FILL
X_1278_ _1344_/B _1278_/B _1278_/C _1279_/B vdd gnd NAND3X1
XFILL_2__923_ vdd gnd FILL
XFILL_2__854_ vdd gnd FILL
XFILL_2__785_ vdd gnd FILL
X_791_ _797_/C _792_/B vdd gnd INVX1
X_860_ _860_/A _965_/B _894_/A _868_/B vdd gnd OAI21X1
XFILL_2__1572_ vdd gnd FILL
XFILL88050x78150 vdd gnd FILL
XFILL_0__1070_ vdd gnd FILL
XFILL_2__1006_ vdd gnd FILL
XFILL_1__941_ vdd gnd FILL
XFILL_1__872_ vdd gnd FILL
X_1201_ _1221_/A _1201_/B _1201_/C _1217_/B vdd gnd NAND3X1
XFILL_3__819_ vdd gnd FILL
X_989_ _999_/B _999_/A _998_/A _996_/B vdd gnd OAI21X1
X_1063_ _965_/B _964_/B _1065_/A _1149_/C vdd gnd OAI21X1
X_1132_ Xin[2] Cin[6] _1139_/C vdd gnd AND2X2
XFILL_3__1115_ vdd gnd FILL
XFILL_3__1046_ vdd gnd FILL
XFILL_0__1406_ vdd gnd FILL
XFILL_0__1268_ vdd gnd FILL
XFILL_0__1337_ vdd gnd FILL
XFILL_0__1199_ vdd gnd FILL
XFILL_1__1446_ vdd gnd FILL
XFILL_1__1515_ vdd gnd FILL
XFILL_1__1377_ vdd gnd FILL
XFILL_2__906_ vdd gnd FILL
XFILL_2__837_ vdd gnd FILL
XFILL_0__890_ vdd gnd FILL
XFILL_2__768_ vdd gnd FILL
X_912_ _912_/A _912_/B _912_/C _916_/A vdd gnd NAND3X1
X_843_ _903_/C _849_/C _850_/C _866_/B vdd gnd NAND3X1
X_774_ _774_/A _795_/C _774_/Y vdd gnd NOR2X1
XFILL_2__1486_ vdd gnd FILL
XFILL_0__1122_ vdd gnd FILL
XFILL_3_BUFX2_insert15 vdd gnd FILL
XFILL_0__1053_ vdd gnd FILL
XFILL_1__924_ vdd gnd FILL
XFILL_1__855_ vdd gnd FILL
XFILL_1__786_ vdd gnd FILL
X_1115_ _1115_/A _1115_/B _1209_/A _1117_/B vdd gnd AOI21X1
X_1046_ Xin[0] Cin[7] _1152_/B _1046_/D _1052_/A vdd gnd AOI22X1
XFILL_1__1231_ vdd gnd FILL
XFILL_1__1300_ vdd gnd FILL
XFILL_1__1093_ vdd gnd FILL
XFILL_3__1029_ vdd gnd FILL
XFILL_1__1162_ vdd gnd FILL
XFILL_2__1340_ vdd gnd FILL
XFILL_4__1069_ vdd gnd FILL
XFILL_0__942_ vdd gnd FILL
XFILL_4__1207_ vdd gnd FILL
XFILL_4__1138_ vdd gnd FILL
XFILL_2__1271_ vdd gnd FILL
XFILL_1__1429_ vdd gnd FILL
XFILL_0__873_ vdd gnd FILL
X_826_ _835_/A _872_/C _835_/B _829_/A vdd gnd OAI21X1
X_757_ Xin[0] _886_/A vdd gnd INVX1
XFILL_3__1380_ vdd gnd FILL
XFILL_2__1469_ vdd gnd FILL
XFILL_0__1105_ vdd gnd FILL
XFILL_0__1036_ vdd gnd FILL
XFILL_1__907_ vdd gnd FILL
XFILL_1__838_ vdd gnd FILL
XFILL_3__1578_ vdd gnd FILL
X_1029_ _1053_/A _1050_/A vdd gnd INVX1
XFILL_1__769_ vdd gnd FILL
XFILL_1__1214_ vdd gnd FILL
XFILL_1__1145_ vdd gnd FILL
XFILL_1__1076_ vdd gnd FILL
XFILL_2__1323_ vdd gnd FILL
XFILL_0__925_ vdd gnd FILL
XFILL_2__1185_ vdd gnd FILL
XFILL_2__1254_ vdd gnd FILL
XFILL_0__787_ vdd gnd FILL
XFILL_0__856_ vdd gnd FILL
X_1380_ _1431_/A _1386_/C vdd gnd INVX1
X_809_ Yin[3] _814_/C vdd gnd INVX1
XFILL_3__998_ vdd gnd FILL
XFILL_3__1432_ vdd gnd FILL
XFILL_3__1501_ vdd gnd FILL
XFILL_3__1363_ vdd gnd FILL
XFILL_4__903_ vdd gnd FILL
XFILL_4__834_ vdd gnd FILL
XFILL_3__1294_ vdd gnd FILL
XFILL_4__765_ vdd gnd FILL
X_1578_ _1578_/A Yout[4] vdd gnd BUFX2
XFILL_0__1019_ vdd gnd FILL
XFILL_1__1128_ vdd gnd FILL
XFILL_3__921_ vdd gnd FILL
XFILL_1__1059_ vdd gnd FILL
XFILL_3__783_ vdd gnd FILL
XFILL_3__852_ vdd gnd FILL
XFILL88950x85950 vdd gnd FILL
XFILL_2__1306_ vdd gnd FILL
XFILL_2__1237_ vdd gnd FILL
XFILL_0__1370_ vdd gnd FILL
XFILL_0__908_ vdd gnd FILL
XFILL_0__839_ vdd gnd FILL
XFILL_2__1099_ vdd gnd FILL
XFILL_2__1168_ vdd gnd FILL
X_1432_ Cin[6] Xin[7] _1470_/C vdd gnd NAND2X1
X_1501_ _1501_/A _1504_/C _1514_/C vdd gnd XNOR2X1
X_1363_ _1364_/B _1423_/A _1554_/D vdd gnd XOR2X1
X_1294_ _1294_/A _1297_/B _1553_/D vdd gnd XNOR2X1
XFILL_3__1346_ vdd gnd FILL
XFILL_3__1415_ vdd gnd FILL
XFILL_2__870_ vdd gnd FILL
XFILL_0__1568_ vdd gnd FILL
XFILL_3__1277_ vdd gnd FILL
XFILL_0__1499_ vdd gnd FILL
XFILL_2__999_ vdd gnd FILL
XFILL_2__1022_ vdd gnd FILL
XFILL88650x15750 vdd gnd FILL
XFILL_3__904_ vdd gnd FILL
XFILL_3__835_ vdd gnd FILL
XFILL_3__766_ vdd gnd FILL
XFILL_3__1200_ vdd gnd FILL
XFILL_3__1062_ vdd gnd FILL
XFILL_3__1131_ vdd gnd FILL
XFILL_0__1353_ vdd gnd FILL
XFILL_0__1422_ vdd gnd FILL
XFILL_0__1284_ vdd gnd FILL
X_1346_ _1406_/B _1406_/A _1354_/B vdd gnd NOR2X1
X_1415_ _1415_/A _1458_/A _1415_/C _1459_/C vdd gnd NAND3X1
XFILL_2__922_ vdd gnd FILL
XFILL_1__1462_ vdd gnd FILL
X_1277_ _1277_/A _1277_/B _1279_/A vdd gnd NAND2X1
XFILL_1__1393_ vdd gnd FILL
XFILL_3__1329_ vdd gnd FILL
XFILL_2__784_ vdd gnd FILL
XFILL_2__853_ vdd gnd FILL
XFILL89250x7950 vdd gnd FILL
X_790_ _803_/B _823_/B vdd gnd INVX1
XFILL_2__1571_ vdd gnd FILL
XFILL_4__1507_ vdd gnd FILL
XFILL_2__1005_ vdd gnd FILL
XFILL_3__818_ vdd gnd FILL
XFILL_1__940_ vdd gnd FILL
X_988_ _992_/B _992_/A _993_/B _993_/A _999_/B vdd gnd AOI22X1
XFILL_1__871_ vdd gnd FILL
X_1200_ _1275_/A _1276_/B _1276_/A _1217_/A vdd gnd NAND3X1
X_1062_ Cin[2] _912_/B _1065_/A vdd gnd NAND2X1
X_1131_ _1145_/C _1146_/C vdd gnd INVX1
XFILL_0__1405_ vdd gnd FILL
XFILL_3__1114_ vdd gnd FILL
XFILL_3__1045_ vdd gnd FILL
XFILL_0__1267_ vdd gnd FILL
XFILL_0__1336_ vdd gnd FILL
XFILL_0__1198_ vdd gnd FILL
XFILL_1__1514_ vdd gnd FILL
X_1329_ Yin[9] _1329_/B _1344_/A vdd gnd NAND2X1
XFILL_2__905_ vdd gnd FILL
XFILL_1__1376_ vdd gnd FILL
XFILL_1__1445_ vdd gnd FILL
XFILL_2__836_ vdd gnd FILL
XFILL_2__767_ vdd gnd FILL
X_911_ Yin[5] _911_/B _916_/B vdd gnd NAND2X1
X_842_ _903_/A _849_/C vdd gnd INVX1
XFILL88650x39150 vdd gnd FILL
X_773_ _773_/A _773_/B _773_/C _774_/A vdd gnd AOI21X1
XFILL_2__1485_ vdd gnd FILL
XFILL_0__1121_ vdd gnd FILL
XFILL_0__1052_ vdd gnd FILL
XFILL_3_BUFX2_insert16 vdd gnd FILL
XFILL_1__923_ vdd gnd FILL
X_1114_ _1114_/A _1114_/B _1114_/C _1117_/C vdd gnd AOI21X1
XFILL_1__785_ vdd gnd FILL
XFILL_1__854_ vdd gnd FILL
X_1045_ _1045_/A _1045_/B _1045_/C _1052_/B vdd gnd AOI21X1
XFILL_1__1230_ vdd gnd FILL
XFILL_1__1161_ vdd gnd FILL
XFILL_1__1092_ vdd gnd FILL
XFILL_3__1028_ vdd gnd FILL
XFILL_0__1319_ vdd gnd FILL
XFILL_2__1270_ vdd gnd FILL
XFILL_0__941_ vdd gnd FILL
XFILL_0__872_ vdd gnd FILL
XFILL_1__1359_ vdd gnd FILL
XFILL_1__1428_ vdd gnd FILL
XFILL_2__819_ vdd gnd FILL
X_825_ _825_/A _825_/B _825_/C _835_/A vdd gnd AOI21X1
X_756_ _814_/A _758_/A vdd gnd INVX1
XFILL_2__1399_ vdd gnd FILL
XFILL_2__1468_ vdd gnd FILL
XFILL_0__1104_ vdd gnd FILL
XFILL_0__1035_ vdd gnd FILL
XFILL_3__1577_ vdd gnd FILL
XFILL_1__906_ vdd gnd FILL
XFILL_1__837_ vdd gnd FILL
XFILL_1__768_ vdd gnd FILL
X_1028_ _951_/B _951_/A _1053_/A vdd gnd NAND2X1
XFILL_1__1144_ vdd gnd FILL
XFILL_1__1213_ vdd gnd FILL
XFILL_1__1075_ vdd gnd FILL
XFILL_2__1322_ vdd gnd FILL
XFILL_2__1253_ vdd gnd FILL
XFILL_0__924_ vdd gnd FILL
XFILL_0__855_ vdd gnd FILL
XFILL_2__1184_ vdd gnd FILL
XFILL_2_BUFX2_insert6 vdd gnd FILL
XFILL_3__997_ vdd gnd FILL
XFILL_0__786_ vdd gnd FILL
XFILL_3__1500_ vdd gnd FILL
X_808_ _912_/A _836_/B Yin[3] _847_/A vdd gnd NAND3X1
XFILL_3__1362_ vdd gnd FILL
XFILL_3__1431_ vdd gnd FILL
XFILL_3__1293_ vdd gnd FILL
XFILL_0__1018_ vdd gnd FILL
X_1577_ _1577_/A Yout[3] vdd gnd BUFX2
XFILL_1__1127_ vdd gnd FILL
XFILL_3__851_ vdd gnd FILL
XFILL_3__920_ vdd gnd FILL
XFILL_1__1058_ vdd gnd FILL
XFILL_3__782_ vdd gnd FILL
XFILL_2__1236_ vdd gnd FILL
XFILL_2__1305_ vdd gnd FILL
XFILL_2__1167_ vdd gnd FILL
XFILL_0__907_ vdd gnd FILL
XFILL_0__838_ vdd gnd FILL
XFILL_2__1098_ vdd gnd FILL
XFILL_0__769_ vdd gnd FILL
X_1500_ _1506_/C _1500_/B _1504_/C vdd gnd XNOR2X1
X_1362_ _1425_/B _1362_/B _1423_/A vdd gnd NAND2X1
X_1431_ _1431_/A _1431_/B _1431_/C _1440_/C vdd gnd OAI21X1
X_1293_ _1296_/C _1295_/A _1297_/B vdd gnd NAND2X1
XFILL_0__1567_ vdd gnd FILL
XFILL_3__1276_ vdd gnd FILL
XFILL_3__1345_ vdd gnd FILL
XFILL_3__1414_ vdd gnd FILL
XFILL_0__1498_ vdd gnd FILL
XFILL_2__1021_ vdd gnd FILL
XFILL_2__998_ vdd gnd FILL
XFILL_3__903_ vdd gnd FILL
XFILL_3__834_ vdd gnd FILL
XFILL_3__765_ vdd gnd FILL
XFILL_3__1130_ vdd gnd FILL
XFILL_0__1421_ vdd gnd FILL
XFILL_3__1061_ vdd gnd FILL
XFILL_2__1219_ vdd gnd FILL
XFILL_0__1352_ vdd gnd FILL
XFILL_0__1283_ vdd gnd FILL
XFILL_0_CLKBUF1_insert0 vdd gnd FILL
X_1276_ _1276_/A _1276_/B _1276_/C _1299_/C vdd gnd AOI21X1
X_1345_ _1345_/A _1345_/B _1406_/B vdd gnd NAND2X1
X_1414_ _1414_/A _1414_/B _1414_/C _1417_/A vdd gnd OAI21X1
XFILL_2__921_ vdd gnd FILL
XFILL_3__1328_ vdd gnd FILL
XFILL_1__1461_ vdd gnd FILL
XFILL_1__1392_ vdd gnd FILL
XFILL_3__1259_ vdd gnd FILL
XFILL_4__1170_ vdd gnd FILL
XFILL_2__783_ vdd gnd FILL
XFILL_2__852_ vdd gnd FILL
XFILL_4__1437_ vdd gnd FILL
XFILL_4__1368_ vdd gnd FILL
XFILL_2__1570_ vdd gnd FILL
XFILL_2__1004_ vdd gnd FILL
XFILL_4__1299_ vdd gnd FILL
XFILL_3__817_ vdd gnd FILL
X_987_ _987_/A _987_/B _987_/C _993_/B vdd gnd OAI21X1
XFILL_1__870_ vdd gnd FILL
X_1130_ Xin[1] Cin[7] _1145_/C vdd gnd NAND2X1
XFILL_3__1113_ vdd gnd FILL
X_1061_ _1065_/B _1239_/A _1143_/C vdd gnd NAND2X1
XFILL_0__1404_ vdd gnd FILL
XFILL_0__1335_ vdd gnd FILL
XFILL_3__1044_ vdd gnd FILL
XFILL_0__1197_ vdd gnd FILL
XFILL_0__1266_ vdd gnd FILL
XFILL_1__999_ vdd gnd FILL
X_1328_ _1367_/B _1349_/B _1370_/A vdd gnd NAND2X1
XFILL_1__1444_ vdd gnd FILL
XFILL_1__1513_ vdd gnd FILL
X_1259_ _1259_/A Yin[9] _1262_/A vdd gnd XNOR2X1
XFILL_2__904_ vdd gnd FILL
XFILL_2__835_ vdd gnd FILL
XFILL_1__1375_ vdd gnd FILL
XFILL_2__766_ vdd gnd FILL
X_910_ _969_/C _917_/C _917_/A _954_/B vdd gnd NAND3X1
X_841_ Cin[1] _961_/A _903_/A vdd gnd NAND2X1
X_772_ _772_/A _795_/C vdd gnd INVX1
XFILL_2__1484_ vdd gnd FILL
XFILL_3_BUFX2_insert17 vdd gnd FILL
XFILL_0__1120_ vdd gnd FILL
XFILL_0__1051_ vdd gnd FILL
XFILL_1__922_ vdd gnd FILL
X_1113_ _1113_/A _1114_/C vdd gnd INVX1
XFILL_1__784_ vdd gnd FILL
XFILL_1__853_ vdd gnd FILL
X_1044_ _1152_/A _1051_/B _1052_/C _1125_/A vdd gnd NAND3X1
XFILL_4__995_ vdd gnd FILL
XFILL_1__1091_ vdd gnd FILL
XFILL_0__1318_ vdd gnd FILL
XFILL_1__1160_ vdd gnd FILL
XFILL_3__1027_ vdd gnd FILL
XFILL_0__1249_ vdd gnd FILL
XFILL_1__1427_ vdd gnd FILL
XFILL_2__818_ vdd gnd FILL
XFILL_0__940_ vdd gnd FILL
XFILL_0__871_ vdd gnd FILL
XFILL_1__1289_ vdd gnd FILL
XFILL_1__1358_ vdd gnd FILL
X_824_ _877_/A _872_/C vdd gnd INVX1
XFILL_2__1467_ vdd gnd FILL
XFILL_2__1398_ vdd gnd FILL
XFILL_0__1103_ vdd gnd FILL
XFILL_0__1034_ vdd gnd FILL
XFILL_1__905_ vdd gnd FILL
XFILL_1__836_ vdd gnd FILL
X_1027_ _996_/C _1027_/B _998_/Y _1208_/C vdd gnd OAI21X1
XFILL_1__767_ vdd gnd FILL
XFILL_3__1576_ vdd gnd FILL
XFILL_1__1143_ vdd gnd FILL
XFILL_1__1212_ vdd gnd FILL
XFILL_1__1074_ vdd gnd FILL
XFILL_2__1252_ vdd gnd FILL
XFILL_2__1321_ vdd gnd FILL
XFILL_2__1183_ vdd gnd FILL
XFILL_0__923_ vdd gnd FILL
XFILL_0__785_ vdd gnd FILL
XFILL_0__854_ vdd gnd FILL
XFILL_2_BUFX2_insert7 vdd gnd FILL
XFILL_3__996_ vdd gnd FILL
XFILL_0__1583_ vdd gnd FILL
XFILL_2__1519_ vdd gnd FILL
X_807_ _837_/A _848_/A vdd gnd INVX1
XFILL_3__1430_ vdd gnd FILL
XFILL_3__1361_ vdd gnd FILL
XFILL_3__1292_ vdd gnd FILL
XFILL_0__1017_ vdd gnd FILL
X_1576_ _1576_/A Yout[2] vdd gnd BUFX2
XFILL_4__1470_ vdd gnd FILL
XFILL_1__819_ vdd gnd FILL
XFILL_1__1057_ vdd gnd FILL
XFILL_1__1126_ vdd gnd FILL
XFILL_3__850_ vdd gnd FILL
XFILL_3__781_ vdd gnd FILL
XFILL_2__1304_ vdd gnd FILL
XFILL_0__906_ vdd gnd FILL
XFILL_2__1235_ vdd gnd FILL
XFILL_2__1166_ vdd gnd FILL
XFILL_0__837_ vdd gnd FILL
XFILL_2__1097_ vdd gnd FILL
XFILL_0__768_ vdd gnd FILL
X_1430_ _1430_/A _1430_/B _1455_/B vdd gnd AND2X2
XFILL_3__979_ vdd gnd FILL
XFILL_3__1413_ vdd gnd FILL
X_1361_ _1361_/A _1361_/B _1361_/C _1425_/B vdd gnd NAND3X1
X_1292_ _1292_/A _1292_/B _1292_/C _1295_/A vdd gnd OAI21X1
XFILL_0__1566_ vdd gnd FILL
XFILL_3__1275_ vdd gnd FILL
XFILL_3__1344_ vdd gnd FILL
XFILL_0__1497_ vdd gnd FILL
XFILL_4__815_ vdd gnd FILL
XFILL89550x11850 vdd gnd FILL
X_1559_ _1559_/D _1559_/CLK _1559_/Q vdd gnd DFFPOSX1
XFILL_2__1020_ vdd gnd FILL
XFILL_2__997_ vdd gnd FILL
XFILL_1__1109_ vdd gnd FILL
XFILL_3__833_ vdd gnd FILL
XFILL_3__902_ vdd gnd FILL
XFILL_3__764_ vdd gnd FILL
XFILL_3__1060_ vdd gnd FILL
XFILL_0__1351_ vdd gnd FILL
XFILL_0__1420_ vdd gnd FILL
XFILL_2__1149_ vdd gnd FILL
XFILL_2__1218_ vdd gnd FILL
XFILL_0__1282_ vdd gnd FILL
XFILL_0_CLKBUF1_insert1 vdd gnd FILL
X_1413_ _1413_/A _1413_/B _1413_/C _1414_/B vdd gnd AOI21X1
X_1275_ _1275_/A _1276_/C vdd gnd INVX1
X_1344_ _1344_/A _1344_/B _1369_/A _1345_/B vdd gnd NAND3X1
XFILL_1__1460_ vdd gnd FILL
XFILL_2__851_ vdd gnd FILL
XFILL_2__920_ vdd gnd FILL
XFILL_1__1391_ vdd gnd FILL
XFILL_3__1327_ vdd gnd FILL
XFILL_3__1258_ vdd gnd FILL
XFILL_3__1189_ vdd gnd FILL
XFILL_2__782_ vdd gnd FILL
XFILL89550x23550 vdd gnd FILL
XFILL89250x58650 vdd gnd FILL
XFILL_2__1003_ vdd gnd FILL
XFILL_3__816_ vdd gnd FILL
X_986_ _986_/A _986_/B _986_/C _993_/A vdd gnd NAND3X1
X_1060_ Cin[2] _1249_/A _1239_/A vdd gnd AND2X2
XFILL_3__1112_ vdd gnd FILL
XFILL_3__1043_ vdd gnd FILL
XFILL_0__1334_ vdd gnd FILL
XFILL_0__1403_ vdd gnd FILL
XFILL_0__1196_ vdd gnd FILL
XFILL_0__1265_ vdd gnd FILL
XFILL_1__998_ vdd gnd FILL
XFILL_4__1152_ vdd gnd FILL
XFILL_4__1221_ vdd gnd FILL
XFILL_1__1443_ vdd gnd FILL
XFILL_1__1512_ vdd gnd FILL
X_1327_ _1327_/A _1327_/B _1327_/C _1349_/B vdd gnd NAND3X1
X_1258_ _1316_/A _1258_/B _1258_/C _1261_/B vdd gnd NAND3X1
X_1189_ _1248_/C _1266_/B _1266_/A _1220_/A vdd gnd NAND3X1
XFILL_2__903_ vdd gnd FILL
XFILL_2__834_ vdd gnd FILL
XFILL_4__1083_ vdd gnd FILL
XFILL89550x35250 vdd gnd FILL
XFILL_1__1374_ vdd gnd FILL
XFILL_2__765_ vdd gnd FILL
X_840_ _903_/B _850_/C vdd gnd INVX1
X_771_ _773_/A _773_/B _773_/C _772_/A vdd gnd NAND3X1
XFILL_2__1483_ vdd gnd FILL
XFILL_4__1419_ vdd gnd FILL
XFILL_0__1050_ vdd gnd FILL
XFILL_1__921_ vdd gnd FILL
XFILL_1__852_ vdd gnd FILL
X_969_ _969_/A _969_/B _969_/C _986_/A vdd gnd OAI21X1
XFILL_1__783_ vdd gnd FILL
X_1112_ _1112_/A _1112_/B _1112_/C _1121_/A vdd gnd NAND3X1
X_1043_ _966_/A _1043_/B _963_/C _1052_/C vdd gnd OAI21X1
XFILL_3__1026_ vdd gnd FILL
XFILL_1__1090_ vdd gnd FILL
XFILL_0__1317_ vdd gnd FILL
XFILL_0__1248_ vdd gnd FILL
XFILL_0__1179_ vdd gnd FILL
XFILL_1__1426_ vdd gnd FILL
XFILL_1__1357_ vdd gnd FILL
XFILL_2__817_ vdd gnd FILL
XFILL_0__870_ vdd gnd FILL
XFILL_1__1288_ vdd gnd FILL
X_823_ _856_/C _823_/B _823_/C _835_/B vdd gnd OAI21X1
XFILL_2__1466_ vdd gnd FILL
XFILL_0__1102_ vdd gnd FILL
XFILL_2__1397_ vdd gnd FILL
XFILL_0__999_ vdd gnd FILL
XFILL_0__1033_ vdd gnd FILL
XFILL_1__904_ vdd gnd FILL
XFILL_1__835_ vdd gnd FILL
XFILL_3__1575_ vdd gnd FILL
X_1026_ _998_/C _998_/B _998_/A _1027_/B vdd gnd AOI21X1
XFILL_1__766_ vdd gnd FILL
XFILL_1__1211_ vdd gnd FILL
XFILL_3__1009_ vdd gnd FILL
XFILL_1__1142_ vdd gnd FILL
XFILL_1__1073_ vdd gnd FILL
XFILL_2__1320_ vdd gnd FILL
XFILL_0__922_ vdd gnd FILL
XFILL_1__1409_ vdd gnd FILL
XFILL_2__1251_ vdd gnd FILL
XFILL_2__1182_ vdd gnd FILL
XFILL_0__784_ vdd gnd FILL
XFILL_0__853_ vdd gnd FILL
XFILL_2_BUFX2_insert8 vdd gnd FILL
XFILL88050x74250 vdd gnd FILL
XFILL_3__995_ vdd gnd FILL
X_806_ Cin[1] Xin[2] _837_/A vdd gnd NAND2X1
XFILL_2__1518_ vdd gnd FILL
XFILL_0__1582_ vdd gnd FILL
XFILL_2__1449_ vdd gnd FILL
XFILL_3__1360_ vdd gnd FILL
XFILL_3__1291_ vdd gnd FILL
XFILL_0__1016_ vdd gnd FILL
X_1575_ _1575_/A Yout[15] vdd gnd BUFX2
XFILL_1__818_ vdd gnd FILL
X_1009_ _1022_/A _1022_/B _948_/Y _1113_/A vdd gnd NAND3X1
XFILL_3__1489_ vdd gnd FILL
XFILL_1__1056_ vdd gnd FILL
XFILL_1__1125_ vdd gnd FILL
XFILL_3__780_ vdd gnd FILL
XFILL_2__1303_ vdd gnd FILL
XFILL_0__905_ vdd gnd FILL
XFILL_2__1096_ vdd gnd FILL
XFILL_2__1165_ vdd gnd FILL
XFILL_2__1234_ vdd gnd FILL
XFILL_0__836_ vdd gnd FILL
XFILL_0__767_ vdd gnd FILL
X_1360_ _1414_/A _1360_/B _1360_/C _1361_/B vdd gnd NAND3X1
XFILL_3__978_ vdd gnd FILL
XFILL_3__1343_ vdd gnd FILL
XFILL_3__1412_ vdd gnd FILL
X_1291_ _1300_/B _1358_/C _1300_/A _1292_/B vdd gnd AOI21X1
XFILL_0__1565_ vdd gnd FILL
XFILL_3__1274_ vdd gnd FILL
XFILL_0__1496_ vdd gnd FILL
X_1489_ _1513_/B _1513_/A _1489_/C _1489_/D _1505_/B vdd gnd AOI22X1
X_1558_ _1558_/D _1559_/CLK _1558_/Q vdd gnd DFFPOSX1
XFILL_2__996_ vdd gnd FILL
XFILL_1__1108_ vdd gnd FILL
XFILL_3__901_ vdd gnd FILL
XFILL_1__1039_ vdd gnd FILL
XFILL_3__832_ vdd gnd FILL
XFILL_3__763_ vdd gnd FILL
XFILL_2__1217_ vdd gnd FILL
XFILL_0__1350_ vdd gnd FILL
XFILL_0__1281_ vdd gnd FILL
XFILL_0_CLKBUF1_insert2 vdd gnd FILL
XFILL_0__819_ vdd gnd FILL
XFILL_2__1148_ vdd gnd FILL
XFILL_2__1079_ vdd gnd FILL
X_1343_ _1343_/A _1396_/A _1369_/A vdd gnd AND2X2
X_1412_ _1412_/A _1412_/B _1412_/C _1511_/A vdd gnd OAI21X1
X_1274_ _1357_/C _1357_/B _1357_/A _1358_/C vdd gnd NAND3X1
XFILL_1__1390_ vdd gnd FILL
XFILL_3__1326_ vdd gnd FILL
XFILL_2__850_ vdd gnd FILL
XFILL_2__781_ vdd gnd FILL
XFILL_0__1479_ vdd gnd FILL
XFILL_3__1257_ vdd gnd FILL
XFILL_3__1188_ vdd gnd FILL
XFILL_2__979_ vdd gnd FILL
XFILL_2__1002_ vdd gnd FILL
X_985_ _994_/B _994_/C _994_/A _999_/A vdd gnd AOI21X1
XFILL_3__815_ vdd gnd FILL
XFILL_3__1111_ vdd gnd FILL
XFILL_3__1042_ vdd gnd FILL
XFILL_0__1264_ vdd gnd FILL
XFILL_0__1402_ vdd gnd FILL
XFILL_0__1333_ vdd gnd FILL
XFILL_0__1195_ vdd gnd FILL
XFILL_1__997_ vdd gnd FILL
XFILL_1__1511_ vdd gnd FILL
X_1326_ _1326_/A _1326_/B _1326_/C _1327_/C vdd gnd OAI21X1
XFILL_1__1373_ vdd gnd FILL
XFILL_1__1442_ vdd gnd FILL
XFILL_3__1309_ vdd gnd FILL
X_1257_ _965_/B _1470_/A _1320_/B _1258_/C vdd gnd OAI21X1
X_1188_ _1188_/A _1188_/B _1266_/A vdd gnd AND2X2
XFILL_2__833_ vdd gnd FILL
XFILL_2__902_ vdd gnd FILL
XFILL_2__764_ vdd gnd FILL
X_770_ _777_/B _770_/B _777_/A _773_/B vdd gnd OAI21X1
XFILL_2__1482_ vdd gnd FILL
X_968_ _977_/A _970_/B Yin[5] _969_/B vdd gnd AOI21X1
XFILL_1__851_ vdd gnd FILL
XFILL_1__920_ vdd gnd FILL
X_899_ Cin[2] _961_/A _952_/B vdd gnd NAND2X1
XFILL_1__782_ vdd gnd FILL
X_1111_ _1209_/A _1115_/B _1115_/A _1112_/C vdd gnd NAND3X1
X_1042_ _962_/C _1047_/B _1043_/B vdd gnd AND2X2
XFILL_3__1025_ vdd gnd FILL
XFILL_0__1316_ vdd gnd FILL
XFILL_0__1247_ vdd gnd FILL
XFILL_0__1178_ vdd gnd FILL
X_1309_ _1371_/B _1319_/C _1371_/A _1325_/B vdd gnd OAI21X1
XFILL_4__1203_ vdd gnd FILL
XFILL_1__1425_ vdd gnd FILL
XFILL_1__1356_ vdd gnd FILL
XFILL_1__1287_ vdd gnd FILL
XFILL_2__816_ vdd gnd FILL
X_822_ Xin[1] Cin[3] _856_/C vdd gnd NAND2X1
XFILL_2__1396_ vdd gnd FILL
XFILL_2__1465_ vdd gnd FILL
XFILL_0__998_ vdd gnd FILL
XFILL_0__1101_ vdd gnd FILL
XFILL_0__1032_ vdd gnd FILL
XFILL_1__903_ vdd gnd FILL
XFILL_1__834_ vdd gnd FILL
XFILL_1__765_ vdd gnd FILL
XFILL_3__1574_ vdd gnd FILL
XFILL_4__976_ vdd gnd FILL
X_1025_ _1209_/A _1124_/A vdd gnd INVX1
XFILL_1__1141_ vdd gnd FILL
XFILL_1__1210_ vdd gnd FILL
XFILL_3__1008_ vdd gnd FILL
XFILL_1__1072_ vdd gnd FILL
XFILL_2__1250_ vdd gnd FILL
XFILL_2__1181_ vdd gnd FILL
XFILL_0__921_ vdd gnd FILL
XFILL_0__852_ vdd gnd FILL
XFILL_1__1339_ vdd gnd FILL
XFILL_1__1408_ vdd gnd FILL
XFILL88650x23550 vdd gnd FILL
XFILL_0__783_ vdd gnd FILL
XFILL_2_BUFX2_insert9 vdd gnd FILL
XFILL_3__994_ vdd gnd FILL
X_805_ _805_/A _805_/B _805_/C _825_/C vdd gnd OAI21X1
XFILL_0__1581_ vdd gnd FILL
XFILL_2__1448_ vdd gnd FILL
XFILL_2__1517_ vdd gnd FILL
XFILL_3__1290_ vdd gnd FILL
XFILL_2__1379_ vdd gnd FILL
XFILL_0__1015_ vdd gnd FILL
X_1574_ _1574_/A Yout[14] vdd gnd BUFX2
XFILL_1__817_ vdd gnd FILL
XFILL_3__1488_ vdd gnd FILL
X_1008_ _946_/Y _1114_/A vdd gnd INVX1
XFILL_1__1124_ vdd gnd FILL
XFILL_1__1055_ vdd gnd FILL
XFILL88650x35250 vdd gnd FILL
XFILL_2__1233_ vdd gnd FILL
XFILL_2__1302_ vdd gnd FILL
XFILL_0__904_ vdd gnd FILL
XFILL_0__835_ vdd gnd FILL
XFILL_2__1095_ vdd gnd FILL
XFILL_2__1164_ vdd gnd FILL
XFILL_3__977_ vdd gnd FILL
XFILL_0__766_ vdd gnd FILL
XFILL_0__1564_ vdd gnd FILL
XFILL_3__1342_ vdd gnd FILL
XFILL_3__1411_ vdd gnd FILL
X_1290_ _1290_/A _1290_/B _1358_/A _1292_/A vdd gnd AOI21X1
XFILL_3__1273_ vdd gnd FILL
XFILL_0__1495_ vdd gnd FILL
XFILL_2_BUFX2_insert10 vdd gnd FILL
X_1557_ _1557_/D _1557_/CLK _1557_/Q vdd gnd DFFPOSX1
XFILL_4__1451_ vdd gnd FILL
X_1488_ _1488_/A _1488_/B _1488_/C _1513_/A vdd gnd OAI21X1
XFILL_4__1382_ vdd gnd FILL
XFILL_2__995_ vdd gnd FILL
XFILL_1__1107_ vdd gnd FILL
XFILL_3__831_ vdd gnd FILL
XFILL_3__900_ vdd gnd FILL
XFILL_1__1038_ vdd gnd FILL
XFILL_3__762_ vdd gnd FILL
XFILL_2__1216_ vdd gnd FILL
XFILL_0__1280_ vdd gnd FILL
XFILL_0__818_ vdd gnd FILL
XFILL_0_CLKBUF1_insert3 vdd gnd FILL
XFILL_2__1078_ vdd gnd FILL
XFILL_2__1147_ vdd gnd FILL
X_1273_ _1303_/A _1348_/C _1303_/B _1357_/A vdd gnd OAI21X1
X_1342_ _1342_/A _1369_/B _1345_/A vdd gnd NAND2X1
X_1411_ _1415_/C _1458_/A _1415_/A _1412_/B vdd gnd AOI21X1
XFILL_3__1325_ vdd gnd FILL
XFILL_3__1256_ vdd gnd FILL
XFILL_2__780_ vdd gnd FILL
XFILL_3__1187_ vdd gnd FILL
XFILL_0__1478_ vdd gnd FILL
XFILL_2__1001_ vdd gnd FILL
XFILL_2__978_ vdd gnd FILL
XFILL_3__814_ vdd gnd FILL
X_984_ _986_/B _986_/C _987_/C _994_/C vdd gnd NAND3X1
XFILL_3__1110_ vdd gnd FILL
XFILL_0__1401_ vdd gnd FILL
XFILL_3__1041_ vdd gnd FILL
XFILL_0__1194_ vdd gnd FILL
XFILL_0__1263_ vdd gnd FILL
XFILL_0__1332_ vdd gnd FILL
XFILL_1__996_ vdd gnd FILL
XFILL_1__1510_ vdd gnd FILL
X_1325_ _1325_/A _1325_/B _1325_/C _1327_/B vdd gnd NAND3X1
X_1256_ _964_/A _1468_/A _1336_/A _1258_/B vdd gnd OAI21X1
XFILL_2__901_ vdd gnd FILL
X_1187_ _1187_/A _1187_/B _1187_/C _1195_/C vdd gnd AOI21X1
XFILL_3__1308_ vdd gnd FILL
XFILL_1__1441_ vdd gnd FILL
XFILL_1__1372_ vdd gnd FILL
XFILL_3__1239_ vdd gnd FILL
XFILL_2__832_ vdd gnd FILL
XFILL_2__763_ vdd gnd FILL
XFILL_2__1481_ vdd gnd FILL
XFILL_1__850_ vdd gnd FILL
X_967_ _992_/B _992_/A _994_/A vdd gnd NAND2X1
X_898_ Cin[2] _961_/A _952_/A _901_/B vdd gnd NAND3X1
XFILL_1__781_ vdd gnd FILL
X_1110_ _1208_/A _1208_/B _1110_/C _1115_/A vdd gnd NAND3X1
X_1041_ Cin[2] Xin[4] _1047_/B vdd gnd NAND2X1
XFILL_0__1177_ vdd gnd FILL
XFILL_3__1024_ vdd gnd FILL
XFILL_0__1246_ vdd gnd FILL
XFILL_0__1315_ vdd gnd FILL
XFILL_1__979_ vdd gnd FILL
X_1308_ _1436_/A Cin[5] Xin[4] Cin[6] _1371_/B vdd gnd AOI22X1
XFILL_1__1424_ vdd gnd FILL
X_1239_ _1239_/A _1336_/A _1239_/C _1239_/D _1243_/B vdd gnd AOI22X1
XFILL_2__815_ vdd gnd FILL
XFILL_4__1064_ vdd gnd FILL
XFILL_4__1133_ vdd gnd FILL
XFILL_1__1355_ vdd gnd FILL
XFILL_1__1286_ vdd gnd FILL
X_821_ _877_/A _872_/B _872_/A _877_/B vdd gnd NAND3X1
XFILL_2__1395_ vdd gnd FILL
XFILL_2__1464_ vdd gnd FILL
XFILL_0__997_ vdd gnd FILL
XFILL_0__1100_ vdd gnd FILL
XFILL_0__1031_ vdd gnd FILL
XFILL_1__902_ vdd gnd FILL
XFILL_1__833_ vdd gnd FILL
X_1024_ _997_/B _997_/A _1209_/A vdd gnd NAND2X1
XFILL_1__764_ vdd gnd FILL
XFILL_3__1573_ vdd gnd FILL
XFILL_1__1140_ vdd gnd FILL
XFILL_3__1007_ vdd gnd FILL
XFILL_1__1071_ vdd gnd FILL
XFILL_0__1229_ vdd gnd FILL
XFILL_1__1407_ vdd gnd FILL
XFILL_2__1180_ vdd gnd FILL
XFILL_0__851_ vdd gnd FILL
XFILL_0__920_ vdd gnd FILL
XFILL_0__782_ vdd gnd FILL
XFILL_1__1338_ vdd gnd FILL
XFILL_1__1269_ vdd gnd FILL
XFILL_3__993_ vdd gnd FILL
XFILL_0__1580_ vdd gnd FILL
X_804_ _884_/A _823_/C _872_/A vdd gnd AND2X2
XFILL_2__1516_ vdd gnd FILL
XFILL_4__760_ vdd gnd FILL
XFILL_2__1447_ vdd gnd FILL
XFILL_2__1378_ vdd gnd FILL
XFILL_0__1014_ vdd gnd FILL
X_1573_ _1573_/A Yout[13] vdd gnd BUFX2
X_1007_ _1015_/C _1015_/B _946_/Y _1012_/B vdd gnd AOI21X1
XFILL_1__816_ vdd gnd FILL
XFILL_3__1487_ vdd gnd FILL
XFILL_4__889_ vdd gnd FILL
XFILL_1__1123_ vdd gnd FILL
XFILL_1__1054_ vdd gnd FILL
XFILL_4__958_ vdd gnd FILL
XFILL_2__1232_ vdd gnd FILL
XFILL88950x19650 vdd gnd FILL
XFILL_2__1163_ vdd gnd FILL
XFILL_2__1301_ vdd gnd FILL
XFILL_0__903_ vdd gnd FILL
XFILL_0__834_ vdd gnd FILL
XFILL_2__1094_ vdd gnd FILL
XFILL_0__765_ vdd gnd FILL
XFILL_3__976_ vdd gnd FILL
XFILL_0__1563_ vdd gnd FILL
XFILL_3__1272_ vdd gnd FILL
XFILL_3__1341_ vdd gnd FILL
XFILL_3__1410_ vdd gnd FILL
XFILL_0__1494_ vdd gnd FILL
XFILL_2_BUFX2_insert11 vdd gnd FILL
X_1556_ _1556_/D _1559_/CLK _1556_/Q vdd gnd DFFPOSX1
X_1487_ _1512_/C _1489_/D vdd gnd INVX1
XFILL_2__994_ vdd gnd FILL
XFILL_1__1106_ vdd gnd FILL
XFILL_1__1037_ vdd gnd FILL
XFILL_3__830_ vdd gnd FILL
XFILL_3__761_ vdd gnd FILL
XFILL_4__1579_ vdd gnd FILL
XFILL_2__1146_ vdd gnd FILL
XFILL_2__1215_ vdd gnd FILL
XFILL_0__817_ vdd gnd FILL
XFILL_0_CLKBUF1_insert4 vdd gnd FILL
XFILL_2__1077_ vdd gnd FILL
X_1410_ _1459_/A _1459_/B _1415_/C vdd gnd NAND2X1
XFILL_3__959_ vdd gnd FILL
X_1272_ _1344_/B _1278_/B _1277_/A _1303_/A vdd gnd AOI21X1
X_1341_ _1367_/B _1349_/B _1406_/A vdd gnd AND2X2
XFILL_0__1477_ vdd gnd FILL
XFILL_3__1255_ vdd gnd FILL
XFILL_3__1324_ vdd gnd FILL
XFILL_3__1186_ vdd gnd FILL
X_1539_ _1555_/Q _1557_/CLK _1571_/A vdd gnd DFFPOSX1
XFILL_4__1502_ vdd gnd FILL
XFILL_4__1433_ vdd gnd FILL
XFILL_4__1364_ vdd gnd FILL
XFILL_4__1295_ vdd gnd FILL
XFILL_2__977_ vdd gnd FILL
XFILL_2__1000_ vdd gnd FILL
XFILL_3__813_ vdd gnd FILL
X_983_ _983_/A _983_/B _983_/C _986_/C vdd gnd NAND3X1
XFILL_3__1040_ vdd gnd FILL
XFILL_0__1400_ vdd gnd FILL
XFILL_0__1331_ vdd gnd FILL
XFILL_2__1129_ vdd gnd FILL
XFILL_0__1193_ vdd gnd FILL
XFILL_0__1262_ vdd gnd FILL
XFILL_1__995_ vdd gnd FILL
X_1186_ _1186_/A _1187_/C vdd gnd INVX1
X_1255_ _1321_/A _1321_/B _1316_/C _1261_/A vdd gnd NAND3X1
XFILL_1__1440_ vdd gnd FILL
X_1324_ _1324_/A _1327_/A vdd gnd INVX1
XFILL_2__831_ vdd gnd FILL
XFILL_2__900_ vdd gnd FILL
XFILL_3__1238_ vdd gnd FILL
XFILL_1__1371_ vdd gnd FILL
XFILL_3__1307_ vdd gnd FILL
XFILL_3__1169_ vdd gnd FILL
XFILL_2__762_ vdd gnd FILL
XFILL_1__1569_ vdd gnd FILL
XFILL_2__1480_ vdd gnd FILL
XFILL_1__780_ vdd gnd FILL
X_897_ _897_/A _897_/B _897_/C _952_/C vdd gnd NAND3X1
X_966_ _966_/A _966_/B _966_/C _992_/A vdd gnd NAND3X1
X_1040_ _1045_/C _1045_/A _1045_/B _1051_/B vdd gnd NAND3X1
XFILL_3__1023_ vdd gnd FILL
XFILL_0__1314_ vdd gnd FILL
XFILL_0__1245_ vdd gnd FILL
XFILL_0__1176_ vdd gnd FILL
XFILL_1__978_ vdd gnd FILL
X_1238_ _1304_/A _1304_/B _1238_/C _1244_/B vdd gnd NOR3X1
XFILL_1__1423_ vdd gnd FILL
X_1307_ _1307_/A _1381_/A _1319_/C vdd gnd NOR2X1
X_1169_ _1235_/A _1169_/B _1169_/C _1188_/B vdd gnd NAND3X1
XFILL_2__814_ vdd gnd FILL
XFILL_1__1354_ vdd gnd FILL
XFILL_1__1285_ vdd gnd FILL
X_820_ _820_/A _820_/B _820_/C _872_/B vdd gnd OAI21X1
XFILL_2__1463_ vdd gnd FILL
XFILL_2__1394_ vdd gnd FILL
XFILL_0__996_ vdd gnd FILL
XFILL_0__1030_ vdd gnd FILL
XFILL_1__832_ vdd gnd FILL
XFILL_1__901_ vdd gnd FILL
XFILL_3__1572_ vdd gnd FILL
X_1023_ _946_/Y _1023_/B _1113_/A _1112_/A vdd gnd OAI21X1
X_949_ Xin[1] Cin[6] _951_/B vdd gnd AND2X2
XFILL_1__763_ vdd gnd FILL
XFILL_1__1070_ vdd gnd FILL
XFILL_3__1006_ vdd gnd FILL
XFILL_0__1228_ vdd gnd FILL
XFILL_0__1159_ vdd gnd FILL
XFILL_4__1115_ vdd gnd FILL
XFILL89250x54750 vdd gnd FILL
XFILL_1__1406_ vdd gnd FILL
XFILL_1__1337_ vdd gnd FILL
XFILL_0__850_ vdd gnd FILL
XFILL_0__781_ vdd gnd FILL
XFILL_1__1199_ vdd gnd FILL
XFILL_4__1046_ vdd gnd FILL
XFILL_1__1268_ vdd gnd FILL
XFILL_3__992_ vdd gnd FILL
X_803_ _861_/C _803_/B _884_/A vdd gnd NAND2X1
XFILL_2__1446_ vdd gnd FILL
XFILL_2__1515_ vdd gnd FILL
XFILL_2__1377_ vdd gnd FILL
XFILL_0__979_ vdd gnd FILL
XFILL_0__1013_ vdd gnd FILL
X_1572_ _1572_/A Yout[12] vdd gnd BUFX2
XFILL_1__815_ vdd gnd FILL
X_1006_ _1022_/A _1022_/B _1010_/C _1015_/C vdd gnd NAND3X1
XFILL_3__1486_ vdd gnd FILL
XFILL_1__1122_ vdd gnd FILL
XFILL_1__1053_ vdd gnd FILL
XFILL89550x31350 vdd gnd FILL
XFILL_2__1300_ vdd gnd FILL
XFILL_0__902_ vdd gnd FILL
XFILL_2__1093_ vdd gnd FILL
XFILL_2__1231_ vdd gnd FILL
XFILL_2__1162_ vdd gnd FILL
XFILL_0__833_ vdd gnd FILL
XFILL_0__764_ vdd gnd FILL
XFILL_3__975_ vdd gnd FILL
XFILL_0__1562_ vdd gnd FILL
XFILL_3__1271_ vdd gnd FILL
XFILL_3__1340_ vdd gnd FILL
XFILL_2__1429_ vdd gnd FILL
XFILL_0__1493_ vdd gnd FILL
XFILL_4__811_ vdd gnd FILL
XFILL_2_BUFX2_insert12 vdd gnd FILL
X_1555_ _1555_/D _1557_/CLK _1555_/Q vdd gnd DFFPOSX1
X_1486_ _1486_/A _1488_/C _1486_/C _1512_/C vdd gnd NAND3X1
XFILL_2__993_ vdd gnd FILL
XFILL89550x43050 vdd gnd FILL
XFILL_3__1469_ vdd gnd FILL
XFILL89250x78150 vdd gnd FILL
XFILL_1__1105_ vdd gnd FILL
XFILL_1__1036_ vdd gnd FILL
XFILL_3__760_ vdd gnd FILL
XFILL_2__1145_ vdd gnd FILL
XFILL_2__1076_ vdd gnd FILL
XFILL_2__1214_ vdd gnd FILL
XFILL_0_CLKBUF1_insert5 vdd gnd FILL
XFILL_0__816_ vdd gnd FILL
X_1340_ _1370_/A _1370_/B _1354_/A vdd gnd NOR2X1
XFILL_3__889_ vdd gnd FILL
XFILL_3__958_ vdd gnd FILL
X_1271_ _1278_/C _1277_/B _1348_/C vdd gnd NOR2X1
XFILL_3__1185_ vdd gnd FILL
XFILL_0__1476_ vdd gnd FILL
XFILL_3__1323_ vdd gnd FILL
XFILL_3__1254_ vdd gnd FILL
X_1538_ _1554_/Q _1557_/CLK _1570_/A vdd gnd DFFPOSX1
X_1469_ _1507_/B _1507_/C _1471_/A vdd gnd NAND2X1
XFILL_2__976_ vdd gnd FILL
XFILL_1__1019_ vdd gnd FILL
XFILL_3__812_ vdd gnd FILL
X_982_ _982_/A _982_/B _982_/C _986_/B vdd gnd NAND3X1
XFILL_0__1330_ vdd gnd FILL
XFILL_0__1261_ vdd gnd FILL
XFILL_2__1128_ vdd gnd FILL
XFILL_2__1059_ vdd gnd FILL
XFILL_0__1192_ vdd gnd FILL
XFILL_1__994_ vdd gnd FILL
X_1323_ _1324_/A _1367_/A _1323_/C _1367_/B vdd gnd NAND3X1
XFILL_3__1306_ vdd gnd FILL
X_1185_ _1195_/B _1195_/A _1220_/C _1201_/B vdd gnd OAI21X1
XFILL_1__1370_ vdd gnd FILL
X_1254_ _964_/A _1468_/A _965_/B _1470_/A _1321_/B vdd gnd OAI22X1
XFILL_2__830_ vdd gnd FILL
XFILL_2__761_ vdd gnd FILL
XFILL_3__1237_ vdd gnd FILL
XFILL_0__1459_ vdd gnd FILL
XFILL_3__1168_ vdd gnd FILL
XFILL_3__1099_ vdd gnd FILL
XFILL_1__1568_ vdd gnd FILL
XFILL_1__1499_ vdd gnd FILL
XFILL_2__959_ vdd gnd FILL
X_965_ _965_/A _965_/B _965_/C _966_/C vdd gnd OAI21X1
X_896_ _964_/A _965_/A _952_/A _897_/B vdd gnd OAI21X1
XFILL_4__990_ vdd gnd FILL
XFILL_3__1022_ vdd gnd FILL
XFILL_0__1244_ vdd gnd FILL
XFILL_0__1313_ vdd gnd FILL
XFILL_0__1175_ vdd gnd FILL
XFILL_1__977_ vdd gnd FILL
X_1306_ _1436_/A Cin[5] _1381_/A vdd gnd NAND2X1
X_1099_ _1099_/A _1099_/B _1127_/C _1105_/B vdd gnd OAI21X1
X_1237_ _1304_/C _1237_/B _1237_/C _1244_/A vdd gnd AOI21X1
XFILL_1__1353_ vdd gnd FILL
XFILL_1__1422_ vdd gnd FILL
X_1168_ Cin[2] Xin[6] _1234_/A _1169_/C vdd gnd NAND3X1
XFILL_2__813_ vdd gnd FILL
XFILL_1__1284_ vdd gnd FILL
XFILL_2__1462_ vdd gnd FILL
XFILL_2__1393_ vdd gnd FILL
XFILL_0__995_ vdd gnd FILL
XFILL_1__831_ vdd gnd FILL
X_948_ _948_/A _948_/B _948_/C _948_/Y vdd gnd OAI21X1
XFILL_1__900_ vdd gnd FILL
XFILL_3__1571_ vdd gnd FILL
X_879_ _936_/C _884_/B _884_/A _882_/C vdd gnd OAI21X1
X_1022_ _1022_/A _1022_/B _948_/Y _1023_/B vdd gnd AOI21X1
XFILL_1__762_ vdd gnd FILL
XFILL_3__1005_ vdd gnd FILL
XFILL_0__1227_ vdd gnd FILL
XFILL_0__1089_ vdd gnd FILL
XFILL_0__1158_ vdd gnd FILL
XFILL_1__1405_ vdd gnd FILL
XFILL_1__1336_ vdd gnd FILL
XFILL_0__780_ vdd gnd FILL
XFILL_1__1198_ vdd gnd FILL
XFILL_1__1267_ vdd gnd FILL
XFILL_3__991_ vdd gnd FILL
X_802_ Xin[1] Cin[3] _861_/C vdd gnd AND2X2
XFILL_2__1376_ vdd gnd FILL
XFILL_2__1445_ vdd gnd FILL
XFILL_2__1514_ vdd gnd FILL
XFILL_0__978_ vdd gnd FILL
XFILL_0__1012_ vdd gnd FILL
X_1571_ _1571_/A Yout[11] vdd gnd BUFX2
XFILL_1__814_ vdd gnd FILL
XFILL_3__1485_ vdd gnd FILL
X_1005_ _996_/C _996_/B _996_/A _1022_/B vdd gnd NAND3X1
XFILL_1__1121_ vdd gnd FILL
XFILL_1__1052_ vdd gnd FILL
XFILL_2__1230_ vdd gnd FILL
XFILL_0__832_ vdd gnd FILL
XFILL_2__1092_ vdd gnd FILL
XFILL_0__901_ vdd gnd FILL
XFILL_4__1028_ vdd gnd FILL
XFILL_1__1319_ vdd gnd FILL
XFILL_2__1161_ vdd gnd FILL
XFILL_0__763_ vdd gnd FILL
XFILL_3__974_ vdd gnd FILL
XFILL_0__1561_ vdd gnd FILL
XFILL_2__1359_ vdd gnd FILL
XFILL_2__1428_ vdd gnd FILL
XFILL_3__1270_ vdd gnd FILL
XFILL_0__1492_ vdd gnd FILL
XFILL_2_BUFX2_insert13 vdd gnd FILL
X_1485_ _1488_/A _1488_/B _1513_/B vdd gnd NAND2X1
X_1554_ _1554_/D _1557_/CLK _1554_/Q vdd gnd DFFPOSX1
.ends


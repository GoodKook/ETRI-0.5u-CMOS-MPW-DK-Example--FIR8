/* Verilog module written by vlog2Verilog (qflow) */
/* With bit-blasted vectors */
/* With power connections converted to binary 1, 0 */

module fir_pe(
    input [7:0] Cin,
    input [7:0] Xin,
    output [7:0] Xout,
    input [15:0] Yin,
    output [15:0] Yout,
    input clk
);

wire [15:0] y ;
wire _588_ ;
wire _168_ ;
wire _60_ ;
wire _397_ ;
wire _703_ ;
wire _19_ ;
wire _512_ ;
wire _741_ ;
wire _321_ ;
wire _57_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _415_ ;
wire _95_ ;
wire _644_ ;
wire _224_ ;
wire _453_ ;
wire _509_ ;
wire _682_ ;
wire _262_ ;
wire _738_ ;
wire _318_ ;
wire _491_ ;
wire _547_ ;
wire _127_ ;
wire _356_ ;
wire _585_ ;
wire _165_ ;
wire _394_ ;
wire _679_ ;
wire _259_ ;
wire _488_ ;
wire _700_ ;
wire _297_ ;
wire _16_ ;
wire _54_ ;
wire _603_ ;
wire _412_ ;
wire _92_ ;
wire _641_ ;
wire _221_ ;
wire _450_ ;
wire _506_ ;
wire _735_ ;
wire _315_ ;
wire _544_ ;
wire _124_ ;
wire _353_ ;
wire _409_ ;
wire _89_ ;
wire _582_ ;
wire _162_ ;
wire _638_ ;
wire _218_ ;
wire _391_ ;
wire _447_ ;
wire _676_ ;
wire _256_ ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire _388_ ;
wire _600_ ;
wire _197_ ;
wire _7_ ;
wire _503_ ;
wire _732_ ;
wire _312_ ;
wire _48_ ;
wire _541_ ;
wire _121_ ;
wire _350_ ;
wire _406_ ;
wire _86_ ;
wire _635_ ;
wire _215_ ;
wire _444_ ;
wire _673_ ;
wire _253_ ;
wire _729_ ;
wire _309_ ;
wire _482_ ;
wire _538_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _347_ ;
wire _576_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire _479_ ;
wire _288_ ;
wire _4_ ;
wire _500_ ;
wire _45_ ;
wire _403_ ;
wire _83_ ;
wire _632_ ;
wire _212_ ;
wire _441_ ;
wire _670_ ;
wire _250_ ;
wire _726_ ;
wire _306_ ;
wire _535_ ;
wire _115_ ;
wire _344_ ;
wire _573_ ;
wire _153_ ;
wire _629_ ;
wire _209_ ;
wire Xin_5_bF$buf0 ;
wire Xin_5_bF$buf1 ;
wire Xin_5_bF$buf2 ;
wire Xin_5_bF$buf3 ;
wire _382_ ;
wire _438_ ;
wire _191_ ;
wire _667_ ;
wire _247_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire _285_ ;
wire _1_ ;
wire _42_ ;
wire _379_ ;
wire _188_ ;
wire _400_ ;
wire _80_ ;
wire _723_ ;
wire _303_ ;
wire _39_ ;
wire _532_ ;
wire _112_ ;
wire _341_ ;
wire clk ;
wire _77_ ;
wire _570_ ;
wire _150_ ;
wire _626_ ;
wire _206_ ;
wire _435_ ;
wire _664_ ;
wire _244_ ;
wire _473_ ;
wire _529_ ;
wire _109_ ;
wire _282_ ;
wire _338_ ;
wire _567_ ;
wire _147_ ;
wire _376_ ;
wire _185_ ;
wire _699_ ;
wire _279_ ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire _74_ ;
wire _623_ ;
wire _203_ ;
wire _432_ ;
wire _661_ ;
wire _241_ ;
wire _717_ ;
wire _470_ ;
wire _526_ ;
wire _106_ ;
wire [15:0] _755_ ;
wire _335_ ;
wire _564_ ;
wire _144_ ;
wire _373_ ;
wire _429_ ;
wire _182_ ;
wire _658_ ;
wire _238_ ;
wire _467_ ;
wire _696_ ;
wire _276_ ;
wire _33_ ;
wire _599_ ;
wire _179_ ;
wire _71_ ;
wire _620_ ;
wire _200_ ;
wire _714_ ;
wire _523_ ;
wire _103_ ;
wire [4:4] _752_ ;
wire _332_ ;
wire _68_ ;
wire _561_ ;
wire _141_ ;
wire _617_ ;
wire _370_ ;
wire _426_ ;
wire _655_ ;
wire _235_ ;
wire _464_ ;
wire _693_ ;
wire _273_ ;
wire [1:1] _749_ ;
wire _329_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _367_ ;
wire _596_ ;
wire _176_ ;
wire _499_ ;
wire _711_ ;
wire _27_ ;
wire _520_ ;
wire _100_ ;
wire _65_ ;
wire _614_ ;
wire _423_ ;
wire _652_ ;
wire _232_ ;
wire _708_ ;
wire _461_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _746_ ;
wire _326_ ;
wire _555_ ;
wire _135_ ;
wire _364_ ;
wire _593_ ;
wire _173_ ;
wire _649_ ;
wire _229_ ;
wire _458_ ;
wire _687_ ;
wire _267_ ;
wire _496_ ;
wire _24_ ;
wire _62_ ;
wire _399_ ;
wire _611_ ;
wire _420_ ;
wire _705_ ;
wire _514_ ;
wire _743_ ;
wire _323_ ;
wire _59_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _361_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _646_ ;
wire _226_ ;
wire _455_ ;
wire _684_ ;
wire _264_ ;
wire _493_ ;
wire _549_ ;
wire _129_ ;
wire _21_ ;
wire _358_ ;
wire _587_ ;
wire _167_ ;
wire _396_ ;
wire _702_ ;
wire _299_ ;
wire _18_ ;
wire _511_ ;
wire _740_ ;
wire _320_ ;
wire _56_ ;
wire _605_ ;
wire _414_ ;
wire _94_ ;
wire _643_ ;
wire _223_ ;
wire _452_ ;
wire _508_ ;
wire _681_ ;
wire _261_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _546_ ;
wire _126_ ;
wire _355_ ;
wire _584_ ;
wire _164_ ;
wire _393_ ;
wire _449_ ;
wire _678_ ;
wire _258_ ;
wire _487_ ;
wire _296_ ;
wire _15_ ;
wire _53_ ;
wire _602_ ;
wire _199_ ;
wire _411_ ;
wire _91_ ;
wire _640_ ;
wire _220_ ;
wire _9_ ;
wire _505_ ;
wire _734_ ;
wire _314_ ;
wire _543_ ;
wire _123_ ;
wire _352_ ;
wire _408_ ;
wire _88_ ;
wire _581_ ;
wire _161_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _446_ ;
wire [15:0] Yin ;
wire _675_ ;
wire _255_ ;
wire _484_ ;
wire _293_ ;
wire _12_ ;
wire _349_ ;
wire _578_ ;
wire _158_ ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire _6_ ;
wire _502_ ;
wire _731_ ;
wire _311_ ;
wire _47_ ;
wire _540_ ;
wire _120_ ;
wire _405_ ;
wire _85_ ;
wire _634_ ;
wire _214_ ;
wire _443_ ;
wire _672_ ;
wire _252_ ;
wire _728_ ;
wire _308_ ;
wire _481_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _346_ ;
wire _575_ ;
wire _155_ ;
wire _384_ ;
wire _193_ ;
wire _669_ ;
wire _249_ ;
wire _478_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _402_ ;
wire _82_ ;
wire _631_ ;
wire _211_ ;
wire _440_ ;
wire _725_ ;
wire _305_ ;
wire _534_ ;
wire _114_ ;
wire _343_ ;
wire _79_ ;
wire _572_ ;
wire _152_ ;
wire _628_ ;
wire _208_ ;
wire _381_ ;
wire _437_ ;
wire _190_ ;
wire _666_ ;
wire _246_ ;
wire _475_ ;
wire _284_ ;
wire _0_ ;
wire _569_ ;
wire _149_ ;
wire _41_ ;
wire _378_ ;
wire _187_ ;
wire [15:0] Yout ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _531_ ;
wire _111_ ;
wire _340_ ;
wire _76_ ;
wire _625_ ;
wire _205_ ;
wire _434_ ;
wire _663_ ;
wire _243_ ;
wire _719_ ;
wire _472_ ;
wire _528_ ;
wire _108_ ;
wire _281_ ;
wire _337_ ;
wire _566_ ;
wire _146_ ;
wire _375_ ;
wire _184_ ;
wire _469_ ;
wire _698_ ;
wire _278_ ;
wire _35_ ;
wire [7:0] Xout ;
wire _73_ ;
wire _622_ ;
wire _202_ ;
wire _431_ ;
wire _660_ ;
wire _240_ ;
wire _716_ ;
wire _525_ ;
wire _105_ ;
wire [7:0] _754_ ;
wire _334_ ;
wire _563_ ;
wire _143_ ;
wire _619_ ;
wire _372_ ;
wire _428_ ;
wire _181_ ;
wire _657_ ;
wire _237_ ;
wire _466_ ;
wire _695_ ;
wire _275_ ;
wire _32_ ;
wire _369_ ;
wire _598_ ;
wire _178_ ;
wire _70_ ;
wire _713_ ;
wire _29_ ;
wire _522_ ;
wire _102_ ;
wire [3:3] _751_ ;
wire _331_ ;
wire _67_ ;
wire _560_ ;
wire _140_ ;
wire _616_ ;
wire _425_ ;
wire _654_ ;
wire _234_ ;
wire _463_ ;
wire _519_ ;
wire _692_ ;
wire _272_ ;
wire [0:0] _748_ ;
wire _328_ ;
wire _557_ ;
wire _137_ ;
wire _366_ ;
wire _595_ ;
wire _175_ ;
wire _689_ ;
wire _269_ ;
wire _498_ ;
wire _710_ ;
wire _26_ ;
wire Cin_0_bF$buf0 ;
wire Cin_0_bF$buf1 ;
wire Cin_0_bF$buf2 ;
wire Cin_0_bF$buf3 ;
wire _64_ ;
wire _613_ ;
wire _422_ ;
wire _651_ ;
wire _231_ ;
wire _707_ ;
wire _460_ ;
wire _516_ ;
wire _745_ ;
wire _325_ ;
wire _554_ ;
wire _134_ ;
wire _363_ ;
wire _419_ ;
wire _99_ ;
wire _592_ ;
wire _172_ ;
wire _648_ ;
wire _228_ ;
wire _457_ ;
wire _686_ ;
wire _266_ ;
wire _495_ ;
wire _23_ ;
wire _589_ ;
wire _169_ ;
wire _61_ ;
wire _398_ ;
wire _610_ ;
wire _704_ ;
wire _513_ ;
wire _742_ ;
wire _322_ ;
wire _58_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _360_ ;
wire _416_ ;
wire _96_ ;
wire [7:0] Cin ;
wire _645_ ;
wire _225_ ;
wire _454_ ;
wire _683_ ;
wire _263_ ;
wire _739_ ;
wire _319_ ;
wire _492_ ;
wire _548_ ;
wire _128_ ;
wire _20_ ;
wire _357_ ;
wire _586_ ;
wire _166_ ;
wire _395_ ;
wire _489_ ;
wire _701_ ;
wire _298_ ;
wire _17_ ;
wire _510_ ;
wire _55_ ;
wire _604_ ;
wire _413_ ;
wire _93_ ;
wire _642_ ;
wire _222_ ;
wire _451_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _736_ ;
wire _316_ ;
wire _545_ ;
wire _125_ ;
wire _354_ ;
wire _583_ ;
wire _163_ ;
wire _639_ ;
wire _219_ ;
wire _392_ ;
wire _448_ ;
wire _677_ ;
wire _257_ ;
wire _486_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _601_ ;
wire _198_ ;
wire _410_ ;
wire _90_ ;
wire _8_ ;
wire _504_ ;
wire _733_ ;
wire _313_ ;
wire _49_ ;
wire _542_ ;
wire _122_ ;
wire _351_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _636_ ;
wire _216_ ;
wire _445_ ;
wire _674_ ;
wire _254_ ;
wire _483_ ;
wire _539_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _348_ ;
wire _577_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire _289_ ;
wire _5_ ;
wire _501_ ;
wire _730_ ;
wire _310_ ;
wire _46_ ;
wire _404_ ;
wire _84_ ;
wire _633_ ;
wire _213_ ;
wire _442_ ;
wire _671_ ;
wire _251_ ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire _536_ ;
wire _116_ ;
wire _345_ ;
wire _574_ ;
wire _154_ ;
wire _383_ ;
wire _439_ ;
wire _192_ ;
wire _668_ ;
wire _248_ ;
wire _477_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire _189_ ;
wire _401_ ;
wire _81_ ;
wire _630_ ;
wire _210_ ;
wire _724_ ;
wire _304_ ;
wire _533_ ;
wire _113_ ;
wire _342_ ;
wire _78_ ;
wire _571_ ;
wire _151_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _436_ ;
wire [7:0] Xin ;
wire _665_ ;
wire _245_ ;
wire _474_ ;
wire _283_ ;
wire _339_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire _377_ ;
wire _186_ ;
wire _721_ ;
wire _301_ ;
wire _37_ ;
wire _530_ ;
wire _110_ ;
wire _75_ ;
wire _624_ ;
wire _204_ ;
wire _433_ ;
wire _662_ ;
wire _242_ ;
wire _718_ ;
wire _471_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _336_ ;
wire _565_ ;
wire _145_ ;
wire _374_ ;
wire _183_ ;
wire _659_ ;
wire _239_ ;
wire _468_ ;
wire _697_ ;
wire _277_ ;
wire _34_ ;
wire _72_ ;
wire _621_ ;
wire _201_ ;
wire _430_ ;
wire _715_ ;
wire _524_ ;
wire _104_ ;
wire [15:5] _753_ ;
wire _333_ ;
wire _69_ ;
wire _562_ ;
wire _142_ ;
wire _618_ ;
wire _371_ ;
wire _427_ ;
wire _180_ ;
wire _656_ ;
wire _236_ ;
wire _465_ ;
wire _694_ ;
wire _274_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _368_ ;
wire _597_ ;
wire _177_ ;
wire _712_ ;
wire _28_ ;
wire _521_ ;
wire _101_ ;
wire [2:2] _750_ ;
wire _330_ ;
wire _66_ ;
wire _615_ ;
wire _424_ ;
wire _653_ ;
wire _233_ ;
wire _709_ ;
wire _462_ ;
wire _518_ ;
wire _691_ ;
wire _271_ ;
wire _747_ ;
wire _327_ ;
wire _556_ ;
wire _136_ ;
wire _365_ ;
wire _594_ ;
wire _174_ ;
wire _459_ ;
wire _688_ ;
wire _268_ ;
wire _497_ ;
wire Xin_3_bF$buf0 ;
wire Xin_3_bF$buf1 ;
wire Xin_3_bF$buf2 ;
wire Xin_3_bF$buf3 ;
wire _25_ ;
wire _63_ ;
wire _612_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire _706_ ;
wire _515_ ;
wire _744_ ;
wire _324_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _362_ ;
wire _418_ ;
wire _98_ ;
wire _591_ ;
wire _171_ ;
wire _647_ ;
wire _227_ ;
wire _456_ ;
wire _685_ ;
wire _265_ ;
wire _494_ ;
wire _22_ ;
wire _359_ ;

FILL FILL_0__1241_ (
);

FILL FILL_2__1259_ (
);

FILL FILL_2__770_ (
);

FILL FILL_1__1402_ (
);

FILL FILL_3__1328_ (
);

OAI21X1 _1257_ (
    .A(_740_),
    .B(_352_),
    .C(_445_),
    .Y(_451_)
);

FILL FILL_3__1081_ (
);

FILL FILL_1__792_ (
);

FILL FILL_2__826_ (
);

FILL FILL_4__1570_ (
);

FILL FILL_0__1470_ (
);

FILL FILL_2__1488_ (
);

FILL FILL_0__1050_ (
);

FILL FILL_2__1068_ (
);

FILL FILL_3__941_ (
);

NAND2X1 _800_ (
    .A(Xin[1]),
    .B(Cin[2]),
    .Y(_741_)
);

FILL FILL_1__1211_ (
);

FILL FILL_3__1137_ (
);

NAND3X1 _1486_ (
    .A(_668_),
    .B(_670_),
    .C(_694_),
    .Y(_696_)
);

OAI21X1 _1066_ (
    .A(_740_),
    .B(_151_),
    .C(_250_),
    .Y(_256_)
);

FILL FILL_1__848_ (
);

FILL FILL_0__1106_ (
);

FILL FILL_2__1297_ (
);

FILL FILL_1__1440_ (
);

FILL FILL_1__1020_ (
);

FILL FILL_3__1366_ (
);

INVX1 _1295_ (
    .A(_489_),
    .Y(_491_)
);

FILL FILL_0__1335_ (
);

FILL FILL_2__864_ (
);

FILL FILL_3__806_ (
);

FILL FILL_3__1175_ (
);

FILL FILL_1__886_ (
);

FILL FILL_4__1244_ (
);

FILL FILL_0__1564_ (
);

FILL FILL_0__1144_ (
);

FILL FILL_1__1305_ (
);

FILL FILL_0__1373_ (
);

FILL FILL_3__844_ (
);

FILL FILL_1__1114_ (
);

NAND3X1 _1389_ (
    .A(_574_),
    .B(_587_),
    .C(_592_),
    .Y(_593_)
);

FILL FILL_0__1429_ (
);

FILL FILL_0__1009_ (
);

FILL FILL_2__958_ (
);

FILL FILL_0__1182_ (
);

OAI21X1 _932_ (
    .A(_119_),
    .B(_118_),
    .C(_82_),
    .Y(_124_)
);

FILL FILL_1__1343_ (
);

FILL FILL_3__1269_ (
);

INVX1 _1198_ (
    .A(_281_),
    .Y(_388_)
);

FILL FILL_2__1412_ (
);

FILL FILL_0__1238_ (
);

FILL FILL_2__767_ (
);

FILL FILL89250x74250 (
);

NAND2X1 _1410_ (
    .A(_611_),
    .B(_608_),
    .Y(_616_)
);

FILL FILL_3__882_ (
);

FILL FILL_1__1572_ (
);

FILL FILL_1__1152_ (
);

FILL FILL_3__1498_ (
);

FILL FILL_3__1078_ (
);

FILL FILL_1__789_ (
);

FILL FILL_2__1221_ (
);

FILL FILL_4__1147_ (
);

FILL FILL_0__1467_ (
);

FILL FILL_0__1047_ (
);

FILL FILL_2__996_ (
);

FILL FILL_3__938_ (
);

FILL FILL88950x19650 (
);

FILL FILL_1__1208_ (
);

NAND2X1 _970_ (
    .A(Cin[1]),
    .B(Xin_5_bF$buf0),
    .Y(_161_)
);

FILL FILL_1__1381_ (
);

FILL FILL_2__1450_ (
);

FILL FILL_2__1030_ (
);

FILL FILL_0__1276_ (
);

FILL FILL_1__1437_ (
);

FILL FILL_1__1017_ (
);

FILL FILL_1__810_ (
);

FILL FILL_1__1190_ (
);

FILL FILL_2__1506_ (
);

FILL FILL_0__1085_ (
);

OAI21X1 _1504_ (
    .A(_686_),
    .B(_701_),
    .C(_712_),
    .Y(_715_)
);

FILL FILL_0__832_ (
);

FILL FILL_3__976_ (
);

OAI21X1 _835_ (
    .A(_18_),
    .B(_16_),
    .C(_9_),
    .Y(_27_)
);

FILL FILL_1__1246_ (
);

FILL FILL_2__1315_ (
);

INVX1 _1313_ (
    .A(_506_),
    .Y(_511_)
);

FILL FILL_3__785_ (
);

FILL FILL_1__1475_ (
);

FILL FILL_1__1055_ (
);

FILL FILL_2__1124_ (
);

FILL FILL_2__899_ (
);

DFFPOSX1 _1542_ (
    .D(y[14]),
    .CLK(clk_bF$buf2),
    .Q(_755_[14])
);

OAI22X1 _1122_ (
    .A(_309_),
    .B(_310_),
    .C(_308_),
    .D(_208_),
    .Y(_311_)
);

FILL FILL_0__870_ (
);

FILL FILL_1__904_ (
);

OAI21X1 _873_ (
    .A(_57_),
    .B(_58_),
    .C(_55_),
    .Y(_65_)
);

FILL FILL_1__1284_ (
);

FILL FILL_2__1353_ (
);

FILL FILL_0__1179_ (
);

FILL FILL_0__926_ (
);

FILL FILL_3__1422_ (
);

FILL FILL_3__1002_ (
);

NAND3X1 _929_ (
    .A(_81_),
    .B(_116_),
    .C(_120_),
    .Y(_121_)
);

NAND3X1 _1351_ (
    .A(_551_),
    .B(_552_),
    .C(_550_),
    .Y(_553_)
);

FILL FILL89550x7950 (
);

FILL FILL_4__857_ (
);

FILL FILL_1__1093_ (
);

FILL FILL_2__1409_ (
);

FILL FILL_2__920_ (
);

FILL FILL_2__1582_ (
);

FILL FILL_2__1162_ (
);

NAND3X1 _1407_ (
    .A(_604_),
    .B(_607_),
    .C(_611_),
    .Y(_613_)
);

FILL FILL_3__879_ (
);

FILL FILL_3__1231_ (
);

FILL FILL_1__1569_ (
);

FILL FILL_1__1149_ (
);

BUFX2 _1580_ (
    .A(_755_[6]),
    .Y(Yout[6])
);

INVX1 _1160_ (
    .A(_348_),
    .Y(_349_)
);

FILL FILL_1__942_ (
);

FILL FILL_0__1200_ (
);

FILL FILL_2__1218_ (
);

FILL FILL_2__1391_ (
);

OAI21X1 _1216_ (
    .A(_404_),
    .B(_405_),
    .C(_403_),
    .Y(_406_)
);

FILL FILL_0__964_ (
);

FILL FILL_3__1460_ (
);

FILL FILL_3__1040_ (
);

NAND2X1 _967_ (
    .A(_154_),
    .B(_157_),
    .Y(_158_)
);

FILL FILL_1__1378_ (
);

FILL FILL_2__1447_ (
);

FILL FILL_2__1027_ (
);

FILL FILL_3__900_ (
);

FILL FILL_3__1516_ (
);

NAND2X1 _1445_ (
    .A(_650_),
    .B(_651_),
    .Y(_653_)
);

INVX1 _1025_ (
    .A(_214_),
    .Y(_215_)
);

FILL FILL_0__773_ (
);

FILL FILL_1__807_ (
);

NOR2X1 _776_ (
    .A(_397_),
    .B(_590_),
    .Y(_601_)
);

FILL FILL_1__1187_ (
);

FILL FILL_1__980_ (
);

FILL FILL_2__1256_ (
);

FILL FILL_0__829_ (
);

FILL FILL_3__1325_ (
);

OAI22X1 _1254_ (
    .A(_590_),
    .B(_447_),
    .C(_740_),
    .D(_352_),
    .Y(_448_)
);

FILL FILL_2__823_ (
);

FILL FILL_2__1485_ (
);

FILL FILL_2__1065_ (
);

FILL FILL_3__1134_ (
);

XOR2X1 _1483_ (
    .A(_693_),
    .B(_674_),
    .Y(_694_)
);

OAI21X1 _1063_ (
    .A(_740_),
    .B(_151_),
    .C(_252_),
    .Y(_253_)
);

FILL FILL_1__845_ (
);

FILL FILL_4__1203_ (
);

FILL FILL_0__1103_ (
);

FILL FILL_2__1294_ (
);

DFFPOSX1 _1539_ (
    .D(y[11]),
    .CLK(clk_bF$buf5),
    .Q(_755_[11])
);

XNOR2X1 _1119_ (
    .A(_211_),
    .B(_308_),
    .Y(_753_[7])
);

FILL FILL_0__867_ (
);

FILL FILL_3__1363_ (
);

OAI21X1 _1292_ (
    .A(_487_),
    .B(_488_),
    .C(_486_),
    .Y(_489_)
);

FILL FILL_0__1332_ (
);

FILL FILL_2__861_ (
);

FILL FILL_3__803_ (
);

FILL FILL_3__1419_ (
);

AOI21X1 _1348_ (
    .A(_439_),
    .B(_463_),
    .C(_466_),
    .Y(_550_)
);

FILL FILL_3__1172_ (
);

FILL FILL_1__883_ (
);

FILL FILL_2__917_ (
);

FILL FILL_2__1579_ (
);

FILL FILL_0__1561_ (
);

FILL FILL_0__1141_ (
);

FILL FILL_2__1159_ (
);

FILL FILL89250x39150 (
);

FILL FILL_1__1302_ (
);

FILL FILL_3__1228_ (
);

BUFX2 _1577_ (
    .A(_755_[3]),
    .Y(Yout[3])
);

AOI21X1 _1157_ (
    .A(_270_),
    .B(_267_),
    .C(_260_),
    .Y(_346_)
);

FILL FILL_1__939_ (
);

FILL FILL_4__1470_ (
);

FILL FILL_2__1388_ (
);

FILL FILL_0__1370_ (
);

FILL FILL_3__841_ (
);

FILL FILL_1__1111_ (
);

FILL FILL_3__1457_ (
);

FILL FILL_3__1037_ (
);

AOI21X1 _1386_ (
    .A(_585_),
    .B(_579_),
    .C(_583_),
    .Y(_589_)
);

FILL FILL_4__1106_ (
);

FILL FILL_0__1426_ (
);

FILL FILL_0__1006_ (
);

FILL FILL_2__955_ (
);

FILL FILL_2__1197_ (
);

FILL FILL_1__1340_ (
);

FILL FILL_3__1266_ (
);

OAI21X1 _1195_ (
    .A(_368_),
    .B(_373_),
    .C(_376_),
    .Y(_384_)
);

FILL FILL_1__977_ (
);

FILL FILL_0__1235_ (
);

FILL FILL_2__764_ (
);

FILL FILL89550x78150 (
);

FILL FILL_0__999_ (
);

FILL FILL_3__1495_ (
);

FILL FILL_3__1075_ (
);

FILL FILL_1__786_ (
);

FILL FILL_0__1464_ (
);

FILL FILL_0__1044_ (
);

FILL FILL_2__993_ (
);

FILL FILL_3__935_ (
);

FILL FILL_1__1205_ (
);

FILL FILL_4__1373_ (
);

FILL FILL_0__1273_ (
);

FILL FILL_1__1434_ (
);

FILL FILL_1__1014_ (
);

AOI21X1 _1289_ (
    .A(_314_),
    .B(_395_),
    .C(_485_),
    .Y(_486_)
);

FILL FILL_2__1503_ (
);

FILL FILL_4__1009_ (
);

FILL FILL_0__1329_ (
);

FILL FILL_2__858_ (
);

FILL FILL_0__1082_ (
);

XNOR2X1 _1501_ (
    .A(_702_),
    .B(_712_),
    .Y(_713_)
);

FILL FILL_3__973_ (
);

OAI21X1 _832_ (
    .A(_22_),
    .B(_21_),
    .C(_735_),
    .Y(_25_)
);

FILL FILL_1__1243_ (
);

FILL FILL_3__1169_ (
);

FILL FILL_4__760_ (
);

NAND2X1 _1098_ (
    .A(_240_),
    .B(_243_),
    .Y(_288_)
);

FILL FILL_2__1312_ (
);

FILL FILL_0__1138_ (
);

INVX1 _1310_ (
    .A(_502_),
    .Y(_508_)
);

FILL FILL_3__782_ (
);

FILL FILL_1__1472_ (
);

FILL FILL_1__1052_ (
);

FILL FILL_3__1398_ (
);

FILL FILL_2__1121_ (
);

FILL FILL_0__1367_ (
);

FILL FILL_2__896_ (
);

FILL FILL_3__838_ (
);

FILL FILL_1__1108_ (
);

FILL FILL_1__901_ (
);

OAI21X1 _870_ (
    .A(_57_),
    .B(_58_),
    .C(_61_),
    .Y(_62_)
);

FILL FILL_1__1281_ (
);

FILL FILL_2__1350_ (
);

FILL FILL_4__1276_ (
);

FILL FILL_0__1176_ (
);

FILL FILL89250x27450 (
);

FILL FILL_0__923_ (
);

AOI21X1 _926_ (
    .A(_113_),
    .B(_114_),
    .C(_112_),
    .Y(_118_)
);

FILL FILL_1__1337_ (
);

FILL FILL_1__1090_ (
);

FILL FILL_2__1406_ (
);

NAND2X1 _1404_ (
    .A(_573_),
    .B(_608_),
    .Y(_609_)
);

FILL FILL_3__876_ (
);

FILL FILL_1__1566_ (
);

FILL FILL_1__1146_ (
);

FILL FILL_2__1215_ (
);

NAND2X1 _1213_ (
    .A(_403_),
    .B(_398_),
    .Y(_404_)
);

FILL FILL_0__961_ (
);

OAI21X1 _964_ (
    .A(_590_),
    .B(_151_),
    .C(_85_),
    .Y(_155_)
);

FILL FILL_1__1375_ (
);

FILL FILL_2__1444_ (
);

FILL FILL_2__1024_ (
);

FILL FILL89550x66450 (
);

FILL FILL_2__799_ (
);

FILL FILL_3__1513_ (
);

INVX1 _1442_ (
    .A(Yin[12]),
    .Y(_650_)
);

AOI21X1 _1022_ (
    .A(_195_),
    .B(_196_),
    .C(_139_),
    .Y(_212_)
);

FILL FILL_0__770_ (
);

FILL FILL_1__804_ (
);

AOI21X1 _773_ (
    .A(_515_),
    .B(_537_),
    .C(_429_),
    .Y(_569_)
);

FILL FILL_1__1184_ (
);

FILL FILL_2__1253_ (
);

FILL FILL_0__1499_ (
);

FILL FILL_0__1079_ (
);

FILL FILL_0__826_ (
);

FILL FILL_3__1322_ (
);

AOI21X1 _829_ (
    .A(_19_),
    .B(_14_),
    .C(_738_),
    .Y(_22_)
);

AND2X2 _1251_ (
    .A(Cin[2]),
    .B(Xin[7]),
    .Y(_445_)
);

FILL FILL_2__1309_ (
);

FILL FILL_2__820_ (
);

FILL FILL_2__1482_ (
);

FILL FILL_2__1062_ (
);

NOR2X1 _1307_ (
    .A(_417_),
    .B(_503_),
    .Y(_505_)
);

FILL FILL_3__779_ (
);

FILL FILL_3__1131_ (
);

FILL FILL_1__1469_ (
);

FILL FILL_1__1049_ (
);

NAND2X1 _1480_ (
    .A(_689_),
    .B(_690_),
    .Y(_691_)
);

AND2X2 _1060_ (
    .A(Cin[2]),
    .B(Xin_5_bF$buf1),
    .Y(_250_)
);

FILL FILL_1__842_ (
);

FILL FILL_4__986_ (
);

FILL FILL_2__1118_ (
);

FILL FILL_0__1100_ (
);

FILL FILL_2__1291_ (
);

DFFPOSX1 _1536_ (
    .D(y[8]),
    .CLK(clk_bF$buf1),
    .Q(_755_[8])
);

AOI21X1 _1116_ (
    .A(_297_),
    .B(_292_),
    .C(_215_),
    .Y(_306_)
);

FILL FILL_0__864_ (
);

FILL FILL_3__1360_ (
);

NAND3X1 _867_ (
    .A(_48_),
    .B(_50_),
    .C(_46_),
    .Y(_59_)
);

FILL FILL_1__1278_ (
);

FILL FILL_2__1347_ (
);

FILL FILL_3__800_ (
);

FILL FILL_3__1416_ (
);

NAND2X1 _1345_ (
    .A(_543_),
    .B(_545_),
    .Y(_546_)
);

FILL FILL_1__1087_ (
);

FILL FILL_1__880_ (
);

FILL FILL_2__914_ (
);

FILL FILL_2__1576_ (
);

FILL FILL_2__1156_ (
);

FILL FILL_3__1225_ (
);

BUFX2 _1574_ (
    .A(_755_[14]),
    .Y(Yout[14])
);

OAI21X1 _1154_ (
    .A(_335_),
    .B(_334_),
    .C(_332_),
    .Y(_343_)
);

FILL FILL_1__936_ (
);

FILL FILL89250x15750 (
);

FILL FILL_2__1385_ (
);

FILL FILL_0__958_ (
);

FILL FILL_3__1454_ (
);

FILL FILL_3__1034_ (
);

NAND3X1 _1383_ (
    .A(_583_),
    .B(_579_),
    .C(_585_),
    .Y(_586_)
);

FILL FILL_4__889_ (
);

FILL FILL_0__1423_ (
);

FILL FILL_0__1003_ (
);

FILL FILL_2__952_ (
);

FILL FILL_2__1194_ (
);

INVX1 _1439_ (
    .A(_646_),
    .Y(_647_)
);

AOI21X1 _1019_ (
    .A(_203_),
    .B(_207_),
    .C(_136_),
    .Y(_210_)
);

FILL FILL_0__767_ (
);

FILL FILL_3__1263_ (
);

FILL FILL88950x4050 (
);

AOI21X1 _1192_ (
    .A(_380_),
    .B(_374_),
    .C(_345_),
    .Y(_381_)
);

FILL FILL_1__974_ (
);

FILL FILL_4__1332_ (
);

FILL FILL_0__1232_ (
);

FILL FILL_2__761_ (
);

FILL FILL_3__1319_ (
);

OAI21X1 _1248_ (
    .A(_359_),
    .B(_441_),
    .C(_369_),
    .Y(_442_)
);

FILL FILL_0__996_ (
);

FILL FILL_3__1492_ (
);

FILL FILL_3__1072_ (
);

OAI21X1 _999_ (
    .A(_176_),
    .B(_179_),
    .C(_182_),
    .Y(_190_)
);

FILL FILL_1__783_ (
);

FILL FILL_2__817_ (
);

FILL FILL_2__1479_ (
);

FILL FILL_0__1461_ (
);

FILL FILL_0__1041_ (
);

FILL FILL_2__1059_ (
);

FILL FILL89550x54750 (
);

FILL FILL_2__990_ (
);

FILL FILL_3__932_ (
);

FILL FILL_1__1202_ (
);

FILL FILL_3__1128_ (
);

OAI21X1 _1477_ (
    .A(_686_),
    .B(_685_),
    .C(_646_),
    .Y(_688_)
);

NAND2X1 _1057_ (
    .A(Xin_3_bF$buf1),
    .B(Cin[4]),
    .Y(_247_)
);

FILL FILL_1__839_ (
);

FILL FILL_0__1517_ (
);

FILL FILL_2__1288_ (
);

FILL FILL_0__1270_ (
);

FILL FILL_1__1431_ (
);

FILL FILL_1__1011_ (
);

FILL FILL_3__1357_ (
);

NAND3X1 _1286_ (
    .A(_479_),
    .B(_480_),
    .C(_481_),
    .Y(_482_)
);

FILL FILL_2__1500_ (
);

FILL FILL_0__1326_ (
);

FILL FILL_2__855_ (
);

FILL FILL_2__1097_ (
);

FILL FILL_3__970_ (
);

FILL FILL_1__1240_ (
);

FILL FILL_3__1166_ (
);

AOI22X1 _1095_ (
    .A(_254_),
    .B(_257_),
    .C(_275_),
    .D(_271_),
    .Y(_285_)
);

FILL FILL_1__877_ (
);

FILL FILL_4__1235_ (
);

FILL FILL_0__1135_ (
);

FILL FILL_0__899_ (
);

FILL FILL_3__1395_ (
);

FILL FILL_0__1364_ (
);

FILL FILL_2__893_ (
);

FILL FILL_3__835_ (
);

FILL FILL_1__1105_ (
);

FILL FILL_2__949_ (
);

FILL FILL_0__1173_ (
);

FILL FILL_0__920_ (
);

NAND3X1 _923_ (
    .A(_112_),
    .B(_114_),
    .C(_113_),
    .Y(_115_)
);

FILL FILL_1__1334_ (
);

NAND3X1 _1189_ (
    .A(_369_),
    .B(_372_),
    .C(_377_),
    .Y(_378_)
);

FILL FILL_2__1403_ (
);

FILL FILL_0__1229_ (
);

FILL FILL_2__758_ (
);

AOI21X1 _1401_ (
    .A(_592_),
    .B(_587_),
    .C(_574_),
    .Y(_606_)
);

FILL FILL_3__873_ (
);

FILL FILL_4__907_ (
);

FILL FILL_1__1563_ (
);

FILL FILL_1__1143_ (
);

FILL FILL_3__1489_ (
);

FILL FILL_3__1069_ (
);

FILL FILL_2__1212_ (
);

FILL FILL_4__1138_ (
);

FILL FILL_0__1458_ (
);

FILL FILL_0__1038_ (
);

FILL FILL_2__987_ (
);

FILL FILL_3__929_ (
);

NAND3X1 _1210_ (
    .A(_314_),
    .B(_394_),
    .C(_395_),
    .Y(_401_)
);

NAND2X1 _961_ (
    .A(Xin_3_bF$buf2),
    .B(Cin[3]),
    .Y(_152_)
);

FILL FILL_1__1372_ (
);

FILL FILL_3__1298_ (
);

FILL FILL_2__1441_ (
);

FILL FILL_2__1021_ (
);

FILL FILL_0__1267_ (
);

FILL FILL_2__796_ (
);

FILL FILL_3__1510_ (
);

FILL FILL_1__1428_ (
);

FILL FILL_1__1008_ (
);

FILL FILL_1__801_ (
);

OAI21X1 _770_ (
    .A(_493_),
    .B(_526_),
    .C(_461_),
    .Y(_537_)
);

FILL FILL_1__1181_ (
);

FILL FILL_2__1250_ (
);

FILL FILL_0__1496_ (
);

FILL FILL_0__1076_ (
);

FILL FILL_0__823_ (
);

FILL FILL_3__967_ (
);

FILL FILL_1_BUFX2_insert6 (
);

FILL FILL_1_BUFX2_insert7 (
);

FILL FILL_1_BUFX2_insert8 (
);

FILL FILL_1_BUFX2_insert9 (
);

OAI21X1 _826_ (
    .A(_18_),
    .B(_17_),
    .C(_16_),
    .Y(_19_)
);

FILL FILL_1__1237_ (
);

FILL FILL_2__1306_ (
);

OAI21X1 _1304_ (
    .A(_415_),
    .B(_416_),
    .C(_424_),
    .Y(_501_)
);

FILL FILL_3__776_ (
);

FILL FILL_1__1466_ (
);

FILL FILL_1__1046_ (
);

FILL FILL_2__1115_ (
);

DFFPOSX1 _1533_ (
    .D(y[5]),
    .CLK(clk_bF$buf3),
    .Q(_755_[5])
);

INVX1 _1113_ (
    .A(_200_),
    .Y(_303_)
);

FILL FILL_0__861_ (
);

NAND3X1 _864_ (
    .A(_38_),
    .B(_55_),
    .C(_43_),
    .Y(_56_)
);

FILL FILL_1__1275_ (
);

FILL FILL_4__792_ (
);

FILL FILL_2__1344_ (
);

FILL FILL_0__917_ (
);

FILL FILL_3__1413_ (
);

NAND2X1 _1342_ (
    .A(_539_),
    .B(_530_),
    .Y(_543_)
);

FILL FILL_4__848_ (
);

FILL FILL_1__1084_ (
);

FILL FILL_2__911_ (
);

FILL FILL_2__1573_ (
);

FILL FILL_2__1153_ (
);

FILL FILL_0__1399_ (
);

FILL FILL_3__1222_ (
);

FILL FILL_3_BUFX2_insert6 (
);

FILL FILL_3_BUFX2_insert7 (
);

FILL FILL_3_BUFX2_insert8 (
);

FILL FILL_3_BUFX2_insert9 (
);

BUFX2 _1571_ (
    .A(_755_[11]),
    .Y(Yout[11])
);

NAND3X1 _1151_ (
    .A(_318_),
    .B(_333_),
    .C(_339_),
    .Y(_340_)
);

FILL FILL_1__933_ (
);

FILL FILL_2__1209_ (
);

FILL FILL89550x19650 (
);

FILL FILL_2__1382_ (
);

OAI21X1 _1207_ (
    .A(_396_),
    .B(_393_),
    .C(_313_),
    .Y(_398_)
);

FILL FILL_0__955_ (
);

FILL FILL_3__1451_ (
);

FILL FILL_3__1031_ (
);

AND2X2 _958_ (
    .A(Cin[2]),
    .B(Xin[4]),
    .Y(_149_)
);

FILL FILL_1__1369_ (
);

INVX1 _1380_ (
    .A(_582_),
    .Y(_583_)
);

FILL FILL_2__1438_ (
);

FILL FILL_0__1420_ (
);

FILL FILL_0__1000_ (
);

FILL FILL_2__1018_ (
);

FILL FILL_2__1191_ (
);

FILL FILL_3__1507_ (
);

NAND2X1 _1436_ (
    .A(Xin_5_bF$buf3),
    .B(Cin[7]),
    .Y(_643_)
);

NAND3X1 _1016_ (
    .A(_204_),
    .B(_205_),
    .C(_206_),
    .Y(_207_)
);

FILL FILL_0__764_ (
);

FILL FILL_3__1260_ (
);

INVX1 _767_ (
    .A(_493_),
    .Y(_504_)
);

FILL FILL_1__1178_ (
);

FILL FILL_1__971_ (
);

FILL FILL_2__1247_ (
);

FILL FILL_3__1316_ (
);

NAND3X1 _1245_ (
    .A(_435_),
    .B(_436_),
    .C(_437_),
    .Y(_438_)
);

FILL FILL_0__993_ (
);

AOI21X1 _996_ (
    .A(_186_),
    .B(_180_),
    .C(_144_),
    .Y(_187_)
);

FILL FILL_1__780_ (
);

FILL FILL_2__814_ (
);

FILL FILL_2__1476_ (
);

FILL FILL_2__1056_ (
);

FILL FILL_3__1125_ (
);

NAND3X1 _1474_ (
    .A(_652_),
    .B(_657_),
    .C(_683_),
    .Y(_684_)
);

AND2X2 _1054_ (
    .A(_240_),
    .B(_243_),
    .Y(_244_)
);

FILL FILL_1__836_ (
);

FILL FILL_0__1514_ (
);

FILL FILL_2__1285_ (
);

FILL FILL_0__858_ (
);

FILL FILL_3__1354_ (
);

INVX1 _1283_ (
    .A(_410_),
    .Y(_479_)
);

FILL FILL_0__1323_ (
);

FILL FILL_2__852_ (
);

FILL FILL_2__1094_ (
);

XOR2X1 _1339_ (
    .A(_530_),
    .B(_539_),
    .Y(_540_)
);

FILL FILL_3__1583_ (
);

FILL FILL_3__1163_ (
);

INVX1 _1092_ (
    .A(_177_),
    .Y(_282_)
);

FILL FILL_1__874_ (
);

FILL FILL_2__908_ (
);

FILL FILL_0__1132_ (
);

FILL FILL_3__1219_ (
);

BUFX2 _1568_ (
    .A(_755_[0]),
    .Y(Yout[0])
);

INVX1 _1148_ (
    .A(_336_),
    .Y(_337_)
);

FILL FILL_0__896_ (
);

FILL FILL_3__1392_ (
);

NAND2X1 _899_ (
    .A(Cin[2]),
    .B(Xin_3_bF$buf2),
    .Y(_91_)
);

FILL FILL_4__1041_ (
);

FILL FILL_2__1379_ (
);

FILL FILL_0__1361_ (
);

FILL FILL_2__890_ (
);

FILL FILL_3__832_ (
);

FILL FILL_1__1102_ (
);

FILL FILL_3__1448_ (
);

FILL FILL_3__1028_ (
);

OAI21X1 _1377_ (
    .A(_503_),
    .B(_576_),
    .C(_579_),
    .Y(_580_)
);

FILL FILL_0__1417_ (
);

FILL FILL_2__946_ (
);

FILL FILL_0__1170_ (
);

FILL FILL_2__1188_ (
);

NAND2X1 _920_ (
    .A(_93_),
    .B(_89_),
    .Y(_112_)
);

FILL FILL_1__1331_ (
);

FILL FILL_3__1257_ (
);

INVX1 _1186_ (
    .A(_271_),
    .Y(_375_)
);

FILL FILL_1__968_ (
);

FILL FILL_2__1400_ (
);

FILL FILL_0__1226_ (
);

FILL FILL_3__870_ (
);

FILL FILL_1__1560_ (
);

FILL FILL_1__1140_ (
);

FILL FILL_3__1486_ (
);

FILL FILL_3__1066_ (
);

FILL FILL_1__777_ (
);

FILL FILL_0__1455_ (
);

FILL FILL_0__1035_ (
);

FILL FILL_2__984_ (
);

FILL FILL_3__926_ (
);

FILL FILL_0__799_ (
);

FILL FILL_3__1295_ (
);

FILL FILL_4__1364_ (
);

FILL FILL_0__1264_ (
);

FILL FILL_2__793_ (
);

FILL FILL_1__1425_ (
);

FILL FILL_1__1005_ (
);

FILL FILL_2__849_ (
);

FILL FILL_0__1493_ (
);

FILL FILL_0__1073_ (
);

FILL FILL_0__820_ (
);

FILL FILL_3__964_ (
);

OAI21X1 _823_ (
    .A(_15_),
    .B(_732_),
    .C(_742_),
    .Y(_16_)
);

FILL FILL_1__1234_ (
);

NAND3X1 _1089_ (
    .A(_267_),
    .B(_270_),
    .C(_272_),
    .Y(_279_)
);

FILL FILL_2__1303_ (
);

FILL FILL_0__1129_ (
);

NAND2X1 _1301_ (
    .A(_428_),
    .B(_434_),
    .Y(_498_)
);

FILL FILL_3__773_ (
);

FILL FILL_1__1463_ (
);

FILL FILL_1__1043_ (
);

FILL FILL_3__1389_ (
);

FILL FILL_2__1112_ (
);

FILL FILL_0__1358_ (
);

FILL FILL_2__887_ (
);

FILL FILL_3__829_ (
);

FILL FILL_1__1519_ (
);

DFFPOSX1 _1530_ (
    .D(y[2]),
    .CLK(clk_bF$buf1),
    .Q(_755_[2])
);

NAND3X1 _1110_ (
    .A(_287_),
    .B(_291_),
    .C(_294_),
    .Y(_300_)
);

OAI21X1 _861_ (
    .A(_47_),
    .B(_590_),
    .C(_743_),
    .Y(_53_)
);

FILL FILL_1__1272_ (
);

FILL FILL_3__1198_ (
);

FILL FILL_2__1341_ (
);

FILL FILL_4__1267_ (
);

FILL FILL_0__1167_ (
);

FILL FILL_0__914_ (
);

FILL FILL_3__1410_ (
);

AOI21X1 _917_ (
    .A(_101_),
    .B(_98_),
    .C(_97_),
    .Y(_109_)
);

FILL FILL_1__1328_ (
);

FILL FILL_1__1081_ (
);

FILL FILL_2__1570_ (
);

FILL FILL_2__1150_ (
);

FILL FILL_0__1396_ (
);

FILL FILL_3__867_ (
);

FILL FILL_1__1137_ (
);

FILL FILL_1__930_ (
);

FILL FILL_2__1206_ (
);

NAND3X1 _1204_ (
    .A(_391_),
    .B(_317_),
    .C(_390_),
    .Y(_394_)
);

FILL FILL_0__952_ (
);

OAI21X1 _955_ (
    .A(_112_),
    .B(_145_),
    .C(_106_),
    .Y(_146_)
);

FILL FILL_1__1366_ (
);

FILL FILL_2__1435_ (
);

FILL FILL_2__1015_ (
);

FILL FILL_3__1504_ (
);

OAI21X1 _1433_ (
    .A(_77_),
    .B(_447_),
    .C(_576_),
    .Y(_640_)
);

INVX1 _1013_ (
    .A(_127_),
    .Y(_204_)
);

FILL FILL_0__761_ (
);

INVX1 _764_ (
    .A(_461_),
    .Y(_472_)
);

FILL FILL_1__1175_ (
);

FILL FILL_2__1244_ (
);

FILL FILL_0__817_ (
);

FILL FILL_3__1313_ (
);

AND2X2 _1242_ (
    .A(_327_),
    .B(_323_),
    .Y(_435_)
);

FILL FILL_0__990_ (
);

NAND3X1 _993_ (
    .A(_177_),
    .B(_178_),
    .C(_183_),
    .Y(_184_)
);

FILL FILL_2__811_ (
);

FILL FILL_2__1473_ (
);

FILL FILL_2__1053_ (
);

FILL FILL_0__1299_ (
);

FILL FILL_3__1122_ (
);

AND2X2 _1471_ (
    .A(_679_),
    .B(_680_),
    .Y(_681_)
);

NAND3X1 _1051_ (
    .A(_226_),
    .B(_230_),
    .C(_238_),
    .Y(_241_)
);

FILL FILL_1__833_ (
);

FILL FILL_0__1511_ (
);

FILL FILL_2__1109_ (
);

FILL FILL_2__1282_ (
);

DFFPOSX1 _1527_ (
    .D(Xin[7]),
    .CLK(clk_bF$buf2),
    .Q(_754_[7])
);

OAI21X1 _1107_ (
    .A(_295_),
    .B(_296_),
    .C(_294_),
    .Y(_297_)
);

FILL FILL_0__855_ (
);

FILL FILL_3__999_ (
);

FILL FILL_3__1351_ (
);

INVX1 _858_ (
    .A(_44_),
    .Y(_50_)
);

FILL FILL_1__1269_ (
);

AOI22X1 _1280_ (
    .A(_434_),
    .B(_438_),
    .C(_463_),
    .D(_458_),
    .Y(_476_)
);

FILL FILL_4__1000_ (
);

FILL FILL_0__1320_ (
);

FILL FILL_2__1338_ (
);

FILL FILL_2__1091_ (
);

FILL FILL_3__1407_ (
);

AND2X2 _1336_ (
    .A(_350_),
    .B(_532_),
    .Y(_536_)
);

FILL FILL_3__1580_ (
);

FILL FILL_3__1160_ (
);

FILL FILL_1__1498_ (
);

FILL FILL_1__1078_ (
);

FILL FILL_1__871_ (
);

FILL FILL_2__905_ (
);

FILL FILL_2__1567_ (
);

FILL FILL_2__1147_ (
);

FILL FILL_3__1216_ (
);

FILL FILL88050x35250 (
);

BUFX2 _1565_ (
    .A(_754_[5]),
    .Y(Xout[5])
);

AOI21X1 _1145_ (
    .A(_328_),
    .B(_329_),
    .C(_319_),
    .Y(_334_)
);

FILL FILL_0__893_ (
);

FILL FILL_1__927_ (
);

OAI21X1 _896_ (
    .A(_590_),
    .B(_87_),
    .C(_79_),
    .Y(_88_)
);

FILL FILL_2__1376_ (
);

FILL FILL_0__949_ (
);

FILL FILL_3__1445_ (
);

FILL FILL_3__1025_ (
);

INVX1 _1374_ (
    .A(Xin_5_bF$buf3),
    .Y(_577_)
);

FILL FILL_0__1414_ (
);

FILL FILL_2__943_ (
);

FILL FILL_2__1185_ (
);

FILL FILL_0__758_ (
);

FILL FILL_3__1254_ (
);

NAND3X1 _1183_ (
    .A(_263_),
    .B(_267_),
    .C(_371_),
    .Y(_372_)
);

FILL FILL_1__965_ (
);

FILL FILL_0__1223_ (
);

AOI22X1 _1239_ (
    .A(_250_),
    .B(_350_),
    .C(_353_),
    .D(_349_),
    .Y(_432_)
);

FILL FILL88350x74250 (
);

FILL FILL_0__987_ (
);

FILL FILL_3__1483_ (
);

FILL FILL_3__1063_ (
);

FILL FILL_1__774_ (
);

FILL FILL_2__808_ (
);

FILL FILL_0__1452_ (
);

FILL FILL_0__1032_ (
);

FILL FILL_2__981_ (
);

FILL FILL_3__923_ (
);

FILL FILL_3__1119_ (
);

NOR2X1 _1468_ (
    .A(_447_),
    .B(_575_),
    .Y(_678_)
);

AOI21X1 _1048_ (
    .A(_148_),
    .B(_153_),
    .C(_237_),
    .Y(_238_)
);

FILL FILL_0__796_ (
);

FILL FILL_3__1292_ (
);

INVX2 _799_ (
    .A(Cin[3]),
    .Y(_740_)
);

FILL FILL_0__1508_ (
);

FILL FILL_0__1261_ (
);

FILL FILL_2__1279_ (
);

FILL FILL_2__790_ (
);

FILL FILL_1__1422_ (
);

FILL FILL_1__1002_ (
);

FILL FILL_3__1348_ (
);

NAND2X1 _1277_ (
    .A(_442_),
    .B(_462_),
    .Y(_473_)
);

FILL FILL_0__1317_ (
);

FILL FILL_2__846_ (
);

FILL FILL_4__1170_ (
);

FILL FILL_0__1490_ (
);

FILL FILL_0__1070_ (
);

FILL FILL_2__1088_ (
);

FILL FILL_3__961_ (
);

OAI21X1 _820_ (
    .A(_12_),
    .B(_11_),
    .C(_10_),
    .Y(_13_)
);

FILL FILL_1__1231_ (
);

FILL FILL_3__1577_ (
);

FILL FILL_3__1157_ (
);

NAND3X1 _1086_ (
    .A(_271_),
    .B(_275_),
    .C(_258_),
    .Y(_276_)
);

FILL FILL_1__868_ (
);

FILL FILL_2__1300_ (
);

FILL FILL_4__1226_ (
);

FILL FILL_0__1126_ (
);

FILL FILL_3__770_ (
);

FILL FILL_1__1460_ (
);

FILL FILL_1__1040_ (
);

FILL FILL_3__1386_ (
);

FILL FILL_0__1355_ (
);

FILL FILL_2__884_ (
);

FILL FILL_3__826_ (
);

FILL FILL_1__1516_ (
);

FILL FILL_3__1195_ (
);

FILL FILL_0__1164_ (
);

FILL FILL_0__911_ (
);

NAND3X1 _914_ (
    .A(_95_),
    .B(_102_),
    .C(_105_),
    .Y(_106_)
);

FILL FILL_1__1325_ (
);

FILL FILL_4__1493_ (
);

FILL FILL_0__1393_ (
);

FILL FILL_3__864_ (
);

FILL FILL_1__1134_ (
);

FILL FILL88950x7950 (
);

FILL FILL_2__1203_ (
);

FILL FILL_4__1129_ (
);

FILL FILL_0__1449_ (
);

FILL FILL_0__1029_ (
);

FILL FILL_2__978_ (
);

NAND3X1 _1201_ (
    .A(_345_),
    .B(_374_),
    .C(_380_),
    .Y(_391_)
);

OAI21X1 _952_ (
    .A(_79_),
    .B(_91_),
    .C(_89_),
    .Y(_143_)
);

FILL FILL_1__1363_ (
);

FILL FILL_3__1289_ (
);

FILL FILL88350x4050 (
);

FILL FILL_4__880_ (
);

FILL FILL_2__1432_ (
);

FILL FILL_2__1012_ (
);

FILL FILL_0__1258_ (
);

FILL FILL_2__787_ (
);

FILL FILL_3__1501_ (
);

FILL FILL_1__1419_ (
);

AND2X2 _1430_ (
    .A(_604_),
    .B(_600_),
    .Y(_637_)
);

OAI21X1 _1010_ (
    .A(_187_),
    .B(_191_),
    .C(_194_),
    .Y(_201_)
);

NOR2X1 _761_ (
    .A(Yin[0]),
    .B(_407_),
    .Y(_440_)
);

FILL FILL_1__1172_ (
);

FILL FILL_3__1098_ (
);

FILL FILL_2__1241_ (
);

FILL FILL_0__1487_ (
);

FILL FILL_0__1067_ (
);

FILL FILL_0__814_ (
);

FILL FILL_3__958_ (
);

FILL FILL_3__1310_ (
);

INVX1 _817_ (
    .A(_746_),
    .Y(_10_)
);

FILL FILL_1__1228_ (
);

INVX1 _990_ (
    .A(_106_),
    .Y(_181_)
);

FILL FILL_2__1470_ (
);

FILL FILL_2__1050_ (
);

FILL FILL_4__1396_ (
);

FILL FILL_0__1296_ (
);

FILL FILL_3__767_ (
);

FILL FILL_1__1457_ (
);

FILL FILL_1__1037_ (
);

FILL FILL_1__830_ (
);

FILL FILL_2__1106_ (
);

DFFPOSX1 _1524_ (
    .D(Xin[4]),
    .CLK(clk_bF$buf1),
    .Q(_754_[4])
);

AOI21X1 _1104_ (
    .A(_188_),
    .B(_190_),
    .C(_293_),
    .Y(_294_)
);

FILL FILL_0__852_ (
);

FILL FILL_3__996_ (
);

INVX2 _855_ (
    .A(Xin[2]),
    .Y(_47_)
);

FILL FILL_1__1266_ (
);

FILL FILL_4__783_ (
);

FILL FILL_2__1335_ (
);

FILL FILL_0__908_ (
);

FILL FILL_3__1404_ (
);

AOI21X1 _1333_ (
    .A(_350_),
    .B(_532_),
    .C(_531_),
    .Y(_533_)
);

FILL FILL_1__1495_ (
);

FILL FILL_1__1075_ (
);

FILL FILL_2__902_ (
);

FILL FILL_2__1564_ (
);

FILL FILL_2__1144_ (
);

FILL FILL_3__1213_ (
);

BUFX2 _1562_ (
    .A(_754_[2]),
    .Y(Xout[2])
);

AOI22X1 _1142_ (
    .A(Cin[2]),
    .B(Xin_5_bF$buf2),
    .C(Cin[3]),
    .D(Xin[4]),
    .Y(_331_)
);

FILL FILL_0__890_ (
);

FILL FILL_1__924_ (
);

AND2X2 _893_ (
    .A(Xin_3_bF$buf1),
    .B(Cin[3]),
    .Y(_85_)
);

FILL FILL_2__1373_ (
);

FILL FILL_4__1299_ (
);

FILL FILL_0__1199_ (
);

FILL FILL_0__946_ (
);

FILL FILL_3__1442_ (
);

FILL FILL_3__1022_ (
);

AND2X2 _949_ (
    .A(Xin[1]),
    .B(Cin[6]),
    .Y(_140_)
);

OAI21X1 _1371_ (
    .A(_502_),
    .B(_506_),
    .C(_510_),
    .Y(_574_)
);

FILL FILL_4__1511_ (
);

FILL FILL_0__1411_ (
);

FILL FILL_2__1429_ (
);

FILL FILL_2__1009_ (
);

FILL FILL_2__940_ (
);

FILL FILL_2__1182_ (
);

NAND3X1 _1427_ (
    .A(_630_),
    .B(_632_),
    .C(_628_),
    .Y(_634_)
);

AOI21X1 _1007_ (
    .A(_197_),
    .B(_192_),
    .C(_137_),
    .Y(_198_)
);

FILL FILL_3__899_ (
);

FILL FILL_3__1251_ (
);

NOR2X1 _758_ (
    .A(_386_),
    .B(_397_),
    .Y(_407_)
);

FILL FILL_1__1169_ (
);

NAND2X1 _1180_ (
    .A(_361_),
    .B(_366_),
    .Y(_369_)
);

FILL FILL_1__962_ (
);

FILL FILL_0__1220_ (
);

FILL FILL_2__1238_ (
);

FILL FILL_3__1307_ (
);

FILL FILL88650x78150 (
);

NAND3X1 _1236_ (
    .A(_425_),
    .B(_420_),
    .C(_427_),
    .Y(_428_)
);

FILL FILL_0__984_ (
);

FILL FILL_3__1480_ (
);

FILL FILL_3__1060_ (
);

OAI21X1 _987_ (
    .A(_170_),
    .B(_166_),
    .C(_172_),
    .Y(_178_)
);

FILL FILL_1__1398_ (
);

FILL FILL_1__771_ (
);

FILL FILL_2__805_ (
);

FILL FILL_2__1467_ (
);

FILL FILL_2__1047_ (
);

FILL FILL_3__920_ (
);

FILL FILL_3_CLKBUF1_insert0 (
);

FILL FILL_3_CLKBUF1_insert1 (
);

FILL FILL_3_CLKBUF1_insert2 (
);

FILL FILL_3_CLKBUF1_insert3 (
);

FILL FILL_3__1116_ (
);

FILL FILL_3_CLKBUF1_insert4 (
);

FILL FILL_3_CLKBUF1_insert5 (
);

AOI21X1 _1465_ (
    .A(_635_),
    .B(_660_),
    .C(_662_),
    .Y(_674_)
);

AOI21X1 _1045_ (
    .A(_228_),
    .B(_229_),
    .C(_220_),
    .Y(_235_)
);

FILL FILL_0__793_ (
);

FILL FILL_1__827_ (
);

NOR2X1 _796_ (
    .A(_737_),
    .B(_736_),
    .Y(_750_[2])
);

FILL FILL_0__1505_ (
);

FILL FILL_2__1276_ (
);

FILL FILL_0__849_ (
);

FILL FILL_3__1345_ (
);

NAND3X1 _1274_ (
    .A(_412_),
    .B(_464_),
    .C(_468_),
    .Y(_469_)
);

FILL FILL_4__1414_ (
);

FILL FILL_0__1314_ (
);

FILL FILL_2__843_ (
);

FILL FILL_2__1085_ (
);

FILL FILL_3__1574_ (
);

FILL FILL_3__1154_ (
);

AOI21X1 _1083_ (
    .A(_269_),
    .B(_268_),
    .C(_261_),
    .Y(_273_)
);

FILL FILL_1__865_ (
);

FILL FILL88950x31350 (
);

FILL FILL_0__1123_ (
);

FILL FILL_4__801_ (
);

DFFPOSX1 _1559_ (
    .D(_753_[15]),
    .CLK(clk_bF$buf2),
    .Q(y[15])
);

OAI21X1 _1139_ (
    .A(_87_),
    .B(_77_),
    .C(_321_),
    .Y(_328_)
);

FILL FILL_0__887_ (
);

FILL FILL_3__1383_ (
);

FILL FILL_4__1032_ (
);

FILL FILL_0__1352_ (
);

FILL FILL_2__881_ (
);

FILL FILL_3__823_ (
);

FILL FILL_1__1513_ (
);

FILL FILL_3__1439_ (
);

FILL FILL_3__1019_ (
);

INVX1 _1368_ (
    .A(_570_),
    .Y(_571_)
);

FILL FILL_3__1192_ (
);

FILL FILL_0__1408_ (
);

FILL FILL_2__937_ (
);

FILL FILL_0__1581_ (
);

FILL FILL_2__1179_ (
);

FILL FILL_0__1161_ (
);

NAND2X1 _911_ (
    .A(Yin[5]),
    .B(_100_),
    .Y(_103_)
);

FILL FILL_1__1322_ (
);

FILL FILL_3__1248_ (
);

NOR2X1 _1177_ (
    .A(_364_),
    .B(_363_),
    .Y(_366_)
);

FILL FILL_1__959_ (
);

FILL FILL_0__1217_ (
);

FILL FILL_0__1390_ (
);

FILL FILL_3__861_ (
);

FILL FILL_1__1131_ (
);

FILL FILL_3__1477_ (
);

FILL FILL_3__1057_ (
);

FILL FILL_1__768_ (
);

FILL FILL_2__1200_ (
);

FILL FILL_0__1446_ (
);

FILL FILL_0__1026_ (
);

FILL FILL_2__975_ (
);

FILL FILL_3__917_ (
);

FILL FILL_1__1360_ (
);

FILL FILL_3__1286_ (
);

FILL FILL_1__997_ (
);

FILL FILL_4__1355_ (
);

FILL FILL_0__1255_ (
);

FILL FILL_2__784_ (
);

FILL FILL_1__1416_ (
);

FILL FILL_3__1095_ (
);

FILL FILL_0__1484_ (
);

FILL FILL_0__1064_ (
);

FILL FILL_0__811_ (
);

FILL FILL_3__955_ (
);

NAND3X1 _814_ (
    .A(Cin_0_bF$buf1),
    .B(Xin_3_bF$buf0),
    .C(_2_),
    .Y(_7_)
);

FILL FILL_1__1225_ (
);

FILL FILL_0__1293_ (
);

FILL FILL_3__764_ (
);

FILL FILL_1__1454_ (
);

FILL FILL_1__1034_ (
);

FILL FILL_2__1103_ (
);

FILL FILL_0__1349_ (
);

FILL FILL_2__878_ (
);

DFFPOSX1 _1521_ (
    .D(Xin[1]),
    .CLK(clk_bF$buf1),
    .Q(_754_[1])
);

NAND3X1 _1101_ (
    .A(_288_),
    .B(_289_),
    .C(_290_),
    .Y(_291_)
);

FILL FILL_3__993_ (
);

NAND2X1 _852_ (
    .A(Xin[0]),
    .B(Cin[4]),
    .Y(_44_)
);

FILL FILL_1__1263_ (
);

FILL FILL_3__1189_ (
);

FILL FILL_2__1332_ (
);

FILL FILL_4__1258_ (
);

FILL FILL_0__1578_ (
);

FILL FILL_0__1158_ (
);

FILL FILL_0__905_ (
);

FILL FILL_3__1401_ (
);

NAND2X1 _908_ (
    .A(Cin_0_bF$buf3),
    .B(Xin_5_bF$buf0),
    .Y(_100_)
);

FILL FILL_1__1319_ (
);

NAND2X1 _1330_ (
    .A(_529_),
    .B(_454_),
    .Y(_530_)
);

FILL FILL_1__1492_ (
);

FILL FILL_1__1072_ (
);

FILL FILL_2__1561_ (
);

FILL FILL_2__1141_ (
);

FILL FILL_0__1387_ (
);

FILL FILL_3__858_ (
);

FILL FILL_3__1210_ (
);

FILL FILL_1__1128_ (
);

FILL FILL_1__921_ (
);

OAI21X1 _890_ (
    .A(_61_),
    .B(_58_),
    .C(_38_),
    .Y(_82_)
);

FILL FILL_2__1370_ (
);

FILL FILL_0__1196_ (
);

FILL FILL88350x15750 (
);

FILL FILL_0__943_ (
);

NAND2X1 _946_ (
    .A(_78_),
    .B(_80_),
    .Y(_137_)
);

FILL FILL_1__1357_ (
);

FILL FILL_2__1426_ (
);

FILL FILL_2__1006_ (
);

NAND3X1 _1424_ (
    .A(_626_),
    .B(_629_),
    .C(_492_),
    .Y(_630_)
);

NAND3X1 _1004_ (
    .A(_188_),
    .B(_189_),
    .C(_190_),
    .Y(_195_)
);

FILL FILL_3__896_ (
);

FILL FILL_1__1166_ (
);

FILL FILL_2__1235_ (
);

FILL FILL_0__808_ (
);

FILL FILL_3__1304_ (
);

NAND3X1 _1233_ (
    .A(_421_),
    .B(_422_),
    .C(_424_),
    .Y(_425_)
);

FILL FILL_0__981_ (
);

NAND3X1 _984_ (
    .A(_173_),
    .B(_174_),
    .C(_172_),
    .Y(_175_)
);

FILL FILL_1__1395_ (
);

FILL FILL_2__802_ (
);

FILL FILL_2__1464_ (
);

FILL FILL_2__1044_ (
);

FILL FILL88650x54750 (
);

FILL FILL_3__1113_ (
);

XNOR2X1 _1462_ (
    .A(_634_),
    .B(_671_),
    .Y(_753_[12])
);

AND2X2 _1042_ (
    .A(_152_),
    .B(_231_),
    .Y(_232_)
);

FILL FILL_0__790_ (
);

FILL FILL_1__824_ (
);

NAND3X1 _793_ (
    .A(_559_),
    .B(_734_),
    .C(_731_),
    .Y(_735_)
);

FILL FILL_0__1502_ (
);

FILL FILL_2__1273_ (
);

FILL FILL_0__1099_ (
);

OAI21X1 _1518_ (
    .A(_739_),
    .B(_20_),
    .C(_24_),
    .Y(_730_)
);

FILL FILL_0__846_ (
);

FILL FILL_3__1342_ (
);

OAI21X1 _849_ (
    .A(_31_),
    .B(_36_),
    .C(_34_),
    .Y(_41_)
);

NOR2X1 _1271_ (
    .A(_460_),
    .B(_462_),
    .Y(_466_)
);

FILL FILL_0__1311_ (
);

FILL FILL_2__1329_ (
);

FILL FILL_2__840_ (
);

FILL FILL_2__1082_ (
);

NAND3X1 _1327_ (
    .A(_523_),
    .B(_524_),
    .C(_525_),
    .Y(_527_)
);

FILL FILL_3__799_ (
);

FILL FILL_3__1571_ (
);

FILL FILL_3__1151_ (
);

FILL FILL_1__1489_ (
);

FILL FILL_1__1069_ (
);

NAND3X1 _1080_ (
    .A(_261_),
    .B(_268_),
    .C(_269_),
    .Y(_270_)
);

FILL FILL_1__862_ (
);

FILL FILL_0__1120_ (
);

FILL FILL_2__1138_ (
);

FILL FILL_3__1207_ (
);

DFFPOSX1 _1556_ (
    .D(_753_[12]),
    .CLK(clk_bF$buf2),
    .Q(y[12])
);

NAND2X1 _1136_ (
    .A(Xin_3_bF$buf3),
    .B(Cin[5]),
    .Y(_325_)
);

FILL FILL_0__884_ (
);

FILL FILL_1__918_ (
);

FILL FILL_3__1380_ (
);

NAND2X1 _887_ (
    .A(Xin[2]),
    .B(Cin[3]),
    .Y(_79_)
);

FILL FILL_1__1298_ (
);

FILL FILL_2__1367_ (
);

FILL FILL_3__820_ (
);

FILL FILL_1__1510_ (
);

FILL FILL_3__1436_ (
);

FILL FILL_3__1016_ (
);

INVX1 _1365_ (
    .A(_555_),
    .Y(_567_)
);

FILL FILL_0__1405_ (
);

FILL FILL_2__934_ (
);

FILL FILL_2__1176_ (
);

FILL FILL_3__1245_ (
);

INVX1 _1174_ (
    .A(_362_),
    .Y(_363_)
);

FILL FILL_1__956_ (
);

FILL FILL_0__1214_ (
);

FILL FILL_0__978_ (
);

FILL FILL_3__1474_ (
);

FILL FILL_3__1054_ (
);

FILL FILL_1__765_ (
);

FILL FILL_0__1443_ (
);

FILL FILL_0__1023_ (
);

FILL FILL_2__972_ (
);

FILL FILL_3__914_ (
);

OAI21X1 _1459_ (
    .A(_611_),
    .B(_608_),
    .C(_621_),
    .Y(_669_)
);

NAND2X1 _1039_ (
    .A(_224_),
    .B(_222_),
    .Y(_229_)
);

FILL FILL_0__787_ (
);

FILL FILL_3__1283_ (
);

FILL FILL_1__994_ (
);

FILL FILL_0__1252_ (
);

FILL FILL_2__781_ (
);

FILL FILL_1__1413_ (
);

FILL FILL_3__1339_ (
);

FILL FILL_4__930_ (
);

NAND2X1 _1268_ (
    .A(_460_),
    .B(_462_),
    .Y(_463_)
);

FILL FILL_3__1092_ (
);

FILL FILL_0__1308_ (
);

FILL FILL_2__837_ (
);

FILL FILL_4__1161_ (
);

FILL FILL_2__1499_ (
);

FILL FILL_0__1481_ (
);

FILL FILL_0__1061_ (
);

FILL FILL_2__1079_ (
);

FILL FILL_3__952_ (
);

NAND2X1 _811_ (
    .A(_2_),
    .B(_3_),
    .Y(_4_)
);

FILL FILL_1__1222_ (
);

FILL FILL_3__1568_ (
);

FILL FILL_3__1148_ (
);

NAND2X1 _1497_ (
    .A(_675_),
    .B(_681_),
    .Y(_709_)
);

NAND3X1 _1077_ (
    .A(_263_),
    .B(_262_),
    .C(_266_),
    .Y(_267_)
);

FILL FILL_1__859_ (
);

FILL FILL_0__1117_ (
);

FILL FILL_0__1290_ (
);

FILL FILL_3__761_ (
);

FILL FILL_1__1451_ (
);

FILL FILL_1__1031_ (
);

FILL FILL_3__1377_ (
);

FILL FILL_2__1100_ (
);

FILL FILL_0__1346_ (
);

FILL FILL_2__875_ (
);

FILL FILL_3__817_ (
);

FILL FILL_1__1507_ (
);

FILL FILL_3__990_ (
);

FILL FILL_1__1260_ (
);

FILL FILL_3__1186_ (
);

FILL FILL_1__897_ (
);

FILL FILL_0__1575_ (
);

FILL FILL_0__1155_ (
);

FILL FILL_0__902_ (
);

INVX1 _905_ (
    .A(_96_),
    .Y(_97_)
);

FILL FILL_1__1316_ (
);

FILL FILL_4__1484_ (
);

FILL FILL_4__1064_ (
);

FILL FILL_0__1384_ (
);

FILL FILL_3__855_ (
);

FILL FILL_1__1125_ (
);

FILL FILL_2__969_ (
);

FILL FILL_0__1193_ (
);

FILL FILL88650x19650 (
);

FILL FILL_0__940_ (
);

NAND2X1 _943_ (
    .A(_132_),
    .B(_134_),
    .Y(_135_)
);

FILL FILL_1__1354_ (
);

FILL FILL_4__871_ (
);

FILL FILL_2__1423_ (
);

FILL FILL_2__1003_ (
);

FILL FILL_0__1249_ (
);

FILL FILL_2__778_ (
);

NOR2X1 _1421_ (
    .A(_625_),
    .B(_565_),
    .Y(_627_)
);

OAI21X1 _1001_ (
    .A(_191_),
    .B(_187_),
    .C(_139_),
    .Y(_192_)
);

FILL FILL_3__893_ (
);

FILL FILL_1__1583_ (
);

FILL FILL_1__1163_ (
);

FILL FILL_3__1089_ (
);

FILL FILL_2__1232_ (
);

FILL FILL_0__1478_ (
);

FILL FILL_0__1058_ (
);

FILL FILL_0__805_ (
);

FILL FILL_3__949_ (
);

FILL FILL_3__1301_ (
);

NAND3X1 _808_ (
    .A(Cin_0_bF$buf2),
    .B(Xin_3_bF$buf0),
    .C(Yin[3]),
    .Y(_1_)
);

FILL FILL_1__1219_ (
);

INVX1 _1230_ (
    .A(_416_),
    .Y(_422_)
);

INVX1 _981_ (
    .A(_160_),
    .Y(_172_)
);

FILL FILL_1__1392_ (
);

FILL FILL_2__1461_ (
);

FILL FILL_2__1041_ (
);

FILL FILL_4__1387_ (
);

FILL FILL_0__1287_ (
);

FILL FILL88950x58650 (
);

FILL FILL_3__758_ (
);

FILL FILL_3__1110_ (
);

FILL FILL_1__1448_ (
);

FILL FILL_1__1028_ (
);

FILL FILL_1__821_ (
);

INVX1 _790_ (
    .A(_601_),
    .Y(_732_)
);

FILL FILL_2__1517_ (
);

FILL FILL_2__1270_ (
);

FILL FILL_0__1096_ (
);

INVX1 _1515_ (
    .A(_721_),
    .Y(_727_)
);

FILL FILL_0__843_ (
);

FILL FILL_3__987_ (
);

NAND3X1 _846_ (
    .A(_29_),
    .B(_35_),
    .C(_37_),
    .Y(_38_)
);

FILL FILL_1__1257_ (
);

FILL FILL_4__774_ (
);

FILL FILL_2__1326_ (
);

INVX1 _1324_ (
    .A(_501_),
    .Y(_523_)
);

FILL FILL_3__796_ (
);

FILL FILL_1__1486_ (
);

FILL FILL_1__1066_ (
);

FILL FILL_2__1135_ (
);

FILL FILL_3__1204_ (
);

DFFPOSX1 _1553_ (
    .D(_753_[9]),
    .CLK(clk_bF$buf5),
    .Q(y[9])
);

AND2X2 _1133_ (
    .A(Xin_3_bF$buf3),
    .B(Cin[5]),
    .Y(_322_)
);

FILL FILL_0__881_ (
);

FILL FILL_1__915_ (
);

OAI21X1 _884_ (
    .A(_744_),
    .B(_70_),
    .C(_63_),
    .Y(_76_)
);

FILL FILL_1__1295_ (
);

FILL FILL_2__1364_ (
);

FILL FILL_1_CLKBUF1_insert0 (
);

FILL FILL_1_CLKBUF1_insert1 (
);

FILL FILL_1_CLKBUF1_insert2 (
);

FILL FILL_1_CLKBUF1_insert3 (
);

FILL FILL_1_CLKBUF1_insert4 (
);

FILL FILL_1_CLKBUF1_insert5 (
);

FILL FILL_0__937_ (
);

FILL FILL_3__1433_ (
);

FILL FILL_3__1013_ (
);

NAND2X1 _1362_ (
    .A(_564_),
    .B(_558_),
    .Y(_565_)
);

FILL FILL_4__1502_ (
);

FILL FILL_0__1402_ (
);

FILL FILL_2__931_ (
);

FILL FILL_2__1173_ (
);

NAND2X1 _1418_ (
    .A(_624_),
    .B(_618_),
    .Y(_625_)
);

FILL FILL_3__1242_ (
);

AOI21X1 _1171_ (
    .A(Cin_0_bF$buf0),
    .B(Xin[7]),
    .C(Yin[7]),
    .Y(_360_)
);

FILL FILL_1__953_ (
);

FILL FILL_0__1211_ (
);

FILL FILL_2__1229_ (
);

FILL FILL88350x7950 (
);

NOR2X1 _1227_ (
    .A(_325_),
    .B(_417_),
    .Y(_419_)
);

FILL FILL_0__975_ (
);

FILL FILL_3__1471_ (
);

FILL FILL_3__1051_ (
);

NAND2X1 _978_ (
    .A(_164_),
    .B(_162_),
    .Y(_169_)
);

FILL FILL_1__1389_ (
);

FILL FILL_1__762_ (
);

FILL FILL_4__1120_ (
);

FILL FILL_0__1440_ (
);

FILL FILL_2__1458_ (
);

FILL FILL_0__1020_ (
);

FILL FILL_2__1038_ (
);

FILL FILL_3__911_ (
);

FILL FILL_3__1107_ (
);

NAND3X1 _1456_ (
    .A(_635_),
    .B(_660_),
    .C(_664_),
    .Y(_665_)
);

NAND3X1 _1036_ (
    .A(_225_),
    .B(_221_),
    .C(_223_),
    .Y(_226_)
);

FILL FILL_0__784_ (
);

FILL FILL_1__818_ (
);

FILL FILL89550x43050 (
);

FILL FILL_3__1280_ (
);

AOI21X1 _787_ (
    .A(_697_),
    .B(_676_),
    .C(_612_),
    .Y(_718_)
);

FILL FILL_1__1198_ (
);

FILL FILL_1__991_ (
);

FILL FILL_2__1267_ (
);

FILL FILL_1__1410_ (
);

FILL FILL_3__1336_ (
);

AOI21X1 _1265_ (
    .A(_263_),
    .B(_267_),
    .C(_371_),
    .Y(_459_)
);

FILL FILL_4__1405_ (
);

FILL FILL_0__1305_ (
);

FILL FILL_2__834_ (
);

FILL FILL_2__1496_ (
);

FILL FILL_2__1076_ (
);

FILL FILL_3__1565_ (
);

FILL FILL_3__1145_ (
);

INVX1 _1494_ (
    .A(_678_),
    .Y(_705_)
);

INVX1 _1074_ (
    .A(Yin[7]),
    .Y(_264_)
);

FILL FILL_1__856_ (
);

FILL FILL_0__1114_ (
);

FILL FILL_0__878_ (
);

FILL FILL_3__1374_ (
);

BUFX2 BUFX2_insert6 (
    .A(Cin[0]),
    .Y(Cin_0_bF$buf3)
);

BUFX2 BUFX2_insert7 (
    .A(Cin[0]),
    .Y(Cin_0_bF$buf2)
);

BUFX2 BUFX2_insert8 (
    .A(Cin[0]),
    .Y(Cin_0_bF$buf1)
);

BUFX2 BUFX2_insert9 (
    .A(Cin[0]),
    .Y(Cin_0_bF$buf0)
);

FILL FILL_4__1023_ (
);

FILL FILL_0__1343_ (
);

FILL FILL_2__872_ (
);

FILL FILL_3__814_ (
);

FILL FILL_1__1504_ (
);

NAND3X1 _1359_ (
    .A(_555_),
    .B(_498_),
    .C(_556_),
    .Y(_562_)
);

FILL FILL_3__1183_ (
);

FILL FILL_1__894_ (
);

FILL FILL_2__928_ (
);

FILL FILL_0__1572_ (
);

FILL FILL_0__1152_ (
);

AND2X2 _902_ (
    .A(_89_),
    .B(_93_),
    .Y(_94_)
);

FILL FILL_1__1313_ (
);

FILL FILL_3__1239_ (
);

NAND3X1 _1168_ (
    .A(Cin[2]),
    .B(Xin[6]),
    .C(_336_),
    .Y(_357_)
);

FILL FILL_0__1208_ (
);

FILL FILL89250x78150 (
);

FILL FILL_0__1381_ (
);

FILL FILL_2__1399_ (
);

FILL FILL_3__852_ (
);

FILL FILL_1__1122_ (
);

FILL FILL_3__1468_ (
);

FILL FILL_3__1048_ (
);

NAND2X1 _1397_ (
    .A(_599_),
    .B(_600_),
    .Y(_602_)
);

FILL FILL_1__759_ (
);

FILL FILL_0__1437_ (
);

FILL FILL_0__1017_ (
);

FILL FILL_2__966_ (
);

FILL FILL_3__908_ (
);

FILL FILL_4__1290_ (
);

FILL FILL_0__1190_ (
);

NAND3X1 _940_ (
    .A(_127_),
    .B(_131_),
    .C(_75_),
    .Y(_132_)
);

FILL FILL_1__1351_ (
);

FILL FILL_3__1277_ (
);

FILL FILL_1__988_ (
);

FILL FILL_2__1420_ (
);

FILL FILL_2__1000_ (
);

FILL FILL_0__1246_ (
);

FILL FILL_2__775_ (
);

FILL FILL_1__1407_ (
);

FILL FILL_3__890_ (
);

FILL FILL_1__1580_ (
);

FILL FILL_1__1160_ (
);

FILL FILL_3__1086_ (
);

FILL FILL_1__797_ (
);

FILL FILL_0__1475_ (
);

FILL FILL_0__1055_ (
);

FILL FILL_0__802_ (
);

FILL FILL_3__946_ (
);

OAI21X1 _805_ (
    .A(_623_),
    .B(_655_),
    .C(_644_),
    .Y(_746_)
);

FILL FILL_1__1216_ (
);

FILL FILL89550x31350 (
);

FILL FILL_0__1284_ (
);

FILL FILL_1__1445_ (
);

FILL FILL_1__1025_ (
);

FILL FILL_2__1514_ (
);

FILL FILL_2__869_ (
);

FILL FILL_4__1193_ (
);

FILL FILL_0__1093_ (
);

AOI21X1 _1512_ (
    .A(_723_),
    .B(_628_),
    .C(_696_),
    .Y(_724_)
);

FILL FILL_0__840_ (
);

FILL FILL_3__984_ (
);

NAND3X1 _843_ (
    .A(_30_),
    .B(_34_),
    .C(_32_),
    .Y(_35_)
);

FILL FILL_1__1254_ (
);

FILL FILL_2__1323_ (
);

FILL FILL_4__1249_ (
);

FILL FILL_0__1569_ (
);

FILL FILL_0__1149_ (
);

AOI21X1 _1321_ (
    .A(_444_),
    .B(_448_),
    .C(_519_),
    .Y(_520_)
);

FILL FILL_3__793_ (
);

FILL FILL_1__1483_ (
);

FILL FILL_1__1063_ (
);

FILL FILL_2__1132_ (
);

FILL FILL_0__1378_ (
);

FILL FILL_3__849_ (
);

FILL FILL_3__1201_ (
);

FILL FILL_1__1119_ (
);

DFFPOSX1 _1550_ (
    .D(_753_[6]),
    .CLK(clk_bF$buf0),
    .Q(y[6])
);

NAND2X1 _1130_ (
    .A(Xin[1]),
    .B(Cin[7]),
    .Y(_319_)
);

FILL FILL_1__912_ (
);

NAND2X1 _881_ (
    .A(_72_),
    .B(_23_),
    .Y(_73_)
);

FILL FILL_1__1292_ (
);

FILL FILL_2__1361_ (
);

FILL FILL_0__1187_ (
);

FILL FILL_0__934_ (
);

FILL FILL_3__1430_ (
);

FILL FILL_3__1010_ (
);

AOI21X1 _937_ (
    .A(_124_),
    .B(_125_),
    .C(_123_),
    .Y(_129_)
);

FILL FILL_1__1348_ (
);

FILL FILL_2__1417_ (
);

FILL FILL_2__1170_ (
);

NAND3X1 _1415_ (
    .A(_570_),
    .B(_615_),
    .C(_616_),
    .Y(_621_)
);

FILL FILL_3__887_ (
);

FILL FILL_1__1577_ (
);

FILL FILL_1__1157_ (
);

FILL FILL_1__950_ (
);

FILL FILL_2__1226_ (
);

NAND2X1 _1224_ (
    .A(Xin[2]),
    .B(Cin[7]),
    .Y(_415_)
);

FILL FILL_0__972_ (
);

AOI21X1 _975_ (
    .A(_165_),
    .B(_163_),
    .C(_161_),
    .Y(_166_)
);

FILL FILL_1__1386_ (
);

FILL FILL_2__1455_ (
);

FILL FILL_2__1035_ (
);

FILL FILL_3__1104_ (
);

NOR2X1 _1453_ (
    .A(_637_),
    .B(_659_),
    .Y(_662_)
);

NAND2X1 _1033_ (
    .A(_140_),
    .B(_222_),
    .Y(_223_)
);

FILL FILL_0__781_ (
);

FILL FILL_1__815_ (
);

INVX1 _784_ (
    .A(_644_),
    .Y(_687_)
);

FILL FILL_1__1195_ (
);

FILL FILL_2__1264_ (
);

XOR2X1 _1509_ (
    .A(_717_),
    .B(_720_),
    .Y(_721_)
);

FILL FILL_0__837_ (
);

FILL FILL_3__1333_ (
);

INVX1 _1262_ (
    .A(_453_),
    .Y(_456_)
);

FILL FILL_0__1302_ (
);

FILL FILL_2__831_ (
);

FILL FILL_2__1493_ (
);

FILL FILL_2__1073_ (
);

AOI21X1 _1318_ (
    .A(_510_),
    .B(_511_),
    .C(_508_),
    .Y(_517_)
);

FILL FILL_3__1562_ (
);

FILL FILL_3__1142_ (
);

NOR2X1 _1491_ (
    .A(_686_),
    .B(_701_),
    .Y(_702_)
);

NAND2X1 _1071_ (
    .A(Cin[1]),
    .B(Xin[6]),
    .Y(_261_)
);

FILL FILL_1__853_ (
);

FILL FILL_0__1111_ (
);

FILL FILL_2__1129_ (
);

DFFPOSX1 _1547_ (
    .D(_751_[3]),
    .CLK(clk_bF$buf3),
    .Q(y[3])
);

AOI21X1 _1127_ (
    .A(_276_),
    .B(_280_),
    .C(_246_),
    .Y(_316_)
);

FILL FILL_0__875_ (
);

FILL FILL_1__909_ (
);

FILL FILL_3__1371_ (
);

AOI21X1 _878_ (
    .A(_62_),
    .B(_56_),
    .C(_27_),
    .Y(_70_)
);

FILL FILL_1__1289_ (
);

FILL FILL_2__1358_ (
);

FILL FILL_0__1340_ (
);

FILL FILL_3__811_ (
);

FILL FILL_1__1501_ (
);

FILL FILL_3__1427_ (
);

FILL FILL_3__1007_ (
);

OAI21X1 _1356_ (
    .A(_554_),
    .B(_557_),
    .C(_497_),
    .Y(_558_)
);

FILL FILL_3__1180_ (
);

FILL FILL_1__1098_ (
);

FILL FILL_1__891_ (
);

FILL FILL_2__925_ (
);

FILL FILL_2__1167_ (
);

FILL FILL_1__1310_ (
);

FILL FILL_3__1236_ (
);

NAND3X1 _1165_ (
    .A(_353_),
    .B(_349_),
    .C(_351_),
    .Y(_354_)
);

FILL FILL_1__947_ (
);

FILL FILL_0__1205_ (
);

FILL FILL_2__1396_ (
);

FILL FILL_0__969_ (
);

FILL FILL_3__1465_ (
);

FILL FILL_3__1045_ (
);

XNOR2X1 _1394_ (
    .A(_532_),
    .B(Yin[11]),
    .Y(_598_)
);

FILL FILL_1__756_ (
);

FILL FILL_0__1434_ (
);

FILL FILL_0__1014_ (
);

FILL FILL89250x54750 (
);

FILL FILL_2__963_ (
);

FILL FILL_3__905_ (
);

FILL FILL_0__778_ (
);

FILL FILL_3__1274_ (
);

FILL FILL_1__985_ (
);

FILL FILL_0__1243_ (
);

FILL FILL_2__772_ (
);

FILL FILL_1__1404_ (
);

FILL FILL_4__921_ (
);

XNOR2X1 _1259_ (
    .A(_362_),
    .B(Yin[9]),
    .Y(_453_)
);

FILL FILL_3__1083_ (
);

FILL FILL_1__794_ (
);

FILL FILL_2__828_ (
);

FILL FILL_4__1152_ (
);

FILL FILL_0__1472_ (
);

FILL FILL_0__1052_ (
);

FILL FILL_3__943_ (
);

AND2X2 _802_ (
    .A(Xin[1]),
    .B(Cin[3]),
    .Y(_743_)
);

FILL FILL_1__1213_ (
);

FILL FILL_3__1139_ (
);

OAI21X1 _1488_ (
    .A(_674_),
    .B(_693_),
    .C(_670_),
    .Y(_699_)
);

AND2X2 _1068_ (
    .A(_257_),
    .B(_254_),
    .Y(_258_)
);

FILL FILL_0__1108_ (
);

FILL FILL_0__1281_ (
);

FILL FILL_2__1299_ (
);

FILL FILL_1__1442_ (
);

FILL FILL_1__1022_ (
);

FILL FILL_3__1368_ (
);

NOR2X1 _1297_ (
    .A(_404_),
    .B(_490_),
    .Y(_494_)
);

FILL FILL_2__1511_ (
);

FILL FILL_4__1437_ (
);

FILL FILL_0__1337_ (
);

FILL FILL_2__866_ (
);

FILL FILL_3__808_ (
);

FILL FILL_0__1090_ (
);

FILL FILL_3__981_ (
);

INVX1 _840_ (
    .A(_31_),
    .Y(_32_)
);

FILL FILL_1__1251_ (
);

FILL FILL_3__1177_ (
);

FILL FILL_1__888_ (
);

FILL FILL_2__1320_ (
);

FILL FILL_0__1566_ (
);

FILL FILL_0__1146_ (
);

FILL FILL_1__1307_ (
);

FILL FILL_3__790_ (
);

FILL FILL_4__824_ (
);

FILL FILL_1__1480_ (
);

FILL FILL_1__1060_ (
);

FILL FILL_4__1055_ (
);

FILL FILL_0__1375_ (
);

FILL FILL_3__846_ (
);

FILL FILL_1__1116_ (
);

FILL FILL_0__1184_ (
);

FILL FILL_0__931_ (
);

NAND3X1 _934_ (
    .A(_123_),
    .B(_125_),
    .C(_124_),
    .Y(_126_)
);

FILL FILL_1__1345_ (
);

FILL FILL_2__1414_ (
);

FILL FILL_2__769_ (
);

OAI21X1 _1412_ (
    .A(_614_),
    .B(_617_),
    .C(_568_),
    .Y(_618_)
);

FILL FILL_3__884_ (
);

FILL FILL_1__1574_ (
);

FILL FILL_1__1154_ (
);

FILL FILL89250x4050 (
);

FILL FILL_2__1223_ (
);

FILL FILL_0__1469_ (
);

FILL FILL_0__1049_ (
);

FILL FILL_2__998_ (
);

OAI21X1 _1221_ (
    .A(_345_),
    .B(_411_),
    .C(_383_),
    .Y(_412_)
);

NAND2X1 _972_ (
    .A(Yin[6]),
    .B(_162_),
    .Y(_163_)
);

FILL FILL_1__1383_ (
);

FILL FILL_2__1452_ (
);

FILL FILL_2__1032_ (
);

FILL FILL_4__1378_ (
);

FILL FILL_0__1278_ (
);

FILL FILL_3__1101_ (
);

FILL FILL_1__1439_ (
);

FILL FILL_1__1019_ (
);

NAND2X1 _1450_ (
    .A(_658_),
    .B(_657_),
    .Y(_659_)
);

NAND2X1 _1030_ (
    .A(Xin[0]),
    .B(Cin[7]),
    .Y(_220_)
);

FILL FILL_1__812_ (
);

AOI21X1 _781_ (
    .A(Cin_0_bF$buf1),
    .B(Xin[2]),
    .C(Yin[2]),
    .Y(_655_)
);

FILL FILL_1__1192_ (
);

FILL FILL_2__1508_ (
);

FILL FILL_2__1261_ (
);

FILL FILL_0__1087_ (
);

NAND3X1 _1506_ (
    .A(_703_),
    .B(_706_),
    .C(_711_),
    .Y(_717_)
);

FILL FILL_0__834_ (
);

FILL FILL_3__978_ (
);

FILL FILL_3__1330_ (
);

OAI21X1 _837_ (
    .A(_747_),
    .B(_28_),
    .C(_1_),
    .Y(_29_)
);

FILL FILL_1__1248_ (
);

FILL FILL_4__765_ (
);

FILL FILL_2__1317_ (
);

FILL FILL_2__1490_ (
);

FILL FILL_2__1070_ (
);

NOR2X1 _1315_ (
    .A(_350_),
    .B(_445_),
    .Y(_513_)
);

FILL FILL_3__787_ (
);

FILL FILL_1__1477_ (
);

FILL FILL_1__1057_ (
);

FILL FILL_1__850_ (
);

FILL FILL_2__1126_ (
);

DFFPOSX1 _1544_ (
    .D(_748_[0]),
    .CLK(clk_bF$buf4),
    .Q(y[0])
);

AOI21X1 _1124_ (
    .A(_215_),
    .B(_297_),
    .C(_312_),
    .Y(_313_)
);

FILL FILL_0__872_ (
);

FILL FILL_1__906_ (
);

NAND3X1 _875_ (
    .A(_65_),
    .B(_66_),
    .C(_64_),
    .Y(_67_)
);

FILL FILL_1__1286_ (
);

FILL FILL89250x19650 (
);

FILL FILL_2__1355_ (
);

FILL FILL_0__928_ (
);

FILL FILL_3__1424_ (
);

FILL FILL_3__1004_ (
);

NAND3X1 _1353_ (
    .A(_551_),
    .B(_552_),
    .C(_500_),
    .Y(_555_)
);

FILL FILL_1__1095_ (
);

FILL FILL_2__922_ (
);

FILL FILL_2__1164_ (
);

NAND3X1 _1409_ (
    .A(_604_),
    .B(_607_),
    .C(_573_),
    .Y(_615_)
);

FILL FILL_3__1233_ (
);

BUFX2 _1582_ (
    .A(_755_[8]),
    .Y(Yout[8])
);

NAND2X1 _1162_ (
    .A(_250_),
    .B(_350_),
    .Y(_351_)
);

FILL FILL_1__944_ (
);

FILL FILL_0__1202_ (
);

FILL FILL_2__1393_ (
);

OAI21X1 _1218_ (
    .A(_315_),
    .B(_408_),
    .C(_394_),
    .Y(_409_)
);

FILL FILL_0__966_ (
);

FILL FILL_3__1462_ (
);

FILL FILL_3__1042_ (
);

OAI21X1 _969_ (
    .A(_96_),
    .B(_159_),
    .C(_98_),
    .Y(_160_)
);

NAND3X1 _1391_ (
    .A(_588_),
    .B(_581_),
    .C(_586_),
    .Y(_595_)
);

FILL FILL_0__1431_ (
);

FILL FILL_2__1449_ (
);

FILL FILL_0__1011_ (
);

FILL FILL_2__1029_ (
);

FILL FILL89550x58650 (
);

FILL FILL_2__960_ (
);

FILL FILL_3__902_ (
);

FILL FILL_3__1518_ (
);

INVX1 _1447_ (
    .A(_654_),
    .Y(_656_)
);

OAI21X1 _1027_ (
    .A(_144_),
    .B(_216_),
    .C(_189_),
    .Y(_217_)
);

FILL FILL_0__775_ (
);

FILL FILL_1__809_ (
);

FILL FILL_3__1271_ (
);

NAND2X1 _778_ (
    .A(Xin[1]),
    .B(Cin[1]),
    .Y(_623_)
);

FILL FILL_1__1189_ (
);

FILL FILL_1__982_ (
);

FILL FILL_0__1240_ (
);

FILL FILL_2__1258_ (
);

FILL FILL_1__1401_ (
);

FILL FILL_3__1327_ (
);

OAI21X1 _1256_ (
    .A(_590_),
    .B(_447_),
    .C(_350_),
    .Y(_450_)
);

FILL FILL_3__1080_ (
);

FILL FILL_1__791_ (
);

FILL FILL_2__825_ (
);

FILL FILL_2__1487_ (
);

FILL FILL_2__1067_ (
);

FILL FILL_3__940_ (
);

FILL FILL_1__1210_ (
);

FILL FILL_3__1136_ (
);

NAND2X1 _1485_ (
    .A(_674_),
    .B(_693_),
    .Y(_695_)
);

NAND2X1 _1065_ (
    .A(_252_),
    .B(_249_),
    .Y(_255_)
);

FILL FILL_1__847_ (
);

FILL FILL_0__1105_ (
);

FILL FILL_2__1296_ (
);

FILL FILL_0__869_ (
);

FILL FILL_3__1365_ (
);

XNOR2X1 _1294_ (
    .A(_406_),
    .B(_490_),
    .Y(_753_[9])
);

FILL FILL_4__1014_ (
);

FILL FILL_0__1334_ (
);

FILL FILL_2__863_ (
);

FILL FILL_3__805_ (
);

FILL FILL_3__1174_ (
);

FILL FILL_1__885_ (
);

FILL FILL_2__919_ (
);

FILL FILL_0__1563_ (
);

FILL FILL_0__1143_ (
);

FILL FILL_1__1304_ (
);

FILL FILL_0_BUFX2_insert10 (
);

FILL FILL_0_BUFX2_insert11 (
);

FILL FILL_0_BUFX2_insert12 (
);

FILL FILL_0_BUFX2_insert13 (
);

BUFX2 _1579_ (
    .A(_755_[5]),
    .Y(Yout[5])
);

FILL FILL_0_BUFX2_insert14 (
);

FILL FILL_0_BUFX2_insert15 (
);

NAND2X1 _1159_ (
    .A(Xin[4]),
    .B(Cin[4]),
    .Y(_348_)
);

FILL FILL_0_BUFX2_insert16 (
);

FILL FILL_0_BUFX2_insert17 (
);

FILL FILL_0__1372_ (
);

FILL FILL_3__843_ (
);

FILL FILL_1__1113_ (
);

FILL FILL_3__1459_ (
);

FILL FILL_3__1039_ (
);

OAI21X1 _1388_ (
    .A(_591_),
    .B(_589_),
    .C(_588_),
    .Y(_592_)
);

FILL FILL_0__1428_ (
);

FILL FILL_0__1008_ (
);

FILL FILL_2__957_ (
);

FILL FILL_4__1281_ (
);

FILL FILL_0__1181_ (
);

FILL FILL_2__1199_ (
);

XOR2X1 _931_ (
    .A(_80_),
    .B(_122_),
    .Y(_123_)
);

FILL FILL_1__1342_ (
);

FILL FILL_3__1268_ (
);

OAI21X1 _1197_ (
    .A(_381_),
    .B(_385_),
    .C(_317_),
    .Y(_387_)
);

FILL FILL_1__979_ (
);

FILL FILL_2__1411_ (
);

FILL FILL_0__1237_ (
);

FILL FILL_2__766_ (
);

FILL FILL_3__881_ (
);

FILL FILL_1__1571_ (
);

FILL FILL_1__1151_ (
);

FILL FILL_3__1497_ (
);

FILL FILL_3__1077_ (
);

FILL FILL_1__788_ (
);

FILL FILL89550x46950 (
);

FILL FILL_2__1220_ (
);

FILL FILL_0__1466_ (
);

FILL FILL_0__1046_ (
);

FILL FILL_2__995_ (
);

FILL FILL_3__937_ (
);

FILL FILL_1__1207_ (
);

FILL FILL_1__1380_ (
);

FILL FILL_0__1275_ (
);

FILL FILL_1__1436_ (
);

FILL FILL_1__1016_ (
);

FILL FILL_4__953_ (
);

FILL FILL_2__1505_ (
);

FILL FILL_4__1184_ (
);

FILL FILL_0__1084_ (
);

XOR2X1 _1503_ (
    .A(_700_),
    .B(_714_),
    .Y(_753_[14])
);

FILL FILL_0__831_ (
);

FILL FILL_3__975_ (
);

INVX1 _834_ (
    .A(_744_),
    .Y(_26_)
);

FILL FILL_1__1245_ (
);

FILL FILL_2__1314_ (
);

NAND2X1 _1312_ (
    .A(_423_),
    .B(_509_),
    .Y(_510_)
);

FILL FILL_3__784_ (
);

FILL FILL_1__1474_ (
);

FILL FILL_1__1054_ (
);

FILL FILL_2__1123_ (
);

FILL FILL_0__1369_ (
);

FILL FILL_2__898_ (
);

DFFPOSX1 _1541_ (
    .D(y[13]),
    .CLK(clk_bF$buf5),
    .Q(_755_[13])
);

AND2X2 _1121_ (
    .A(_302_),
    .B(_207_),
    .Y(_310_)
);

FILL FILL_1__903_ (
);

AOI21X1 _872_ (
    .A(_745_),
    .B(_13_),
    .C(_17_),
    .Y(_64_)
);

FILL FILL_1__1283_ (
);

FILL FILL_2__1352_ (
);

FILL FILL_0__1178_ (
);

FILL FILL_0__925_ (
);

FILL FILL_3__1421_ (
);

FILL FILL_3__1001_ (
);

OAI21X1 _928_ (
    .A(_119_),
    .B(_118_),
    .C(_117_),
    .Y(_120_)
);

FILL FILL_1__1339_ (
);

NAND2X1 _1350_ (
    .A(_528_),
    .B(_540_),
    .Y(_552_)
);

FILL FILL_1__1092_ (
);

FILL FILL_2__1408_ (
);

FILL FILL_2__1581_ (
);

FILL FILL_2__1161_ (
);

FILL FILL_4__1087_ (
);

AOI21X1 _1406_ (
    .A(_542_),
    .B(_546_),
    .C(_610_),
    .Y(_611_)
);

FILL FILL_3__878_ (
);

FILL FILL_3__1230_ (
);

FILL FILL_1__1568_ (
);

FILL FILL_1__1148_ (
);

FILL FILL_1__941_ (
);

FILL FILL_2__1217_ (
);

FILL FILL_2__1390_ (
);

INVX1 _1215_ (
    .A(_311_),
    .Y(_405_)
);

FILL FILL_0__963_ (
);

NAND3X1 _966_ (
    .A(_147_),
    .B(_155_),
    .C(_156_),
    .Y(_157_)
);

FILL FILL_1__1377_ (
);

FILL FILL_4__894_ (
);

FILL FILL_2__1446_ (
);

FILL FILL_2__1026_ (
);

FILL FILL_3__1515_ (
);

OR2X2 _1444_ (
    .A(_651_),
    .B(_650_),
    .Y(_652_)
);

NAND2X1 _1024_ (
    .A(_142_),
    .B(_143_),
    .Y(_214_)
);

FILL FILL_0__772_ (
);

FILL FILL_1__806_ (
);

INVX2 _775_ (
    .A(Cin[2]),
    .Y(_590_)
);

FILL FILL_1__1186_ (
);

FILL FILL_2__1255_ (
);

FILL FILL_0__828_ (
);

FILL FILL_3__1324_ (
);

INVX1 _1253_ (
    .A(Xin[7]),
    .Y(_447_)
);

FILL FILL_2__822_ (
);

FILL FILL_2__1484_ (
);

FILL FILL_2__1064_ (
);

OAI21X1 _1309_ (
    .A(_506_),
    .B(_505_),
    .C(_502_),
    .Y(_507_)
);

FILL FILL_3__1133_ (
);

NAND2X1 _1482_ (
    .A(_692_),
    .B(_688_),
    .Y(_693_)
);

NAND2X1 _1062_ (
    .A(Cin[2]),
    .B(Xin_5_bF$buf2),
    .Y(_252_)
);

FILL FILL_1__844_ (
);

FILL FILL_0__1102_ (
);

FILL FILL_2__1293_ (
);

DFFPOSX1 _1538_ (
    .D(y[10]),
    .CLK(clk_bF$buf5),
    .Q(_755_[10])
);

NAND2X1 _1118_ (
    .A(_302_),
    .B(_307_),
    .Y(_308_)
);

FILL FILL_0__866_ (
);

FILL FILL_3__1362_ (
);

NAND2X1 _869_ (
    .A(_59_),
    .B(_60_),
    .Y(_61_)
);

AOI21X1 _1291_ (
    .A(_477_),
    .B(_469_),
    .C(_410_),
    .Y(_488_)
);

FILL FILL_4__797_ (
);

FILL FILL_0__1331_ (
);

FILL FILL_2__1349_ (
);

FILL FILL_2__860_ (
);

FILL FILL_3__802_ (
);

FILL FILL_3__1418_ (
);

OAI21X1 _1347_ (
    .A(_541_),
    .B(_547_),
    .C(_500_),
    .Y(_549_)
);

FILL FILL_3__1171_ (
);

FILL FILL_1__1089_ (
);

FILL FILL_1__882_ (
);

FILL FILL_2__916_ (
);

FILL FILL_2__1578_ (
);

FILL FILL_0__1560_ (
);

FILL FILL_2__1158_ (
);

FILL FILL_0__1140_ (
);

FILL FILL_1__1301_ (
);

FILL FILL_3__1227_ (
);

BUFX2 _1576_ (
    .A(_755_[2]),
    .Y(Yout[2])
);

NAND2X1 _1156_ (
    .A(_340_),
    .B(_344_),
    .Y(_345_)
);

FILL FILL_1__938_ (
);

FILL FILL_2__1387_ (
);

FILL FILL_3__840_ (
);

FILL FILL88050x74250 (
);

FILL FILL_1__1110_ (
);

FILL FILL_3__1456_ (
);

FILL FILL_3__1036_ (
);

INVX1 _1385_ (
    .A(_536_),
    .Y(_588_)
);

FILL FILL_0__1425_ (
);

FILL FILL_0__1005_ (
);

FILL FILL_2__954_ (
);

FILL FILL_2__1196_ (
);

FILL FILL_0__769_ (
);

FILL FILL_3__1265_ (
);

NAND3X1 _1194_ (
    .A(_379_),
    .B(_347_),
    .C(_378_),
    .Y(_383_)
);

FILL FILL_1__976_ (
);

FILL FILL_0__1234_ (
);

FILL FILL_2__763_ (
);

FILL FILL_4__912_ (
);

FILL FILL_0__998_ (
);

FILL FILL_3__1494_ (
);

FILL FILL_3__1074_ (
);

FILL FILL_1__785_ (
);

FILL FILL_2__819_ (
);

FILL FILL_4__1143_ (
);

FILL FILL_0__1463_ (
);

FILL FILL_0__1043_ (
);

FILL FILL_2__992_ (
);

FILL FILL_3__934_ (
);

FILL FILL_1__1204_ (
);

INVX1 _1479_ (
    .A(_683_),
    .Y(_690_)
);

AND2X2 _1059_ (
    .A(Cin[3]),
    .B(Xin[4]),
    .Y(_249_)
);

FILL FILL_0__1519_ (
);

FILL FILL_0__1272_ (
);

FILL FILL_1__1433_ (
);

FILL FILL_1__1013_ (
);

FILL FILL_3__1359_ (
);

INVX1 _1288_ (
    .A(_394_),
    .Y(_485_)
);

FILL FILL_2__1502_ (
);

FILL FILL_4__1428_ (
);

FILL FILL_0__1328_ (
);

FILL FILL_2__857_ (
);

FILL FILL_2__1099_ (
);

FILL FILL_0__1081_ (
);

XNOR2X1 _1500_ (
    .A(_711_),
    .B(_707_),
    .Y(_712_)
);

FILL FILL_3__972_ (
);

INVX1 _831_ (
    .A(_23_),
    .Y(_24_)
);

FILL FILL_1__1242_ (
);

FILL FILL_3__1168_ (
);

NAND3X1 _1097_ (
    .A(_281_),
    .B(_286_),
    .C(_244_),
    .Y(_287_)
);

FILL FILL_1__879_ (
);

FILL FILL_2__1311_ (
);

FILL FILL_0__1137_ (
);

FILL FILL_3__781_ (
);

FILL FILL_4__815_ (
);

FILL FILL_1__1471_ (
);

FILL FILL_1__1051_ (
);

FILL FILL_3__1397_ (
);

FILL FILL_2__1120_ (
);

FILL FILL_4__1046_ (
);

FILL FILL_0__1366_ (
);

FILL FILL_2__895_ (
);

FILL FILL_3__837_ (
);

FILL FILL_1__1107_ (
);

FILL FILL_1__900_ (
);

FILL FILL_1__1280_ (
);

FILL FILL_0__1175_ (
);

FILL FILL_0__922_ (
);

AOI21X1 _925_ (
    .A(_43_),
    .B(_55_),
    .C(_57_),
    .Y(_117_)
);

FILL FILL_1__1336_ (
);

FILL FILL_2__1405_ (
);

NAND2X1 _1403_ (
    .A(_604_),
    .B(_607_),
    .Y(_608_)
);

FILL FILL_3__875_ (
);

FILL FILL_1__1565_ (
);

FILL FILL_1__1145_ (
);

FILL FILL_2__1214_ (
);

FILL FILL_2__989_ (
);

NAND3X1 _1212_ (
    .A(_400_),
    .B(_401_),
    .C(_402_),
    .Y(_403_)
);

FILL FILL_0__960_ (
);

NAND3X1 _963_ (
    .A(_153_),
    .B(_148_),
    .C(_150_),
    .Y(_154_)
);

FILL FILL_1__1374_ (
);

FILL FILL_2__1443_ (
);

FILL FILL_2__1023_ (
);

FILL FILL_0__1269_ (
);

FILL FILL_2__798_ (
);

FILL FILL_3__1512_ (
);

NOR2X1 _1441_ (
    .A(_648_),
    .B(_647_),
    .Y(_649_)
);

NAND2X1 _1021_ (
    .A(_207_),
    .B(_208_),
    .Y(_211_)
);

FILL FILL_1__803_ (
);

INVX1 _772_ (
    .A(_548_),
    .Y(_559_)
);

FILL FILL_1__1183_ (
);

FILL FILL_2__1252_ (
);

FILL FILL_0__1498_ (
);

FILL FILL_0__1078_ (
);

FILL FILL_0__825_ (
);

FILL FILL_3__969_ (
);

FILL FILL_3__1321_ (
);

NOR2X1 _828_ (
    .A(_739_),
    .B(_20_),
    .Y(_21_)
);

FILL FILL_1__1239_ (
);

INVX1 _1250_ (
    .A(_443_),
    .Y(_444_)
);

FILL FILL_2__1308_ (
);

FILL FILL_2__1481_ (
);

FILL FILL_2__1061_ (
);

NAND2X1 _1306_ (
    .A(Xin_5_bF$buf3),
    .B(Cin[5]),
    .Y(_503_)
);

FILL FILL_3__778_ (
);

FILL FILL_3__1130_ (
);

FILL FILL_1__1468_ (
);

FILL FILL_1__1048_ (
);

FILL FILL_1__841_ (
);

FILL FILL_2__1117_ (
);

FILL FILL_2__1290_ (
);

DFFPOSX1 _1535_ (
    .D(y[7]),
    .CLK(clk_bF$buf0),
    .Q(_755_[7])
);

AOI21X1 _1115_ (
    .A(_300_),
    .B(_299_),
    .C(_214_),
    .Y(_305_)
);

FILL FILL_0__863_ (
);

AOI21X1 _866_ (
    .A(_37_),
    .B(_35_),
    .C(_29_),
    .Y(_58_)
);

FILL FILL_1__1277_ (
);

FILL FILL_2__1346_ (
);

FILL FILL_0__919_ (
);

FILL FILL_3__1415_ (
);

NAND3X1 _1344_ (
    .A(_529_),
    .B(_454_),
    .C(_544_),
    .Y(_545_)
);

FILL FILL_1__1086_ (
);

FILL FILL_2__913_ (
);

FILL FILL_2__1575_ (
);

FILL FILL_2__1155_ (
);

FILL FILL_3__1224_ (
);

BUFX2 _1573_ (
    .A(_755_[13]),
    .Y(Yout[13])
);

NAND3X1 _1153_ (
    .A(_327_),
    .B(_338_),
    .C(_330_),
    .Y(_342_)
);

FILL FILL_1__935_ (
);

FILL FILL_2__1384_ (
);

OAI21X1 _1209_ (
    .A(_214_),
    .B(_399_),
    .C(_292_),
    .Y(_400_)
);

FILL FILL88350x78150 (
);

FILL FILL_0__957_ (
);

FILL FILL_3__1453_ (
);

FILL FILL_3__1033_ (
);

INVX1 _1382_ (
    .A(_584_),
    .Y(_585_)
);

FILL FILL_0__1422_ (
);

FILL FILL_0__1002_ (
);

FILL FILL_2__951_ (
);

FILL FILL89250x7950 (
);

FILL FILL_2__1193_ (
);

FILL FILL_3__1509_ (
);

NAND3X1 _1438_ (
    .A(_638_),
    .B(_642_),
    .C(_645_),
    .Y(_646_)
);

INVX1 _1018_ (
    .A(_208_),
    .Y(_209_)
);

FILL FILL_0__766_ (
);

FILL FILL_3__1262_ (
);

INVX1 _769_ (
    .A(_483_),
    .Y(_526_)
);

NAND3X1 _1191_ (
    .A(_378_),
    .B(_379_),
    .C(_376_),
    .Y(_380_)
);

FILL FILL_1__973_ (
);

FILL FILL_0__1231_ (
);

FILL FILL_2__1249_ (
);

FILL FILL_2__760_ (
);

FILL FILL_3__1318_ (
);

NOR2X1 _1247_ (
    .A(_361_),
    .B(_366_),
    .Y(_441_)
);

FILL FILL_0__995_ (
);

FILL FILL_3__1491_ (
);

FILL FILL_3__1071_ (
);

NAND3X1 _998_ (
    .A(_146_),
    .B(_185_),
    .C(_184_),
    .Y(_189_)
);

FILL FILL_1__782_ (
);

FILL FILL_2__816_ (
);

FILL FILL_4__1560_ (
);

FILL FILL_0__1460_ (
);

FILL FILL_2__1478_ (
);

FILL FILL_0__1040_ (
);

FILL FILL_2__1058_ (
);

FILL FILL_3__931_ (
);

FILL FILL_1__1201_ (
);

FILL FILL_3__1127_ (
);

AOI21X1 _1476_ (
    .A(_652_),
    .B(_657_),
    .C(_683_),
    .Y(_686_)
);

OAI21X1 _1056_ (
    .A(_245_),
    .B(_158_),
    .C(_177_),
    .Y(_246_)
);

FILL FILL_1__838_ (
);

FILL FILL_0__1516_ (
);

FILL FILL_2__1287_ (
);

FILL FILL_1__1430_ (
);

FILL FILL_1__1010_ (
);

FILL FILL_3__1356_ (
);

NAND3X1 _1285_ (
    .A(_464_),
    .B(_468_),
    .C(_471_),
    .Y(_481_)
);

FILL FILL_4__1005_ (
);

FILL FILL_0__1325_ (
);

FILL FILL_2__854_ (
);

FILL FILL_2__1096_ (
);

FILL FILL_3__1165_ (
);

AOI21X1 _1094_ (
    .A(_278_),
    .B(_279_),
    .C(_277_),
    .Y(_284_)
);

FILL FILL_1__876_ (
);

FILL FILL_0__1134_ (
);

FILL FILL_0__898_ (
);

FILL FILL_3__1394_ (
);

FILL FILL_0__1363_ (
);

FILL FILL_2__892_ (
);

FILL FILL_3__834_ (
);

FILL FILL_1__1104_ (
);

NAND2X1 _1379_ (
    .A(Xin[4]),
    .B(Cin[7]),
    .Y(_582_)
);

FILL FILL_0__1419_ (
);

FILL FILL_2__948_ (
);

FILL FILL_4__1272_ (
);

FILL FILL_0__1172_ (
);

NAND3X1 _922_ (
    .A(_102_),
    .B(_105_),
    .C(_107_),
    .Y(_114_)
);

FILL FILL_1__1333_ (
);

FILL FILL_3__1259_ (
);

AND2X2 _1188_ (
    .A(_354_),
    .B(_358_),
    .Y(_377_)
);

FILL FILL_2__1402_ (
);

FILL FILL_0__1228_ (
);

FILL FILL_2__757_ (
);

AOI21X1 _1400_ (
    .A(_596_),
    .B(_595_),
    .C(_594_),
    .Y(_605_)
);

FILL FILL_3__872_ (
);

FILL FILL_1__1562_ (
);

FILL FILL_1__1142_ (
);

FILL FILL_3__1488_ (
);

FILL FILL_3__1068_ (
);

FILL FILL_1__779_ (
);

FILL FILL_2__1211_ (
);

FILL FILL_0__1457_ (
);

FILL FILL_0__1037_ (
);

FILL FILL_2__986_ (
);

FILL FILL_3__928_ (
);

INVX2 _960_ (
    .A(Xin[4]),
    .Y(_151_)
);

FILL FILL_1__1371_ (
);

FILL FILL_3__1297_ (
);

FILL FILL_2__1440_ (
);

FILL FILL_2__1020_ (
);

FILL FILL_0__1266_ (
);

FILL FILL_2__795_ (
);

FILL FILL_1__1427_ (
);

FILL FILL_1__1007_ (
);

FILL FILL_1__800_ (
);

FILL FILL_4__944_ (
);

FILL FILL_1__1180_ (
);

FILL FILL_4__1175_ (
);

FILL FILL_0__1495_ (
);

FILL FILL_0__1075_ (
);

FILL FILL_0__822_ (
);

FILL FILL_3__966_ (
);

AOI21X1 _825_ (
    .A(_8_),
    .B(_5_),
    .C(_746_),
    .Y(_18_)
);

FILL FILL_1__1236_ (
);

FILL FILL_2__1305_ (
);

OAI21X1 _1303_ (
    .A(_467_),
    .B(_465_),
    .C(_458_),
    .Y(_500_)
);

FILL FILL_3__775_ (
);

FILL FILL_1__1465_ (
);

FILL FILL_1__1045_ (
);

FILL FILL_2__1114_ (
);

FILL FILL_2__889_ (
);

DFFPOSX1 _1532_ (
    .D(y[4]),
    .CLK(clk_bF$buf3),
    .Q(_755_[4])
);

NAND3X1 _1112_ (
    .A(_213_),
    .B(_298_),
    .C(_301_),
    .Y(_302_)
);

FILL FILL_0__860_ (
);

NAND2X1 _863_ (
    .A(_49_),
    .B(_54_),
    .Y(_55_)
);

FILL FILL_1__1274_ (
);

FILL FILL_2__1343_ (
);

FILL FILL_0__1169_ (
);

FILL FILL_0__916_ (
);

FILL FILL_3__1412_ (
);

NAND3X1 _919_ (
    .A(_106_),
    .B(_110_),
    .C(_94_),
    .Y(_111_)
);

AND2X2 _1341_ (
    .A(_522_),
    .B(_527_),
    .Y(_542_)
);

FILL FILL_1__1083_ (
);

FILL FILL_2__910_ (
);

FILL FILL_2__1572_ (
);

FILL FILL_2__1152_ (
);

FILL FILL_4__1078_ (
);

FILL FILL_0__1398_ (
);

FILL FILL_3__869_ (
);

FILL FILL_3__1221_ (
);

FILL FILL_1__1139_ (
);

BUFX2 _1570_ (
    .A(_755_[10]),
    .Y(Yout[10])
);

OAI21X1 _1150_ (
    .A(_335_),
    .B(_334_),
    .C(_338_),
    .Y(_339_)
);

FILL FILL_1__932_ (
);

FILL FILL_2__1208_ (
);

FILL FILL_2__1381_ (
);

AOI21X1 _1206_ (
    .A(_395_),
    .B(_394_),
    .C(_314_),
    .Y(_396_)
);

FILL FILL_0__954_ (
);

FILL FILL_3__1450_ (
);

FILL FILL_3__1030_ (
);

INVX1 _957_ (
    .A(_147_),
    .Y(_148_)
);

FILL FILL_1__1368_ (
);

FILL FILL_2__1437_ (
);

FILL FILL_2__1017_ (
);

FILL FILL_2__1190_ (
);

FILL FILL88350x54750 (
);

FILL FILL_3__1506_ (
);

OAI21X1 _1435_ (
    .A(_577_),
    .B(_575_),
    .C(_641_),
    .Y(_642_)
);

NAND3X1 _1015_ (
    .A(_137_),
    .B(_192_),
    .C(_197_),
    .Y(_206_)
);

FILL FILL_0__763_ (
);

AOI21X1 _766_ (
    .A(Cin_0_bF$buf1),
    .B(Xin[1]),
    .C(Yin[1]),
    .Y(_493_)
);

FILL FILL_1__1177_ (
);

FILL FILL_1__970_ (
);

FILL FILL_2__1246_ (
);

FILL FILL_0__819_ (
);

FILL FILL_3__1315_ (
);

OAI21X1 _1244_ (
    .A(_430_),
    .B(_431_),
    .C(_427_),
    .Y(_437_)
);

FILL FILL_0__992_ (
);

NAND3X1 _995_ (
    .A(_184_),
    .B(_185_),
    .C(_182_),
    .Y(_186_)
);

FILL FILL_2__813_ (
);

FILL FILL_2__1475_ (
);

FILL FILL_2__1055_ (
);

FILL FILL_3__1124_ (
);

XNOR2X1 _1473_ (
    .A(_682_),
    .B(Yin[13]),
    .Y(_683_)
);

NAND3X1 _1053_ (
    .A(_218_),
    .B(_241_),
    .C(_242_),
    .Y(_243_)
);

FILL FILL_1__835_ (
);

FILL FILL88950x35250 (
);

FILL FILL_0__1513_ (
);

FILL FILL_2__1284_ (
);

DFFPOSX1 _1529_ (
    .D(y[1]),
    .CLK(clk_bF$buf4),
    .Q(_755_[1])
);

OAI21X1 _1109_ (
    .A(_295_),
    .B(_296_),
    .C(_217_),
    .Y(_299_)
);

FILL FILL_0__857_ (
);

FILL FILL_3__1353_ (
);

NAND3X1 _1282_ (
    .A(_410_),
    .B(_469_),
    .C(_477_),
    .Y(_478_)
);

FILL FILL_4__788_ (
);

FILL FILL_0__1322_ (
);

FILL FILL_2__851_ (
);

FILL FILL_2__1093_ (
);

FILL FILL_3__1409_ (
);

NAND2X1 _1338_ (
    .A(_534_),
    .B(_538_),
    .Y(_539_)
);

FILL FILL_3__1582_ (
);

FILL FILL_3__1162_ (
);

NAND3X1 _1091_ (
    .A(_280_),
    .B(_246_),
    .C(_276_),
    .Y(_281_)
);

FILL FILL_1__873_ (
);

FILL FILL_2__907_ (
);

FILL FILL_2__1569_ (
);

FILL FILL_2__1149_ (
);

FILL FILL_0__1131_ (
);

FILL FILL_3__1218_ (
);

BUFX2 _1567_ (
    .A(_754_[7]),
    .Y(Xout[7])
);

NAND2X1 _1147_ (
    .A(Cin[3]),
    .B(Xin_5_bF$buf1),
    .Y(_336_)
);

FILL FILL_0__895_ (
);

FILL FILL_1__929_ (
);

FILL FILL_3__1391_ (
);

NAND3X1 _898_ (
    .A(Cin[2]),
    .B(Xin_3_bF$buf2),
    .C(_79_),
    .Y(_90_)
);

FILL FILL_4__1460_ (
);

FILL FILL_2__1378_ (
);

FILL FILL_0__1360_ (
);

FILL FILL_3__831_ (
);

FILL FILL_1__1101_ (
);

FILL FILL_3__1447_ (
);

FILL FILL_3__1027_ (
);

OAI21X1 _1376_ (
    .A(_577_),
    .B(_324_),
    .C(_578_),
    .Y(_579_)
);

FILL FILL_4__1516_ (
);

FILL FILL_0__1416_ (
);

FILL FILL_2__945_ (
);

FILL FILL_2__1187_ (
);

FILL FILL_1__1330_ (
);

FILL FILL_3__1256_ (
);

OAI21X1 _1185_ (
    .A(_373_),
    .B(_368_),
    .C(_347_),
    .Y(_374_)
);

FILL FILL_1__967_ (
);

FILL FILL_0__1225_ (
);

FILL FILL_4__903_ (
);

FILL FILL_0__989_ (
);

FILL FILL_3__1485_ (
);

FILL FILL_3__1065_ (
);

FILL FILL_1__776_ (
);

FILL FILL_0__1454_ (
);

FILL FILL_0__1034_ (
);

FILL FILL_2__983_ (
);

FILL FILL_3__925_ (
);

FILL FILL_0__798_ (
);

FILL FILL_3__1294_ (
);

FILL FILL_0__1263_ (
);

FILL FILL_2__792_ (
);

FILL FILL_1__1424_ (
);

FILL FILL_1__1004_ (
);

AOI21X1 _1279_ (
    .A(_473_),
    .B(_474_),
    .C(_465_),
    .Y(_475_)
);

FILL FILL_4__1419_ (
);

FILL FILL_0__1319_ (
);

FILL FILL_2__848_ (
);

FILL FILL_0__1492_ (
);

FILL FILL_0__1072_ (
);

FILL FILL_3__963_ (
);

NAND2X1 _822_ (
    .A(Xin[1]),
    .B(Cin[3]),
    .Y(_15_)
);

FILL FILL_1__1233_ (
);

FILL FILL_3__1579_ (
);

FILL FILL_3__1159_ (
);

FILL FILL88950x23550 (
);

OAI21X1 _1088_ (
    .A(_274_),
    .B(_273_),
    .C(_260_),
    .Y(_278_)
);

FILL FILL_2__1302_ (
);

FILL FILL_0__1128_ (
);

AOI21X1 _1300_ (
    .A(_410_),
    .B(_477_),
    .C(_496_),
    .Y(_497_)
);

FILL FILL_3__772_ (
);

FILL FILL_4__806_ (
);

FILL FILL_1__1462_ (
);

FILL FILL_1__1042_ (
);

FILL FILL_3__1388_ (
);

FILL FILL_2__1111_ (
);

FILL FILL_4__1037_ (
);

FILL FILL_0__1357_ (
);

FILL FILL_2__886_ (
);

FILL FILL_3__828_ (
);

FILL FILL_1__1518_ (
);

OAI21X1 _860_ (
    .A(_51_),
    .B(_740_),
    .C(_45_),
    .Y(_52_)
);

FILL FILL_1__1271_ (
);

FILL FILL_3__1197_ (
);

FILL FILL_2__1340_ (
);

FILL FILL_0__1166_ (
);

FILL FILL88350x19650 (
);

FILL FILL_0__913_ (
);

AOI21X1 _916_ (
    .A(_104_),
    .B(_103_),
    .C(_96_),
    .Y(_108_)
);

FILL FILL_1__1327_ (
);

FILL FILL_1__1080_ (
);

FILL FILL_0__1395_ (
);

FILL FILL_3__866_ (
);

FILL FILL_1__1136_ (
);

FILL FILL_2__1205_ (
);

AOI21X1 _1203_ (
    .A(_392_),
    .B(_387_),
    .C(_315_),
    .Y(_393_)
);

FILL FILL_0__951_ (
);

AOI21X1 _954_ (
    .A(_105_),
    .B(_102_),
    .C(_95_),
    .Y(_145_)
);

FILL FILL_1__1365_ (
);

FILL FILL_2__1434_ (
);

FILL FILL_2__1014_ (
);

FILL FILL_2__789_ (
);

FILL FILL88650x58650 (
);

FILL FILL_3__1503_ (
);

NAND2X1 _1432_ (
    .A(Cin[6]),
    .B(Xin[7]),
    .Y(_639_)
);

OAI21X1 _1012_ (
    .A(_202_),
    .B(_198_),
    .C(_127_),
    .Y(_203_)
);

FILL FILL_0__760_ (
);

NAND2X1 _763_ (
    .A(Xin[0]),
    .B(Cin[1]),
    .Y(_461_)
);

FILL FILL_1__1174_ (
);

FILL FILL_2__1243_ (
);

FILL FILL_0__1489_ (
);

FILL FILL_0__1069_ (
);

FILL FILL_0__816_ (
);

FILL FILL_3__1312_ (
);

AOI21X1 _819_ (
    .A(_4_),
    .B(_1_),
    .C(_0_),
    .Y(_12_)
);

NAND3X1 _1241_ (
    .A(_414_),
    .B(_428_),
    .C(_433_),
    .Y(_434_)
);

AND2X2 _992_ (
    .A(_157_),
    .B(_154_),
    .Y(_183_)
);

FILL FILL_2__810_ (
);

FILL FILL_2__1472_ (
);

FILL FILL_2__1052_ (
);

FILL FILL_0__1298_ (
);

FILL FILL_3__769_ (
);

FILL FILL_3__1121_ (
);

FILL FILL_1__1459_ (
);

FILL FILL_1__1039_ (
);

OAI21X1 _1470_ (
    .A(_352_),
    .B(_575_),
    .C(_639_),
    .Y(_680_)
);

NAND3X1 _1050_ (
    .A(_219_),
    .B(_234_),
    .C(_239_),
    .Y(_240_)
);

FILL FILL_1__832_ (
);

FILL FILL_4__976_ (
);

FILL FILL_0__1510_ (
);

FILL FILL_2__1108_ (
);

FILL FILL_2__1281_ (
);

DFFPOSX1 _1526_ (
    .D(Xin[6]),
    .CLK(clk_bF$buf3),
    .Q(_754_[6])
);

AOI21X1 _1106_ (
    .A(_281_),
    .B(_286_),
    .C(_244_),
    .Y(_296_)
);

FILL FILL_0__854_ (
);

FILL FILL_3__998_ (
);

FILL FILL_3__1350_ (
);

NAND3X1 _857_ (
    .A(_44_),
    .B(_48_),
    .C(_46_),
    .Y(_49_)
);

FILL FILL_1__1268_ (
);

FILL FILL_2__1337_ (
);

FILL FILL_2__1090_ (
);

FILL FILL_3__1406_ (
);

INVX1 _1335_ (
    .A(Yin[10]),
    .Y(_535_)
);

FILL FILL_1__1497_ (
);

FILL FILL_1__1077_ (
);

FILL FILL_1__870_ (
);

FILL FILL_2__904_ (
);

FILL FILL_2__1566_ (
);

FILL FILL_2__1146_ (
);

FILL FILL_3__1215_ (
);

BUFX2 _1564_ (
    .A(_754_[4]),
    .Y(Xout[4])
);

NAND3X1 _1144_ (
    .A(_332_),
    .B(_327_),
    .C(_330_),
    .Y(_333_)
);

FILL FILL_0__892_ (
);

FILL FILL_1__926_ (
);

INVX1 _895_ (
    .A(Xin_3_bF$buf1),
    .Y(_87_)
);

FILL FILL_2__1375_ (
);

FILL FILL_0__948_ (
);

FILL FILL_3__1444_ (
);

FILL FILL_3__1024_ (
);

FILL FILL_2_BUFX2_insert10 (
);

FILL FILL_2_BUFX2_insert11 (
);

FILL FILL_2_BUFX2_insert12 (
);

FILL FILL_2_BUFX2_insert13 (
);

FILL FILL_2_BUFX2_insert14 (
);

FILL FILL_2_BUFX2_insert15 (
);

FILL FILL_2_BUFX2_insert16 (
);

FILL FILL_2_BUFX2_insert17 (
);

NAND2X1 _1373_ (
    .A(Xin[6]),
    .B(Cin[6]),
    .Y(_576_)
);

FILL FILL_0__1413_ (
);

FILL FILL_2__942_ (
);

FILL FILL_2__1184_ (
);

INVX1 _1429_ (
    .A(_635_),
    .Y(_636_)
);

NAND3X1 _1009_ (
    .A(_195_),
    .B(_196_),
    .C(_139_),
    .Y(_200_)
);

FILL FILL_0__757_ (
);

FILL FILL_3__1253_ (
);

NAND2X1 _1182_ (
    .A(_362_),
    .B(_370_),
    .Y(_371_)
);

FILL FILL_1__964_ (
);

FILL FILL_4__1322_ (
);

FILL FILL_0__1222_ (
);

FILL FILL_3__1309_ (
);

NOR3X1 _1238_ (
    .A(_415_),
    .B(_416_),
    .C(_419_),
    .Y(_431_)
);

FILL FILL_0__986_ (
);

FILL FILL_3__1482_ (
);

FILL FILL_3__1062_ (
);

OAI21X1 _989_ (
    .A(_179_),
    .B(_176_),
    .C(_146_),
    .Y(_180_)
);

FILL FILL_1__773_ (
);

FILL FILL_2__807_ (
);

FILL FILL_4_CLKBUF1_insert4 (
);

FILL FILL_2__1469_ (
);

FILL FILL_0__1451_ (
);

FILL FILL_2__1049_ (
);

FILL FILL_0__1031_ (
);

FILL FILL_2__980_ (
);

FILL FILL_3__922_ (
);

FILL FILL_3__1118_ (
);

INVX1 _1467_ (
    .A(_576_),
    .Y(_677_)
);

NOR2X1 _1047_ (
    .A(_152_),
    .B(_231_),
    .Y(_237_)
);

FILL FILL_0__795_ (
);

FILL FILL_1__829_ (
);

FILL FILL_3__1291_ (
);

INVX1 _798_ (
    .A(_738_),
    .Y(_739_)
);

FILL FILL_0__1507_ (
);

FILL FILL_0__1260_ (
);

FILL FILL_2__1278_ (
);

FILL FILL_1__1421_ (
);

FILL FILL_1__1001_ (
);

FILL FILL_3__1347_ (
);

AOI21X1 _1276_ (
    .A(_382_),
    .B(_384_),
    .C(_470_),
    .Y(_471_)
);

FILL FILL_0__1316_ (
);

FILL FILL_2__845_ (
);

FILL FILL_2__1087_ (
);

FILL FILL_3__960_ (
);

FILL FILL_1__1230_ (
);

FILL FILL_3__1576_ (
);

FILL FILL_3__1156_ (
);

OAI21X1 _1085_ (
    .A(_274_),
    .B(_273_),
    .C(_272_),
    .Y(_275_)
);

FILL FILL_1__867_ (
);

FILL FILL_0__1125_ (
);

FILL FILL88950x85950 (
);

FILL FILL_0__889_ (
);

FILL FILL_3__1385_ (
);

FILL FILL_0__1354_ (
);

FILL FILL_2__883_ (
);

FILL FILL_3__825_ (
);

FILL FILL_1__1515_ (
);

FILL FILL_3__1194_ (
);

FILL FILL_2__939_ (
);

FILL FILL_0__1583_ (
);

FILL FILL_0__1163_ (
);

FILL FILL_0__910_ (
);

NAND3X1 _913_ (
    .A(_96_),
    .B(_103_),
    .C(_104_),
    .Y(_105_)
);

FILL FILL_1__1324_ (
);

AOI21X1 _1179_ (
    .A(_367_),
    .B(_365_),
    .C(_359_),
    .Y(_368_)
);

FILL FILL_0__1219_ (
);

FILL FILL_0__1392_ (
);

FILL FILL_3__863_ (
);

FILL FILL_1__1133_ (
);

FILL FILL_3__1479_ (
);

FILL FILL_3__1059_ (
);

FILL FILL_2__1202_ (
);

FILL FILL_0__1448_ (
);

FILL FILL_0__1028_ (
);

FILL FILL_2__977_ (
);

FILL FILL_3__919_ (
);

NAND3X1 _1200_ (
    .A(_383_),
    .B(_384_),
    .C(_382_),
    .Y(_390_)
);

FILL FILL89250x31350 (
);

AOI21X1 _951_ (
    .A(_78_),
    .B(_140_),
    .C(_141_),
    .Y(_142_)
);

FILL FILL_1__1362_ (
);

FILL FILL_3__1288_ (
);

FILL FILL_1__999_ (
);

FILL FILL_2__1431_ (
);

FILL FILL_2__1011_ (
);

FILL FILL_0__1257_ (
);

FILL FILL_2__786_ (
);

FILL FILL_3__1500_ (
);

FILL FILL_1__1418_ (
);

FILL FILL_4__935_ (
);

INVX1 _760_ (
    .A(_418_),
    .Y(_429_)
);

FILL FILL_1__1171_ (
);

FILL FILL_3__1097_ (
);

FILL FILL_2__1240_ (
);

FILL FILL_4__1166_ (
);

FILL FILL_0__1486_ (
);

FILL FILL_0__1066_ (
);

FILL FILL_0__813_ (
);

FILL FILL_3__957_ (
);

NAND3X1 _816_ (
    .A(_746_),
    .B(_5_),
    .C(_8_),
    .Y(_9_)
);

FILL FILL_1__1227_ (
);

FILL FILL_0__1295_ (
);

FILL FILL_3__766_ (
);

FILL FILL_1__1456_ (
);

FILL FILL_1__1036_ (
);

FILL FILL_2__1105_ (
);

DFFPOSX1 _1523_ (
    .D(Xin_3_bF$buf1),
    .CLK(clk_bF$buf4),
    .Q(_754_[3])
);

INVX1 _1103_ (
    .A(_189_),
    .Y(_293_)
);

FILL FILL_0__851_ (
);

FILL FILL_3__995_ (
);

NAND2X1 _854_ (
    .A(_743_),
    .B(_45_),
    .Y(_46_)
);

FILL FILL_1__1265_ (
);

FILL FILL_2__1334_ (
);

FILL FILL_0__907_ (
);

FILL FILL_3__1403_ (
);

AND2X2 _1332_ (
    .A(Cin[4]),
    .B(Xin[7]),
    .Y(_532_)
);

FILL FILL_4__838_ (
);

FILL FILL_1__1494_ (
);

FILL FILL_1__1074_ (
);

FILL FILL_2__901_ (
);

FILL FILL_2__1563_ (
);

FILL FILL_2__1143_ (
);

FILL FILL_4__1069_ (
);

FILL FILL_0__1389_ (
);

FILL FILL_3__1212_ (
);

BUFX2 _1561_ (
    .A(_754_[1]),
    .Y(Xout[1])
);

NAND3X1 _1141_ (
    .A(_319_),
    .B(_328_),
    .C(_329_),
    .Y(_330_)
);

FILL FILL_1__923_ (
);

INVX1 _892_ (
    .A(_83_),
    .Y(_84_)
);

FILL FILL_2__1372_ (
);

FILL FILL_0__1198_ (
);

FILL FILL_0__945_ (
);

FILL FILL_3__1441_ (
);

FILL FILL_3__1021_ (
);

OAI21X1 _948_ (
    .A(_123_),
    .B(_138_),
    .C(_116_),
    .Y(_139_)
);

FILL FILL_1__1359_ (
);

OAI21X1 _1370_ (
    .A(_528_),
    .B(_540_),
    .C(_572_),
    .Y(_573_)
);

FILL FILL_2__1428_ (
);

FILL FILL_0__1410_ (
);

FILL FILL_2__1008_ (
);

FILL FILL_2__1181_ (
);

NAND2X1 _1426_ (
    .A(_618_),
    .B(_631_),
    .Y(_632_)
);

NAND3X1 _1006_ (
    .A(_195_),
    .B(_196_),
    .C(_194_),
    .Y(_197_)
);

FILL FILL_3__898_ (
);

FILL FILL_3__1250_ (
);

INVX1 _757_ (
    .A(Xin[0]),
    .Y(_397_)
);

FILL FILL_1__1168_ (
);

FILL FILL_1__961_ (
);

FILL FILL_2__1237_ (
);

FILL FILL_3__1306_ (
);

OAI21X1 _1235_ (
    .A(_348_),
    .B(_426_),
    .C(_351_),
    .Y(_427_)
);

FILL FILL_0__983_ (
);

NAND3X1 _986_ (
    .A(_160_),
    .B(_173_),
    .C(_174_),
    .Y(_177_)
);

FILL FILL_1__1397_ (
);

FILL FILL_1__770_ (
);

FILL FILL_2__804_ (
);

FILL FILL_2__1466_ (
);

FILL FILL_2__1046_ (
);

FILL FILL_3__1115_ (
);

OAI21X1 _1464_ (
    .A(_671_),
    .B(_672_),
    .C(_670_),
    .Y(_673_)
);

NAND3X1 _1044_ (
    .A(_226_),
    .B(_230_),
    .C(_233_),
    .Y(_234_)
);

FILL FILL_0__792_ (
);

FILL FILL_1__826_ (
);

AOI21X1 _795_ (
    .A(_731_),
    .B(_734_),
    .C(_559_),
    .Y(_737_)
);

FILL FILL_0__1504_ (
);

FILL FILL_2__1275_ (
);

FILL FILL_0__848_ (
);

FILL FILL_3__1344_ (
);

OAI21X1 _1273_ (
    .A(_467_),
    .B(_466_),
    .C(_465_),
    .Y(_468_)
);

FILL FILL_0__1313_ (
);

FILL FILL_2__842_ (
);

FILL FILL_2__1084_ (
);

NAND2X1 _1329_ (
    .A(Yin[9]),
    .B(_363_),
    .Y(_529_)
);

FILL FILL_3__1573_ (
);

FILL FILL_3__1153_ (
);

INVX1 _1082_ (
    .A(_260_),
    .Y(_272_)
);

FILL FILL_1__864_ (
);

FILL FILL_0__1122_ (
);

FILL FILL_3__1209_ (
);

DFFPOSX1 _1558_ (
    .D(_753_[14]),
    .CLK(clk_bF$buf2),
    .Q(y[14])
);

NAND3X1 _1138_ (
    .A(_326_),
    .B(_320_),
    .C(_323_),
    .Y(_327_)
);

FILL FILL_0__886_ (
);

FILL FILL_3__1382_ (
);

XOR2X1 _889_ (
    .A(_80_),
    .B(_78_),
    .Y(_81_)
);

FILL FILL_4__1451_ (
);

FILL FILL_0__1351_ (
);

FILL FILL_2__1369_ (
);

FILL FILL_2__880_ (
);

FILL FILL_3__822_ (
);

FILL FILL_1__1512_ (
);

FILL FILL_3__1438_ (
);

FILL FILL_3__1018_ (
);

NAND2X1 _1367_ (
    .A(_516_),
    .B(_522_),
    .Y(_570_)
);

FILL FILL_3__1191_ (
);

FILL FILL_4__1507_ (
);

FILL FILL_0__1407_ (
);

FILL FILL_2__936_ (
);

FILL FILL_0__1580_ (
);

FILL FILL_2__1178_ (
);

FILL FILL_0__1160_ (
);

NAND3X1 _910_ (
    .A(_98_),
    .B(_97_),
    .C(_101_),
    .Y(_102_)
);

FILL FILL_1__1321_ (
);

FILL FILL_3__1247_ (
);

OAI21X1 _1176_ (
    .A(_363_),
    .B(_364_),
    .C(_361_),
    .Y(_365_)
);

FILL FILL_1__958_ (
);

FILL FILL_0__1216_ (
);

FILL FILL_3__860_ (
);

FILL FILL_1__1130_ (
);

FILL FILL_3__1476_ (
);

FILL FILL_3__1056_ (
);

FILL FILL_1__767_ (
);

FILL FILL_0__1445_ (
);

FILL FILL_0__1025_ (
);

FILL FILL_2__974_ (
);

FILL FILL_3__916_ (
);

FILL FILL89550x35250 (
);

FILL FILL_0__789_ (
);

FILL FILL_3__1285_ (
);

FILL FILL_1__996_ (
);

FILL FILL_0__1254_ (
);

FILL FILL_2__783_ (
);

FILL FILL_1__1415_ (
);

FILL FILL_3__1094_ (
);

FILL FILL_2__839_ (
);

FILL FILL_4__1583_ (
);

FILL FILL_0__1483_ (
);

FILL FILL_0__1063_ (
);

FILL FILL_0__810_ (
);

FILL FILL_3__954_ (
);

NAND2X1 _813_ (
    .A(Yin[3]),
    .B(_3_),
    .Y(_6_)
);

FILL FILL_1__1224_ (
);

NAND2X1 _1499_ (
    .A(_709_),
    .B(_710_),
    .Y(_711_)
);

NAND3X1 _1079_ (
    .A(Cin_0_bF$buf0),
    .B(Xin[7]),
    .C(_264_),
    .Y(_269_)
);

FILL FILL_0__1119_ (
);

FILL FILL_0__1292_ (
);

FILL FILL_3__763_ (
);

FILL FILL_1__1453_ (
);

FILL FILL_1__1033_ (
);

FILL FILL_3__1379_ (
);

FILL FILL_2__1102_ (
);

FILL FILL_4__1028_ (
);

FILL FILL_0__1348_ (
);

FILL FILL_2__877_ (
);

FILL FILL_3__819_ (
);

FILL FILL_1__1509_ (
);

DFFPOSX1 _1520_ (
    .D(Xin[0]),
    .CLK(clk_bF$buf1),
    .Q(_754_[0])
);

NAND3X1 _1100_ (
    .A(_276_),
    .B(_280_),
    .C(_283_),
    .Y(_290_)
);

FILL FILL_3__992_ (
);

NAND3X1 _851_ (
    .A(_42_),
    .B(_41_),
    .C(_40_),
    .Y(_43_)
);

FILL FILL_1__1262_ (
);

FILL FILL_3__1188_ (
);

FILL FILL_1__899_ (
);

FILL FILL_2__1331_ (
);

FILL FILL_0__1577_ (
);

FILL FILL_0__1157_ (
);

FILL FILL_0__904_ (
);

FILL FILL_3__1400_ (
);

INVX1 _907_ (
    .A(Yin[5]),
    .Y(_99_)
);

FILL FILL_1__1318_ (
);

FILL FILL_1__1491_ (
);

FILL FILL_1__1071_ (
);

FILL FILL_2__1560_ (
);

FILL FILL_2__1140_ (
);

FILL FILL_0__1386_ (
);

FILL FILL_3__857_ (
);

FILL FILL_1__1127_ (
);

FILL FILL_1__920_ (
);

FILL FILL_4__1295_ (
);

FILL FILL_0__1195_ (
);

FILL FILL_0__942_ (
);

OAI21X1 _945_ (
    .A(_73_),
    .B(_133_),
    .C(_132_),
    .Y(_136_)
);

FILL FILL_1__1356_ (
);

FILL FILL_2__1425_ (
);

FILL FILL_2__1005_ (
);

INVX1 _1423_ (
    .A(_565_),
    .Y(_629_)
);

AOI21X1 _1003_ (
    .A(_81_),
    .B(_120_),
    .C(_193_),
    .Y(_194_)
);

FILL FILL_3__895_ (
);

FILL FILL_1__1165_ (
);

FILL FILL_2__1234_ (
);

FILL FILL_0__807_ (
);

FILL FILL_3__1303_ (
);

FILL FILL89550x23550 (
);

NAND2X1 _1232_ (
    .A(_322_),
    .B(_423_),
    .Y(_424_)
);

FILL FILL_0__980_ (
);

NAND3X1 _983_ (
    .A(_161_),
    .B(_163_),
    .C(_165_),
    .Y(_174_)
);

FILL FILL_1__1394_ (
);

FILL FILL_2__801_ (
);

FILL FILL_2__1463_ (
);

FILL FILL_2__1043_ (
);

FILL FILL_0__1289_ (
);

FILL FILL_3__1112_ (
);

NAND2X1 _1461_ (
    .A(_670_),
    .B(_668_),
    .Y(_671_)
);

NAND2X1 _1041_ (
    .A(Cin[2]),
    .B(Xin[4]),
    .Y(_231_)
);

FILL FILL_1__823_ (
);

FILL FILL_4__967_ (
);

OAI21X1 _792_ (
    .A(_718_),
    .B(_733_),
    .C(_732_),
    .Y(_734_)
);

FILL FILL_2__1519_ (
);

FILL FILL_0__1501_ (
);

FILL FILL_2__1272_ (
);

FILL FILL_4__1198_ (
);

FILL FILL_0__1098_ (
);

NAND2X1 _1517_ (
    .A(_728_),
    .B(_722_),
    .Y(_753_[15])
);

FILL FILL_0__845_ (
);

FILL FILL_3__989_ (
);

FILL FILL_3__1341_ (
);

AOI21X1 _848_ (
    .A(_0_),
    .B(_4_),
    .C(_39_),
    .Y(_40_)
);

FILL FILL_1__1259_ (
);

NAND2X1 _1270_ (
    .A(_434_),
    .B(_438_),
    .Y(_465_)
);

FILL FILL_4__1410_ (
);

FILL FILL_0__1310_ (
);

FILL FILL_2__1328_ (
);

FILL FILL_2__1081_ (
);

OAI21X1 _1326_ (
    .A(_517_),
    .B(_518_),
    .C(_514_),
    .Y(_525_)
);

FILL FILL_3__798_ (
);

FILL FILL_3__1570_ (
);

FILL FILL_3__1150_ (
);

FILL FILL_1__1488_ (
);

FILL FILL_1__1068_ (
);

FILL FILL_1__861_ (
);

FILL FILL_2__1137_ (
);

FILL FILL_3__1206_ (
);

DFFPOSX1 _1555_ (
    .D(_753_[11]),
    .CLK(clk_bF$buf5),
    .Q(y[11])
);

INVX1 _1135_ (
    .A(Cin[6]),
    .Y(_324_)
);

FILL FILL_0__883_ (
);

FILL FILL_1__917_ (
);

NOR2X1 _886_ (
    .A(_397_),
    .B(_77_),
    .Y(_78_)
);

FILL FILL_1__1297_ (
);

FILL FILL_2_CLKBUF1_insert0 (
);

FILL FILL_2_CLKBUF1_insert1 (
);

FILL FILL_2_CLKBUF1_insert2 (
);

FILL FILL_2_CLKBUF1_insert3 (
);

FILL FILL_2_CLKBUF1_insert4 (
);

FILL FILL_2_CLKBUF1_insert5 (
);

FILL FILL_2__1366_ (
);

FILL FILL_0__939_ (
);

FILL FILL_3__1435_ (
);

FILL FILL_3__1015_ (
);

OAI21X1 _1364_ (
    .A(_565_),
    .B(_495_),
    .C(_564_),
    .Y(_566_)
);

FILL FILL_0__1404_ (
);

FILL FILL89250x58650 (
);

FILL FILL_2__933_ (
);

FILL FILL_2__1175_ (
);

FILL FILL_3__1244_ (
);

NAND3X1 _1173_ (
    .A(Cin[1]),
    .B(Xin[7]),
    .C(Yin[8]),
    .Y(_362_)
);

FILL FILL_1__955_ (
);

FILL FILL_4__1313_ (
);

FILL FILL_0__1213_ (
);

INVX1 _1229_ (
    .A(_415_),
    .Y(_421_)
);

FILL FILL_0__977_ (
);

FILL FILL_3__1473_ (
);

FILL FILL_3__1053_ (
);

FILL FILL_1__764_ (
);

FILL FILL_0__1442_ (
);

FILL FILL_0__1022_ (
);

FILL FILL_2__971_ (
);

FILL FILL_3__913_ (
);

FILL FILL_3__1109_ (
);

NAND3X1 _1458_ (
    .A(_615_),
    .B(_621_),
    .C(_667_),
    .Y(_668_)
);

NAND2X1 _1038_ (
    .A(_227_),
    .B(_140_),
    .Y(_228_)
);

FILL FILL_0__786_ (
);

FILL FILL_3__1282_ (
);

NAND3X1 _789_ (
    .A(_601_),
    .B(_708_),
    .C(_729_),
    .Y(_731_)
);

FILL FILL_1__993_ (
);

FILL FILL_0__1251_ (
);

FILL FILL_2__1269_ (
);

FILL FILL_2__780_ (
);

FILL FILL89550x11850 (
);

FILL FILL_1__1412_ (
);

FILL FILL_3__1338_ (
);

NAND2X1 _1267_ (
    .A(_454_),
    .B(_457_),
    .Y(_462_)
);

FILL FILL_3__1091_ (
);

FILL FILL_0__1307_ (
);

FILL FILL_2__836_ (
);

FILL FILL_2__1498_ (
);

FILL FILL_0__1480_ (
);

FILL FILL_2__1078_ (
);

FILL FILL_0__1060_ (
);

FILL FILL_3__951_ (
);

NAND2X1 _810_ (
    .A(Cin_0_bF$buf2),
    .B(Xin_3_bF$buf0),
    .Y(_3_)
);

FILL FILL_1__1221_ (
);

FILL FILL_3__1567_ (
);

FILL FILL_3__1147_ (
);

NAND2X1 _1496_ (
    .A(_703_),
    .B(_706_),
    .Y(_707_)
);

NAND2X1 _1076_ (
    .A(_264_),
    .B(_265_),
    .Y(_266_)
);

FILL FILL_1__858_ (
);

FILL FILL_4__1216_ (
);

FILL FILL_0__1116_ (
);

FILL FILL_3__760_ (
);

FILL FILL_1__1450_ (
);

FILL FILL_1__1030_ (
);

FILL FILL_3__1376_ (
);

FILL FILL_0__1345_ (
);

FILL FILL_2__874_ (
);

FILL FILL_3__816_ (
);

FILL FILL_1__1506_ (
);

FILL FILL_3__1185_ (
);

FILL FILL_1__896_ (
);

FILL FILL_0__1574_ (
);

FILL FILL_0__1154_ (
);

FILL FILL_0__901_ (
);

NAND2X1 _904_ (
    .A(Cin[1]),
    .B(Xin[4]),
    .Y(_96_)
);

FILL FILL_1__1315_ (
);

FILL FILL_0__1383_ (
);

FILL FILL_3__854_ (
);

FILL FILL_1__1124_ (
);

NAND3X1 _1399_ (
    .A(_593_),
    .B(_597_),
    .C(_603_),
    .Y(_604_)
);

FILL FILL_0__1439_ (
);

FILL FILL_0__1019_ (
);

FILL FILL_2__968_ (
);

FILL FILL_0__1192_ (
);

INVX1 _942_ (
    .A(_133_),
    .Y(_134_)
);

FILL FILL_1__1353_ (
);

FILL FILL_3__1279_ (
);

FILL FILL_2__1422_ (
);

FILL FILL_2__1002_ (
);

FILL FILL_0__1248_ (
);

FILL FILL_2__777_ (
);

FILL FILL_1__1409_ (
);

XOR2X1 _1420_ (
    .A(_566_),
    .B(_626_),
    .Y(_753_[11])
);

AOI21X1 _1000_ (
    .A(_190_),
    .B(_189_),
    .C(_188_),
    .Y(_191_)
);

FILL FILL_3__892_ (
);

FILL FILL_4__926_ (
);

FILL FILL_1__1582_ (
);

FILL FILL_1__1162_ (
);

FILL FILL_3__1088_ (
);

FILL FILL_1__799_ (
);

FILL FILL_2__1231_ (
);

FILL FILL_4__1157_ (
);

FILL FILL_0__1477_ (
);

FILL FILL_0__1057_ (
);

FILL FILL_0__804_ (
);

FILL FILL_3__948_ (
);

FILL FILL_3__1300_ (
);

INVX1 _807_ (
    .A(_747_),
    .Y(_0_)
);

FILL FILL_1__1218_ (
);

OAI21X1 _980_ (
    .A(_170_),
    .B(_166_),
    .C(_160_),
    .Y(_171_)
);

FILL FILL_1__1391_ (
);

FILL FILL89550x85950 (
);

FILL FILL_2__1460_ (
);

FILL FILL_2__1040_ (
);

FILL FILL_0__1286_ (
);

FILL FILL_3__757_ (
);

FILL FILL_1__1447_ (
);

FILL FILL_1__1027_ (
);

FILL FILL_1__820_ (
);

FILL FILL_2__1516_ (
);

FILL FILL_0__1095_ (
);

OAI21X1 _1514_ (
    .A(_725_),
    .B(_724_),
    .C(_713_),
    .Y(_726_)
);

FILL FILL_0__842_ (
);

FILL FILL_3__986_ (
);

OAI21X1 _845_ (
    .A(_31_),
    .B(_36_),
    .C(_33_),
    .Y(_37_)
);

FILL FILL_1__1256_ (
);

FILL FILL_2__1325_ (
);

NAND3X1 _1323_ (
    .A(_501_),
    .B(_516_),
    .C(_521_),
    .Y(_522_)
);

FILL FILL_3__795_ (
);

FILL FILL_4__829_ (
);

FILL FILL_1__1485_ (
);

FILL FILL_1__1065_ (
);

FILL FILL_2__1134_ (
);

FILL FILL_3__1203_ (
);

DFFPOSX1 _1552_ (
    .D(_753_[8]),
    .CLK(clk_bF$buf1),
    .Q(y[8])
);

AND2X2 _1132_ (
    .A(Xin[2]),
    .B(Cin[6]),
    .Y(_321_)
);

FILL FILL_0__880_ (
);

FILL FILL_1__914_ (
);

INVX1 _883_ (
    .A(_74_),
    .Y(_75_)
);

FILL FILL_1__1294_ (
);

FILL FILL_2__1363_ (
);

FILL FILL_0__1189_ (
);

FILL FILL_0__936_ (
);

FILL FILL_3__1432_ (
);

FILL FILL_3__1012_ (
);

OAI21X1 _939_ (
    .A(_129_),
    .B(_130_),
    .C(_128_),
    .Y(_131_)
);

NAND3X1 _1361_ (
    .A(_562_),
    .B(_563_),
    .C(_561_),
    .Y(_564_)
);

FILL FILL_2__1419_ (
);

FILL FILL_0__1401_ (
);

FILL FILL_2__930_ (
);

FILL FILL_2__1172_ (
);

NAND3X1 _1417_ (
    .A(_620_),
    .B(_621_),
    .C(_622_),
    .Y(_624_)
);

FILL FILL_3__889_ (
);

FILL FILL_3__1241_ (
);

FILL FILL_1__1579_ (
);

FILL FILL_1__1159_ (
);

NAND2X1 _1170_ (
    .A(_358_),
    .B(_354_),
    .Y(_359_)
);

FILL FILL_1__952_ (
);

FILL FILL_0__1210_ (
);

FILL FILL_2__1228_ (
);

NAND2X1 _1226_ (
    .A(Xin[4]),
    .B(Cin[6]),
    .Y(_417_)
);

FILL FILL_0__974_ (
);

FILL FILL_3__1470_ (
);

FILL FILL_3__1050_ (
);

NAND3X1 _977_ (
    .A(Cin_0_bF$buf3),
    .B(Xin[6]),
    .C(Yin[6]),
    .Y(_168_)
);

FILL FILL_1__1388_ (
);

FILL FILL_1__761_ (
);

FILL FILL_2__1457_ (
);

FILL FILL_2__1037_ (
);

FILL FILL_3__910_ (
);

FILL FILL_3__1106_ (
);

OR2X2 _1455_ (
    .A(_659_),
    .B(_637_),
    .Y(_664_)
);

OAI21X1 _1035_ (
    .A(_47_),
    .B(_77_),
    .C(_224_),
    .Y(_225_)
);

FILL FILL_0__783_ (
);

FILL FILL_1__817_ (
);

NAND3X1 _786_ (
    .A(_612_),
    .B(_676_),
    .C(_697_),
    .Y(_708_)
);

FILL FILL_1__1197_ (
);

FILL FILL_1__990_ (
);

FILL FILL_2__1266_ (
);

FILL FILL_0__839_ (
);

FILL FILL_3__1335_ (
);

NAND3X1 _1264_ (
    .A(_454_),
    .B(_457_),
    .C(_442_),
    .Y(_458_)
);

FILL FILL_0__1304_ (
);

FILL FILL_2__833_ (
);

FILL FILL_2__1495_ (
);

FILL FILL_2__1075_ (
);

FILL FILL_3__1564_ (
);

FILL FILL_3__1144_ (
);

INVX1 _1493_ (
    .A(Yin[14]),
    .Y(_704_)
);

NAND3X1 _1073_ (
    .A(Cin_0_bF$buf0),
    .B(Xin[7]),
    .C(Yin[7]),
    .Y(_263_)
);

FILL FILL_1__855_ (
);

FILL FILL_4__999_ (
);

FILL FILL_0__1113_ (
);

DFFPOSX1 _1549_ (
    .D(_753_[5]),
    .CLK(clk_bF$buf3),
    .Q(y[5])
);

OAI21X1 _1129_ (
    .A(_224_),
    .B(_227_),
    .C(_226_),
    .Y(_318_)
);

FILL FILL_0__877_ (
);

FILL FILL_3__1373_ (
);

FILL FILL_4__1442_ (
);

FILL FILL_0__1342_ (
);

FILL FILL_2__871_ (
);

FILL FILL_3__813_ (
);

FILL FILL_1__1503_ (
);

FILL FILL_3__1429_ (
);

FILL FILL_3__1009_ (
);

OAI21X1 _1358_ (
    .A(_479_),
    .B(_560_),
    .C(_469_),
    .Y(_561_)
);

FILL FILL_3__1182_ (
);

FILL FILL_1__893_ (
);

FILL FILL_2__927_ (
);

FILL FILL_0__1571_ (
);

FILL FILL_0__1151_ (
);

FILL FILL_2__1169_ (
);

NAND3X1 _901_ (
    .A(_83_),
    .B(_90_),
    .C(_92_),
    .Y(_93_)
);

FILL FILL_1__1312_ (
);

FILL FILL_3__1238_ (
);

NAND3X1 _1167_ (
    .A(Cin[3]),
    .B(Xin_5_bF$buf1),
    .C(_355_),
    .Y(_356_)
);

FILL FILL_1__949_ (
);

FILL FILL_0__1207_ (
);

FILL FILL_4__1060_ (
);

FILL FILL_0__1380_ (
);

FILL FILL_2__1398_ (
);

FILL FILL_3__851_ (
);

FILL FILL_1__1121_ (
);

FILL FILL_3__1467_ (
);

FILL FILL_3__1047_ (
);

OR2X2 _1396_ (
    .A(_534_),
    .B(_598_),
    .Y(_600_)
);

FILL FILL_1__758_ (
);

FILL FILL_0__1436_ (
);

FILL FILL_0__1016_ (
);

FILL FILL_2__965_ (
);

FILL FILL_3__907_ (
);

FILL FILL_1__1350_ (
);

FILL FILL_3__1276_ (
);

FILL FILL_1__987_ (
);

FILL FILL_4__1345_ (
);

FILL FILL_0__1245_ (
);

FILL FILL_2__774_ (
);

FILL FILL_1__1406_ (
);

FILL FILL_3__1085_ (
);

FILL FILL_1__796_ (
);

FILL FILL_4__1574_ (
);

FILL FILL_0__1474_ (
);

FILL FILL_0__1054_ (
);

FILL FILL_0__801_ (
);

FILL FILL_3__945_ (
);

AND2X2 _804_ (
    .A(_744_),
    .B(_742_),
    .Y(_745_)
);

FILL FILL_1__1215_ (
);

FILL FILL_0__1283_ (
);

FILL FILL_1__1444_ (
);

FILL FILL_1__1024_ (
);

NOR3X1 _1299_ (
    .A(_475_),
    .B(_476_),
    .C(_471_),
    .Y(_496_)
);

FILL FILL_2__1513_ (
);

FILL FILL_0__1339_ (
);

FILL FILL_2__868_ (
);

FILL FILL_0__1092_ (
);

AOI22X1 _1511_ (
    .A(_618_),
    .B(_631_),
    .C(_627_),
    .D(_492_),
    .Y(_723_)
);

FILL FILL_3__983_ (
);

INVX1 _842_ (
    .A(_33_),
    .Y(_34_)
);

FILL FILL_1__1253_ (
);

FILL FILL_3__1179_ (
);

FILL FILL_2__1322_ (
);

FILL FILL_0__1568_ (
);

FILL FILL_0__1148_ (
);

FILL FILL_1__1309_ (
);

AND2X2 _1320_ (
    .A(_350_),
    .B(_445_),
    .Y(_519_)
);

FILL FILL_3__792_ (
);

FILL FILL_1__1482_ (
);

FILL FILL_1__1062_ (
);

FILL FILL_2__1131_ (
);

FILL FILL_0__1377_ (
);

FILL FILL_3__848_ (
);

FILL FILL_3__1200_ (
);

FILL FILL_1__1118_ (
);

FILL FILL_1__911_ (
);

AND2X2 _880_ (
    .A(_71_),
    .B(_68_),
    .Y(_72_)
);

FILL FILL_1__1291_ (
);

FILL FILL_2__1360_ (
);

FILL FILL_0__1186_ (
);

FILL FILL_0__933_ (
);

AOI21X1 _936_ (
    .A(_67_),
    .B(_26_),
    .C(_69_),
    .Y(_128_)
);

FILL FILL_1__1347_ (
);

FILL FILL_2__1416_ (
);

OAI21X1 _1414_ (
    .A(_499_),
    .B(_619_),
    .C(_555_),
    .Y(_620_)
);

FILL FILL_3__886_ (
);

FILL FILL_4_BUFX2_insert13 (
);

FILL FILL_4_BUFX2_insert17 (
);

FILL FILL_1__1576_ (
);

FILL FILL_1__1156_ (
);

FILL FILL_2__1225_ (
);

OAI21X1 _1223_ (
    .A(_227_),
    .B(_413_),
    .C(_327_),
    .Y(_414_)
);

FILL FILL_0__971_ (
);

NAND3X1 _974_ (
    .A(Cin_0_bF$buf3),
    .B(Xin[6]),
    .C(_164_),
    .Y(_165_)
);

FILL FILL_1__1385_ (
);

FILL FILL_2__1454_ (
);

FILL FILL_2__1034_ (
);

FILL FILL_3__1103_ (
);

INVX1 _1452_ (
    .A(_660_),
    .Y(_661_)
);

AND2X2 _1032_ (
    .A(Xin[2]),
    .B(Cin[5]),
    .Y(_222_)
);

FILL FILL_0__780_ (
);

FILL FILL_1__814_ (
);

FILL FILL_0_CLKBUF1_insert0 (
);

FILL FILL_0_CLKBUF1_insert1 (
);

FILL FILL_0_CLKBUF1_insert2 (
);

FILL FILL_0_CLKBUF1_insert3 (
);

FILL FILL_4__958_ (
);

FILL FILL_0_CLKBUF1_insert4 (
);

FILL FILL_0_CLKBUF1_insert5 (
);

NAND3X1 _783_ (
    .A(_633_),
    .B(_644_),
    .C(_666_),
    .Y(_676_)
);

FILL FILL_1__1194_ (
);

FILL FILL_2__1263_ (
);

FILL FILL_4__1189_ (
);

FILL FILL_0__1089_ (
);

XNOR2X1 _1508_ (
    .A(_719_),
    .B(Yin[15]),
    .Y(_720_)
);

FILL FILL_0__836_ (
);

FILL FILL_3__1332_ (
);

AOI21X1 _839_ (
    .A(Cin_0_bF$buf2),
    .B(Xin[4]),
    .C(Yin[4]),
    .Y(_31_)
);

NAND2X1 _1261_ (
    .A(_449_),
    .B(_452_),
    .Y(_455_)
);

FILL FILL_4__1401_ (
);

FILL FILL_0__1301_ (
);

FILL FILL_2__1319_ (
);

FILL FILL_2__830_ (
);

FILL FILL_2__1492_ (
);

FILL FILL_2__1072_ (
);

NAND3X1 _1317_ (
    .A(_507_),
    .B(_512_),
    .C(_514_),
    .Y(_516_)
);

FILL FILL_3__789_ (
);

FILL FILL_3__1561_ (
);

FILL FILL_3__1141_ (
);

FILL FILL_1__1479_ (
);

FILL FILL_1__1059_ (
);

INVX1 _1490_ (
    .A(_692_),
    .Y(_701_)
);

OAI21X1 _1070_ (
    .A(_161_),
    .B(_259_),
    .C(_168_),
    .Y(_260_)
);

FILL FILL_1__852_ (
);

FILL FILL_0__1110_ (
);

FILL FILL_2__1128_ (
);

DFFPOSX1 _1546_ (
    .D(_750_[2]),
    .CLK(clk_bF$buf4),
    .Q(y[2])
);

INVX1 _1126_ (
    .A(_314_),
    .Y(_315_)
);

FILL FILL_0__874_ (
);

FILL FILL_1__908_ (
);

FILL FILL_3__1370_ (
);

AOI22X1 _877_ (
    .A(_9_),
    .B(_14_),
    .C(_65_),
    .D(_66_),
    .Y(_69_)
);

FILL FILL_1__1288_ (
);

FILL FILL_2__1357_ (
);

FILL FILL_3__810_ (
);

FILL FILL88050x78150 (
);

FILL FILL_1__1500_ (
);

FILL FILL_3__1426_ (
);

FILL FILL_3__1006_ (
);

AOI21X1 _1355_ (
    .A(_556_),
    .B(_555_),
    .C(_498_),
    .Y(_557_)
);

FILL FILL_1__1097_ (
);

FILL FILL_1__890_ (
);

FILL FILL_2__924_ (
);

FILL FILL_2__1166_ (
);

FILL FILL_3__1235_ (
);

OAI21X1 _1164_ (
    .A(_590_),
    .B(_352_),
    .C(_336_),
    .Y(_353_)
);

FILL FILL_1__946_ (
);

FILL FILL_4__1304_ (
);

FILL FILL_0__1204_ (
);

FILL FILL_2__1395_ (
);

FILL FILL_0__968_ (
);

FILL FILL_3__1464_ (
);

FILL FILL_3__1044_ (
);

NAND3X1 _1393_ (
    .A(_594_),
    .B(_595_),
    .C(_596_),
    .Y(_597_)
);

FILL FILL_0__1433_ (
);

FILL FILL_0__1013_ (
);

FILL FILL_2__962_ (
);

FILL FILL_3__904_ (
);

OAI21X1 _1449_ (
    .A(_648_),
    .B(_647_),
    .C(_654_),
    .Y(_658_)
);

INVX1 _1029_ (
    .A(_218_),
    .Y(_219_)
);

FILL FILL_0__777_ (
);

FILL FILL_3__1273_ (
);

FILL FILL_1__984_ (
);

FILL FILL_0__1242_ (
);

FILL FILL_2__771_ (
);

FILL FILL_1__1403_ (
);

FILL FILL_3__1329_ (
);

NAND3X1 _1258_ (
    .A(_443_),
    .B(_450_),
    .C(_451_),
    .Y(_452_)
);

FILL FILL_3__1082_ (
);

FILL FILL_1__793_ (
);

FILL FILL_2__827_ (
);

FILL FILL_0__1471_ (
);

FILL FILL_2__1489_ (
);

FILL FILL_2__1069_ (
);

FILL FILL_0__1051_ (
);

FILL FILL_3__942_ (
);

OAI21X1 _801_ (
    .A(_397_),
    .B(_740_),
    .C(_741_),
    .Y(_742_)
);

FILL FILL_1__1212_ (
);

FILL FILL_3__1138_ (
);

INVX1 _1487_ (
    .A(_696_),
    .Y(_698_)
);

NAND3X1 _1067_ (
    .A(_247_),
    .B(_255_),
    .C(_256_),
    .Y(_257_)
);

FILL FILL_1__849_ (
);

FILL FILL_4__1207_ (
);

FILL FILL_0__1107_ (
);

FILL FILL_2__1298_ (
);

FILL FILL_0__1280_ (
);

FILL FILL_1__1441_ (
);

FILL FILL_1__1021_ (
);

FILL FILL_3__1367_ (
);

OAI21X1 _1296_ (
    .A(_403_),
    .B(_491_),
    .C(_484_),
    .Y(_492_)
);

FILL FILL_2__1510_ (
);

FILL FILL_0__1336_ (
);

FILL FILL_2__865_ (
);

FILL FILL_3__807_ (
);

FILL FILL_3__980_ (
);

FILL FILL_1__1250_ (
);

FILL FILL_3__1176_ (
);

FILL FILL_1__887_ (
);

FILL FILL_0__1565_ (
);

FILL FILL_0__1145_ (
);

FILL FILL_1__1306_ (
);

FILL FILL_4__1474_ (
);

FILL FILL_0__1374_ (
);

FILL FILL_3__845_ (
);

FILL FILL_1__1115_ (
);

FILL FILL_2__959_ (
);

FILL FILL_0__1183_ (
);

FILL FILL_0__930_ (
);

NAND3X1 _933_ (
    .A(_115_),
    .B(_111_),
    .C(_117_),
    .Y(_125_)
);

FILL FILL_1__1344_ (
);

FILL FILL_4__861_ (
);

AOI21X1 _1199_ (
    .A(_244_),
    .B(_286_),
    .C(_388_),
    .Y(_389_)
);

FILL FILL_2__1413_ (
);

FILL FILL_0__1239_ (
);

FILL FILL_2__768_ (
);

FILL FILL_4__1092_ (
);

AOI21X1 _1411_ (
    .A(_616_),
    .B(_615_),
    .C(_570_),
    .Y(_617_)
);

FILL FILL_3__883_ (
);

FILL FILL_4__917_ (
);

FILL FILL_1__1573_ (
);

FILL FILL_1__1153_ (
);

FILL FILL_3__1499_ (
);

FILL FILL_3__1079_ (
);

FILL FILL_2__1222_ (
);

FILL FILL_0__1468_ (
);

FILL FILL_0__1048_ (
);

FILL FILL_2__997_ (
);

FILL FILL_3__939_ (
);

FILL FILL_1__1209_ (
);

AOI21X1 _1220_ (
    .A(_378_),
    .B(_379_),
    .C(_347_),
    .Y(_411_)
);

NAND2X1 _971_ (
    .A(Cin_0_bF$buf3),
    .B(Xin[6]),
    .Y(_162_)
);

FILL FILL_1__1382_ (
);

FILL FILL_2__1451_ (
);

FILL FILL_2__1031_ (
);

FILL FILL_0__1277_ (
);

FILL FILL_3__1100_ (
);

FILL FILL_1__1438_ (
);

FILL FILL_1__1018_ (
);

FILL FILL_1__811_ (
);

NAND3X1 _780_ (
    .A(Cin_0_bF$buf1),
    .B(Xin[2]),
    .C(Yin[2]),
    .Y(_644_)
);

FILL FILL_1__1191_ (
);

FILL FILL_2__1507_ (
);

FILL FILL_2__1260_ (
);

FILL FILL_0__1086_ (
);

OAI21X1 _1505_ (
    .A(_714_),
    .B(_700_),
    .C(_715_),
    .Y(_716_)
);

FILL FILL_0__833_ (
);

FILL FILL_3__977_ (
);

AOI21X1 _836_ (
    .A(Cin_0_bF$buf2),
    .B(Xin_3_bF$buf0),
    .C(Yin[3]),
    .Y(_28_)
);

FILL FILL_1__1247_ (
);

FILL FILL_2__1316_ (
);

FILL FILL89250x150 (
);

NAND3X1 _1314_ (
    .A(_508_),
    .B(_511_),
    .C(_510_),
    .Y(_512_)
);

FILL FILL_3__786_ (
);

FILL FILL_1__1476_ (
);

FILL FILL_1__1056_ (
);

FILL FILL_2__1125_ (
);

DFFPOSX1 _1543_ (
    .D(y[15]),
    .CLK(clk_bF$buf2),
    .Q(_755_[15])
);

INVX1 _1123_ (
    .A(_292_),
    .Y(_312_)
);

FILL FILL_0__871_ (
);

FILL FILL_1__905_ (
);

NAND3X1 _874_ (
    .A(_38_),
    .B(_61_),
    .C(_43_),
    .Y(_66_)
);

FILL FILL_1__1285_ (
);

FILL FILL_2__1354_ (
);

FILL FILL_0__927_ (
);

FILL FILL_3__1423_ (
);

FILL FILL_3__1003_ (
);

AOI21X1 _1352_ (
    .A(_549_),
    .B(_553_),
    .C(_499_),
    .Y(_554_)
);

FILL FILL_1__1094_ (
);

FILL FILL_2__921_ (
);

FILL FILL_2__1583_ (
);

FILL FILL_2__1163_ (
);

FILL FILL88050x54750 (
);

AOI21X1 _1408_ (
    .A(_609_),
    .B(_613_),
    .C(_571_),
    .Y(_614_)
);

FILL FILL_3__1232_ (
);

BUFX2 _1581_ (
    .A(_755_[7]),
    .Y(Yout[7])
);

AND2X2 _1161_ (
    .A(Cin[3]),
    .B(Xin[6]),
    .Y(_350_)
);

FILL FILL_1__943_ (
);

FILL FILL_0__1201_ (
);

FILL FILL_2__1219_ (
);

FILL FILL_2__1392_ (
);

AOI21X1 _1217_ (
    .A(_390_),
    .B(_391_),
    .C(_317_),
    .Y(_408_)
);

FILL FILL_0__965_ (
);

FILL FILL_3__1461_ (
);

FILL FILL_3__1041_ (
);

AOI21X1 _968_ (
    .A(Cin_0_bF$buf3),
    .B(Xin_5_bF$buf0),
    .C(Yin[5]),
    .Y(_159_)
);

FILL FILL_1__1379_ (
);

INVX1 _1390_ (
    .A(_574_),
    .Y(_594_)
);

FILL FILL_4__1110_ (
);

FILL FILL_2__1448_ (
);

FILL FILL_0__1430_ (
);

FILL FILL_0__1010_ (
);

FILL FILL_2__1028_ (
);

FILL FILL_3__901_ (
);

FILL FILL_3__1517_ (
);

NAND2X1 _1446_ (
    .A(_653_),
    .B(_652_),
    .Y(_654_)
);

AOI21X1 _1026_ (
    .A(_184_),
    .B(_185_),
    .C(_146_),
    .Y(_216_)
);

FILL FILL_0__774_ (
);

FILL FILL_1__808_ (
);

FILL FILL_3__1270_ (
);

OAI21X1 _777_ (
    .A(_461_),
    .B(_493_),
    .C(_483_),
    .Y(_612_)
);

FILL FILL88650x35250 (
);

FILL FILL_1__1188_ (
);

FILL FILL_1__981_ (
);

FILL FILL_2__1257_ (
);

FILL FILL_1__1400_ (
);

FILL FILL_3__1326_ (
);

NAND3X1 _1255_ (
    .A(_444_),
    .B(_448_),
    .C(_446_),
    .Y(_449_)
);

FILL FILL_1__790_ (
);

FILL FILL_2__824_ (
);

FILL FILL_2__1486_ (
);

FILL FILL_2__1066_ (
);

FILL FILL_3__1135_ (
);

XOR2X1 _1484_ (
    .A(_673_),
    .B(_694_),
    .Y(_753_[13])
);

NAND3X1 _1064_ (
    .A(_253_),
    .B(_248_),
    .C(_251_),
    .Y(_254_)
);

FILL FILL_1__846_ (
);

FILL FILL_0__1104_ (
);

FILL FILL_2__1295_ (
);

FILL FILL_0__868_ (
);

FILL FILL_3__1364_ (
);

FILL FILL88950x74250 (
);

NAND2X1 _1293_ (
    .A(_484_),
    .B(_489_),
    .Y(_490_)
);

FILL FILL_4__1433_ (
);

FILL FILL_0__1333_ (
);

FILL FILL_2__862_ (
);

FILL FILL_3__804_ (
);

NAND3X1 _1349_ (
    .A(_522_),
    .B(_527_),
    .C(_546_),
    .Y(_551_)
);

FILL FILL_3__1173_ (
);

FILL FILL_1__884_ (
);

FILL FILL_2__918_ (
);

FILL FILL_0__1562_ (
);

FILL FILL_0__1142_ (
);

FILL FILL_1__1303_ (
);

FILL FILL_3__1229_ (
);

FILL FILL_4__820_ (
);

BUFX2 _1578_ (
    .A(_755_[4]),
    .Y(Yout[4])
);

OAI21X1 _1158_ (
    .A(_346_),
    .B(_277_),
    .C(_271_),
    .Y(_347_)
);

FILL FILL_4__1051_ (
);

FILL FILL_0__1371_ (
);

FILL FILL_2__1389_ (
);

FILL FILL_3__842_ (
);

FILL FILL_1__1112_ (
);

FILL FILL_3__1458_ (
);

FILL FILL_3__1038_ (
);

NOR2X1 _1387_ (
    .A(_582_),
    .B(_580_),
    .Y(_591_)
);

FILL FILL_0__1427_ (
);

FILL FILL_0__1007_ (
);

FILL FILL_2__956_ (
);

FILL FILL_2__1198_ (
);

FILL FILL_0__1180_ (
);

INVX1 _930_ (
    .A(_78_),
    .Y(_122_)
);

FILL FILL_1__1341_ (
);

FILL FILL_3__1267_ (
);

AOI21X1 _1196_ (
    .A(_383_),
    .B(_384_),
    .C(_382_),
    .Y(_385_)
);

FILL FILL_1__978_ (
);

FILL FILL_2__1410_ (
);

FILL FILL_4__1336_ (
);

FILL FILL_0__1236_ (
);

FILL FILL_2__765_ (
);

FILL FILL_3__880_ (
);

FILL FILL_1__1570_ (
);

FILL FILL_1__1150_ (
);

FILL FILL_3__1496_ (
);

FILL FILL_3__1076_ (
);

BUFX2 BUFX2_insert10 (
    .A(Xin[3]),
    .Y(Xin_3_bF$buf3)
);

BUFX2 BUFX2_insert11 (
    .A(Xin[3]),
    .Y(Xin_3_bF$buf2)
);

BUFX2 BUFX2_insert12 (
    .A(Xin[3]),
    .Y(Xin_3_bF$buf1)
);

BUFX2 BUFX2_insert13 (
    .A(Xin[3]),
    .Y(Xin_3_bF$buf0)
);

BUFX2 BUFX2_insert14 (
    .A(Xin[5]),
    .Y(Xin_5_bF$buf3)
);

BUFX2 BUFX2_insert15 (
    .A(Xin[5]),
    .Y(Xin_5_bF$buf2)
);

BUFX2 BUFX2_insert16 (
    .A(Xin[5]),
    .Y(Xin_5_bF$buf1)
);

BUFX2 BUFX2_insert17 (
    .A(Xin[5]),
    .Y(Xin_5_bF$buf0)
);

FILL FILL_1__787_ (
);

FILL FILL_4__1565_ (
);

FILL FILL_0__1465_ (
);

FILL FILL_0__1045_ (
);

FILL FILL_2__994_ (
);

FILL FILL_3__936_ (
);

FILL FILL_1__1206_ (
);

FILL FILL88650x23550 (
);

FILL FILL_0__1274_ (
);

FILL FILL_1__1435_ (
);

FILL FILL_1__1015_ (
);

FILL FILL_2__1504_ (
);

FILL FILL_2__859_ (
);

FILL FILL_0__1083_ (
);

INVX1 _1502_ (
    .A(_713_),
    .Y(_714_)
);

FILL FILL_0__830_ (
);

FILL FILL_3__974_ (
);

AND2X2 _833_ (
    .A(_24_),
    .B(_25_),
    .Y(_751_[3])
);

FILL FILL_1__1244_ (
);

OAI21X1 _1099_ (
    .A(_285_),
    .B(_284_),
    .C(_246_),
    .Y(_289_)
);

FILL FILL_2__1313_ (
);

FILL FILL_4__1239_ (
);

FILL FILL_0__1139_ (
);

FILL FILL88050x19650 (
);

AND2X2 _1311_ (
    .A(Xin_5_bF$buf3),
    .B(Cin[5]),
    .Y(_509_)
);

FILL FILL_3__783_ (
);

FILL FILL_1__1473_ (
);

FILL FILL_1__1053_ (
);

FILL FILL_3__1399_ (
);

FILL FILL_4__990_ (
);

FILL FILL_2__1122_ (
);

FILL FILL_0__1368_ (
);

FILL FILL_2__897_ (
);

FILL FILL_3__839_ (
);

FILL FILL_1__1109_ (
);

DFFPOSX1 _1540_ (
    .D(y[12]),
    .CLK(clk_bF$buf2),
    .Q(_755_[12])
);

INVX1 _1120_ (
    .A(_307_),
    .Y(_309_)
);

FILL FILL_1__902_ (
);

NAND3X1 _871_ (
    .A(_27_),
    .B(_56_),
    .C(_62_),
    .Y(_63_)
);

FILL FILL_1__1282_ (
);

FILL FILL_2__1351_ (
);

FILL FILL_0__1177_ (
);

FILL FILL_0__924_ (
);

FILL FILL_3__1420_ (
);

FILL FILL_3__1000_ (
);

AOI22X1 _927_ (
    .A(_89_),
    .B(_93_),
    .C(_110_),
    .D(_106_),
    .Y(_119_)
);

FILL FILL_1__1338_ (
);

FILL FILL_1__1091_ (
);

FILL FILL_2__1407_ (
);

FILL FILL_2__1580_ (
);

FILL FILL_2__1160_ (
);

INVX1 _1405_ (
    .A(_572_),
    .Y(_610_)
);

FILL FILL_3__877_ (
);

FILL FILL_1__1567_ (
);

FILL FILL_1__1147_ (
);

FILL FILL_1__940_ (
);

FILL FILL_2__1216_ (
);

XNOR2X1 _1214_ (
    .A(_311_),
    .B(_404_),
    .Y(_753_[8])
);

FILL FILL_0__962_ (
);

OAI21X1 _965_ (
    .A(_87_),
    .B(_740_),
    .C(_149_),
    .Y(_156_)
);

FILL FILL_1__1376_ (
);

FILL FILL_2__1445_ (
);

FILL FILL_2__1025_ (
);

FILL FILL_3__1514_ (
);

NAND2X1 _1443_ (
    .A(Yin[11]),
    .B(_532_),
    .Y(_651_)
);

OAI21X1 _1023_ (
    .A(_137_),
    .B(_212_),
    .C(_200_),
    .Y(_213_)
);

FILL FILL_0__771_ (
);

FILL FILL_1__805_ (
);

FILL FILL_4__949_ (
);

FILL FILL88950x39150 (
);

NOR2X1 _774_ (
    .A(_569_),
    .B(_559_),
    .Y(_749_[1])
);

FILL FILL_1__1185_ (
);

FILL FILL_2__1254_ (
);

FILL FILL_0__827_ (
);

FILL FILL_3__1323_ (
);

NAND2X1 _1252_ (
    .A(_350_),
    .B(_445_),
    .Y(_446_)
);

FILL FILL_2__821_ (
);

FILL FILL_2__1483_ (
);

FILL FILL_2__1063_ (
);

AOI22X1 _1308_ (
    .A(Xin_5_bF$buf3),
    .B(Cin[5]),
    .C(Xin[4]),
    .D(Cin[6]),
    .Y(_506_)
);

FILL FILL_3__1132_ (
);

NAND3X1 _1481_ (
    .A(_647_),
    .B(_684_),
    .C(_691_),
    .Y(_692_)
);

NAND2X1 _1061_ (
    .A(_249_),
    .B(_250_),
    .Y(_251_)
);

FILL FILL_1__843_ (
);

FILL FILL_2__1119_ (
);

FILL FILL_0__1101_ (
);

FILL FILL_2__1292_ (
);

DFFPOSX1 _1537_ (
    .D(y[9]),
    .CLK(clk_bF$buf0),
    .Q(_755_[9])
);

OAI21X1 _1117_ (
    .A(_306_),
    .B(_305_),
    .C(_304_),
    .Y(_307_)
);

FILL FILL_0__865_ (
);

FILL FILL_3__1361_ (
);

NAND3X1 _868_ (
    .A(_44_),
    .B(_52_),
    .C(_53_),
    .Y(_60_)
);

FILL FILL_1__1279_ (
);

AOI21X1 _1290_ (
    .A(_481_),
    .B(_480_),
    .C(_479_),
    .Y(_487_)
);

FILL FILL_2__1348_ (
);

FILL FILL_0__1330_ (
);

FILL FILL_3__801_ (
);

FILL FILL_3__1417_ (
);

NOR2X1 _1346_ (
    .A(_546_),
    .B(_542_),
    .Y(_547_)
);

FILL FILL_3__1170_ (
);

FILL FILL_1__1088_ (
);

FILL FILL_1__881_ (
);

FILL FILL_2__915_ (
);

FILL FILL_2__1577_ (
);

FILL FILL_2__1157_ (
);

FILL FILL_1__1300_ (
);

FILL FILL_3__1226_ (
);

BUFX2 _1575_ (
    .A(_755_[15]),
    .Y(Yout[15])
);

NAND3X1 _1155_ (
    .A(_341_),
    .B(_342_),
    .C(_343_),
    .Y(_344_)
);

FILL FILL_1__937_ (
);

FILL FILL_2__1386_ (
);

FILL FILL_0__959_ (
);

FILL FILL_3__1455_ (
);

FILL FILL_3__1035_ (
);

NAND3X1 _1384_ (
    .A(_536_),
    .B(_581_),
    .C(_586_),
    .Y(_587_)
);

FILL FILL_0__1424_ (
);

FILL FILL_0__1004_ (
);

FILL FILL_2__953_ (
);

FILL FILL_2__1195_ (
);

FILL FILL_0__768_ (
);

FILL FILL_3__1264_ (
);

AND2X2 _1193_ (
    .A(_340_),
    .B(_344_),
    .Y(_382_)
);

FILL FILL_1__975_ (
);

FILL FILL_0__1233_ (
);

FILL FILL_2__762_ (
);

NAND2X1 _1249_ (
    .A(Xin_5_bF$buf1),
    .B(Cin[4]),
    .Y(_443_)
);

FILL FILL_0__997_ (
);

FILL FILL_3__1493_ (
);

FILL FILL_3__1073_ (
);

FILL FILL_1__784_ (
);

FILL FILL_2__818_ (
);

FILL FILL_0__1462_ (
);

FILL FILL_0__1042_ (
);

FILL FILL_2__991_ (
);

FILL FILL_3__933_ (
);

FILL FILL_1__1203_ (
);

FILL FILL_3__1129_ (
);

FILL FILL88950x27450 (
);

OAI21X1 _1478_ (
    .A(_650_),
    .B(_651_),
    .C(_657_),
    .Y(_689_)
);

INVX1 _1058_ (
    .A(_247_),
    .Y(_248_)
);

FILL FILL_0__1518_ (
);

FILL FILL88650x85950 (
);

FILL FILL_2__1289_ (
);

FILL FILL_0__1271_ (
);

FILL FILL_1__1432_ (
);

FILL FILL_1__1012_ (
);

FILL FILL_3__1358_ (
);

NAND3X1 _1287_ (
    .A(_409_),
    .B(_478_),
    .C(_482_),
    .Y(_484_)
);

FILL FILL_2__1501_ (
);

FILL FILL_0__1327_ (
);

FILL FILL_2__856_ (
);

FILL FILL_4__1180_ (
);

FILL FILL_2__1098_ (
);

FILL FILL_0__1080_ (
);

FILL FILL_3__971_ (
);

NOR3X1 _830_ (
    .A(_735_),
    .B(_22_),
    .C(_21_),
    .Y(_23_)
);

FILL FILL_1__1241_ (
);

FILL FILL_3__1167_ (
);

OAI21X1 _1096_ (
    .A(_284_),
    .B(_285_),
    .C(_283_),
    .Y(_286_)
);

FILL FILL_1__878_ (
);

FILL FILL_2__1310_ (
);

FILL FILL_0__1136_ (
);

FILL FILL_3__780_ (
);

FILL FILL_1__1470_ (
);

FILL FILL_1__1050_ (
);

FILL FILL_3__1396_ (
);

FILL FILL_4__1465_ (
);

FILL FILL_0__1365_ (
);

FILL FILL_2__894_ (
);

FILL FILL_3__836_ (
);

FILL FILL_1__1106_ (
);

FILL FILL_0__1174_ (
);

FILL FILL_0__921_ (
);

NAND3X1 _924_ (
    .A(_115_),
    .B(_111_),
    .C(_82_),
    .Y(_116_)
);

FILL FILL_1__1335_ (
);

FILL FILL_4__852_ (
);

FILL FILL_2__1404_ (
);

FILL FILL_2__759_ (
);

FILL FILL_4__1083_ (
);

OAI21X1 _1402_ (
    .A(_605_),
    .B(_606_),
    .C(_602_),
    .Y(_607_)
);

FILL FILL_3__874_ (
);

FILL FILL_1__1564_ (
);

FILL FILL_1__1144_ (
);

FILL FILL_2__1213_ (
);

FILL FILL_0__1459_ (
);

FILL FILL_0__1039_ (
);

FILL FILL_2__988_ (
);

NAND3X1 _1211_ (
    .A(_315_),
    .B(_387_),
    .C(_392_),
    .Y(_402_)
);

OAI21X1 _962_ (
    .A(_590_),
    .B(_151_),
    .C(_152_),
    .Y(_153_)
);

FILL FILL_1__1373_ (
);

FILL FILL_3__1299_ (
);

FILL FILL_2__1442_ (
);

FILL FILL_2__1022_ (
);

FILL FILL_4__1368_ (
);

FILL FILL_0__1268_ (
);

FILL FILL_2__797_ (
);

FILL FILL_3__1511_ (
);

FILL FILL_1__1429_ (
);

FILL FILL_1__1009_ (
);

AOI21X1 _1440_ (
    .A(_645_),
    .B(_642_),
    .C(_638_),
    .Y(_648_)
);

NOR2X1 _1020_ (
    .A(_210_),
    .B(_209_),
    .Y(_753_[6])
);

FILL FILL_1__802_ (
);

NAND3X1 _771_ (
    .A(_515_),
    .B(_537_),
    .C(_429_),
    .Y(_548_)
);

FILL FILL_1__1182_ (
);

FILL FILL_2__1251_ (
);

FILL FILL_0__1497_ (
);

FILL FILL_0__1077_ (
);

FILL FILL_0__824_ (
);

FILL FILL_3__968_ (
);

FILL FILL_3__1320_ (
);

NAND2X1 _827_ (
    .A(_14_),
    .B(_19_),
    .Y(_20_)
);

FILL FILL_1__1238_ (
);

FILL FILL88950x15750 (
);

FILL FILL_2__1307_ (
);

FILL FILL_2__1480_ (
);

FILL FILL_2__1060_ (
);

NAND2X1 _1305_ (
    .A(Xin_3_bF$buf3),
    .B(Cin[7]),
    .Y(_502_)
);

FILL FILL_3__777_ (
);

FILL FILL_1__1467_ (
);

FILL FILL_1__1047_ (
);

FILL FILL_1__840_ (
);

FILL FILL_2__1116_ (
);

DFFPOSX1 _1534_ (
    .D(y[6]),
    .CLK(clk_bF$buf0),
    .Q(_755_[6])
);

AOI21X1 _1114_ (
    .A(_199_),
    .B(_201_),
    .C(_303_),
    .Y(_304_)
);

FILL FILL_0__862_ (
);

AOI21X1 _865_ (
    .A(_41_),
    .B(_42_),
    .C(_40_),
    .Y(_57_)
);

FILL FILL_1__1276_ (
);

FILL FILL_2__1345_ (
);

FILL FILL_0__918_ (
);

FILL FILL_3__1414_ (
);

AND2X2 _1343_ (
    .A(_538_),
    .B(_534_),
    .Y(_544_)
);

FILL FILL_1__1085_ (
);

FILL FILL_2__912_ (
);

FILL FILL_2__1574_ (
);

FILL FILL_2__1154_ (
);

FILL FILL_3__1223_ (
);

BUFX2 _1572_ (
    .A(_755_[12]),
    .Y(Yout[12])
);

AND2X2 _1152_ (
    .A(_226_),
    .B(_223_),
    .Y(_341_)
);

FILL FILL_1__934_ (
);

FILL FILL_2__1383_ (
);

AOI21X1 _1208_ (
    .A(_287_),
    .B(_291_),
    .C(_217_),
    .Y(_399_)
);

FILL FILL_0__956_ (
);

FILL FILL_3__1452_ (
);

FILL FILL_3__1032_ (
);

NAND2X1 _959_ (
    .A(_85_),
    .B(_149_),
    .Y(_150_)
);

NOR2X1 _1381_ (
    .A(_503_),
    .B(_576_),
    .Y(_584_)
);

FILL FILL_4__1101_ (
);

FILL FILL_0__1421_ (
);

FILL FILL_2__1439_ (
);

FILL FILL_2__1019_ (
);

FILL FILL_0__1001_ (
);

FILL FILL_2__950_ (
);

FILL FILL_2__1192_ (
);

FILL FILL_3__1508_ (
);

OR2X2 _1437_ (
    .A(_641_),
    .B(_643_),
    .Y(_645_)
);

NAND3X1 _1017_ (
    .A(_136_),
    .B(_207_),
    .C(_203_),
    .Y(_208_)
);

FILL FILL_0__765_ (
);

FILL FILL_3__1261_ (
);

NAND3X1 _768_ (
    .A(_472_),
    .B(_483_),
    .C(_504_),
    .Y(_515_)
);

FILL FILL_1__1179_ (
);

NAND3X1 _1190_ (
    .A(_365_),
    .B(_359_),
    .C(_367_),
    .Y(_379_)
);

FILL FILL_1__972_ (
);

FILL FILL_0__1230_ (
);

FILL FILL_2__1248_ (
);

FILL FILL_3__1317_ (
);

AND2X2 _1246_ (
    .A(_434_),
    .B(_438_),
    .Y(_439_)
);

FILL FILL_0__994_ (
);

FILL FILL_3__1490_ (
);

FILL FILL_3__1070_ (
);

XOR2X1 _997_ (
    .A(_143_),
    .B(_142_),
    .Y(_188_)
);

FILL FILL_1__781_ (
);

FILL FILL_2__815_ (
);

FILL FILL_2__1477_ (
);

FILL FILL_2__1057_ (
);

FILL FILL_3__930_ (
);

FILL FILL_1__1200_ (
);

FILL FILL_3__1126_ (
);

INVX1 _1475_ (
    .A(_684_),
    .Y(_685_)
);

AOI21X1 _1055_ (
    .A(_174_),
    .B(_173_),
    .C(_160_),
    .Y(_245_)
);

FILL FILL_1__837_ (
);

FILL FILL_0__1515_ (
);

FILL FILL_2__1286_ (
);

FILL FILL_0__859_ (
);

FILL FILL_3__1355_ (
);

OAI21X1 _1284_ (
    .A(_476_),
    .B(_475_),
    .C(_412_),
    .Y(_480_)
);

FILL FILL_4__1424_ (
);

FILL FILL_0__1324_ (
);

FILL FILL_1_BUFX2_insert10 (
);

FILL FILL_1_BUFX2_insert11 (
);

FILL FILL_1_BUFX2_insert12 (
);

FILL FILL_1_BUFX2_insert13 (
);

FILL FILL_1_BUFX2_insert14 (
);

FILL FILL_1_BUFX2_insert15 (
);

FILL FILL_2__853_ (
);

FILL FILL_1_BUFX2_insert16 (
);

FILL FILL_1_BUFX2_insert17 (
);

FILL FILL_2__1095_ (
);

FILL FILL_3__1164_ (
);

AOI21X1 _1093_ (
    .A(_183_),
    .B(_178_),
    .C(_282_),
    .Y(_283_)
);

FILL FILL_1__875_ (
);

FILL FILL_2__909_ (
);

FILL FILL_0__1133_ (
);

FILL FILL_4__811_ (
);

BUFX2 _1569_ (
    .A(_755_[1]),
    .Y(Yout[1])
);

AOI22X1 _1149_ (
    .A(_149_),
    .B(_337_),
    .C(_253_),
    .D(_248_),
    .Y(_338_)
);

FILL FILL_0__897_ (
);

FILL FILL_3__1393_ (
);

FILL FILL_0__1362_ (
);

FILL FILL_2__891_ (
);

FILL FILL_3__833_ (
);

FILL FILL_1__1103_ (
);

FILL FILL_3__1449_ (
);

FILL FILL_3__1029_ (
);

OAI21X1 _1378_ (
    .A(_151_),
    .B(_575_),
    .C(_580_),
    .Y(_581_)
);

FILL FILL_0__1418_ (
);

FILL FILL_2__947_ (
);

FILL FILL89550x150 (
);

FILL FILL88650x4050 (
);

FILL FILL_0__1171_ (
);

FILL FILL_2__1189_ (
);

FILL FILL89250x35250 (
);

OAI21X1 _921_ (
    .A(_109_),
    .B(_108_),
    .C(_95_),
    .Y(_113_)
);

FILL FILL_1__1332_ (
);

FILL FILL_3__1258_ (
);

AOI21X1 _1187_ (
    .A(_258_),
    .B(_275_),
    .C(_375_),
    .Y(_376_)
);

FILL FILL_1__969_ (
);

FILL FILL_2__1401_ (
);

FILL FILL_4__1327_ (
);

FILL FILL_0__1227_ (
);

FILL FILL_2__756_ (
);

FILL FILL_3__871_ (
);

FILL FILL_1__1561_ (
);

FILL FILL_1__1141_ (
);

FILL FILL_3__1487_ (
);

FILL FILL_3__1067_ (
);

FILL FILL_1__778_ (
);

FILL FILL_2__1210_ (
);

FILL FILL_0__1456_ (
);

FILL FILL_0__1036_ (
);

FILL FILL_2__985_ (
);

FILL FILL_3__927_ (
);

FILL FILL_1__1370_ (
);

FILL FILL_3__1296_ (
);

FILL FILL_0__1265_ (
);

FILL FILL_2__794_ (
);

FILL FILL89550x74250 (
);

FILL FILL_1__1426_ (
);

FILL FILL_1__1006_ (
);

FILL FILL_0__1494_ (
);

FILL FILL_0__1074_ (
);

FILL FILL_0__821_ (
);

FILL FILL_3__965_ (
);

INVX1 _824_ (
    .A(_9_),
    .Y(_17_)
);

FILL FILL_1__1235_ (
);

FILL FILL_2__1304_ (
);

INVX1 _1302_ (
    .A(_498_),
    .Y(_499_)
);

FILL FILL_3__774_ (
);

FILL FILL_1__1464_ (
);

FILL FILL_1__1044_ (
);

FILL FILL_4__981_ (
);

FILL FILL_2__1113_ (
);

FILL FILL_0__1359_ (
);

FILL FILL_2__888_ (
);

DFFPOSX1 _1531_ (
    .D(y[3]),
    .CLK(clk_bF$buf3),
    .Q(_755_[3])
);

NAND3X1 _1111_ (
    .A(_214_),
    .B(_299_),
    .C(_300_),
    .Y(_301_)
);

NAND3X1 _862_ (
    .A(_50_),
    .B(_52_),
    .C(_53_),
    .Y(_54_)
);

FILL FILL_1__1273_ (
);

FILL FILL_3__1199_ (
);

FILL FILL_2__1342_ (
);

FILL FILL_0__1168_ (
);

FILL FILL_0__915_ (
);

FILL FILL_3__1411_ (
);

OAI21X1 _918_ (
    .A(_109_),
    .B(_108_),
    .C(_107_),
    .Y(_110_)
);

FILL FILL_1__1329_ (
);

NOR2X1 _1340_ (
    .A(_528_),
    .B(_540_),
    .Y(_541_)
);

FILL FILL_1__1082_ (
);

FILL FILL_2__1571_ (
);

FILL FILL_2__1151_ (
);

FILL FILL_4__1497_ (
);

FILL FILL_0__1397_ (
);

FILL FILL_3__868_ (
);

FILL FILL_3__1220_ (
);

FILL FILL_1__1138_ (
);

FILL FILL_1__931_ (
);

FILL FILL_2__1207_ (
);

FILL FILL_2__1380_ (
);

FILL FILL89250x23550 (
);

OAI21X1 _1205_ (
    .A(_381_),
    .B(_385_),
    .C(_389_),
    .Y(_395_)
);

FILL FILL_0__953_ (
);

NAND2X1 _956_ (
    .A(Xin[2]),
    .B(Cin[4]),
    .Y(_147_)
);

FILL FILL_1__1367_ (
);

FILL FILL_4__884_ (
);

FILL FILL_2__1436_ (
);

FILL FILL_2__1016_ (
);

FILL FILL_3__1505_ (
);

OAI21X1 _1434_ (
    .A(_578_),
    .B(_639_),
    .C(_640_),
    .Y(_641_)
);

NAND3X1 _1014_ (
    .A(_199_),
    .B(_200_),
    .C(_201_),
    .Y(_205_)
);

FILL FILL_0__762_ (
);

NAND3X1 _765_ (
    .A(Cin_0_bF$buf1),
    .B(Xin[1]),
    .C(Yin[1]),
    .Y(_483_)
);

FILL FILL_1__1176_ (
);

FILL FILL_2__1245_ (
);

FILL FILL_0__818_ (
);

FILL FILL_3__1314_ (
);

NAND3X1 _1243_ (
    .A(_425_),
    .B(_432_),
    .C(_420_),
    .Y(_436_)
);

FILL FILL_0__991_ (
);

NAND3X1 _994_ (
    .A(_158_),
    .B(_171_),
    .C(_175_),
    .Y(_185_)
);

FILL FILL_2__812_ (
);

FILL FILL_2__1474_ (
);

FILL FILL_2__1054_ (
);

FILL FILL_3__1123_ (
);

XOR2X1 _1472_ (
    .A(_681_),
    .B(_675_),
    .Y(_682_)
);

OAI21X1 _1052_ (
    .A(_236_),
    .B(_235_),
    .C(_233_),
    .Y(_242_)
);

FILL FILL_1__834_ (
);

FILL FILL_0__1512_ (
);

FILL FILL_2__1283_ (
);

DFFPOSX1 _1528_ (
    .D(y[0]),
    .CLK(clk_bF$buf4),
    .Q(_755_[0])
);

NAND3X1 _1108_ (
    .A(_215_),
    .B(_292_),
    .C(_297_),
    .Y(_298_)
);

FILL FILL_0__856_ (
);

FILL FILL_3__1352_ (
);

INVX1 _859_ (
    .A(Xin[1]),
    .Y(_51_)
);

OAI21X1 _1281_ (
    .A(_475_),
    .B(_476_),
    .C(_471_),
    .Y(_477_)
);

FILL FILL_0__1321_ (
);

FILL FILL_2__1339_ (
);

FILL FILL_2__850_ (
);

FILL FILL_2__1092_ (
);

FILL FILL_3__1408_ (
);

OAI21X1 _1337_ (
    .A(_531_),
    .B(_536_),
    .C(_535_),
    .Y(_538_)
);

FILL FILL_3__1581_ (
);

FILL FILL_3__1161_ (
);

FILL FILL_1__1499_ (
);

FILL FILL_1__1079_ (
);

NAND3X1 _1090_ (
    .A(_277_),
    .B(_279_),
    .C(_278_),
    .Y(_280_)
);

FILL FILL_1__872_ (
);

FILL FILL_2__906_ (
);

FILL FILL_4__1230_ (
);

FILL FILL_2__1568_ (
);

FILL FILL_2__1148_ (
);

FILL FILL_0__1130_ (
);

FILL FILL_3__1217_ (
);

BUFX2 _1566_ (
    .A(_754_[6]),
    .Y(Xout[6])
);

AOI21X1 _1146_ (
    .A(_323_),
    .B(_326_),
    .C(_320_),
    .Y(_335_)
);

FILL FILL_0__894_ (
);

FILL FILL_1__928_ (
);

FILL FILL_3__1390_ (
);

NAND3X1 _897_ (
    .A(_84_),
    .B(_88_),
    .C(_86_),
    .Y(_89_)
);

FILL FILL_2__1377_ (
);

FILL FILL_3__830_ (
);

FILL FILL_1__1100_ (
);

FILL FILL_3__1446_ (
);

FILL FILL_3__1026_ (
);

NAND2X1 _1375_ (
    .A(Cin[5]),
    .B(Xin[6]),
    .Y(_578_)
);

FILL FILL_0__1415_ (
);

FILL FILL_2__944_ (
);

FILL FILL_2__1186_ (
);

FILL FILL89550x39150 (
);

FILL FILL_0__759_ (
);

FILL FILL_3__1255_ (
);

AOI22X1 _1184_ (
    .A(_354_),
    .B(_358_),
    .C(_369_),
    .D(_372_),
    .Y(_373_)
);

FILL FILL_1__966_ (
);

FILL FILL_0__1224_ (
);

FILL FILL89250x11850 (
);

FILL FILL_0__988_ (
);

FILL FILL_3__1484_ (
);

FILL FILL_3__1064_ (
);

FILL FILL_1__775_ (
);

FILL FILL_2__809_ (
);

FILL FILL_4__1133_ (
);

FILL FILL_0__1453_ (
);

FILL FILL_0__1033_ (
);

FILL FILL_2__982_ (
);

FILL FILL_3__924_ (
);

NAND2X1 _1469_ (
    .A(_677_),
    .B(_678_),
    .Y(_679_)
);

OAI21X1 _1049_ (
    .A(_236_),
    .B(_235_),
    .C(_238_),
    .Y(_239_)
);

FILL FILL_0__797_ (
);

FILL FILL_3__1293_ (
);

FILL FILL_0__1509_ (
);

FILL FILL_0__1262_ (
);

FILL FILL_2__791_ (
);

FILL FILL_1__1423_ (
);

FILL FILL_1__1003_ (
);

FILL FILL_3__1349_ (
);

FILL FILL_4__940_ (
);

NAND3X1 _1278_ (
    .A(_454_),
    .B(_457_),
    .C(_460_),
    .Y(_474_)
);

FILL FILL_0__1318_ (
);

FILL FILL_2__847_ (
);

FILL FILL_0__1491_ (
);

FILL FILL_2__1089_ (
);

FILL FILL_0__1071_ (
);

FILL FILL_3__962_ (
);

NAND3X1 _821_ (
    .A(_9_),
    .B(_13_),
    .C(_745_),
    .Y(_14_)
);

FILL FILL_1__1232_ (
);

FILL FILL_3__1578_ (
);

FILL FILL_3__1158_ (
);

NAND2X1 _1087_ (
    .A(_254_),
    .B(_257_),
    .Y(_277_)
);

FILL FILL_1__869_ (
);

FILL FILL_2__1301_ (
);

FILL FILL_0__1127_ (
);

FILL FILL_3__771_ (
);

FILL FILL_1__1461_ (
);

FILL FILL_1__1041_ (
);

FILL FILL_3__1387_ (
);

FILL FILL_2__1110_ (
);

FILL FILL_4__1456_ (
);

FILL FILL_0__1356_ (
);

FILL FILL_2__885_ (
);

FILL FILL_3__827_ (
);

FILL FILL_1__1517_ (
);

FILL FILL_1__1270_ (
);

FILL FILL_3__1196_ (
);

FILL FILL_0__1165_ (
);

FILL FILL_0__912_ (
);

INVX1 _915_ (
    .A(_95_),
    .Y(_107_)
);

FILL FILL_1__1326_ (
);

FILL FILL_4__843_ (
);

FILL FILL_4__1074_ (
);

FILL FILL_0__1394_ (
);

FILL FILL_3__865_ (
);

FILL FILL_1__1135_ (
);

FILL FILL_2__1204_ (
);

FILL FILL_2__979_ (
);

FILL FILL89550x27450 (
);

NAND3X1 _1202_ (
    .A(_390_),
    .B(_391_),
    .C(_389_),
    .Y(_392_)
);

FILL FILL_0__950_ (
);

XNOR2X1 _953_ (
    .A(_143_),
    .B(_142_),
    .Y(_144_)
);

FILL FILL_1__1364_ (
);

FILL FILL89250x85950 (
);

FILL FILL_2__1433_ (
);

FILL FILL_2__1013_ (
);

FILL FILL_4__1359_ (
);

FILL FILL_0__1259_ (
);

FILL FILL_2__788_ (
);

FILL FILL_3__1502_ (
);

OAI21X1 _1431_ (
    .A(_582_),
    .B(_580_),
    .C(_585_),
    .Y(_638_)
);

AOI21X1 _1011_ (
    .A(_201_),
    .B(_200_),
    .C(_199_),
    .Y(_202_)
);

NOR2X1 _762_ (
    .A(_440_),
    .B(_429_),
    .Y(_748_[0])
);

FILL FILL_1__1173_ (
);

FILL FILL_3__1099_ (
);

FILL FILL_2__1242_ (
);

FILL FILL_0__1488_ (
);

FILL FILL_0__1068_ (
);

FILL FILL_0__815_ (
);

FILL FILL_3__959_ (
);

FILL FILL_3__1311_ (
);

AOI21X1 _818_ (
    .A(_7_),
    .B(_6_),
    .C(_747_),
    .Y(_11_)
);

FILL FILL_1__1229_ (
);

OAI21X1 _1240_ (
    .A(_430_),
    .B(_431_),
    .C(_432_),
    .Y(_433_)
);

AOI21X1 _991_ (
    .A(_94_),
    .B(_110_),
    .C(_181_),
    .Y(_182_)
);

FILL FILL_2__1471_ (
);

FILL FILL_2__1051_ (
);

FILL FILL_0__1297_ (
);

FILL FILL_3__768_ (
);

FILL FILL_3__1120_ (
);

FILL FILL_1__1458_ (
);

FILL FILL_1__1038_ (
);

FILL FILL_1__831_ (
);

FILL FILL_2__1107_ (
);

FILL FILL_2__1280_ (
);

DFFPOSX1 _1525_ (
    .D(Xin_5_bF$buf2),
    .CLK(clk_bF$buf0),
    .Q(_754_[5])
);

AOI21X1 _1105_ (
    .A(_290_),
    .B(_289_),
    .C(_288_),
    .Y(_295_)
);

FILL FILL_0__853_ (
);

FILL FILL_3__997_ (
);

OAI21X1 _856_ (
    .A(_47_),
    .B(_590_),
    .C(_15_),
    .Y(_48_)
);

FILL FILL_1__1267_ (
);

FILL FILL_2__1336_ (
);

FILL FILL_0__909_ (
);

FILL FILL_3__1405_ (
);

NAND2X1 _1334_ (
    .A(Yin[10]),
    .B(_533_),
    .Y(_534_)
);

FILL FILL_1__1496_ (
);

FILL FILL_1__1076_ (
);

FILL FILL_2__903_ (
);

FILL FILL_2__1565_ (
);

FILL FILL_2__1145_ (
);

FILL FILL_3__1214_ (
);

BUFX2 _1563_ (
    .A(_754_[3]),
    .Y(Xout[3])
);

OAI21X1 _1143_ (
    .A(_247_),
    .B(_331_),
    .C(_251_),
    .Y(_332_)
);

FILL FILL_0__891_ (
);

FILL FILL_1__925_ (
);

NAND2X1 _894_ (
    .A(_45_),
    .B(_85_),
    .Y(_86_)
);

FILL FILL_2__1374_ (
);

FILL FILL_0__947_ (
);

FILL FILL_3__1443_ (
);

FILL FILL_3__1023_ (
);

INVX1 _1372_ (
    .A(Cin[7]),
    .Y(_575_)
);

FILL FILL_0__1412_ (
);

FILL FILL_2__941_ (
);

FILL FILL_2__1183_ (
);

NAND2X1 _1428_ (
    .A(_587_),
    .B(_593_),
    .Y(_635_)
);

INVX1 _1008_ (
    .A(_137_),
    .Y(_199_)
);

FILL FILL_0__756_ (
);

FILL FILL_3__1252_ (
);

NAND2X1 _759_ (
    .A(Yin[0]),
    .B(_407_),
    .Y(_418_)
);

INVX1 _1181_ (
    .A(_364_),
    .Y(_370_)
);

FILL FILL_1__963_ (
);

FILL FILL_0__1221_ (
);

FILL FILL_2__1239_ (
);

FILL FILL89550x15750 (
);

FILL FILL_3__1308_ (
);

AOI21X1 _1237_ (
    .A(_424_),
    .B(_422_),
    .C(_421_),
    .Y(_430_)
);

FILL FILL_0__985_ (
);

FILL FILL_3__1481_ (
);

FILL FILL_3__1061_ (
);

AOI22X1 _988_ (
    .A(_154_),
    .B(_157_),
    .C(_178_),
    .D(_177_),
    .Y(_179_)
);

FILL FILL_1__1399_ (
);

FILL FILL_1__772_ (
);

FILL FILL_2__806_ (
);

FILL FILL_2__1468_ (
);

FILL FILL_0__1450_ (
);

FILL FILL_2__1048_ (
);

FILL FILL_0__1030_ (
);

FILL FILL_3__921_ (
);

FILL FILL_3__1117_ (
);

OAI22X1 _1466_ (
    .A(_578_),
    .B(_639_),
    .C(_643_),
    .D(_641_),
    .Y(_675_)
);

AOI22X1 _1046_ (
    .A(Xin[0]),
    .B(Cin[7]),
    .C(_223_),
    .D(_225_),
    .Y(_236_)
);

FILL FILL_0__794_ (
);

FILL FILL_1__828_ (
);

FILL FILL_3__1290_ (
);

OAI21X1 _797_ (
    .A(_732_),
    .B(_718_),
    .C(_708_),
    .Y(_738_)
);

FILL FILL_0__1506_ (
);

FILL FILL_2__1277_ (
);

FILL FILL_1__1420_ (
);

FILL FILL_1__1000_ (
);

FILL FILL_3__1346_ (
);

INVX1 _1275_ (
    .A(_383_),
    .Y(_470_)
);

FILL FILL_0__1315_ (
);

FILL FILL_2__844_ (
);

FILL FILL_2__1086_ (
);

FILL FILL_3__1575_ (
);

FILL FILL_3__1155_ (
);

AOI21X1 _1084_ (
    .A(_266_),
    .B(_263_),
    .C(_262_),
    .Y(_274_)
);

FILL FILL_1__866_ (
);

FILL FILL_0__1124_ (
);

FILL FILL_0__888_ (
);

FILL FILL_3__1384_ (
);

FILL FILL_0__1353_ (
);

FILL FILL_2__882_ (
);

FILL FILL_3__824_ (
);

FILL FILL_1__1514_ (
);

NAND2X1 _1369_ (
    .A(_544_),
    .B(_530_),
    .Y(_572_)
);

FILL FILL_3__1193_ (
);

FILL FILL_0__1409_ (
);

FILL FILL_2__938_ (
);

FILL FILL_4__1262_ (
);

FILL FILL_0__1582_ (
);

FILL FILL_0__1162_ (
);

NAND3X1 _912_ (
    .A(Cin_0_bF$buf2),
    .B(Xin_5_bF$buf2),
    .C(_99_),
    .Y(_104_)
);

FILL FILL_1__1323_ (
);

FILL FILL_3__1249_ (
);

NAND3X1 _1178_ (
    .A(_263_),
    .B(_267_),
    .C(_366_),
    .Y(_367_)
);

FILL FILL_4__1318_ (
);

FILL FILL_0__1218_ (
);

FILL FILL_0__1391_ (
);

FILL FILL_3__862_ (
);

FILL FILL_1__1132_ (
);

FILL FILL_3__1478_ (
);

FILL FILL_3__1058_ (
);

FILL FILL_1__769_ (
);

FILL FILL_2__1201_ (
);

FILL FILL_0__1447_ (
);

FILL FILL_0__1027_ (
);

FILL FILL_2__976_ (
);

FILL FILL_3__918_ (
);

AOI22X1 _950_ (
    .A(Xin[0]),
    .B(Cin[6]),
    .C(Xin[1]),
    .D(Cin[5]),
    .Y(_141_)
);

FILL FILL_1__1361_ (
);

FILL FILL_3__1287_ (
);

FILL FILL_1__998_ (
);

FILL FILL_2__1430_ (
);

FILL FILL_2__1010_ (
);

FILL FILL_0__1256_ (
);

FILL FILL_2__785_ (
);

FILL FILL_1__1417_ (
);

FILL FILL_1__1170_ (
);

FILL FILL_3__1096_ (
);

FILL FILL_0__1485_ (
);

FILL FILL_0__1065_ (
);

FILL FILL_0__812_ (
);

FILL FILL_3__956_ (
);

NAND3X1 _815_ (
    .A(_747_),
    .B(_6_),
    .C(_7_),
    .Y(_8_)
);

FILL FILL_1__1226_ (
);

FILL FILL_0__1294_ (
);

FILL FILL_3__765_ (
);

FILL FILL_1__1455_ (
);

FILL FILL_1__1035_ (
);

FILL FILL_4__972_ (
);

FILL FILL_2__1104_ (
);

FILL FILL_2__879_ (
);

DFFPOSX1 _1522_ (
    .D(Xin[2]),
    .CLK(clk_bF$buf4),
    .Q(_754_[2])
);

NAND3X1 _1102_ (
    .A(_291_),
    .B(_287_),
    .C(_217_),
    .Y(_292_)
);

FILL FILL_0__850_ (
);

FILL FILL_3__994_ (
);

AND2X2 _853_ (
    .A(Xin[2]),
    .B(Cin[2]),
    .Y(_45_)
);

FILL FILL_1__1264_ (
);

FILL FILL_2__1333_ (
);

FILL FILL_0__1579_ (
);

FILL FILL_0__1159_ (
);

FILL FILL_0__906_ (
);

FILL FILL_3__1402_ (
);

NAND2X1 _909_ (
    .A(_99_),
    .B(_100_),
    .Y(_101_)
);

AOI22X1 _1331_ (
    .A(Cin[3]),
    .B(Xin[7]),
    .C(Cin[4]),
    .D(Xin[6]),
    .Y(_531_)
);

FILL FILL_1__1493_ (
);

FILL FILL_1__1073_ (
);

FILL FILL_2__900_ (
);

FILL FILL_2__1562_ (
);

FILL FILL_2__1142_ (
);

FILL FILL_4__1488_ (
);

FILL FILL_0__1388_ (
);

FILL FILL_3__859_ (
);

FILL FILL_3__1211_ (
);

FILL FILL88650x7950 (
);

FILL FILL_1__1129_ (
);

BUFX2 _1560_ (
    .A(_754_[0]),
    .Y(Xout[0])
);

OAI21X1 _1140_ (
    .A(_47_),
    .B(_324_),
    .C(_322_),
    .Y(_329_)
);

FILL FILL_1__922_ (
);

NAND2X1 _891_ (
    .A(Xin[1]),
    .B(Cin[4]),
    .Y(_83_)
);

FILL FILL_2__1371_ (
);

FILL FILL_0__1197_ (
);

FILL FILL_0__944_ (
);

FILL FILL_3__1440_ (
);

FILL FILL_3__1020_ (
);

AOI21X1 _947_ (
    .A(_111_),
    .B(_115_),
    .C(_82_),
    .Y(_138_)
);

FILL FILL_1__1358_ (
);

FILL FILL_4__875_ (
);

FILL FILL_2__1427_ (
);

FILL FILL_2__1007_ (
);

FILL FILL_2__1180_ (
);

NAND2X1 _1425_ (
    .A(_624_),
    .B(_564_),
    .Y(_631_)
);

NAND3X1 _1005_ (
    .A(_144_),
    .B(_180_),
    .C(_186_),
    .Y(_196_)
);

FILL FILL_3__897_ (
);

INVX1 _756_ (
    .A(Cin_0_bF$buf1),
    .Y(_386_)
);

FILL FILL_1__1167_ (
);

FILL FILL_1__960_ (
);

FILL FILL_2__1236_ (
);

FILL FILL_0__809_ (
);

FILL FILL_3__1305_ (
);

AND2X2 _1234_ (
    .A(_336_),
    .B(_355_),
    .Y(_426_)
);

FILL FILL_0__982_ (
);

AOI21X1 _985_ (
    .A(_171_),
    .B(_175_),
    .C(_158_),
    .Y(_176_)
);

FILL FILL_1__1396_ (
);

FILL FILL_2__803_ (
);

FILL FILL_2__1465_ (
);

FILL FILL_2__1045_ (
);

FILL FILL_3__1114_ (
);

INVX1 _1463_ (
    .A(_634_),
    .Y(_672_)
);

OAI21X1 _1043_ (
    .A(_147_),
    .B(_232_),
    .C(_150_),
    .Y(_233_)
);

FILL FILL_0__791_ (
);

FILL FILL_1__825_ (
);

INVX1 _794_ (
    .A(_735_),
    .Y(_736_)
);

FILL FILL_0__1503_ (
);

FILL FILL_2__1274_ (
);

XOR2X1 _1519_ (
    .A(_730_),
    .B(_72_),
    .Y(_752_[4])
);

FILL FILL_0__847_ (
);

FILL FILL_3__1343_ (
);

AOI21X1 _1272_ (
    .A(_454_),
    .B(_457_),
    .C(_442_),
    .Y(_467_)
);

FILL FILL_4__778_ (
);

FILL FILL_0__1312_ (
);

FILL FILL_2__841_ (
);

FILL FILL_2__1083_ (
);

NAND2X1 _1328_ (
    .A(_522_),
    .B(_527_),
    .Y(_528_)
);

FILL FILL_3__1572_ (
);

FILL FILL_3__1152_ (
);

NAND3X1 _1081_ (
    .A(_260_),
    .B(_267_),
    .C(_270_),
    .Y(_271_)
);

FILL FILL_1__863_ (
);

FILL FILL_4__1221_ (
);

FILL FILL_0__1121_ (
);

FILL FILL_2__1139_ (
);

FILL FILL_3__1208_ (
);

DFFPOSX1 _1557_ (
    .D(_753_[13]),
    .CLK(clk_bF$buf5),
    .Q(y[13])
);

OAI21X1 _1137_ (
    .A(_47_),
    .B(_324_),
    .C(_325_),
    .Y(_326_)
);

FILL FILL_0__885_ (
);

FILL FILL_1__919_ (
);

FILL FILL_3__1381_ (
);

OAI21X1 _888_ (
    .A(_741_),
    .B(_79_),
    .C(_59_),
    .Y(_80_)
);

FILL FILL_1__1299_ (
);

FILL FILL_2__1368_ (
);

FILL FILL_0__1350_ (
);

FILL FILL_3__821_ (
);

FILL FILL_1__1511_ (
);

FILL FILL_3__1437_ (
);

FILL FILL_3__1017_ (
);

AOI21X1 _1366_ (
    .A(_498_),
    .B(_556_),
    .C(_567_),
    .Y(_568_)
);

FILL FILL_3__1190_ (
);

FILL FILL_0__1406_ (
);

FILL FILL_2__935_ (
);

FILL FILL_2__1177_ (
);

FILL FILL_1__1320_ (
);

FILL FILL_3__1246_ (
);

AOI21X1 _1175_ (
    .A(Cin[1]),
    .B(Xin[7]),
    .C(Yin[8]),
    .Y(_364_)
);

FILL FILL_1__957_ (
);

FILL FILL_0__1215_ (
);

FILL FILL_0__979_ (
);

FILL FILL_3__1475_ (
);

FILL FILL_3__1055_ (
);

FILL FILL_1__766_ (
);

FILL FILL_4__1124_ (
);

FILL FILL_0__1444_ (
);

FILL FILL_0__1024_ (
);

FILL FILL_2__973_ (
);

FILL FILL_3__915_ (
);

FILL FILL_0__788_ (
);

FILL FILL_3__1284_ (
);

FILL FILL_1__995_ (
);

FILL FILL_0__1253_ (
);

FILL FILL_2__782_ (
);

FILL FILL_1__1414_ (
);

NAND3X1 _1269_ (
    .A(_458_),
    .B(_463_),
    .C(_439_),
    .Y(_464_)
);

FILL FILL_3__1093_ (
);

FILL FILL_0__1309_ (
);

FILL FILL_2__838_ (
);

FILL FILL_0__1482_ (
);

FILL FILL_0__1062_ (
);

FILL FILL_3__953_ (
);

NAND3X1 _812_ (
    .A(_1_),
    .B(_0_),
    .C(_4_),
    .Y(_5_)
);

FILL FILL_1__1223_ (
);

FILL FILL_3__1569_ (
);

FILL FILL_3__1149_ (
);

NAND2X1 _1498_ (
    .A(Yin[13]),
    .B(_682_),
    .Y(_710_)
);

NAND2X1 _1078_ (
    .A(Yin[7]),
    .B(_265_),
    .Y(_268_)
);

FILL FILL_0__1118_ (
);

FILL FILL_4__1391_ (
);

FILL FILL_0__1291_ (
);

FILL FILL_3__762_ (
);

FILL FILL_1__1452_ (
);

FILL FILL_1__1032_ (
);

FILL FILL_3__1378_ (
);

FILL FILL_2__1101_ (
);

FILL FILL_4__1447_ (
);

FILL FILL_0__1347_ (
);

FILL FILL_2__876_ (
);

FILL FILL_3__818_ (
);

FILL FILL_1__1508_ (
);

FILL FILL_3__991_ (
);

NAND3X1 _850_ (
    .A(_30_),
    .B(_33_),
    .C(_32_),
    .Y(_42_)
);

FILL FILL_1__1261_ (
);

FILL FILL_3__1187_ (
);

FILL FILL_1__898_ (
);

FILL FILL_2__1330_ (
);

FILL FILL_0__1576_ (
);

FILL FILL_0__1156_ (
);

FILL FILL_0__903_ (
);

NAND3X1 _906_ (
    .A(Cin_0_bF$buf3),
    .B(Xin_5_bF$buf0),
    .C(Yin[5]),
    .Y(_98_)
);

FILL FILL_1__1317_ (
);

FILL FILL_4__834_ (
);

FILL FILL_1__1490_ (
);

FILL FILL_1__1070_ (
);

FILL FILL_0__1385_ (
);

FILL FILL_3__856_ (
);

FILL FILL_1__1126_ (
);

FILL FILL_0__1194_ (
);

FILL FILL_0__941_ (
);

XOR2X1 _944_ (
    .A(_135_),
    .B(_73_),
    .Y(_753_[5])
);

FILL FILL_1__1355_ (
);

FILL FILL_2__1424_ (
);

FILL FILL_2__1004_ (
);

FILL FILL_2__779_ (
);

NAND3X1 _1422_ (
    .A(_494_),
    .B(_311_),
    .C(_627_),
    .Y(_628_)
);

INVX1 _1002_ (
    .A(_116_),
    .Y(_193_)
);

FILL FILL_3__894_ (
);

FILL FILL_1__1164_ (
);

FILL FILL_2__1233_ (
);

FILL FILL_4__1579_ (
);

FILL FILL_0__1479_ (
);

FILL FILL_0__1059_ (
);

FILL FILL_0__806_ (
);

FILL FILL_3__1302_ (
);

INVX1 _809_ (
    .A(Yin[3]),
    .Y(_2_)
);

AND2X2 _1231_ (
    .A(Xin[4]),
    .B(Cin[6]),
    .Y(_423_)
);

NAND3X1 _982_ (
    .A(_168_),
    .B(_167_),
    .C(_169_),
    .Y(_173_)
);

FILL FILL_1__1393_ (
);

FILL FILL_2__800_ (
);

FILL FILL_2__1462_ (
);

FILL FILL_2__1042_ (
);

FILL FILL_0__1288_ (
);

FILL FILL_3__759_ (
);

FILL FILL_3__1111_ (
);

FILL FILL_1__1449_ (
);

FILL FILL_1__1029_ (
);

NAND3X1 _1460_ (
    .A(_669_),
    .B(_665_),
    .C(_663_),
    .Y(_670_)
);

NAND3X1 _1040_ (
    .A(_220_),
    .B(_228_),
    .C(_229_),
    .Y(_230_)
);

FILL FILL_1__822_ (
);

INVX1 _791_ (
    .A(_708_),
    .Y(_733_)
);

FILL FILL_2__1518_ (
);

FILL FILL_0__1500_ (
);

FILL FILL_2__1271_ (
);

FILL FILL_0__1097_ (
);

NAND3X1 _1516_ (
    .A(_715_),
    .B(_727_),
    .C(_726_),
    .Y(_728_)
);

FILL FILL_0__844_ (
);

FILL FILL_3__988_ (
);

FILL FILL_3__1340_ (
);

INVX1 _847_ (
    .A(_1_),
    .Y(_39_)
);

FILL FILL_1__1258_ (
);

FILL FILL88950x150 (
);

FILL FILL_2__1327_ (
);

FILL FILL_2__1080_ (
);

NAND3X1 _1325_ (
    .A(_512_),
    .B(_507_),
    .C(_520_),
    .Y(_524_)
);

FILL FILL_3__797_ (
);

FILL FILL_1__1487_ (
);

FILL FILL_1__1067_ (
);

FILL FILL_1__860_ (
);

FILL FILL_2__1136_ (
);

FILL FILL_3_BUFX2_insert10 (
);

FILL FILL_3_BUFX2_insert11 (
);

FILL FILL_3_BUFX2_insert12 (
);

FILL FILL_3_BUFX2_insert13 (
);

FILL FILL_3_BUFX2_insert14 (
);

FILL FILL_3_BUFX2_insert15 (
);

FILL FILL_3_BUFX2_insert16 (
);

FILL FILL_3_BUFX2_insert17 (
);

FILL FILL_3__1205_ (
);

DFFPOSX1 _1554_ (
    .D(_753_[10]),
    .CLK(clk_bF$buf5),
    .Q(y[10])
);

NAND2X1 _1134_ (
    .A(_321_),
    .B(_322_),
    .Y(_323_)
);

FILL FILL_0__882_ (
);

FILL FILL_1__916_ (
);

INVX1 _885_ (
    .A(Cin[5]),
    .Y(_77_)
);

FILL FILL_1__1296_ (
);

FILL FILL_2__1365_ (
);

FILL FILL_0__938_ (
);

FILL FILL_3__1434_ (
);

FILL FILL_3__1014_ (
);

XOR2X1 _1363_ (
    .A(_495_),
    .B(_565_),
    .Y(_753_[10])
);

FILL FILL_0__1403_ (
);

FILL FILL_2__932_ (
);

FILL FILL_2__1174_ (
);

INVX1 _1419_ (
    .A(_625_),
    .Y(_626_)
);

FILL FILL_3__1243_ (
);

FILL FILL88350x35250 (
);

OAI21X1 _1172_ (
    .A(_261_),
    .B(_360_),
    .C(_263_),
    .Y(_361_)
);

FILL FILL_1__954_ (
);

FILL FILL_0__1212_ (
);

OAI21X1 _1228_ (
    .A(_416_),
    .B(_419_),
    .C(_415_),
    .Y(_420_)
);

FILL FILL_0__976_ (
);

FILL FILL_3__1472_ (
);

FILL FILL_3__1052_ (
);

AOI21X1 _979_ (
    .A(_169_),
    .B(_168_),
    .C(_167_),
    .Y(_170_)
);

FILL FILL_1__763_ (
);

FILL FILL_2__1459_ (
);

FILL FILL_0__1441_ (
);

FILL FILL_0__1021_ (
);

FILL FILL_2__1039_ (
);

FILL FILL_2__970_ (
);

FILL FILL_3__912_ (
);

FILL FILL_3__1108_ (
);

NAND2X1 _1457_ (
    .A(_665_),
    .B(_663_),
    .Y(_667_)
);

NAND2X1 _1037_ (
    .A(Xin[2]),
    .B(Cin[5]),
    .Y(_227_)
);

FILL FILL_0__785_ (
);

FILL FILL_1__819_ (
);

FILL FILL_3__1281_ (
);

INVX1 _788_ (
    .A(_718_),
    .Y(_729_)
);

FILL FILL_1__1199_ (
);

FILL FILL_1__992_ (
);

FILL FILL_4__1350_ (
);

FILL FILL_0__1250_ (
);

FILL FILL_2__1268_ (
);

FILL FILL_1__1411_ (
);

FILL FILL_3__1337_ (
);

FILL FILL88650x74250 (
);

AOI21X1 _1266_ (
    .A(_377_),
    .B(_372_),
    .C(_459_),
    .Y(_460_)
);

FILL FILL_3__1090_ (
);

FILL FILL_0__1306_ (
);

FILL FILL_2__835_ (
);

FILL FILL_2__1497_ (
);

FILL FILL_2__1077_ (
);

FILL FILL_3__950_ (
);

FILL FILL_1__1220_ (
);

FILL FILL_3__1566_ (
);

FILL FILL_3__1146_ (
);

OAI21X1 _1495_ (
    .A(_677_),
    .B(_705_),
    .C(_704_),
    .Y(_706_)
);

NAND2X1 _1075_ (
    .A(Cin_0_bF$buf0),
    .B(Xin[7]),
    .Y(_265_)
);

FILL FILL_1__857_ (
);

FILL FILL_0__1115_ (
);

FILL FILL_0__879_ (
);

FILL FILL_3__1375_ (
);

FILL FILL_0__1344_ (
);

FILL FILL_2__873_ (
);

FILL FILL_3__815_ (
);

FILL FILL_1__1505_ (
);

FILL FILL_3__1184_ (
);

FILL FILL_1__895_ (
);

FILL FILL_2__929_ (
);

FILL FILL_4__1253_ (
);

FILL FILL_0__1573_ (
);

FILL FILL_0__1153_ (
);

FILL FILL_0__900_ (
);

OAI21X1 _903_ (
    .A(_33_),
    .B(_31_),
    .C(_30_),
    .Y(_95_)
);

FILL FILL_1__1314_ (
);

NAND3X1 _1169_ (
    .A(_348_),
    .B(_356_),
    .C(_357_),
    .Y(_358_)
);

FILL FILL_4__1309_ (
);

FILL FILL_0__1209_ (
);

FILL FILL_0__1382_ (
);

FILL FILL_3__853_ (
);

FILL FILL89550x4050 (
);

FILL FILL_1__1123_ (
);

FILL FILL_3__1469_ (
);

FILL FILL_3__1049_ (
);

INVX1 _1398_ (
    .A(_602_),
    .Y(_603_)
);

FILL FILL_0__1438_ (
);

FILL FILL_0__1018_ (
);

FILL FILL_2__967_ (
);

FILL FILL_3__909_ (
);

FILL FILL_0__1191_ (
);

AOI22X1 _941_ (
    .A(_127_),
    .B(_131_),
    .C(_72_),
    .D(_21_),
    .Y(_133_)
);

FILL FILL88350x23550 (
);

FILL FILL_1__1352_ (
);

FILL FILL_3__1278_ (
);

FILL FILL_1__989_ (
);

FILL FILL_2__1421_ (
);

FILL FILL_2__1001_ (
);

FILL FILL_0__1247_ (
);

FILL FILL_2__776_ (
);

FILL FILL_1__1408_ (
);

FILL FILL_3__891_ (
);

FILL FILL_1__1581_ (
);

FILL FILL_1__1161_ (
);

FILL FILL_3__1087_ (
);

FILL FILL_1__798_ (
);

FILL FILL_2__1230_ (
);

FILL FILL_0__1476_ (
);

FILL FILL_0__1056_ (
);

FILL FILL_0__803_ (
);

FILL FILL_3__947_ (
);

NAND2X1 _806_ (
    .A(Cin[1]),
    .B(Xin[2]),
    .Y(_747_)
);

FILL FILL_1__1217_ (
);

FILL FILL_1__1390_ (
);

FILL FILL_0_BUFX2_insert6 (
);

FILL FILL_0_BUFX2_insert7 (
);

FILL FILL_0_BUFX2_insert8 (
);

FILL FILL_0_BUFX2_insert9 (
);

FILL FILL_0__1285_ (
);

FILL FILL_3__756_ (
);

FILL FILL_1__1446_ (
);

FILL FILL_1__1026_ (
);

FILL FILL_4__963_ (
);

FILL FILL_2__1515_ (
);

FILL FILL_0__1094_ (
);

AND2X2 _1513_ (
    .A(_699_),
    .B(_695_),
    .Y(_725_)
);

FILL FILL_0__841_ (
);

FILL FILL_3__985_ (
);

INVX1 _844_ (
    .A(_30_),
    .Y(_36_)
);

FILL FILL_1__1255_ (
);

FILL FILL_2__1324_ (
);

OAI21X1 _1322_ (
    .A(_517_),
    .B(_518_),
    .C(_520_),
    .Y(_521_)
);

FILL FILL_3__794_ (
);

FILL FILL_1__1484_ (
);

FILL FILL_1__1064_ (
);

FILL FILL_2__1133_ (
);

FILL FILL_4__1479_ (
);

FILL FILL_0__1379_ (
);

FILL FILL_3__1202_ (
);

DFFPOSX1 _1551_ (
    .D(_753_[7]),
    .CLK(clk_bF$buf0),
    .Q(y[7])
);

INVX1 _1131_ (
    .A(_319_),
    .Y(_320_)
);

FILL FILL_1__913_ (
);

NAND3X1 _882_ (
    .A(_68_),
    .B(_21_),
    .C(_71_),
    .Y(_74_)
);

FILL FILL_1__1293_ (
);

FILL FILL_2_BUFX2_insert6 (
);

FILL FILL_2_BUFX2_insert7 (
);

FILL FILL_2_BUFX2_insert8 (
);

FILL FILL_2_BUFX2_insert9 (
);

FILL FILL_2__1362_ (
);

FILL FILL_0__1188_ (
);

FILL FILL_0__935_ (
);

FILL FILL_3__1431_ (
);

FILL FILL_3__1011_ (
);

AOI21X1 _938_ (
    .A(_120_),
    .B(_116_),
    .C(_81_),
    .Y(_130_)
);

FILL FILL_1__1349_ (
);

NAND3X1 _1360_ (
    .A(_499_),
    .B(_553_),
    .C(_549_),
    .Y(_563_)
);

FILL FILL_4__866_ (
);

FILL FILL_0__1400_ (
);

FILL FILL_2__1418_ (
);

FILL FILL_2__1171_ (
);

FILL FILL_4__1097_ (
);

NAND3X1 _1416_ (
    .A(_571_),
    .B(_613_),
    .C(_609_),
    .Y(_622_)
);

FILL FILL_3__888_ (
);

FILL FILL_3__1240_ (
);

FILL FILL88650x39150 (
);

FILL FILL_1__1578_ (
);

FILL FILL_1__1158_ (
);

FILL FILL_1__951_ (
);

FILL FILL_2__1227_ (
);

AOI22X1 _1225_ (
    .A(Xin_3_bF$buf3),
    .B(Cin[6]),
    .C(Xin[4]),
    .D(Cin[5]),
    .Y(_416_)
);

FILL FILL_0__973_ (
);

INVX1 _976_ (
    .A(_161_),
    .Y(_167_)
);

FILL FILL_1__1387_ (
);

FILL FILL_1__760_ (
);

FILL FILL_2__1456_ (
);

FILL FILL_2__1036_ (
);

FILL FILL_3__1105_ (
);

OAI21X1 _1454_ (
    .A(_662_),
    .B(_661_),
    .C(_636_),
    .Y(_663_)
);

NAND2X1 _1034_ (
    .A(Xin[1]),
    .B(Cin[6]),
    .Y(_224_)
);

FILL FILL_0__782_ (
);

FILL FILL_1__816_ (
);

OAI21X1 _785_ (
    .A(_655_),
    .B(_687_),
    .C(_623_),
    .Y(_697_)
);

FILL FILL_1__1196_ (
);

FILL FILL_4_BUFX2_insert8 (
);

FILL FILL_2__1265_ (
);

FILL FILL_0__838_ (
);

FILL FILL_3__1334_ (
);

FILL FILL88950x78150 (
);

NAND2X1 _1263_ (
    .A(_456_),
    .B(_455_),
    .Y(_457_)
);

FILL FILL_4__769_ (
);

FILL FILL_0__1303_ (
);

FILL FILL_2__832_ (
);

FILL FILL_2__1494_ (
);

FILL FILL_2__1074_ (
);

NOR3X1 _1319_ (
    .A(_502_),
    .B(_506_),
    .C(_505_),
    .Y(_518_)
);

FILL FILL_3__1563_ (
);

FILL FILL_3__1143_ (
);

NAND3X1 _1492_ (
    .A(Yin[14]),
    .B(_576_),
    .C(_678_),
    .Y(_703_)
);

INVX1 _1072_ (
    .A(_261_),
    .Y(_262_)
);

FILL FILL_1__854_ (
);

FILL FILL_4__1212_ (
);

FILL FILL_0__1112_ (
);

DFFPOSX1 _1548_ (
    .D(_752_[4]),
    .CLK(clk_bF$buf3),
    .Q(y[4])
);

OAI21X1 _1128_ (
    .A(_288_),
    .B(_316_),
    .C(_281_),
    .Y(_317_)
);

FILL FILL_0__876_ (
);

FILL FILL_3__1372_ (
);

OAI21X1 _879_ (
    .A(_69_),
    .B(_70_),
    .C(_744_),
    .Y(_71_)
);

FILL FILL_2__1359_ (
);

FILL FILL_0__1341_ (
);

FILL FILL_2__870_ (
);

FILL FILL_3__812_ (
);

FILL FILL_1__1502_ (
);

FILL FILL_3__1428_ (
);

FILL FILL_3__1008_ (
);

AOI21X1 _1357_ (
    .A(_468_),
    .B(_464_),
    .C(_412_),
    .Y(_560_)
);

FILL FILL_3__1181_ (
);

FILL FILL_1__1099_ (
);

FILL FILL_1__892_ (
);

FILL FILL_2__926_ (
);

FILL FILL_0__1570_ (
);

FILL FILL_0__1150_ (
);

FILL FILL_2__1168_ (
);

NAND3X1 _900_ (
    .A(Xin[2]),
    .B(Cin[3]),
    .C(_91_),
    .Y(_92_)
);

FILL FILL_1__1311_ (
);

FILL FILL_3__1237_ (
);

FILL FILL88050x7950 (
);

NAND2X1 _1166_ (
    .A(Cin[2]),
    .B(Xin[6]),
    .Y(_355_)
);

FILL FILL_1__948_ (
);

FILL FILL_0__1206_ (
);

FILL FILL_2__1397_ (
);

FILL FILL_3__850_ (
);

FILL FILL_1__1120_ (
);

FILL FILL_3__1466_ (
);

FILL FILL_3__1046_ (
);

CLKBUF1 CLKBUF1_insert0 (
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert1 (
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert2 (
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert3 (
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert4 (
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert5 (
    .A(clk),
    .Y(clk_bF$buf0)
);

NAND2X1 _1395_ (
    .A(_598_),
    .B(_534_),
    .Y(_599_)
);

FILL FILL_1__757_ (
);

FILL FILL_4__1115_ (
);

FILL FILL_0__1435_ (
);

FILL FILL_0__1015_ (
);

FILL FILL_2__964_ (
);

FILL FILL_3__906_ (
);

FILL FILL_0__779_ (
);

FILL FILL_3__1275_ (
);

FILL FILL_1__986_ (
);

FILL FILL88350x85950 (
);

FILL FILL_0__1244_ (
);

FILL FILL_2__773_ (
);

FILL FILL_1__1405_ (
);

FILL FILL_3__1084_ (
);

FILL FILL_1__795_ (
);

FILL FILL_2__829_ (
);

FILL FILL_0__1473_ (
);

FILL FILL_0__1053_ (
);

FILL FILL_0__800_ (
);

FILL FILL_3__944_ (
);

NAND2X1 _803_ (
    .A(_743_),
    .B(_601_),
    .Y(_744_)
);

FILL FILL_1__1214_ (
);

AOI22X1 _1489_ (
    .A(_695_),
    .B(_699_),
    .C(_634_),
    .D(_698_),
    .Y(_700_)
);

AOI21X1 _1069_ (
    .A(Cin_0_bF$buf0),
    .B(Xin[6]),
    .C(Yin[6]),
    .Y(_259_)
);

FILL FILL_0__1109_ (
);

FILL FILL_4__1382_ (
);

FILL FILL_0__1282_ (
);

FILL FILL_1__1443_ (
);

FILL FILL_1__1023_ (
);

FILL FILL_3__1369_ (
);

AOI21X1 _1298_ (
    .A(_311_),
    .B(_494_),
    .C(_492_),
    .Y(_495_)
);

FILL FILL_2__1512_ (
);

FILL FILL_4__1018_ (
);

FILL FILL_0__1338_ (
);

FILL FILL_2__867_ (
);

FILL FILL_3__809_ (
);

FILL FILL_0__1091_ (
);

NAND2X1 _1510_ (
    .A(_721_),
    .B(_716_),
    .Y(_722_)
);

FILL FILL_3__982_ (
);

NAND2X1 _841_ (
    .A(Cin[1]),
    .B(Xin_3_bF$buf2),
    .Y(_33_)
);

FILL FILL_1__1252_ (
);

FILL FILL_3__1178_ (
);

FILL FILL_1__889_ (
);

FILL FILL_2__1321_ (
);

FILL FILL_0__1567_ (
);

FILL FILL_0__1147_ (
);

FILL FILL_1__1308_ (
);

FILL FILL_3__791_ (
);

FILL FILL_1__1481_ (
);

FILL FILL_1__1061_ (
);

FILL FILL_2__1130_ (
);

FILL FILL_0__1376_ (
);

FILL FILL_3__847_ (
);

FILL FILL_1__1117_ (
);

FILL FILL_1__910_ (
);

FILL FILL_1__1290_ (
);

FILL FILL_4__1285_ (
);

FILL FILL_0__1185_ (
);

FILL FILL_0__932_ (
);

NAND3X1 _935_ (
    .A(_121_),
    .B(_126_),
    .C(_76_),
    .Y(_127_)
);

FILL FILL_1__1346_ (
);

FILL FILL_2__1415_ (
);

AOI21X1 _1413_ (
    .A(_552_),
    .B(_551_),
    .C(_500_),
    .Y(_619_)
);

FILL FILL_3__885_ (
);

FILL FILL_1__1575_ (
);

FILL FILL_1__1155_ (
);

FILL FILL_2__1224_ (
);

FILL FILL_2__999_ (
);

FILL FILL88650x15750 (
);

NAND2X1 _1222_ (
    .A(Xin_3_bF$buf3),
    .B(Cin[6]),
    .Y(_413_)
);

FILL FILL_0__970_ (
);

INVX1 _973_ (
    .A(Yin[6]),
    .Y(_164_)
);

FILL FILL_1__1384_ (
);

FILL FILL_2__1453_ (
);

FILL FILL_2__1033_ (
);

FILL FILL_0__1279_ (
);

FILL FILL_3__1102_ (
);

NAND2X1 _1451_ (
    .A(_637_),
    .B(_659_),
    .Y(_660_)
);

INVX1 _1031_ (
    .A(_220_),
    .Y(_221_)
);

FILL FILL_1__813_ (
);

INVX1 _782_ (
    .A(_655_),
    .Y(_666_)
);

FILL FILL_1__1193_ (
);

FILL FILL_2__1509_ (
);

FILL FILL_2__1262_ (
);

FILL FILL_0__1088_ (
);

OAI21X1 _1507_ (
    .A(Yin[14]),
    .B(_677_),
    .C(_678_),
    .Y(_719_)
);

FILL FILL_0__835_ (
);

FILL FILL_3__979_ (
);

FILL FILL_3__1331_ (
);

NAND3X1 _838_ (
    .A(Cin_0_bF$buf2),
    .B(Xin[4]),
    .C(Yin[4]),
    .Y(_30_)
);

FILL FILL_1__1249_ (
);

NAND3X1 _1260_ (
    .A(_453_),
    .B(_449_),
    .C(_452_),
    .Y(_454_)
);

FILL FILL_2__1318_ (
);

FILL FILL_0__1300_ (
);

FILL FILL_2__1491_ (
);

FILL FILL_2__1071_ (
);

FILL FILL88950x54750 (
);

OAI21X1 _1316_ (
    .A(_443_),
    .B(_513_),
    .C(_446_),
    .Y(_514_)
);

FILL FILL_3__788_ (
);

FILL FILL_3__1560_ (
);

FILL FILL_3__1140_ (
);

FILL FILL_1__1478_ (
);

FILL FILL_1__1058_ (
);

FILL FILL_1__851_ (
);

FILL FILL_4__995_ (
);

FILL FILL_2__1127_ (
);

DFFPOSX1 _1545_ (
    .D(_749_[1]),
    .CLK(clk_bF$buf4),
    .Q(y[1])
);

NAND2X1 _1125_ (
    .A(_234_),
    .B(_240_),
    .Y(_314_)
);

FILL FILL_0__873_ (
);

FILL FILL_1__907_ (
);

NAND3X1 _876_ (
    .A(_26_),
    .B(_63_),
    .C(_67_),
    .Y(_68_)
);

FILL FILL_1__1287_ (
);

FILL FILL_2__1356_ (
);

FILL FILL_0__929_ (
);

FILL FILL_3__1425_ (
);

FILL FILL_3__1005_ (
);

OAI21X1 _1354_ (
    .A(_541_),
    .B(_547_),
    .C(_550_),
    .Y(_556_)
);

FILL FILL_1__1096_ (
);

FILL FILL_2__923_ (
);

FILL FILL_2__1165_ (
);

FILL FILL_3__1234_ (
);

BUFX2 _1583_ (
    .A(_755_[9]),
    .Y(Yout[9])
);

INVX1 _1163_ (
    .A(Xin[6]),
    .Y(_352_)
);

FILL FILL_1__945_ (
);

FILL FILL_0__1203_ (
);

FILL FILL_2__1394_ (
);

NAND2X1 _1219_ (
    .A(_333_),
    .B(_340_),
    .Y(_410_)
);

FILL FILL_0__967_ (
);

FILL FILL_3__1463_ (
);

FILL FILL_3__1043_ (
);

OAI21X1 _1392_ (
    .A(_591_),
    .B(_589_),
    .C(_536_),
    .Y(_596_)
);

FILL FILL_4__898_ (
);

FILL FILL_0__1432_ (
);

FILL FILL_0__1012_ (
);

FILL FILL_2__961_ (
);

FILL FILL_3__903_ (
);

FILL FILL_3__1519_ (
);

NAND2X1 _1448_ (
    .A(_656_),
    .B(_649_),
    .Y(_657_)
);

NAND2X1 _1028_ (
    .A(_140_),
    .B(_78_),
    .Y(_218_)
);

FILL FILL_0__776_ (
);

FILL FILL_3__1272_ (
);

INVX1 _779_ (
    .A(_623_),
    .Y(_633_)
);

FILL FILL_1__983_ (
);

FILL FILL_4__1341_ (
);

endmodule

/* Verilog module written by vlog2Verilog (qflow) */
/* With explicit power connections */

module fir_pe(
    inout vdd,
    inout gnd,
    input [7:0] Cin,
    input Rdy,
    output Vld,
    input [3:0] Xin,
    output [3:0] Xout,
    input [3:0] Yin,
    output [3:0] Yout,
    input clk
);

wire [15:0] y ;
wire _588_ ;
wire _168_ ;
wire _800_ ;
wire _60_ ;
wire _397_ ;
wire _703_ ;
wire _19_ ;
wire _512_ ;
wire [4:0] LoadCtl ;
wire _741_ ;
wire _321_ ;
wire _57_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _835_ ;
wire _415_ ;
wire _95_ ;
wire _148__bF$buf0 ;
wire _148__bF$buf1 ;
wire _148__bF$buf2 ;
wire _148__bF$buf3 ;
wire _148__bF$buf4 ;
wire _644_ ;
wire _224_ ;
wire _873_ ;
wire _453_ ;
wire _509_ ;
wire _682_ ;
wire _262_ ;
wire _738_ ;
wire _318_ ;
wire _491_ ;
wire _547_ ;
wire _127_ ;
wire _776_ ;
wire _356_ ;
wire _585_ ;
wire _165_ ;
wire _394_ ;
wire _679_ ;
wire _259_ ;
wire _488_ ;
wire _700_ ;
wire _297_ ;
wire _16_ ;
wire _54_ ;
wire _603_ ;
wire _832_ ;
wire _412_ ;
wire _92_ ;
wire _641_ ;
wire _221_ ;
wire _870_ ;
wire _450_ ;
wire _506_ ;
wire _735_ ;
wire _315_ ;
wire _544_ ;
wire _124_ ;
wire _773_ ;
wire _353_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _582_ ;
wire _162_ ;
wire _638_ ;
wire _218_ ;
wire _391_ ;
wire _867_ ;
wire _447_ ;
wire _676_ ;
wire _256_ ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire _388_ ;
wire _600_ ;
wire Rdy ;
wire _197_ ;
wire _7_ ;
wire _503_ ;
wire _732_ ;
wire _312_ ;
wire _48_ ;
wire _541_ ;
wire _121_ ;
wire _770_ ;
wire _350_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _635_ ;
wire _215_ ;
wire _864_ ;
wire _444_ ;
wire _673_ ;
wire _253_ ;
wire _729_ ;
wire _309_ ;
wire _482_ ;
wire _538_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _767_ ;
wire _347_ ;
wire _576_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire [7:0] XinHL ;
wire _899_ ;
wire _479_ ;
wire _288_ ;
wire _4_ ;
wire [3:0] _920_ ;
wire _500_ ;
wire _45_ ;
wire _823_ ;
wire _403_ ;
wire _83_ ;
wire _632_ ;
wire _212_ ;
wire _861_ ;
wire _441_ ;
wire _917_ ;
wire _670_ ;
wire _250_ ;
wire _726_ ;
wire _306_ ;
wire _535_ ;
wire _115_ ;
wire _764_ ;
wire _344_ ;
wire _573_ ;
wire _153_ ;
wire _629_ ;
wire _209_ ;
wire _382_ ;
wire _858_ ;
wire _438_ ;
wire _191_ ;
wire _667_ ;
wire _247_ ;
wire _896_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire _285_ ;
wire _1_ ;
wire _42_ ;
wire _799_ ;
wire _379_ ;
wire _188_ ;
wire _820_ ;
wire _400_ ;
wire _80_ ;
wire _914_ ;
wire _723_ ;
wire _303_ ;
wire _39_ ;
wire _532_ ;
wire _112_ ;
wire _761_ ;
wire _341_ ;
wire clk ;
wire _817_ ;
wire _77_ ;
wire _570_ ;
wire _150_ ;
wire _626_ ;
wire _206_ ;
wire _855_ ;
wire _435_ ;
wire _664_ ;
wire _244_ ;
wire _893_ ;
wire _473_ ;
wire _529_ ;
wire _109_ ;
wire _282_ ;
wire _758_ ;
wire _338_ ;
wire _567_ ;
wire _147_ ;
wire _796_ ;
wire _376_ ;
wire _185_ ;
wire _699_ ;
wire _279_ ;
wire _911_ ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire _814_ ;
wire _74_ ;
wire _623_ ;
wire _203_ ;
wire _852_ ;
wire _432_ ;
wire _908_ ;
wire _661_ ;
wire _241_ ;
wire _717_ ;
wire _890_ ;
wire _470_ ;
wire _526_ ;
wire _106_ ;
wire _755_ ;
wire _335_ ;
wire _564_ ;
wire _144_ ;
wire _793_ ;
wire _373_ ;
wire _849_ ;
wire _429_ ;
wire _182_ ;
wire LoadCtl_0_bF$buf0 ;
wire LoadCtl_0_bF$buf1 ;
wire LoadCtl_0_bF$buf2 ;
wire LoadCtl_0_bF$buf3 ;
wire LoadCtl_0_bF$buf4 ;
wire _658_ ;
wire _238_ ;
wire _887_ ;
wire _467_ ;
wire _696_ ;
wire _276_ ;
wire _33_ ;
wire _599_ ;
wire _179_ ;
wire _811_ ;
wire _71_ ;
wire _620_ ;
wire _200_ ;
wire _905_ ;
wire _714_ ;
wire _523_ ;
wire _103_ ;
wire _752_ ;
wire _332_ ;
wire _808_ ;
wire _68_ ;
wire _561_ ;
wire _141_ ;
wire _617_ ;
wire _790_ ;
wire _370_ ;
wire _846_ ;
wire _426_ ;
wire _655_ ;
wire _235_ ;
wire _884_ ;
wire _464_ ;
wire _693_ ;
wire _273_ ;
wire _749_ ;
wire _329_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _787_ ;
wire _367_ ;
wire _596_ ;
wire _176_ ;
wire _902_ ;
wire _499_ ;
wire _711_ ;
wire _27_ ;
wire _520_ ;
wire _100_ ;
wire _805_ ;
wire _65_ ;
wire _614_ ;
wire _843_ ;
wire _423_ ;
wire _652_ ;
wire _232_ ;
wire _708_ ;
wire _881_ ;
wire _461_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _746_ ;
wire _326_ ;
wire _555_ ;
wire _135_ ;
wire _784_ ;
wire _364_ ;
wire _593_ ;
wire _173_ ;
wire _649_ ;
wire _229_ ;
wire _878_ ;
wire _458_ ;
wire _687_ ;
wire _267_ ;
wire _496_ ;
wire _24_ ;
wire _802_ ;
wire _62_ ;
wire _399_ ;
wire _611_ ;
wire _840_ ;
wire _420_ ;
wire _705_ ;
wire [15:0] _y ;
wire _514_ ;
wire _743_ ;
wire _323_ ;
wire _59_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _781_ ;
wire _361_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _646_ ;
wire _226_ ;
wire _875_ ;
wire _455_ ;
wire _684_ ;
wire _264_ ;
wire _493_ ;
wire _549_ ;
wire _129_ ;
wire _21_ ;
wire _778_ ;
wire _358_ ;
wire _587_ ;
wire _167_ ;
wire _396_ ;
wire _702_ ;
wire _299_ ;
wire _18_ ;
wire _511_ ;
wire _740_ ;
wire _320_ ;
wire _56_ ;
wire _605_ ;
wire _834_ ;
wire _414_ ;
wire _94_ ;
wire _643_ ;
wire _223_ ;
wire _872_ ;
wire _452_ ;
wire _508_ ;
wire _681_ ;
wire _261_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _546_ ;
wire _126_ ;
wire _775_ ;
wire _355_ ;
wire _584_ ;
wire _164_ ;
wire _393_ ;
wire _869_ ;
wire _449_ ;
wire _678_ ;
wire _258_ ;
wire _487_ ;
wire _296_ ;
wire _15_ ;
wire _53_ ;
wire _602_ ;
wire _199_ ;
wire _831_ ;
wire _411_ ;
wire _91_ ;
wire _640_ ;
wire _220_ ;
wire _9_ ;
wire _505_ ;
wire _734_ ;
wire _314_ ;
wire _543_ ;
wire _123_ ;
wire _772_ ;
wire _352_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _581_ ;
wire _161_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _866_ ;
wire _446_ ;
wire [3:0] Yin ;
wire _675_ ;
wire _255_ ;
wire _484_ ;
wire _293_ ;
wire _12_ ;
wire _769_ ;
wire _349_ ;
wire _578_ ;
wire _158_ ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire _6_ ;
wire _502_ ;
wire _731_ ;
wire _311_ ;
wire _47_ ;
wire _540_ ;
wire _120_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire [3:0] Yin0 ;
wire [3:0] Yin1 ;
wire [3:0] Yin2 ;
wire [3:0] Yin3 ;
wire _634_ ;
wire _214_ ;
wire _863_ ;
wire _443_ ;
wire _919_ ;
wire _672_ ;
wire _252_ ;
wire _728_ ;
wire _308_ ;
wire _481_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _766_ ;
wire _346_ ;
wire _575_ ;
wire _155_ ;
wire _384_ ;
wire _193_ ;
wire _669_ ;
wire _249_ ;
wire _898_ ;
wire _478_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _822_ ;
wire _402_ ;
wire _82_ ;
wire _631_ ;
wire _211_ ;
wire _860_ ;
wire _440_ ;
wire _916_ ;
wire _725_ ;
wire _305_ ;
wire [3:0] XinH ;
wire _534_ ;
wire _114_ ;
wire _763_ ;
wire _343_ ;
wire _819_ ;
wire _79_ ;
wire _572_ ;
wire _152_ ;
wire _628_ ;
wire _208_ ;
wire _381_ ;
wire _857_ ;
wire _437_ ;
wire _190_ ;
wire _666_ ;
wire _246_ ;
wire _895_ ;
wire _475_ ;
wire _284_ ;
wire _0_ ;
wire _569_ ;
wire _149_ ;
wire _41_ ;
wire _798_ ;
wire _378_ ;
wire _187_ ;
wire [3:0] Yout ;
wire _913_ ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _531_ ;
wire _111_ ;
wire _760_ ;
wire _340_ ;
wire _816_ ;
wire _76_ ;
wire _625_ ;
wire _205_ ;
wire _854_ ;
wire _434_ ;
wire _663_ ;
wire _243_ ;
wire _719_ ;
wire _892_ ;
wire _472_ ;
wire _528_ ;
wire _108_ ;
wire _281_ ;
wire _757_ ;
wire _337_ ;
wire _566_ ;
wire _146_ ;
wire _795_ ;
wire _375_ ;
wire _184_ ;
wire _889_ ;
wire _469_ ;
wire _698_ ;
wire _278_ ;
wire _910_ ;
wire _35_ ;
wire [3:0] Xout ;
wire _813_ ;
wire _73_ ;
wire _622_ ;
wire _202_ ;
wire _851_ ;
wire _431_ ;
wire _907_ ;
wire _660_ ;
wire _240_ ;
wire _716_ ;
wire _525_ ;
wire _105_ ;
wire _754_ ;
wire _334_ ;
wire _563_ ;
wire _143_ ;
wire _619_ ;
wire _792_ ;
wire _372_ ;
wire _848_ ;
wire _428_ ;
wire _181_ ;
wire _657_ ;
wire _237_ ;
wire _886_ ;
wire _466_ ;
wire _695_ ;
wire _275_ ;
wire _32_ ;
wire _789_ ;
wire _369_ ;
wire _598_ ;
wire _178_ ;
wire _810_ ;
wire _70_ ;
wire LoadCtl_4_bF$buf0 ;
wire LoadCtl_4_bF$buf1 ;
wire LoadCtl_4_bF$buf2 ;
wire LoadCtl_4_bF$buf3 ;
wire LoadCtl_4_bF$buf4 ;
wire _904_ ;
wire _713_ ;
wire _29_ ;
wire _522_ ;
wire _102_ ;
wire _751_ ;
wire _331_ ;
wire _807_ ;
wire _67_ ;
wire _560_ ;
wire _140_ ;
wire _616_ ;
wire _845_ ;
wire _425_ ;
wire _654_ ;
wire _234_ ;
wire _883_ ;
wire _463_ ;
wire _519_ ;
wire _692_ ;
wire _272_ ;
wire _748_ ;
wire _328_ ;
wire _557_ ;
wire _137_ ;
wire _786_ ;
wire _366_ ;
wire _595_ ;
wire _175_ ;
wire _689_ ;
wire _269_ ;
wire _901_ ;
wire _498_ ;
wire _710_ ;
wire _26_ ;
wire Cin_0_bF$buf0 ;
wire Cin_0_bF$buf1 ;
wire Cin_0_bF$buf2 ;
wire Cin_0_bF$buf3 ;
wire _804_ ;
wire _64_ ;
wire _613_ ;
wire _842_ ;
wire _422_ ;
wire _651_ ;
wire _231_ ;
wire _707_ ;
wire _880_ ;
wire _460_ ;
wire _516_ ;
wire _745_ ;
wire _325_ ;
wire _554_ ;
wire _134_ ;
wire _783_ ;
wire _363_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _592_ ;
wire _172_ ;
wire Vld ;
wire _648_ ;
wire _228_ ;
wire _877_ ;
wire _457_ ;
wire _686_ ;
wire _266_ ;
wire _495_ ;
wire _23_ ;
wire _589_ ;
wire _169_ ;
wire _801_ ;
wire _61_ ;
wire _398_ ;
wire _610_ ;
wire _704_ ;
wire _513_ ;
wire _742_ ;
wire _322_ ;
wire _58_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _780_ ;
wire _360_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire [7:0] Cin ;
wire _645_ ;
wire _225_ ;
wire _874_ ;
wire _454_ ;
wire _683_ ;
wire _263_ ;
wire _739_ ;
wire _319_ ;
wire _492_ ;
wire _548_ ;
wire _128_ ;
wire _20_ ;
wire _777_ ;
wire _357_ ;
wire _586_ ;
wire _166_ ;
wire _395_ ;
wire _489_ ;
wire _701_ ;
wire _298_ ;
wire _17_ ;
wire _510_ ;
wire _55_ ;
wire _604_ ;
wire _833_ ;
wire _413_ ;
wire _93_ ;
wire _642_ ;
wire _222_ ;
wire _871_ ;
wire _451_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _736_ ;
wire _316_ ;
wire _545_ ;
wire _125_ ;
wire _774_ ;
wire _354_ ;
wire _583_ ;
wire _163_ ;
wire _639_ ;
wire _219_ ;
wire _392_ ;
wire _868_ ;
wire _448_ ;
wire _677_ ;
wire _257_ ;
wire _486_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _601_ ;
wire _198_ ;
wire _830_ ;
wire _410_ ;
wire _90_ ;
wire _8_ ;
wire _504_ ;
wire _733_ ;
wire _313_ ;
wire _49_ ;
wire _542_ ;
wire _122_ ;
wire _771_ ;
wire _351_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _636_ ;
wire _216_ ;
wire _865_ ;
wire _445_ ;
wire _674_ ;
wire _254_ ;
wire _483_ ;
wire _539_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _768_ ;
wire _348_ ;
wire _577_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire _289_ ;
wire _5_ ;
wire [3:0] _921_ ;
wire _501_ ;
wire _730_ ;
wire _310_ ;
wire _46_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _633_ ;
wire _213_ ;
wire _862_ ;
wire _442_ ;
wire _918_ ;
wire _671_ ;
wire _251_ ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire _536_ ;
wire _116_ ;
wire _765_ ;
wire _345_ ;
wire _574_ ;
wire _154_ ;
wire _383_ ;
wire _859_ ;
wire _439_ ;
wire _192_ ;
wire _668_ ;
wire _248_ ;
wire _897_ ;
wire _477_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire _189_ ;
wire _821_ ;
wire _401_ ;
wire _81_ ;
wire _630_ ;
wire _210_ ;
wire _915_ ;
wire _724_ ;
wire _304_ ;
wire _533_ ;
wire _113_ ;
wire _762_ ;
wire _342_ ;
wire _818_ ;
wire _78_ ;
wire _571_ ;
wire _151_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _856_ ;
wire _436_ ;
wire [3:0] Xin ;
wire _665_ ;
wire _245_ ;
wire _894_ ;
wire _474_ ;
wire _283_ ;
wire _759_ ;
wire _339_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire _797_ ;
wire _377_ ;
wire _186_ ;
wire _912_ ;
wire _721_ ;
wire _301_ ;
wire _37_ ;
wire _530_ ;
wire _110_ ;
wire _815_ ;
wire _75_ ;
wire _624_ ;
wire _204_ ;
wire _853_ ;
wire _433_ ;
wire _909_ ;
wire _662_ ;
wire _242_ ;
wire _718_ ;
wire _891_ ;
wire _471_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _756_ ;
wire _336_ ;
wire _565_ ;
wire _145_ ;
wire _794_ ;
wire _374_ ;
wire _183_ ;
wire _659_ ;
wire _239_ ;
wire _888_ ;
wire _468_ ;
wire _697_ ;
wire _277_ ;
wire _34_ ;
wire _812_ ;
wire _72_ ;
wire _621_ ;
wire _201_ ;
wire _850_ ;
wire _430_ ;
wire _906_ ;
wire _715_ ;
wire _524_ ;
wire _104_ ;
wire _753_ ;
wire _333_ ;
wire _809_ ;
wire _69_ ;
wire _562_ ;
wire _142_ ;
wire _618_ ;
wire _791_ ;
wire _371_ ;
wire _847_ ;
wire _427_ ;
wire _180_ ;
wire _656_ ;
wire _236_ ;
wire _885_ ;
wire _465_ ;
wire _694_ ;
wire _274_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _788_ ;
wire _368_ ;
wire _597_ ;
wire _177_ ;
wire _903_ ;
wire _712_ ;
wire _28_ ;
wire _521_ ;
wire _101_ ;
wire _750_ ;
wire _330_ ;
wire _806_ ;
wire _66_ ;
wire _615_ ;
wire _844_ ;
wire _424_ ;
wire _653_ ;
wire _233_ ;
wire _709_ ;
wire _882_ ;
wire _462_ ;
wire _518_ ;
wire _691_ ;
wire _271_ ;
wire _747_ ;
wire _327_ ;
wire _556_ ;
wire _136_ ;
wire _785_ ;
wire _365_ ;
wire _594_ ;
wire _174_ ;
wire _879_ ;
wire _459_ ;
wire _688_ ;
wire _268_ ;
wire _900_ ;
wire _497_ ;
wire _25_ ;
wire _803_ ;
wire _63_ ;
wire _612_ ;
wire _841_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire _706_ ;
wire _515_ ;
wire _744_ ;
wire _324_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _782_ ;
wire _362_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _591_ ;
wire _171_ ;
wire _647_ ;
wire _227_ ;
wire _876_ ;
wire _456_ ;
wire _685_ ;
wire _265_ ;
wire _494_ ;
wire _22_ ;
wire _779_ ;
wire _359_ ;

BUFX2 BUFX2_insert25 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_148_),
    .Y(_148__bF$buf0)
);

BUFX2 BUFX2_insert24 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_148_),
    .Y(_148__bF$buf1)
);

BUFX2 BUFX2_insert23 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_148_),
    .Y(_148__bF$buf2)
);

BUFX2 BUFX2_insert22 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_148_),
    .Y(_148__bF$buf3)
);

BUFX2 BUFX2_insert21 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_148_),
    .Y(_148__bF$buf4)
);

BUFX2 BUFX2_insert20 (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf0)
);

BUFX2 BUFX2_insert19 (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf1)
);

BUFX2 BUFX2_insert18 (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf2)
);

BUFX2 BUFX2_insert17 (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf3)
);

BUFX2 BUFX2_insert16 (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf4)
);

BUFX2 BUFX2_insert15 (
    .vdd(vdd),
    .gnd(gnd),
    .A(Cin[0]),
    .Y(Cin_0_bF$buf0)
);

BUFX2 BUFX2_insert14 (
    .vdd(vdd),
    .gnd(gnd),
    .A(Cin[0]),
    .Y(Cin_0_bF$buf1)
);

BUFX2 BUFX2_insert13 (
    .vdd(vdd),
    .gnd(gnd),
    .A(Cin[0]),
    .Y(Cin_0_bF$buf2)
);

BUFX2 BUFX2_insert12 (
    .vdd(vdd),
    .gnd(gnd),
    .A(Cin[0]),
    .Y(Cin_0_bF$buf3)
);

CLKBUF1 CLKBUF1_insert11 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert10 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert9 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert8 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert7 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert6 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert5 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_bF$buf6)
);

BUFX2 BUFX2_insert4 (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf0)
);

BUFX2 BUFX2_insert3 (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf1)
);

BUFX2 BUFX2_insert2 (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf2)
);

BUFX2 BUFX2_insert1 (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf3)
);

BUFX2 BUFX2_insert0 (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf4)
);

NAND2X1 _1000_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf4),
    .B(_y[12]),
    .Y(_158_)
);

OAI21X1 _1001_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf3),
    .B(_157_),
    .C(_158_),
    .Y(_16_)
);

INVX1 _1002_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_y[13]),
    .Y(_159_)
);

NAND2X1 _1003_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(y[13]),
    .B(_148__bF$buf4),
    .Y(_160_)
);

OAI21X1 _1004_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_148__bF$buf3),
    .B(_159_),
    .C(_160_),
    .Y(_17_)
);

INVX1 _1005_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(y[14]),
    .Y(_161_)
);

NAND2X1 _1006_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf2),
    .B(_y[14]),
    .Y(_162_)
);

OAI21X1 _1007_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf1),
    .B(_161_),
    .C(_162_),
    .Y(_18_)
);

INVX1 _1008_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_y[15]),
    .Y(_163_)
);

NAND2X1 _1009_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(y[15]),
    .B(_148__bF$buf2),
    .Y(_164_)
);

OAI21X1 _1010_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_148__bF$buf1),
    .B(_163_),
    .C(_164_),
    .Y(_19_)
);

NAND3X1 _1011_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[0]),
    .B(Cin_0_bF$buf3),
    .C(Yin0[0]),
    .Y(_165_)
);

INVX1 _1012_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[0]),
    .Y(_166_)
);

INVX1 _1013_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Cin_0_bF$buf2),
    .Y(_167_)
);

INVX1 _1014_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin0[0]),
    .Y(_168_)
);

OAI21X1 _1015_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_166_),
    .B(_167_),
    .C(_168_),
    .Y(_169_)
);

NAND2X1 _1016_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_165_),
    .B(_169_),
    .Y(_170_)
);

NAND2X1 _1017_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_y[0]),
    .B(_148__bF$buf0),
    .Y(_171_)
);

OAI21X1 _1018_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_148__bF$buf4),
    .B(_170_),
    .C(_171_),
    .Y(_20_)
);

AOI21X1 _1019_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[1]),
    .B(Cin_0_bF$buf1),
    .C(Yin0[1]),
    .Y(_172_)
);

NAND3X1 _1020_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[1]),
    .B(Cin_0_bF$buf0),
    .C(Yin0[1]),
    .Y(_173_)
);

INVX1 _1021_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_173_),
    .Y(_174_)
);

NAND2X1 _1022_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[0]),
    .B(Cin[1]),
    .Y(_175_)
);

OAI21X1 _1023_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_172_),
    .B(_174_),
    .C(_175_),
    .Y(_176_)
);

INVX1 _1024_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_172_),
    .Y(_177_)
);

INVX1 _1025_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_175_),
    .Y(_178_)
);

NAND3X1 _1026_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_173_),
    .B(_178_),
    .C(_177_),
    .Y(_179_)
);

NAND2X1 _1027_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_179_),
    .B(_176_),
    .Y(_180_)
);

OR2X2 _1028_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_180_),
    .B(_165_),
    .Y(_181_)
);

NAND2X1 _1029_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_165_),
    .B(_180_),
    .Y(_182_)
);

NAND2X1 _1030_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_182_),
    .B(_181_),
    .Y(_183_)
);

NAND2X1 _1031_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_y[1]),
    .B(_148__bF$buf3),
    .Y(_184_)
);

OAI21X1 _1032_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_148__bF$buf2),
    .B(_183_),
    .C(_184_),
    .Y(_21_)
);

NAND2X1 _1033_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_y[2]),
    .B(_148__bF$buf1),
    .Y(_185_)
);

INVX1 _1034_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_181_),
    .Y(_186_)
);

INVX4 _1035_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Cin[2]),
    .Y(_187_)
);

OAI21X1 _1036_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_175_),
    .B(_172_),
    .C(_173_),
    .Y(_188_)
);

INVX1 _1037_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_188_),
    .Y(_189_)
);

INVX1 _1038_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[1]),
    .Y(_190_)
);

INVX1 _1039_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Cin[1]),
    .Y(_191_)
);

AOI21X1 _1040_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[2]),
    .B(Cin_0_bF$buf3),
    .C(Yin0[2]),
    .Y(_192_)
);

NAND3X1 _1041_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[2]),
    .B(Cin_0_bF$buf2),
    .C(Yin0[2]),
    .Y(_193_)
);

INVX1 _1042_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_193_),
    .Y(_194_)
);

NOR2X1 _1043_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_192_),
    .B(_194_),
    .Y(_195_)
);

OAI21X1 _1044_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_190_),
    .B(_191_),
    .C(_195_),
    .Y(_196_)
);

NAND2X1 _1045_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[1]),
    .B(Cin[1]),
    .Y(_197_)
);

INVX1 _1046_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_197_),
    .Y(_198_)
);

OAI21X1 _1047_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_192_),
    .B(_194_),
    .C(_198_),
    .Y(_199_)
);

NAND3X1 _1048_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_189_),
    .B(_199_),
    .C(_196_),
    .Y(_200_)
);

NAND2X1 _1049_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_198_),
    .B(_195_),
    .Y(_201_)
);

OAI21X1 _1050_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_192_),
    .B(_194_),
    .C(_197_),
    .Y(_202_)
);

NAND3X1 _1051_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_188_),
    .B(_202_),
    .C(_201_),
    .Y(_203_)
);

NAND2X1 _1052_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_203_),
    .B(_200_),
    .Y(_204_)
);

OAI21X1 _1053_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_166_),
    .B(_187_),
    .C(_204_),
    .Y(_205_)
);

NAND2X1 _1054_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[0]),
    .B(Cin[2]),
    .Y(_206_)
);

INVX1 _1055_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_206_),
    .Y(_207_)
);

NAND3X1 _1056_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_207_),
    .B(_203_),
    .C(_200_),
    .Y(_208_)
);

AOI21X1 _1057_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_205_),
    .B(_208_),
    .C(_186_),
    .Y(_209_)
);

NAND3X1 _1058_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_186_),
    .B(_208_),
    .C(_205_),
    .Y(_210_)
);

NAND2X1 _1059_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf0),
    .B(_210_),
    .Y(_211_)
);

OAI21X1 _1060_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_209_),
    .B(_211_),
    .C(_185_),
    .Y(_22_)
);

NAND2X1 _1061_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_y[3]),
    .B(_148__bF$buf0),
    .Y(_212_)
);

AOI21X1 _1062_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_201_),
    .B(_202_),
    .C(_188_),
    .Y(_213_)
);

OAI21X1 _1063_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_206_),
    .B(_213_),
    .C(_203_),
    .Y(_214_)
);

NAND2X1 _1064_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[1]),
    .B(Cin[3]),
    .Y(_215_)
);

NOR2X1 _1065_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_206_),
    .B(_215_),
    .Y(_216_)
);

AOI22X1 _1066_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[0]),
    .B(Cin[3]),
    .C(XinHL[1]),
    .D(Cin[2]),
    .Y(_217_)
);

NOR2X1 _1067_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_217_),
    .B(_216_),
    .Y(_218_)
);

OAI21X1 _1068_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_197_),
    .B(_192_),
    .C(_193_),
    .Y(_219_)
);

NAND2X1 _1069_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[2]),
    .B(Cin[1]),
    .Y(_220_)
);

NAND3X1 _1070_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[3]),
    .B(Cin_0_bF$buf1),
    .C(Yin0[3]),
    .Y(_221_)
);

INVX1 _1071_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_221_),
    .Y(_222_)
);

AOI21X1 _1072_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[3]),
    .B(Cin_0_bF$buf0),
    .C(Yin0[3]),
    .Y(_223_)
);

OAI21X1 _1073_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_223_),
    .B(_222_),
    .C(_220_),
    .Y(_224_)
);

INVX1 _1074_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_220_),
    .Y(_225_)
);

INVX1 _1075_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_223_),
    .Y(_226_)
);

NAND3X1 _1076_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_225_),
    .B(_221_),
    .C(_226_),
    .Y(_227_)
);

NAND3X1 _1077_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_219_),
    .B(_227_),
    .C(_224_),
    .Y(_228_)
);

INVX1 _1078_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_228_),
    .Y(_229_)
);

AOI21X1 _1079_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_224_),
    .B(_227_),
    .C(_219_),
    .Y(_230_)
);

OAI21X1 _1080_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_230_),
    .B(_229_),
    .C(_218_),
    .Y(_231_)
);

INVX1 _1081_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_218_),
    .Y(_232_)
);

INVX1 _1082_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_219_),
    .Y(_233_)
);

AOI21X1 _1083_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_226_),
    .B(_221_),
    .C(_225_),
    .Y(_234_)
);

INVX1 _1084_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin0[3]),
    .Y(_235_)
);

NAND3X1 _1085_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[3]),
    .B(Cin_0_bF$buf3),
    .C(_235_),
    .Y(_236_)
);

INVX2 _1086_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[3]),
    .Y(_237_)
);

OAI21X1 _1087_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_237_),
    .B(_167_),
    .C(Yin0[3]),
    .Y(_238_)
);

AOI21X1 _1088_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_238_),
    .B(_236_),
    .C(_220_),
    .Y(_239_)
);

OAI21X1 _1089_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_234_),
    .B(_239_),
    .C(_233_),
    .Y(_240_)
);

NAND3X1 _1090_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_232_),
    .B(_228_),
    .C(_240_),
    .Y(_241_)
);

NAND2X1 _1091_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_241_),
    .B(_231_),
    .Y(_242_)
);

NOR2X1 _1092_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_214_),
    .B(_242_),
    .Y(_243_)
);

AOI22X1 _1093_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_208_),
    .B(_203_),
    .C(_231_),
    .D(_241_),
    .Y(_244_)
);

OAI21X1 _1094_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_244_),
    .B(_243_),
    .C(_210_),
    .Y(_245_)
);

NOR3X1 _1095_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_244_),
    .B(_210_),
    .C(_243_),
    .Y(_246_)
);

INVX1 _1096_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_246_),
    .Y(_247_)
);

NAND2X1 _1097_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_245_),
    .B(_247_),
    .Y(_248_)
);

OAI21X1 _1098_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_148__bF$buf4),
    .B(_248_),
    .C(_212_),
    .Y(_23_)
);

NAND2X1 _1099_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_y[4]),
    .B(_148__bF$buf3),
    .Y(_249_)
);

INVX1 _1100_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_216_),
    .Y(_250_)
);

OAI21X1 _1101_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_232_),
    .B(_230_),
    .C(_228_),
    .Y(_251_)
);

OAI21X1 _1102_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_220_),
    .B(_223_),
    .C(_221_),
    .Y(_252_)
);

INVX1 _1103_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_252_),
    .Y(_253_)
);

AOI21X1 _1104_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[0]),
    .B(Cin_0_bF$buf2),
    .C(Yin1[0]),
    .Y(_254_)
);

INVX1 _1105_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_254_),
    .Y(_255_)
);

NAND3X1 _1106_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[0]),
    .B(Cin_0_bF$buf1),
    .C(Yin1[0]),
    .Y(_256_)
);

NAND2X1 _1107_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[3]),
    .B(Cin[1]),
    .Y(_257_)
);

NAND3X1 _1108_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_256_),
    .B(_257_),
    .C(_255_),
    .Y(_258_)
);

INVX1 _1109_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_256_),
    .Y(_259_)
);

INVX1 _1110_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_257_),
    .Y(_260_)
);

OAI21X1 _1111_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_254_),
    .B(_259_),
    .C(_260_),
    .Y(_261_)
);

NAND3X1 _1112_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_258_),
    .B(_261_),
    .C(_253_),
    .Y(_262_)
);

NAND3X1 _1113_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_256_),
    .B(_260_),
    .C(_255_),
    .Y(_263_)
);

OAI21X1 _1114_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_254_),
    .B(_259_),
    .C(_257_),
    .Y(_264_)
);

NAND3X1 _1115_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_252_),
    .B(_263_),
    .C(_264_),
    .Y(_265_)
);

NAND2X1 _1116_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[0]),
    .B(Cin[4]),
    .Y(_266_)
);

INVX1 _1117_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_266_),
    .Y(_267_)
);

AND2X2 _1118_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[1]),
    .B(Cin[3]),
    .Y(_268_)
);

AND2X2 _1119_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[2]),
    .B(Cin[2]),
    .Y(_269_)
);

NAND2X1 _1120_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_268_),
    .B(_269_),
    .Y(_270_)
);

INVX2 _1121_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[2]),
    .Y(_271_)
);

OAI21X1 _1122_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_271_),
    .B(_187_),
    .C(_215_),
    .Y(_272_)
);

NAND3X1 _1123_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_272_),
    .B(_267_),
    .C(_270_),
    .Y(_273_)
);

OAI21X1 _1124_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_271_),
    .B(_187_),
    .C(_268_),
    .Y(_274_)
);

INVX2 _1125_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Cin[3]),
    .Y(_275_)
);

OAI21X1 _1126_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_190_),
    .B(_275_),
    .C(_269_),
    .Y(_276_)
);

NAND3X1 _1127_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_266_),
    .B(_274_),
    .C(_276_),
    .Y(_277_)
);

AND2X2 _1128_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_277_),
    .B(_273_),
    .Y(_278_)
);

NAND3X1 _1129_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_262_),
    .B(_265_),
    .C(_278_),
    .Y(_279_)
);

AOI21X1 _1130_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_264_),
    .B(_263_),
    .C(_252_),
    .Y(_280_)
);

AOI21X1 _1131_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_258_),
    .B(_261_),
    .C(_253_),
    .Y(_281_)
);

NAND2X1 _1132_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_273_),
    .B(_277_),
    .Y(_282_)
);

OAI21X1 _1133_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_280_),
    .B(_281_),
    .C(_282_),
    .Y(_283_)
);

AOI21X1 _1134_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_283_),
    .B(_279_),
    .C(_251_),
    .Y(_284_)
);

NAND3X1 _1135_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_218_),
    .B(_228_),
    .C(_240_),
    .Y(_285_)
);

NAND3X1 _1136_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_265_),
    .B(_282_),
    .C(_262_),
    .Y(_286_)
);

OAI21X1 _1137_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_280_),
    .B(_281_),
    .C(_278_),
    .Y(_287_)
);

AOI22X1 _1138_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_228_),
    .B(_285_),
    .C(_287_),
    .D(_286_),
    .Y(_288_)
);

OAI21X1 _1139_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_288_),
    .B(_284_),
    .C(_250_),
    .Y(_289_)
);

AOI21X1 _1140_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_218_),
    .B(_240_),
    .C(_229_),
    .Y(_290_)
);

NAND3X1 _1141_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_286_),
    .B(_287_),
    .C(_290_),
    .Y(_291_)
);

NAND3X1 _1142_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_251_),
    .B(_279_),
    .C(_283_),
    .Y(_292_)
);

NAND3X1 _1143_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_216_),
    .B(_292_),
    .C(_291_),
    .Y(_293_)
);

NAND3X1 _1144_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_244_),
    .B(_289_),
    .C(_293_),
    .Y(_294_)
);

INVX1 _1145_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_244_),
    .Y(_295_)
);

NAND2X1 _1146_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_289_),
    .B(_293_),
    .Y(_296_)
);

NAND2X1 _1147_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_295_),
    .B(_296_),
    .Y(_297_)
);

AOI21X1 _1148_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_297_),
    .B(_294_),
    .C(_246_),
    .Y(_298_)
);

NAND3X1 _1149_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_294_),
    .B(_246_),
    .C(_297_),
    .Y(_299_)
);

NAND2X1 _1150_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf4),
    .B(_299_),
    .Y(_300_)
);

OAI21X1 _1151_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_298_),
    .B(_300_),
    .C(_249_),
    .Y(_24_)
);

NAND2X1 _1152_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_y[5]),
    .B(_148__bF$buf2),
    .Y(_301_)
);

INVX1 _1153_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_294_),
    .Y(_302_)
);

OAI21X1 _1154_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_250_),
    .B(_284_),
    .C(_292_),
    .Y(_303_)
);

INVX1 _1155_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Cin[5]),
    .Y(_304_)
);

NOR2X1 _1156_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_166_),
    .B(_304_),
    .Y(_305_)
);

INVX1 _1157_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_305_),
    .Y(_306_)
);

INVX1 _1158_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_269_),
    .Y(_307_)
);

OAI21X1 _1159_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_215_),
    .B(_307_),
    .C(_273_),
    .Y(_308_)
);

XOR2X1 _1160_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_308_),
    .B(_306_),
    .Y(_309_)
);

AOI21X1 _1161_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_278_),
    .B(_262_),
    .C(_281_),
    .Y(_310_)
);

NAND2X1 _1162_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[1]),
    .B(Cin[4]),
    .Y(_311_)
);

AND2X2 _1163_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[2]),
    .B(Cin[3]),
    .Y(_312_)
);

OAI21X1 _1164_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_237_),
    .B(_187_),
    .C(_312_),
    .Y(_313_)
);

AND2X2 _1165_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[3]),
    .B(Cin[2]),
    .Y(_314_)
);

OAI21X1 _1166_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_271_),
    .B(_275_),
    .C(_314_),
    .Y(_315_)
);

NAND3X1 _1167_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_311_),
    .B(_313_),
    .C(_315_),
    .Y(_316_)
);

INVX1 _1168_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_311_),
    .Y(_317_)
);

NAND2X1 _1169_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_312_),
    .B(_314_),
    .Y(_318_)
);

OAI22X1 _1170_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_271_),
    .B(_275_),
    .C(_237_),
    .D(_187_),
    .Y(_319_)
);

NAND3X1 _1171_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_317_),
    .B(_319_),
    .C(_318_),
    .Y(_320_)
);

NAND2X1 _1172_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_320_),
    .B(_316_),
    .Y(_321_)
);

OAI21X1 _1173_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_257_),
    .B(_254_),
    .C(_256_),
    .Y(_322_)
);

INVX1 _1174_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_322_),
    .Y(_323_)
);

NAND2X1 _1175_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[0]),
    .B(Cin[1]),
    .Y(_324_)
);

NAND3X1 _1176_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[1]),
    .B(Cin_0_bF$buf0),
    .C(Yin1[1]),
    .Y(_325_)
);

INVX1 _1177_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_325_),
    .Y(_326_)
);

AOI21X1 _1178_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[1]),
    .B(Cin_0_bF$buf3),
    .C(Yin1[1]),
    .Y(_327_)
);

OAI21X1 _1179_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_327_),
    .B(_326_),
    .C(_324_),
    .Y(_328_)
);

INVX1 _1180_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_324_),
    .Y(_329_)
);

INVX1 _1181_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_327_),
    .Y(_330_)
);

NAND3X1 _1182_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_329_),
    .B(_325_),
    .C(_330_),
    .Y(_331_)
);

NAND3X1 _1183_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_331_),
    .B(_328_),
    .C(_323_),
    .Y(_332_)
);

AOI21X1 _1184_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_330_),
    .B(_325_),
    .C(_329_),
    .Y(_333_)
);

INVX1 _1185_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin1[1]),
    .Y(_334_)
);

NAND3X1 _1186_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[1]),
    .B(Cin_0_bF$buf2),
    .C(_334_),
    .Y(_335_)
);

OAI21X1 _1187_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_126_),
    .B(_167_),
    .C(Yin1[1]),
    .Y(_336_)
);

AOI21X1 _1188_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_336_),
    .B(_335_),
    .C(_324_),
    .Y(_337_)
);

OAI21X1 _1189_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_333_),
    .B(_337_),
    .C(_322_),
    .Y(_338_)
);

NAND3X1 _1190_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_321_),
    .B(_332_),
    .C(_338_),
    .Y(_339_)
);

AND2X2 _1191_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_316_),
    .B(_320_),
    .Y(_340_)
);

NAND3X1 _1192_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_322_),
    .B(_331_),
    .C(_328_),
    .Y(_341_)
);

OAI21X1 _1193_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_333_),
    .B(_337_),
    .C(_323_),
    .Y(_342_)
);

NAND3X1 _1194_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_341_),
    .B(_342_),
    .C(_340_),
    .Y(_343_)
);

NAND3X1 _1195_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_339_),
    .B(_343_),
    .C(_310_),
    .Y(_344_)
);

OAI21X1 _1196_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_282_),
    .B(_280_),
    .C(_265_),
    .Y(_345_)
);

AOI21X1 _1197_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_341_),
    .B(_342_),
    .C(_340_),
    .Y(_346_)
);

AOI21X1 _1198_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_338_),
    .B(_332_),
    .C(_321_),
    .Y(_347_)
);

OAI21X1 _1199_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_347_),
    .B(_346_),
    .C(_345_),
    .Y(_348_)
);

NAND3X1 _1200_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_309_),
    .B(_344_),
    .C(_348_),
    .Y(_349_)
);

INVX1 _1201_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_309_),
    .Y(_350_)
);

NAND3X1 _1202_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_339_),
    .B(_345_),
    .C(_343_),
    .Y(_351_)
);

OAI21X1 _1203_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_347_),
    .B(_346_),
    .C(_310_),
    .Y(_352_)
);

NAND3X1 _1204_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_351_),
    .B(_350_),
    .C(_352_),
    .Y(_353_)
);

NAND3X1 _1205_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_349_),
    .B(_353_),
    .C(_303_),
    .Y(_354_)
);

AOI21X1 _1206_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_291_),
    .B(_216_),
    .C(_288_),
    .Y(_355_)
);

AOI21X1 _1207_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_352_),
    .B(_351_),
    .C(_350_),
    .Y(_356_)
);

AOI21X1 _1208_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_348_),
    .B(_344_),
    .C(_309_),
    .Y(_357_)
);

OAI21X1 _1209_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_356_),
    .B(_357_),
    .C(_355_),
    .Y(_358_)
);

NAND3X1 _1210_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_354_),
    .B(_358_),
    .C(_302_),
    .Y(_359_)
);

INVX1 _1211_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_359_),
    .Y(_360_)
);

AND2X2 _1212_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_293_),
    .B(_289_),
    .Y(_361_)
);

AOI22X1 _1213_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_361_),
    .B(_244_),
    .C(_354_),
    .D(_358_),
    .Y(_362_)
);

NOR2X1 _1214_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_362_),
    .B(_360_),
    .Y(_363_)
);

XOR2X1 _1215_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_363_),
    .B(_299_),
    .Y(_364_)
);

OAI21X1 _1216_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_148__bF$buf1),
    .B(_364_),
    .C(_301_),
    .Y(_25_)
);

OAI21X1 _1217_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_362_),
    .B(_299_),
    .C(_359_),
    .Y(_365_)
);

INVX1 _1218_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_354_),
    .Y(_366_)
);

NAND2X1 _1219_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_305_),
    .B(_308_),
    .Y(_367_)
);

INVX1 _1220_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_351_),
    .Y(_368_)
);

AOI21X1 _1221_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_350_),
    .B(_352_),
    .C(_368_),
    .Y(_369_)
);

AOI22X1 _1222_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[0]),
    .B(Cin[6]),
    .C(XinHL[1]),
    .D(Cin[5]),
    .Y(_370_)
);

AND2X2 _1223_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[1]),
    .B(Cin[6]),
    .Y(_371_)
);

NAND2X1 _1224_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_371_),
    .B(_305_),
    .Y(_372_)
);

INVX1 _1225_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_372_),
    .Y(_373_)
);

NOR2X1 _1226_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_370_),
    .B(_373_),
    .Y(_374_)
);

NAND2X1 _1227_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[3]),
    .B(Cin[3]),
    .Y(_375_)
);

OAI21X1 _1228_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_307_),
    .B(_375_),
    .C(_320_),
    .Y(_376_)
);

XNOR2X1 _1229_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_374_),
    .B(_376_),
    .Y(_377_)
);

INVX1 _1230_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_341_),
    .Y(_378_)
);

AOI21X1 _1231_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_340_),
    .B(_342_),
    .C(_378_),
    .Y(_379_)
);

NAND2X1 _1232_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[2]),
    .B(Cin[4]),
    .Y(_380_)
);

NAND2X1 _1233_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[0]),
    .B(Cin[2]),
    .Y(_381_)
);

NOR2X1 _1234_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_375_),
    .B(_381_),
    .Y(_382_)
);

AND2X2 _1235_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_375_),
    .B(_381_),
    .Y(_383_)
);

OAI21X1 _1236_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_382_),
    .B(_383_),
    .C(_380_),
    .Y(_384_)
);

INVX1 _1237_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_380_),
    .Y(_385_)
);

AND2X2 _1238_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[0]),
    .B(Cin[3]),
    .Y(_386_)
);

NAND2X1 _1239_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_314_),
    .B(_386_),
    .Y(_387_)
);

OAI21X1 _1240_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_124_),
    .B(_187_),
    .C(_375_),
    .Y(_388_)
);

NAND3X1 _1241_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_388_),
    .B(_385_),
    .C(_387_),
    .Y(_389_)
);

NAND2X1 _1242_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_389_),
    .B(_384_),
    .Y(_390_)
);

OAI21X1 _1243_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_324_),
    .B(_327_),
    .C(_325_),
    .Y(_391_)
);

INVX1 _1244_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_391_),
    .Y(_392_)
);

NAND2X1 _1245_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[1]),
    .B(Cin[1]),
    .Y(_393_)
);

NAND3X1 _1246_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[2]),
    .B(Cin_0_bF$buf1),
    .C(Yin1[2]),
    .Y(_394_)
);

INVX1 _1247_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_394_),
    .Y(_395_)
);

AOI21X1 _1248_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[2]),
    .B(Cin_0_bF$buf0),
    .C(Yin1[2]),
    .Y(_396_)
);

OAI21X1 _1249_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_396_),
    .B(_395_),
    .C(_393_),
    .Y(_397_)
);

INVX1 _1250_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_393_),
    .Y(_398_)
);

INVX1 _1251_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_396_),
    .Y(_399_)
);

NAND3X1 _1252_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_398_),
    .B(_394_),
    .C(_399_),
    .Y(_400_)
);

NAND3X1 _1253_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_400_),
    .B(_397_),
    .C(_392_),
    .Y(_401_)
);

AOI21X1 _1254_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_399_),
    .B(_394_),
    .C(_398_),
    .Y(_402_)
);

INVX1 _1255_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin1[2]),
    .Y(_403_)
);

NAND3X1 _1256_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[2]),
    .B(Cin_0_bF$buf3),
    .C(_403_),
    .Y(_404_)
);

OAI21X1 _1257_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_128_),
    .B(_167_),
    .C(Yin1[2]),
    .Y(_405_)
);

AOI21X1 _1258_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_405_),
    .B(_404_),
    .C(_393_),
    .Y(_406_)
);

OAI21X1 _1259_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_402_),
    .B(_406_),
    .C(_391_),
    .Y(_407_)
);

NAND3X1 _1260_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_390_),
    .B(_401_),
    .C(_407_),
    .Y(_408_)
);

AND2X2 _1261_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_384_),
    .B(_389_),
    .Y(_409_)
);

NAND3X1 _1262_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_391_),
    .B(_400_),
    .C(_397_),
    .Y(_410_)
);

OAI21X1 _1263_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_402_),
    .B(_406_),
    .C(_392_),
    .Y(_411_)
);

NAND3X1 _1264_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_410_),
    .B(_411_),
    .C(_409_),
    .Y(_412_)
);

NAND3X1 _1265_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_408_),
    .B(_412_),
    .C(_379_),
    .Y(_413_)
);

AOI21X1 _1266_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_328_),
    .B(_331_),
    .C(_322_),
    .Y(_414_)
);

OAI21X1 _1267_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_321_),
    .B(_414_),
    .C(_341_),
    .Y(_415_)
);

AOI21X1 _1268_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_410_),
    .B(_411_),
    .C(_409_),
    .Y(_416_)
);

AOI21X1 _1269_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_407_),
    .B(_401_),
    .C(_390_),
    .Y(_417_)
);

OAI21X1 _1270_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_417_),
    .B(_416_),
    .C(_415_),
    .Y(_418_)
);

NAND3X1 _1271_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_377_),
    .B(_413_),
    .C(_418_),
    .Y(_419_)
);

XOR2X1 _1272_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_374_),
    .B(_376_),
    .Y(_420_)
);

NAND3X1 _1273_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_408_),
    .B(_415_),
    .C(_412_),
    .Y(_421_)
);

OAI21X1 _1274_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_417_),
    .B(_416_),
    .C(_379_),
    .Y(_422_)
);

NAND3X1 _1275_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_420_),
    .B(_421_),
    .C(_422_),
    .Y(_423_)
);

NAND3X1 _1276_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_419_),
    .B(_423_),
    .C(_369_),
    .Y(_424_)
);

AOI21X1 _1277_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_343_),
    .B(_339_),
    .C(_345_),
    .Y(_425_)
);

OAI21X1 _1278_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_309_),
    .B(_425_),
    .C(_351_),
    .Y(_426_)
);

AOI21X1 _1279_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_422_),
    .B(_421_),
    .C(_420_),
    .Y(_427_)
);

AOI21X1 _1280_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_418_),
    .B(_413_),
    .C(_377_),
    .Y(_428_)
);

OAI21X1 _1281_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_427_),
    .B(_428_),
    .C(_426_),
    .Y(_429_)
);

NAND3X1 _1282_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_367_),
    .B(_429_),
    .C(_424_),
    .Y(_430_)
);

INVX1 _1283_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_367_),
    .Y(_431_)
);

NAND3X1 _1284_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_426_),
    .B(_423_),
    .C(_419_),
    .Y(_432_)
);

OAI21X1 _1285_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_427_),
    .B(_428_),
    .C(_369_),
    .Y(_433_)
);

NAND3X1 _1286_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_431_),
    .B(_432_),
    .C(_433_),
    .Y(_434_)
);

NAND3X1 _1287_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_366_),
    .B(_434_),
    .C(_430_),
    .Y(_435_)
);

AOI21X1 _1288_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_433_),
    .B(_432_),
    .C(_431_),
    .Y(_436_)
);

AOI21X1 _1289_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_424_),
    .B(_429_),
    .C(_367_),
    .Y(_437_)
);

OAI21X1 _1290_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_436_),
    .B(_437_),
    .C(_354_),
    .Y(_438_)
);

AOI21X1 _1291_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_438_),
    .B(_435_),
    .C(_365_),
    .Y(_439_)
);

NAND3X1 _1292_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_435_),
    .B(_365_),
    .C(_438_),
    .Y(_440_)
);

NAND2X1 _1293_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf3),
    .B(_440_),
    .Y(_441_)
);

OAI22X1 _1294_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf2),
    .B(_149_),
    .C(_439_),
    .D(_441_),
    .Y(_26_)
);

INVX1 _1295_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_435_),
    .Y(_442_)
);

INVX1 _1296_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_440_),
    .Y(_443_)
);

INVX1 _1297_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_432_),
    .Y(_444_)
);

AOI21X1 _1298_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_431_),
    .B(_433_),
    .C(_444_),
    .Y(_445_)
);

NAND2X1 _1299_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_376_),
    .B(_374_),
    .Y(_446_)
);

INVX1 _1300_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_421_),
    .Y(_447_)
);

AOI21X1 _1301_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_420_),
    .B(_422_),
    .C(_447_),
    .Y(_448_)
);

NAND2X1 _1302_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[0]),
    .B(Cin[7]),
    .Y(_449_)
);

INVX1 _1303_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_449_),
    .Y(_450_)
);

AND2X2 _1304_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[2]),
    .B(Cin[5]),
    .Y(_451_)
);

NAND2X1 _1305_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_371_),
    .B(_451_),
    .Y(_452_)
);

NAND2X1 _1306_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[1]),
    .B(Cin[6]),
    .Y(_453_)
);

OAI21X1 _1307_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_271_),
    .B(_304_),
    .C(_453_),
    .Y(_454_)
);

AOI21X1 _1308_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_452_),
    .B(_454_),
    .C(_450_),
    .Y(_455_)
);

INVX1 _1309_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Cin[6]),
    .Y(_456_)
);

OAI21X1 _1310_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_190_),
    .B(_456_),
    .C(_451_),
    .Y(_457_)
);

OAI21X1 _1311_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_271_),
    .B(_304_),
    .C(_371_),
    .Y(_458_)
);

AOI21X1 _1312_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_457_),
    .B(_458_),
    .C(_449_),
    .Y(_459_)
);

OAI21X1 _1313_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_380_),
    .B(_383_),
    .C(_387_),
    .Y(_460_)
);

OAI21X1 _1314_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_455_),
    .B(_459_),
    .C(_460_),
    .Y(_461_)
);

NAND3X1 _1315_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_449_),
    .B(_457_),
    .C(_458_),
    .Y(_462_)
);

NAND3X1 _1316_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_454_),
    .B(_450_),
    .C(_452_),
    .Y(_463_)
);

AOI21X1 _1317_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_385_),
    .B(_388_),
    .C(_382_),
    .Y(_464_)
);

NAND3X1 _1318_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_463_),
    .B(_462_),
    .C(_464_),
    .Y(_465_)
);

NAND3X1 _1319_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_372_),
    .B(_465_),
    .C(_461_),
    .Y(_466_)
);

NAND3X1 _1320_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_463_),
    .B(_462_),
    .C(_460_),
    .Y(_467_)
);

OAI21X1 _1321_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_455_),
    .B(_459_),
    .C(_464_),
    .Y(_468_)
);

NAND3X1 _1322_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_373_),
    .B(_467_),
    .C(_468_),
    .Y(_469_)
);

NAND2X1 _1323_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_466_),
    .B(_469_),
    .Y(_470_)
);

INVX1 _1324_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_410_),
    .Y(_471_)
);

AOI21X1 _1325_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_409_),
    .B(_411_),
    .C(_471_),
    .Y(_472_)
);

NAND2X1 _1326_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[3]),
    .B(Cin[4]),
    .Y(_473_)
);

NAND2X1 _1327_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[0]),
    .B(Cin[3]),
    .Y(_474_)
);

NAND3X1 _1328_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[1]),
    .B(Cin[2]),
    .C(_474_),
    .Y(_475_)
);

NAND2X1 _1329_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[1]),
    .B(Cin[2]),
    .Y(_476_)
);

NAND2X1 _1330_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_476_),
    .B(_386_),
    .Y(_477_)
);

NAND3X1 _1331_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_473_),
    .B(_475_),
    .C(_477_),
    .Y(_478_)
);

INVX1 _1332_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_473_),
    .Y(_479_)
);

AND2X2 _1333_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[1]),
    .B(Cin[2]),
    .Y(_480_)
);

NAND2X1 _1334_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_386_),
    .B(_480_),
    .Y(_481_)
);

OAI21X1 _1335_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_126_),
    .B(_187_),
    .C(_474_),
    .Y(_482_)
);

NAND3X1 _1336_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_479_),
    .B(_482_),
    .C(_481_),
    .Y(_483_)
);

NAND2X1 _1337_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_478_),
    .B(_483_),
    .Y(_484_)
);

OAI21X1 _1338_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_393_),
    .B(_396_),
    .C(_394_),
    .Y(_485_)
);

INVX1 _1339_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_485_),
    .Y(_486_)
);

NAND2X1 _1340_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[2]),
    .B(Cin[1]),
    .Y(_487_)
);

INVX1 _1341_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin1[3]),
    .Y(_488_)
);

NAND3X1 _1342_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[3]),
    .B(Cin_0_bF$buf2),
    .C(_488_),
    .Y(_489_)
);

NAND2X1 _1343_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[3]),
    .B(Cin_0_bF$buf1),
    .Y(_490_)
);

NAND2X1 _1344_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin1[3]),
    .B(_490_),
    .Y(_491_)
);

NAND3X1 _1345_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_487_),
    .B(_491_),
    .C(_489_),
    .Y(_492_)
);

INVX1 _1346_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_487_),
    .Y(_493_)
);

NAND3X1 _1347_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[3]),
    .B(Cin_0_bF$buf0),
    .C(Yin1[3]),
    .Y(_494_)
);

NAND2X1 _1348_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_488_),
    .B(_490_),
    .Y(_495_)
);

NAND3X1 _1349_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_494_),
    .B(_493_),
    .C(_495_),
    .Y(_496_)
);

NAND3X1 _1350_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_492_),
    .B(_496_),
    .C(_486_),
    .Y(_497_)
);

AOI21X1 _1351_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_495_),
    .B(_494_),
    .C(_493_),
    .Y(_498_)
);

AOI21X1 _1352_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_489_),
    .B(_491_),
    .C(_487_),
    .Y(_499_)
);

OAI21X1 _1353_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_498_),
    .B(_499_),
    .C(_485_),
    .Y(_500_)
);

NAND3X1 _1354_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_484_),
    .B(_497_),
    .C(_500_),
    .Y(_501_)
);

AND2X2 _1355_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_483_),
    .B(_478_),
    .Y(_502_)
);

NAND3X1 _1356_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_485_),
    .B(_496_),
    .C(_492_),
    .Y(_503_)
);

OAI21X1 _1357_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_498_),
    .B(_499_),
    .C(_486_),
    .Y(_504_)
);

NAND3X1 _1358_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_503_),
    .B(_504_),
    .C(_502_),
    .Y(_505_)
);

NAND3X1 _1359_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_501_),
    .B(_505_),
    .C(_472_),
    .Y(_506_)
);

AOI21X1 _1360_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_397_),
    .B(_400_),
    .C(_391_),
    .Y(_507_)
);

OAI21X1 _1361_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_390_),
    .B(_507_),
    .C(_410_),
    .Y(_508_)
);

AOI21X1 _1362_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_503_),
    .B(_504_),
    .C(_502_),
    .Y(_509_)
);

AOI21X1 _1363_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_500_),
    .B(_497_),
    .C(_484_),
    .Y(_510_)
);

OAI21X1 _1364_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_510_),
    .B(_509_),
    .C(_508_),
    .Y(_511_)
);

NAND3X1 _1365_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_470_),
    .B(_511_),
    .C(_506_),
    .Y(_512_)
);

AND2X2 _1366_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_466_),
    .B(_469_),
    .Y(_513_)
);

NAND3X1 _1367_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_501_),
    .B(_505_),
    .C(_508_),
    .Y(_514_)
);

OAI21X1 _1368_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_510_),
    .B(_509_),
    .C(_472_),
    .Y(_515_)
);

NAND3X1 _1369_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_514_),
    .B(_513_),
    .C(_515_),
    .Y(_516_)
);

NAND3X1 _1370_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_512_),
    .B(_516_),
    .C(_448_),
    .Y(_517_)
);

AOI21X1 _1371_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_412_),
    .B(_408_),
    .C(_415_),
    .Y(_518_)
);

OAI21X1 _1372_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_518_),
    .B(_377_),
    .C(_421_),
    .Y(_519_)
);

AOI21X1 _1373_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_515_),
    .B(_514_),
    .C(_513_),
    .Y(_520_)
);

AOI21X1 _1374_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_506_),
    .B(_511_),
    .C(_470_),
    .Y(_521_)
);

OAI21X1 _1375_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_520_),
    .B(_521_),
    .C(_519_),
    .Y(_522_)
);

AOI21X1 _1376_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_517_),
    .B(_522_),
    .C(_446_),
    .Y(_523_)
);

INVX1 _1377_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_446_),
    .Y(_524_)
);

NAND3X1 _1378_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_516_),
    .B(_512_),
    .C(_519_),
    .Y(_525_)
);

OAI21X1 _1379_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_520_),
    .B(_521_),
    .C(_448_),
    .Y(_526_)
);

AOI21X1 _1380_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_526_),
    .B(_525_),
    .C(_524_),
    .Y(_527_)
);

OAI21X1 _1381_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_527_),
    .B(_523_),
    .C(_445_),
    .Y(_528_)
);

AOI21X1 _1382_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_419_),
    .B(_423_),
    .C(_426_),
    .Y(_529_)
);

OAI21X1 _1383_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_367_),
    .B(_529_),
    .C(_432_),
    .Y(_530_)
);

NAND3X1 _1384_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_524_),
    .B(_525_),
    .C(_526_),
    .Y(_531_)
);

NAND3X1 _1385_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_446_),
    .B(_522_),
    .C(_517_),
    .Y(_532_)
);

NAND3X1 _1386_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_530_),
    .B(_531_),
    .C(_532_),
    .Y(_533_)
);

NAND2X1 _1387_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_533_),
    .B(_528_),
    .Y(_534_)
);

OAI21X1 _1388_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_442_),
    .B(_443_),
    .C(_534_),
    .Y(_535_)
);

NOR2X1 _1389_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_442_),
    .B(_443_),
    .Y(_536_)
);

INVX1 _1390_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_534_),
    .Y(_537_)
);

AOI21X1 _1391_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_536_),
    .B(_537_),
    .C(_148__bF$buf0),
    .Y(_538_)
);

AOI22X1 _1392_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_148__bF$buf4),
    .B(_151_),
    .C(_538_),
    .D(_535_),
    .Y(_27_)
);

NAND2X1 _1393_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_y[8]),
    .B(_148__bF$buf3),
    .Y(_539_)
);

INVX1 _1394_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_528_),
    .Y(_540_)
);

AND2X2 _1395_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_533_),
    .B(_435_),
    .Y(_541_)
);

OAI22X1 _1396_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_540_),
    .B(_541_),
    .C(_534_),
    .D(_440_),
    .Y(_542_)
);

AOI21X1 _1397_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_512_),
    .B(_516_),
    .C(_519_),
    .Y(_543_)
);

OAI21X1 _1398_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_446_),
    .B(_543_),
    .C(_525_),
    .Y(_544_)
);

NAND2X1 _1399_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_467_),
    .B(_469_),
    .Y(_545_)
);

INVX1 _1400_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_545_),
    .Y(_546_)
);

INVX1 _1401_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_514_),
    .Y(_547_)
);

AOI21X1 _1402_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_513_),
    .B(_515_),
    .C(_547_),
    .Y(_548_)
);

AND2X2 _1403_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_463_),
    .B(_452_),
    .Y(_549_)
);

NAND2X1 _1404_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[1]),
    .B(Cin[7]),
    .Y(_550_)
);

INVX1 _1405_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_550_),
    .Y(_551_)
);

AND2X2 _1406_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[2]),
    .B(Cin[6]),
    .Y(_552_)
);

AND2X2 _1407_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[3]),
    .B(Cin[5]),
    .Y(_553_)
);

NAND2X1 _1408_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_552_),
    .B(_553_),
    .Y(_554_)
);

NAND2X1 _1409_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[3]),
    .B(Cin[5]),
    .Y(_555_)
);

OAI21X1 _1410_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_271_),
    .B(_456_),
    .C(_555_),
    .Y(_556_)
);

AOI21X1 _1411_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_554_),
    .B(_556_),
    .C(_551_),
    .Y(_557_)
);

OAI21X1 _1412_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_271_),
    .B(_456_),
    .C(_553_),
    .Y(_558_)
);

OAI21X1 _1413_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_237_),
    .B(_304_),
    .C(_552_),
    .Y(_559_)
);

AOI21X1 _1414_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_558_),
    .B(_559_),
    .C(_550_),
    .Y(_560_)
);

AND2X2 _1415_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_474_),
    .B(_476_),
    .Y(_561_)
);

OAI21X1 _1416_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_473_),
    .B(_561_),
    .C(_481_),
    .Y(_562_)
);

OAI21X1 _1417_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_557_),
    .B(_560_),
    .C(_562_),
    .Y(_563_)
);

NAND3X1 _1418_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_550_),
    .B(_558_),
    .C(_559_),
    .Y(_564_)
);

NAND3X1 _1419_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_556_),
    .B(_551_),
    .C(_554_),
    .Y(_565_)
);

NOR2X1 _1420_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_474_),
    .B(_476_),
    .Y(_566_)
);

AOI21X1 _1421_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_479_),
    .B(_482_),
    .C(_566_),
    .Y(_567_)
);

NAND3X1 _1422_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_565_),
    .B(_564_),
    .C(_567_),
    .Y(_568_)
);

NAND3X1 _1423_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_549_),
    .B(_568_),
    .C(_563_),
    .Y(_569_)
);

INVX1 _1424_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_451_),
    .Y(_570_)
);

OAI21X1 _1425_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_453_),
    .B(_570_),
    .C(_463_),
    .Y(_571_)
);

NAND3X1 _1426_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_565_),
    .B(_564_),
    .C(_562_),
    .Y(_572_)
);

OAI21X1 _1427_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_557_),
    .B(_560_),
    .C(_567_),
    .Y(_573_)
);

NAND3X1 _1428_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_571_),
    .B(_572_),
    .C(_573_),
    .Y(_574_)
);

NAND2X1 _1429_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_569_),
    .B(_574_),
    .Y(_575_)
);

INVX1 _1430_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_503_),
    .Y(_576_)
);

AOI21X1 _1431_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_502_),
    .B(_504_),
    .C(_576_),
    .Y(_577_)
);

NAND2X1 _1432_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[0]),
    .B(Cin[4]),
    .Y(_578_)
);

NAND2X1 _1433_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[1]),
    .B(Cin[3]),
    .Y(_579_)
);

NAND3X1 _1434_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[2]),
    .B(Cin[2]),
    .C(_579_),
    .Y(_580_)
);

NAND2X1 _1435_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[2]),
    .B(Cin[2]),
    .Y(_581_)
);

NAND3X1 _1436_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[1]),
    .B(Cin[3]),
    .C(_581_),
    .Y(_582_)
);

NAND3X1 _1437_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_578_),
    .B(_580_),
    .C(_582_),
    .Y(_583_)
);

INVX1 _1438_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_578_),
    .Y(_584_)
);

AND2X2 _1439_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[2]),
    .B(Cin[3]),
    .Y(_585_)
);

NAND2X1 _1440_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_480_),
    .B(_585_),
    .Y(_586_)
);

OAI21X1 _1441_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_128_),
    .B(_187_),
    .C(_579_),
    .Y(_587_)
);

NAND3X1 _1442_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_584_),
    .B(_587_),
    .C(_586_),
    .Y(_588_)
);

NAND2X1 _1443_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_583_),
    .B(_588_),
    .Y(_589_)
);

AOI21X1 _1444_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[3]),
    .B(Cin[1]),
    .C(Yin2[0]),
    .Y(_590_)
);

NAND3X1 _1445_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[3]),
    .B(Cin[1]),
    .C(Yin2[0]),
    .Y(_591_)
);

INVX1 _1446_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_591_),
    .Y(_592_)
);

NOR2X1 _1447_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_590_),
    .B(_592_),
    .Y(_593_)
);

NAND3X1 _1448_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_494_),
    .B(_496_),
    .C(_593_),
    .Y(_594_)
);

AOI21X1 _1449_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[3]),
    .B(Cin_0_bF$buf3),
    .C(Yin1[3]),
    .Y(_595_)
);

OAI21X1 _1450_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_487_),
    .B(_595_),
    .C(_494_),
    .Y(_596_)
);

OAI21X1 _1451_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_590_),
    .B(_592_),
    .C(_596_),
    .Y(_597_)
);

NAND3X1 _1452_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_597_),
    .B(_589_),
    .C(_594_),
    .Y(_598_)
);

AND2X2 _1453_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_588_),
    .B(_583_),
    .Y(_599_)
);

INVX1 _1454_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_590_),
    .Y(_600_)
);

NAND2X1 _1455_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_591_),
    .B(_600_),
    .Y(_601_)
);

NOR2X1 _1456_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_596_),
    .B(_601_),
    .Y(_602_)
);

INVX1 _1457_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_597_),
    .Y(_603_)
);

OAI21X1 _1458_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_602_),
    .B(_603_),
    .C(_599_),
    .Y(_604_)
);

NAND3X1 _1459_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_598_),
    .B(_604_),
    .C(_577_),
    .Y(_605_)
);

AOI21X1 _1460_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_492_),
    .B(_496_),
    .C(_485_),
    .Y(_606_)
);

OAI21X1 _1461_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_484_),
    .B(_606_),
    .C(_503_),
    .Y(_607_)
);

NAND2X1 _1462_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_596_),
    .B(_593_),
    .Y(_608_)
);

NAND3X1 _1463_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_494_),
    .B(_496_),
    .C(_601_),
    .Y(_609_)
);

AOI21X1 _1464_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_608_),
    .B(_609_),
    .C(_599_),
    .Y(_610_)
);

AOI21X1 _1465_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_594_),
    .B(_597_),
    .C(_589_),
    .Y(_611_)
);

OAI21X1 _1466_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_611_),
    .B(_610_),
    .C(_607_),
    .Y(_612_)
);

NAND3X1 _1467_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_575_),
    .B(_605_),
    .C(_612_),
    .Y(_613_)
);

AND2X2 _1468_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_569_),
    .B(_574_),
    .Y(_614_)
);

NAND3X1 _1469_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_598_),
    .B(_607_),
    .C(_604_),
    .Y(_615_)
);

OAI21X1 _1470_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_611_),
    .B(_610_),
    .C(_577_),
    .Y(_616_)
);

NAND3X1 _1471_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_615_),
    .B(_616_),
    .C(_614_),
    .Y(_617_)
);

NAND3X1 _1472_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_613_),
    .B(_617_),
    .C(_548_),
    .Y(_618_)
);

AOI21X1 _1473_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_505_),
    .B(_501_),
    .C(_508_),
    .Y(_619_)
);

OAI21X1 _1474_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_470_),
    .B(_619_),
    .C(_514_),
    .Y(_620_)
);

AOI21X1 _1475_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_615_),
    .B(_616_),
    .C(_614_),
    .Y(_621_)
);

AOI21X1 _1476_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_612_),
    .B(_605_),
    .C(_575_),
    .Y(_622_)
);

OAI21X1 _1477_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_622_),
    .B(_621_),
    .C(_620_),
    .Y(_623_)
);

NAND3X1 _1478_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_546_),
    .B(_623_),
    .C(_618_),
    .Y(_624_)
);

NAND3X1 _1479_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_613_),
    .B(_617_),
    .C(_620_),
    .Y(_625_)
);

OAI21X1 _1480_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_621_),
    .B(_622_),
    .C(_548_),
    .Y(_626_)
);

NAND3X1 _1481_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_545_),
    .B(_625_),
    .C(_626_),
    .Y(_627_)
);

NAND3X1 _1482_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_627_),
    .B(_624_),
    .C(_544_),
    .Y(_628_)
);

INVX1 _1483_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_525_),
    .Y(_629_)
);

AOI21X1 _1484_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_524_),
    .B(_526_),
    .C(_629_),
    .Y(_630_)
);

AOI21X1 _1485_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_626_),
    .B(_625_),
    .C(_545_),
    .Y(_631_)
);

AOI21X1 _1486_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_618_),
    .B(_623_),
    .C(_546_),
    .Y(_632_)
);

OAI21X1 _1487_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_631_),
    .B(_632_),
    .C(_630_),
    .Y(_633_)
);

NAND2X1 _1488_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_628_),
    .B(_633_),
    .Y(_634_)
);

XOR2X1 _1489_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_542_),
    .B(_634_),
    .Y(_635_)
);

OAI21X1 _1490_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_148__bF$buf2),
    .B(_635_),
    .C(_539_),
    .Y(_28_)
);

INVX1 _1491_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_628_),
    .Y(_636_)
);

AOI21X1 _1492_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_542_),
    .B(_633_),
    .C(_636_),
    .Y(_637_)
);

INVX1 _1493_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_625_),
    .Y(_638_)
);

AOI21X1 _1494_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_545_),
    .B(_626_),
    .C(_638_),
    .Y(_639_)
);

NAND2X1 _1495_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_572_),
    .B(_574_),
    .Y(_640_)
);

INVX1 _1496_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_640_),
    .Y(_641_)
);

INVX1 _1497_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_615_),
    .Y(_642_)
);

AOI21X1 _1498_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_614_),
    .B(_616_),
    .C(_642_),
    .Y(_643_)
);

AND2X2 _1499_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_565_),
    .B(_554_),
    .Y(_644_)
);

NAND2X1 _1500_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[2]),
    .B(Cin[7]),
    .Y(_645_)
);

NAND2X1 _1501_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[0]),
    .B(Cin[6]),
    .Y(_646_)
);

NOR2X1 _1502_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_555_),
    .B(_646_),
    .Y(_647_)
);

AOI22X1 _1503_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[0]),
    .B(Cin[5]),
    .C(XinHL[3]),
    .D(Cin[6]),
    .Y(_648_)
);

NOR3X1 _1504_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_645_),
    .B(_648_),
    .C(_647_),
    .Y(_649_)
);

INVX1 _1505_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_645_),
    .Y(_650_)
);

AND2X2 _1506_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[0]),
    .B(Cin[6]),
    .Y(_651_)
);

NAND2X1 _1507_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_553_),
    .B(_651_),
    .Y(_652_)
);

INVX1 _1508_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_648_),
    .Y(_653_)
);

AOI21X1 _1509_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_652_),
    .B(_653_),
    .C(_650_),
    .Y(_654_)
);

AND2X2 _1510_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_579_),
    .B(_581_),
    .Y(_655_)
);

OAI21X1 _1511_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_578_),
    .B(_655_),
    .C(_586_),
    .Y(_656_)
);

OAI21X1 _1512_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_654_),
    .B(_649_),
    .C(_656_),
    .Y(_657_)
);

NAND3X1 _1513_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_650_),
    .B(_653_),
    .C(_652_),
    .Y(_658_)
);

OAI21X1 _1514_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_648_),
    .B(_647_),
    .C(_645_),
    .Y(_659_)
);

AOI22X1 _1515_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_480_),
    .B(_585_),
    .C(_587_),
    .D(_584_),
    .Y(_660_)
);

NAND3X1 _1516_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_658_),
    .B(_660_),
    .C(_659_),
    .Y(_661_)
);

NAND3X1 _1517_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_644_),
    .B(_661_),
    .C(_657_),
    .Y(_662_)
);

NAND2X1 _1518_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[3]),
    .B(Cin[6]),
    .Y(_663_)
);

OAI21X1 _1519_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_570_),
    .B(_663_),
    .C(_565_),
    .Y(_664_)
);

NAND3X1 _1520_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_658_),
    .B(_659_),
    .C(_656_),
    .Y(_665_)
);

OAI21X1 _1521_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_654_),
    .B(_649_),
    .C(_660_),
    .Y(_666_)
);

NAND3X1 _1522_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_664_),
    .B(_665_),
    .C(_666_),
    .Y(_667_)
);

NAND2X1 _1523_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_662_),
    .B(_667_),
    .Y(_668_)
);

AOI21X1 _1524_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_494_),
    .B(_496_),
    .C(_601_),
    .Y(_669_)
);

AOI21X1 _1525_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_599_),
    .B(_609_),
    .C(_669_),
    .Y(_670_)
);

NAND2X1 _1526_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[1]),
    .B(Cin[4]),
    .Y(_671_)
);

AND2X2 _1527_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[3]),
    .B(Cin[2]),
    .Y(_672_)
);

OAI21X1 _1528_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_128_),
    .B(_275_),
    .C(_672_),
    .Y(_673_)
);

OAI21X1 _1529_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_130_),
    .B(_187_),
    .C(_585_),
    .Y(_674_)
);

NAND3X1 _1530_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_671_),
    .B(_673_),
    .C(_674_),
    .Y(_675_)
);

INVX1 _1531_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_671_),
    .Y(_676_)
);

NAND2X1 _1532_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_585_),
    .B(_672_),
    .Y(_677_)
);

OAI22X1 _1533_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_128_),
    .B(_275_),
    .C(_130_),
    .D(_187_),
    .Y(_678_)
);

NAND3X1 _1534_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_676_),
    .B(_678_),
    .C(_677_),
    .Y(_679_)
);

NAND2X1 _1535_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_679_),
    .B(_675_),
    .Y(_680_)
);

XNOR2X1 _1536_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_591_),
    .B(Yin2[1]),
    .Y(_681_)
);

INVX1 _1537_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_681_),
    .Y(_682_)
);

NAND2X1 _1538_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_682_),
    .B(_680_),
    .Y(_683_)
);

NAND3X1 _1539_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_681_),
    .B(_679_),
    .C(_675_),
    .Y(_684_)
);

NAND2X1 _1540_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_684_),
    .B(_683_),
    .Y(_685_)
);

NOR2X1 _1541_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_670_),
    .B(_685_),
    .Y(_686_)
);

NOR2X1 _1542_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_596_),
    .B(_593_),
    .Y(_687_)
);

OAI21X1 _1543_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_589_),
    .B(_687_),
    .C(_608_),
    .Y(_688_)
);

AOI21X1 _1544_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_683_),
    .B(_684_),
    .C(_688_),
    .Y(_689_)
);

OAI21X1 _1545_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_689_),
    .B(_686_),
    .C(_668_),
    .Y(_690_)
);

AND2X2 _1546_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_662_),
    .B(_667_),
    .Y(_691_)
);

NAND3X1 _1547_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_683_),
    .B(_684_),
    .C(_688_),
    .Y(_692_)
);

NAND2X1 _1548_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_670_),
    .B(_685_),
    .Y(_693_)
);

NAND3X1 _1549_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_692_),
    .B(_693_),
    .C(_691_),
    .Y(_694_)
);

NAND3X1 _1550_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_694_),
    .B(_690_),
    .C(_643_),
    .Y(_695_)
);

AOI21X1 _1551_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_604_),
    .B(_598_),
    .C(_607_),
    .Y(_696_)
);

OAI21X1 _1552_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_575_),
    .B(_696_),
    .C(_615_),
    .Y(_697_)
);

AOI22X1 _1553_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_662_),
    .B(_667_),
    .C(_693_),
    .D(_692_),
    .Y(_698_)
);

NAND3X1 _1554_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_683_),
    .B(_684_),
    .C(_670_),
    .Y(_699_)
);

OAI21X1 _1555_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_669_),
    .B(_611_),
    .C(_685_),
    .Y(_700_)
);

AOI21X1 _1556_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_700_),
    .B(_699_),
    .C(_668_),
    .Y(_701_)
);

OAI21X1 _1557_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_698_),
    .B(_701_),
    .C(_697_),
    .Y(_702_)
);

AOI21X1 _1558_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_695_),
    .B(_702_),
    .C(_641_),
    .Y(_703_)
);

NAND3X1 _1559_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_697_),
    .B(_694_),
    .C(_690_),
    .Y(_704_)
);

OAI21X1 _1560_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_698_),
    .B(_701_),
    .C(_643_),
    .Y(_705_)
);

AOI21X1 _1561_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_705_),
    .B(_704_),
    .C(_640_),
    .Y(_706_)
);

OAI21X1 _1562_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_703_),
    .B(_706_),
    .C(_639_),
    .Y(_707_)
);

AOI21X1 _1563_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_705_),
    .B(_704_),
    .C(_641_),
    .Y(_708_)
);

AOI21X1 _1564_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_695_),
    .B(_702_),
    .C(_640_),
    .Y(_709_)
);

OAI22X1 _1565_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_708_),
    .B(_709_),
    .C(_638_),
    .D(_632_),
    .Y(_710_)
);

NAND2X1 _1566_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_707_),
    .B(_710_),
    .Y(_711_)
);

XNOR2X1 _1567_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_637_),
    .B(_711_),
    .Y(_712_)
);

NAND2X1 _1568_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_y[9]),
    .B(_148__bF$buf1),
    .Y(_713_)
);

OAI21X1 _1569_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_148__bF$buf0),
    .B(_712_),
    .C(_713_),
    .Y(_29_)
);

NAND2X1 _1570_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_y[10]),
    .B(_148__bF$buf4),
    .Y(_714_)
);

OAI21X1 _1571_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_628_),
    .B(_711_),
    .C(_710_),
    .Y(_715_)
);

NOR2X1 _1572_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_711_),
    .B(_634_),
    .Y(_716_)
);

AOI21X1 _1573_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_542_),
    .B(_716_),
    .C(_715_),
    .Y(_717_)
);

AOI21X1 _1574_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_690_),
    .B(_694_),
    .C(_697_),
    .Y(_718_)
);

OAI21X1 _1575_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_641_),
    .B(_718_),
    .C(_704_),
    .Y(_719_)
);

NAND2X1 _1576_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_665_),
    .B(_667_),
    .Y(_720_)
);

INVX1 _1577_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720_),
    .Y(_721_)
);

AOI21X1 _1578_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_691_),
    .B(_693_),
    .C(_686_),
    .Y(_722_)
);

OAI21X1 _1579_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_645_),
    .B(_648_),
    .C(_652_),
    .Y(_723_)
);

INVX1 _1580_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_723_),
    .Y(_724_)
);

NAND2X1 _1581_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinHL[3]),
    .B(Cin[7]),
    .Y(_725_)
);

AOI22X1 _1582_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[0]),
    .B(Cin[6]),
    .C(XinH[1]),
    .D(Cin[5]),
    .Y(_726_)
);

NAND2X1 _1583_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[1]),
    .B(Cin[5]),
    .Y(_727_)
);

NOR2X1 _1584_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_646_),
    .B(_727_),
    .Y(_728_)
);

NOR3X1 _1585_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_725_),
    .B(_726_),
    .C(_728_),
    .Y(_729_)
);

INVX1 _1586_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_725_),
    .Y(_730_)
);

INVX1 _1587_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_726_),
    .Y(_731_)
);

INVX1 _1588_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_727_),
    .Y(_732_)
);

NAND2X1 _1589_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_651_),
    .B(_732_),
    .Y(_733_)
);

AOI21X1 _1590_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_733_),
    .B(_731_),
    .C(_730_),
    .Y(_734_)
);

NOR2X1 _1591_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_585_),
    .B(_672_),
    .Y(_735_)
);

OAI21X1 _1592_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_671_),
    .B(_735_),
    .C(_677_),
    .Y(_736_)
);

OAI21X1 _1593_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_729_),
    .B(_734_),
    .C(_736_),
    .Y(_737_)
);

NAND3X1 _1594_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_731_),
    .B(_730_),
    .C(_733_),
    .Y(_738_)
);

OAI21X1 _1595_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_726_),
    .B(_728_),
    .C(_725_),
    .Y(_739_)
);

AND2X2 _1596_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_585_),
    .B(_672_),
    .Y(_740_)
);

AOI21X1 _1597_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_676_),
    .B(_678_),
    .C(_740_),
    .Y(_741_)
);

NAND3X1 _1598_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_738_),
    .B(_739_),
    .C(_741_),
    .Y(_742_)
);

NAND3X1 _1599_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_724_),
    .B(_742_),
    .C(_737_),
    .Y(_743_)
);

NAND3X1 _1600_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_738_),
    .B(_739_),
    .C(_736_),
    .Y(_744_)
);

OAI21X1 _1601_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_729_),
    .B(_734_),
    .C(_741_),
    .Y(_745_)
);

NAND3X1 _1602_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_723_),
    .B(_744_),
    .C(_745_),
    .Y(_746_)
);

NAND2X1 _1603_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_746_),
    .B(_743_),
    .Y(_747_)
);

INVX1 _1604_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin2[1]),
    .Y(_748_)
);

OAI21X1 _1605_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_748_),
    .B(_591_),
    .C(_684_),
    .Y(_749_)
);

INVX1 _1606_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin2[2]),
    .Y(_750_)
);

AND2X2 _1607_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[3]),
    .B(Cin[4]),
    .Y(_751_)
);

AND2X2 _1608_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_585_),
    .B(_751_),
    .Y(_752_)
);

AOI22X1 _1609_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[2]),
    .B(Cin[4]),
    .C(XinH[3]),
    .D(Cin[3]),
    .Y(_753_)
);

OAI21X1 _1610_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_753_),
    .B(_752_),
    .C(_750_),
    .Y(_754_)
);

AOI21X1 _1611_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_585_),
    .B(_751_),
    .C(_753_),
    .Y(_755_)
);

NAND2X1 _1612_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin2[2]),
    .B(_755_),
    .Y(_756_)
);

AND2X2 _1613_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_754_),
    .B(_756_),
    .Y(_757_)
);

NAND2X1 _1614_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_757_),
    .B(_749_),
    .Y(_758_)
);

NAND2X1 _1615_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin2[1]),
    .B(_592_),
    .Y(_759_)
);

NAND2X1 _1616_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_756_),
    .B(_754_),
    .Y(_760_)
);

NAND3X1 _1617_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_759_),
    .B(_684_),
    .C(_760_),
    .Y(_761_)
);

NAND2X1 _1618_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_761_),
    .B(_758_),
    .Y(_762_)
);

NAND2X1 _1619_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_747_),
    .B(_762_),
    .Y(_763_)
);

NAND3X1 _1620_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_759_),
    .B(_684_),
    .C(_757_),
    .Y(_764_)
);

NAND2X1 _1621_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_760_),
    .B(_749_),
    .Y(_765_)
);

NAND2X1 _1622_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_764_),
    .B(_765_),
    .Y(_766_)
);

NAND3X1 _1623_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_743_),
    .B(_746_),
    .C(_766_),
    .Y(_767_)
);

NAND3X1 _1624_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_763_),
    .B(_767_),
    .C(_722_),
    .Y(_768_)
);

OAI21X1 _1625_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_689_),
    .B(_668_),
    .C(_692_),
    .Y(_769_)
);

AOI21X1 _1626_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_743_),
    .B(_746_),
    .C(_766_),
    .Y(_770_)
);

NOR2X1 _1627_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_747_),
    .B(_762_),
    .Y(_771_)
);

OAI21X1 _1628_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_771_),
    .B(_770_),
    .C(_769_),
    .Y(_772_)
);

NAND3X1 _1629_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_721_),
    .B(_772_),
    .C(_768_),
    .Y(_773_)
);

NAND3X1 _1630_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_763_),
    .B(_767_),
    .C(_769_),
    .Y(_774_)
);

OAI21X1 _1631_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_771_),
    .B(_770_),
    .C(_722_),
    .Y(_775_)
);

NAND3X1 _1632_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_774_),
    .B(_720_),
    .C(_775_),
    .Y(_776_)
);

NAND3X1 _1633_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_773_),
    .B(_776_),
    .C(_719_),
    .Y(_777_)
);

NOR3X1 _1634_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_698_),
    .B(_701_),
    .C(_643_),
    .Y(_778_)
);

AOI21X1 _1635_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_640_),
    .B(_705_),
    .C(_778_),
    .Y(_779_)
);

AOI21X1 _1636_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_775_),
    .B(_774_),
    .C(_720_),
    .Y(_780_)
);

AOI21X1 _1637_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_768_),
    .B(_772_),
    .C(_721_),
    .Y(_781_)
);

OAI21X1 _1638_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_780_),
    .B(_781_),
    .C(_779_),
    .Y(_782_)
);

NAND2X1 _1639_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_777_),
    .B(_782_),
    .Y(_783_)
);

AND2X2 _1640_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_717_),
    .B(_783_),
    .Y(_784_)
);

OAI21X1 _1641_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_783_),
    .B(_717_),
    .C(LoadCtl_4_bF$buf1),
    .Y(_785_)
);

OAI21X1 _1642_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_785_),
    .B(_784_),
    .C(_714_),
    .Y(_30_)
);

INVX1 _1643_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_y[11]),
    .Y(_786_)
);

OAI21X1 _1644_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_783_),
    .B(_717_),
    .C(_777_),
    .Y(_787_)
);

AOI21X1 _1645_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_763_),
    .B(_767_),
    .C(_769_),
    .Y(_788_)
);

OAI21X1 _1646_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_721_),
    .B(_788_),
    .C(_774_),
    .Y(_789_)
);

NAND2X1 _1647_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_744_),
    .B(_746_),
    .Y(_790_)
);

INVX1 _1648_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_790_),
    .Y(_791_)
);

AND2X2 _1649_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_743_),
    .B(_746_),
    .Y(_792_)
);

INVX1 _1650_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_758_),
    .Y(_793_)
);

AOI21X1 _1651_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_792_),
    .B(_761_),
    .C(_793_),
    .Y(_794_)
);

OAI21X1 _1652_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_725_),
    .B(_726_),
    .C(_733_),
    .Y(_795_)
);

NAND2X1 _1653_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[0]),
    .B(Cin[7]),
    .Y(_796_)
);

INVX1 _1654_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_796_),
    .Y(_797_)
);

AOI22X1 _1655_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[1]),
    .B(Cin[6]),
    .C(XinH[2]),
    .D(Cin[5]),
    .Y(_798_)
);

INVX1 _1656_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_798_),
    .Y(_799_)
);

AND2X2 _1657_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[2]),
    .B(Cin[6]),
    .Y(_800_)
);

NAND2X1 _1658_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_800_),
    .B(_732_),
    .Y(_801_)
);

NAND3X1 _1659_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_799_),
    .B(_797_),
    .C(_801_),
    .Y(_802_)
);

NAND2X1 _1660_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[2]),
    .B(Cin[6]),
    .Y(_803_)
);

NOR2X1 _1661_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_727_),
    .B(_803_),
    .Y(_804_)
);

OAI21X1 _1662_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_798_),
    .B(_804_),
    .C(_796_),
    .Y(_805_)
);

NAND3X1 _1663_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_752_),
    .B(_805_),
    .C(_802_),
    .Y(_806_)
);

INVX1 _1664_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_752_),
    .Y(_807_)
);

NOR3X1 _1665_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_796_),
    .B(_798_),
    .C(_804_),
    .Y(_808_)
);

AOI21X1 _1666_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_801_),
    .B(_799_),
    .C(_797_),
    .Y(_809_)
);

OAI21X1 _1667_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_808_),
    .B(_809_),
    .C(_807_),
    .Y(_810_)
);

AOI21X1 _1668_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_810_),
    .B(_806_),
    .C(_795_),
    .Y(_811_)
);

INVX1 _1669_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_795_),
    .Y(_812_)
);

OAI21X1 _1670_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_808_),
    .B(_809_),
    .C(_752_),
    .Y(_813_)
);

NAND3X1 _1671_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_805_),
    .B(_807_),
    .C(_802_),
    .Y(_814_)
);

AOI21X1 _1672_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_813_),
    .B(_814_),
    .C(_812_),
    .Y(_815_)
);

INVX1 _1673_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin2[3]),
    .Y(_816_)
);

XOR2X1 _1674_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_751_),
    .B(_816_),
    .Y(_817_)
);

OR2X2 _1675_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_756_),
    .B(_817_),
    .Y(_818_)
);

NAND2X1 _1676_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_817_),
    .B(_756_),
    .Y(_819_)
);

NAND2X1 _1677_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_819_),
    .B(_818_),
    .Y(_820_)
);

OAI21X1 _1678_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_811_),
    .B(_815_),
    .C(_820_),
    .Y(_821_)
);

NAND3X1 _1679_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_812_),
    .B(_814_),
    .C(_813_),
    .Y(_822_)
);

NAND3X1 _1680_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_795_),
    .B(_806_),
    .C(_810_),
    .Y(_823_)
);

INVX1 _1681_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_820_),
    .Y(_824_)
);

NAND3X1 _1682_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_822_),
    .B(_823_),
    .C(_824_),
    .Y(_825_)
);

NAND3X1 _1683_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_821_),
    .B(_825_),
    .C(_794_),
    .Y(_826_)
);

NAND2X1 _1684_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_821_),
    .B(_825_),
    .Y(_827_)
);

OAI21X1 _1685_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_793_),
    .B(_771_),
    .C(_827_),
    .Y(_828_)
);

NAND3X1 _1686_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_791_),
    .B(_828_),
    .C(_826_),
    .Y(_829_)
);

OAI21X1 _1687_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_747_),
    .B(_762_),
    .C(_758_),
    .Y(_830_)
);

NAND3X1 _1688_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_821_),
    .B(_825_),
    .C(_830_),
    .Y(_831_)
);

NAND2X1 _1689_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_827_),
    .B(_794_),
    .Y(_832_)
);

NAND3X1 _1690_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_790_),
    .B(_831_),
    .C(_832_),
    .Y(_833_)
);

NAND3X1 _1691_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_833_),
    .B(_789_),
    .C(_829_),
    .Y(_834_)
);

INVX1 _1692_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_774_),
    .Y(_835_)
);

AOI21X1 _1693_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720_),
    .B(_775_),
    .C(_835_),
    .Y(_836_)
);

AOI21X1 _1694_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_832_),
    .B(_831_),
    .C(_790_),
    .Y(_837_)
);

AOI21X1 _1695_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_826_),
    .B(_828_),
    .C(_791_),
    .Y(_838_)
);

OAI21X1 _1696_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_837_),
    .B(_838_),
    .C(_836_),
    .Y(_839_)
);

NAND2X1 _1697_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_834_),
    .B(_839_),
    .Y(_840_)
);

AND2X2 _1698_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_787_),
    .B(_840_),
    .Y(_841_)
);

NOR2X1 _1699_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_840_),
    .B(_787_),
    .Y(_842_)
);

OAI21X1 _1700_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_842_),
    .B(_841_),
    .C(LoadCtl_4_bF$buf0),
    .Y(_843_)
);

OAI21X1 _1701_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf4),
    .B(_786_),
    .C(_843_),
    .Y(_31_)
);

NAND2X1 _1702_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_y[12]),
    .B(_148__bF$buf3),
    .Y(_844_)
);

NOR2X1 _1703_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_840_),
    .B(_783_),
    .Y(_845_)
);

NAND3X1 _1704_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_716_),
    .B(_845_),
    .C(_542_),
    .Y(_846_)
);

NAND2X1 _1705_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_834_),
    .B(_777_),
    .Y(_847_)
);

AOI22X1 _1706_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_839_),
    .B(_847_),
    .C(_845_),
    .D(_715_),
    .Y(_848_)
);

NAND2X1 _1707_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_846_),
    .B(_848_),
    .Y(_849_)
);

OAI21X1 _1708_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_794_),
    .B(_827_),
    .C(_833_),
    .Y(_850_)
);

NAND2X1 _1709_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_806_),
    .B(_823_),
    .Y(_851_)
);

OAI21X1 _1710_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_756_),
    .B(_817_),
    .C(_825_),
    .Y(_852_)
);

OAI21X1 _1711_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_796_),
    .B(_798_),
    .C(_801_),
    .Y(_853_)
);

NAND2X1 _1712_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[1]),
    .B(Cin[7]),
    .Y(_854_)
);

AOI21X1 _1713_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[3]),
    .B(Cin[5]),
    .C(_800_),
    .Y(_855_)
);

NAND2X1 _1714_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[2]),
    .B(Cin[5]),
    .Y(_856_)
);

NAND2X1 _1715_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[3]),
    .B(Cin[6]),
    .Y(_857_)
);

NOR2X1 _1716_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_856_),
    .B(_857_),
    .Y(_858_)
);

NOR2X1 _1717_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_858_),
    .B(_855_),
    .Y(_859_)
);

XNOR2X1 _1718_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_859_),
    .B(_854_),
    .Y(_860_)
);

NOR2X1 _1719_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_853_),
    .B(_860_),
    .Y(_861_)
);

OAI21X1 _1720_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_804_),
    .B(_808_),
    .C(_860_),
    .Y(_862_)
);

INVX1 _1721_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_862_),
    .Y(_863_)
);

INVX1 _1722_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin3[0]),
    .Y(_864_)
);

NAND2X1 _1723_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin2[3]),
    .B(_751_),
    .Y(_865_)
);

NAND2X1 _1724_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_864_),
    .B(_865_),
    .Y(_866_)
);

OR2X2 _1725_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_865_),
    .B(_864_),
    .Y(_867_)
);

NAND2X1 _1726_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_866_),
    .B(_867_),
    .Y(_868_)
);

OAI21X1 _1727_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_861_),
    .B(_863_),
    .C(_868_),
    .Y(_869_)
);

OR2X2 _1728_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_860_),
    .B(_853_),
    .Y(_870_)
);

INVX1 _1729_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_868_),
    .Y(_871_)
);

NAND3X1 _1730_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_862_),
    .B(_871_),
    .C(_870_),
    .Y(_872_)
);

NAND3X1 _1731_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_872_),
    .B(_852_),
    .C(_869_),
    .Y(_873_)
);

NAND2X1 _1732_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_872_),
    .B(_869_),
    .Y(_874_)
);

NAND3X1 _1733_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_818_),
    .B(_825_),
    .C(_874_),
    .Y(_875_)
);

NAND3X1 _1734_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_851_),
    .B(_873_),
    .C(_875_),
    .Y(_876_)
);

INVX1 _1735_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_851_),
    .Y(_877_)
);

INVX1 _1736_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_873_),
    .Y(_878_)
);

INVX1 _1737_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_875_),
    .Y(_879_)
);

OAI21X1 _1738_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_878_),
    .B(_879_),
    .C(_877_),
    .Y(_880_)
);

NAND3X1 _1739_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_850_),
    .B(_876_),
    .C(_880_),
    .Y(_881_)
);

INVX1 _1740_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_850_),
    .Y(_882_)
);

NAND2X1 _1741_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_876_),
    .B(_880_),
    .Y(_883_)
);

NAND2X1 _1742_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_882_),
    .B(_883_),
    .Y(_884_)
);

AND2X2 _1743_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_884_),
    .B(_881_),
    .Y(_885_)
);

XNOR2X1 _1744_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_849_),
    .B(_885_),
    .Y(_886_)
);

OAI21X1 _1745_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_148__bF$buf2),
    .B(_886_),
    .C(_844_),
    .Y(_32_)
);

INVX1 _1746_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_881_),
    .Y(_887_)
);

AND2X2 _1747_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_849_),
    .B(_885_),
    .Y(_888_)
);

AOI21X1 _1748_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_875_),
    .B(_851_),
    .C(_878_),
    .Y(_889_)
);

OAI22X1 _1749_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_856_),
    .B(_857_),
    .C(_854_),
    .D(_855_),
    .Y(_890_)
);

INVX1 _1750_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Cin[7]),
    .Y(_891_)
);

OAI21X1 _1751_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_128_),
    .B(_891_),
    .C(_857_),
    .Y(_892_)
);

NOR2X1 _1752_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_130_),
    .B(_891_),
    .Y(_893_)
);

NAND2X1 _1753_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_800_),
    .B(_893_),
    .Y(_894_)
);

AND2X2 _1754_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_894_),
    .B(_892_),
    .Y(_895_)
);

XOR2X1 _1755_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_895_),
    .B(_890_),
    .Y(_896_)
);

XNOR2X1 _1756_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_896_),
    .B(Yin3[1]),
    .Y(_897_)
);

AOI21X1 _1757_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_872_),
    .B(_867_),
    .C(_897_),
    .Y(_898_)
);

INVX1 _1758_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_898_),
    .Y(_899_)
);

NAND3X1 _1759_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_867_),
    .B(_897_),
    .C(_872_),
    .Y(_900_)
);

NAND3X1 _1760_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_863_),
    .B(_900_),
    .C(_899_),
    .Y(_901_)
);

INVX1 _1761_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_900_),
    .Y(_902_)
);

OAI21X1 _1762_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_898_),
    .B(_902_),
    .C(_862_),
    .Y(_903_)
);

NAND2X1 _1763_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_901_),
    .B(_903_),
    .Y(_904_)
);

XOR2X1 _1764_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_904_),
    .B(_889_),
    .Y(_905_)
);

INVX1 _1765_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_905_),
    .Y(_906_)
);

OAI21X1 _1766_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_887_),
    .B(_888_),
    .C(_906_),
    .Y(_907_)
);

NOR2X1 _1767_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_887_),
    .B(_888_),
    .Y(_908_)
);

AOI21X1 _1768_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_908_),
    .B(_905_),
    .C(_148__bF$buf1),
    .Y(_909_)
);

AOI22X1 _1769_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_148__bF$buf0),
    .B(_159_),
    .C(_909_),
    .D(_907_),
    .Y(_33_)
);

NAND2X1 _1770_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_y[14]),
    .B(_148__bF$buf4),
    .Y(_910_)
);

NAND3X1 _1771_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_881_),
    .B(_905_),
    .C(_884_),
    .Y(_911_)
);

AOI21X1 _1772_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_848_),
    .B(_846_),
    .C(_911_),
    .Y(_912_)
);

NAND2X1 _1773_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_905_),
    .B(_887_),
    .Y(_913_)
);

OAI21X1 _1774_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_889_),
    .B(_904_),
    .C(_913_),
    .Y(_914_)
);

NOR2X1 _1775_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914_),
    .B(_912_),
    .Y(_915_)
);

AOI21X1 _1776_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_863_),
    .B(_900_),
    .C(_898_),
    .Y(_916_)
);

NAND2X1 _1777_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_890_),
    .B(_895_),
    .Y(_917_)
);

OAI21X1 _1778_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_128_),
    .B(_456_),
    .C(_893_),
    .Y(_918_)
);

XOR2X1 _1779_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_918_),
    .B(Yin3[2]),
    .Y(_919_)
);

NAND2X1 _1780_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin3[1]),
    .B(_896_),
    .Y(_56_)
);

OR2X2 _1781_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_56_),
    .B(_919_),
    .Y(_57_)
);

NAND2X1 _1782_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_919_),
    .B(_56_),
    .Y(_58_)
);

NAND2X1 _1783_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_58_),
    .B(_57_),
    .Y(_59_)
);

NAND2X1 _1784_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_917_),
    .B(_59_),
    .Y(_60_)
);

OAI21X1 _1785_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_917_),
    .B(_919_),
    .C(_60_),
    .Y(_61_)
);

OR2X2 _1786_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_61_),
    .B(_916_),
    .Y(_62_)
);

NAND2X1 _1787_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_916_),
    .B(_61_),
    .Y(_63_)
);

AND2X2 _1788_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_62_),
    .B(_63_),
    .Y(_64_)
);

XOR2X1 _1789_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_915_),
    .B(_64_),
    .Y(_65_)
);

OAI21X1 _1790_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_148__bF$buf3),
    .B(_65_),
    .C(_910_),
    .Y(_34_)
);

OAI21X1 _1791_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914_),
    .B(_912_),
    .C(_64_),
    .Y(_66_)
);

OAI21X1 _1792_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_916_),
    .B(_61_),
    .C(_66_),
    .Y(_67_)
);

OAI21X1 _1793_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_917_),
    .B(_919_),
    .C(_57_),
    .Y(_68_)
);

OAI21X1 _1794_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin3[2]),
    .B(_800_),
    .C(_893_),
    .Y(_69_)
);

XOR2X1 _1795_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_69_),
    .B(Yin3[3]),
    .Y(_70_)
);

XNOR2X1 _1796_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_68_),
    .B(_70_),
    .Y(_71_)
);

INVX1 _1797_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_71_),
    .Y(_72_)
);

NAND2X1 _1798_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_72_),
    .B(_67_),
    .Y(_73_)
);

NAND3X1 _1799_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_62_),
    .B(_71_),
    .C(_66_),
    .Y(_74_)
);

AND2X2 _1800_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_74_),
    .B(LoadCtl_4_bF$buf3),
    .Y(_75_)
);

AOI22X1 _1801_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_148__bF$buf2),
    .B(_163_),
    .C(_75_),
    .D(_73_),
    .Y(_35_)
);

INVX1 _1802_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin[0]),
    .Y(_76_)
);

INVX1 _1803_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl[2]),
    .Y(_77_)
);

NAND3X1 _1804_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl[3]),
    .B(_77_),
    .C(_104_),
    .Y(_78_)
);

NAND2X1 _1805_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin3[0]),
    .B(_78_),
    .Y(_79_)
);

OAI21X1 _1806_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_76_),
    .B(_78_),
    .C(_79_),
    .Y(_36_)
);

INVX1 _1807_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin[1]),
    .Y(_80_)
);

NAND2X1 _1808_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin3[1]),
    .B(_78_),
    .Y(_81_)
);

OAI21X1 _1809_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_80_),
    .B(_78_),
    .C(_81_),
    .Y(_37_)
);

INVX1 _1810_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin[2]),
    .Y(_82_)
);

NAND2X1 _1811_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin3[2]),
    .B(_78_),
    .Y(_83_)
);

OAI21X1 _1812_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_82_),
    .B(_78_),
    .C(_83_),
    .Y(_38_)
);

INVX1 _1813_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin[3]),
    .Y(_84_)
);

NAND2X1 _1814_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin3[3]),
    .B(_78_),
    .Y(_85_)
);

OAI21X1 _1815_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_84_),
    .B(_78_),
    .C(_85_),
    .Y(_39_)
);

NOR2X1 _1816_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_77_),
    .B(_105_),
    .Y(_86_)
);

NOR2X1 _1817_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin2[0]),
    .B(_86_),
    .Y(_87_)
);

AOI21X1 _1818_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_76_),
    .B(_86_),
    .C(_87_),
    .Y(_40_)
);

NAND2X1 _1819_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin[1]),
    .B(_86_),
    .Y(_88_)
);

OAI21X1 _1820_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_748_),
    .B(_86_),
    .C(_88_),
    .Y(_41_)
);

NAND2X1 _1821_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin[2]),
    .B(_86_),
    .Y(_89_)
);

OAI21X1 _1822_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_750_),
    .B(_86_),
    .C(_89_),
    .Y(_42_)
);

NAND2X1 _1823_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Yin[3]),
    .B(_86_),
    .Y(_90_)
);

OAI21X1 _1824_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_816_),
    .B(_86_),
    .C(_90_),
    .Y(_43_)
);

INVX1 _1825_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_110_),
    .Y(_91_)
);

OAI21X1 _1826_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf4),
    .B(_109_),
    .C(Yin1[0]),
    .Y(_92_)
);

OAI21X1 _1827_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_76_),
    .B(_91_),
    .C(_92_),
    .Y(_44_)
);

OAI21X1 _1828_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf3),
    .B(_109_),
    .C(Yin1[1]),
    .Y(_93_)
);

OAI21X1 _1829_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_80_),
    .B(_91_),
    .C(_93_),
    .Y(_45_)
);

OAI21X1 _1830_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf2),
    .B(_109_),
    .C(Yin1[2]),
    .Y(_94_)
);

OAI21X1 _1831_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_82_),
    .B(_91_),
    .C(_94_),
    .Y(_46_)
);

OAI21X1 _1832_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf1),
    .B(_109_),
    .C(Yin1[3]),
    .Y(_95_)
);

OAI21X1 _1833_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_84_),
    .B(_91_),
    .C(_95_),
    .Y(_47_)
);

NAND2X1 _1834_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf0),
    .B(Yin[0]),
    .Y(_96_)
);

OAI21X1 _1835_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf4),
    .B(_168_),
    .C(_96_),
    .Y(_48_)
);

NOR2X1 _1836_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf3),
    .B(Yin0[1]),
    .Y(_97_)
);

AOI21X1 _1837_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf2),
    .B(_80_),
    .C(_97_),
    .Y(_49_)
);

NOR2X1 _1838_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf1),
    .B(Yin0[2]),
    .Y(_98_)
);

AOI21X1 _1839_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf0),
    .B(_82_),
    .C(_98_),
    .Y(_50_)
);

NAND2X1 _1840_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf4),
    .B(Yin[3]),
    .Y(_99_)
);

OAI21X1 _1841_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf3),
    .B(_235_),
    .C(_99_),
    .Y(_51_)
);

NAND2X1 _1842_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf2),
    .B(Xin[0]),
    .Y(_100_)
);

OAI21X1 _1843_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf1),
    .B(_166_),
    .C(_100_),
    .Y(_52_)
);

NAND2X1 _1844_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf0),
    .B(Xin[1]),
    .Y(_101_)
);

OAI21X1 _1845_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf4),
    .B(_190_),
    .C(_101_),
    .Y(_53_)
);

NAND2X1 _1846_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf3),
    .B(Xin[2]),
    .Y(_102_)
);

OAI21X1 _1847_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf2),
    .B(_271_),
    .C(_102_),
    .Y(_54_)
);

NAND2X1 _1848_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf1),
    .B(Xin[3]),
    .Y(_103_)
);

OAI21X1 _1849_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf0),
    .B(_237_),
    .C(_103_),
    .Y(_55_)
);

DFFPOSX1 _1850_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_0_),
    .Q(XinH[0])
);

DFFPOSX1 _1851_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_1_),
    .Q(XinH[1])
);

DFFPOSX1 _1852_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_2_),
    .Q(XinH[2])
);

DFFPOSX1 _1853_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_3_),
    .Q(XinH[3])
);

DFFPOSX1 _1854_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_4_),
    .Q(y[0])
);

DFFPOSX1 _1855_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_5_),
    .Q(y[1])
);

DFFPOSX1 _1856_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_6_),
    .Q(y[2])
);

DFFPOSX1 _1857_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_7_),
    .Q(y[3])
);

DFFPOSX1 _1858_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_8_),
    .Q(y[4])
);

DFFPOSX1 _1859_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_9_),
    .Q(y[5])
);

DFFPOSX1 _1860_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_10_),
    .Q(y[6])
);

DFFPOSX1 _1861_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_11_),
    .Q(y[7])
);

DFFPOSX1 _1862_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_12_),
    .Q(y[8])
);

DFFPOSX1 _1863_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_13_),
    .Q(y[9])
);

DFFPOSX1 _1864_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_14_),
    .Q(y[10])
);

DFFPOSX1 _1865_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_15_),
    .Q(y[11])
);

DFFPOSX1 _1866_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_16_),
    .Q(y[12])
);

DFFPOSX1 _1867_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_17_),
    .Q(y[13])
);

DFFPOSX1 _1868_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_18_),
    .Q(y[14])
);

DFFPOSX1 _1869_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_19_),
    .Q(y[15])
);

DFFPOSX1 _1870_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_20_),
    .Q(_y[0])
);

DFFPOSX1 _1871_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_21_),
    .Q(_y[1])
);

DFFPOSX1 _1872_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_22_),
    .Q(_y[2])
);

DFFPOSX1 _1873_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_23_),
    .Q(_y[3])
);

DFFPOSX1 _1874_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_24_),
    .Q(_y[4])
);

DFFPOSX1 _1875_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_25_),
    .Q(_y[5])
);

DFFPOSX1 _1876_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_26_),
    .Q(_y[6])
);

DFFPOSX1 _1877_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_27_),
    .Q(_y[7])
);

DFFPOSX1 _1878_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_28_),
    .Q(_y[8])
);

DFFPOSX1 _1879_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_29_),
    .Q(_y[9])
);

DFFPOSX1 _1880_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_30_),
    .Q(_y[10])
);

DFFPOSX1 _1881_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_31_),
    .Q(_y[11])
);

DFFPOSX1 _1882_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_32_),
    .Q(_y[12])
);

DFFPOSX1 _1883_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_33_),
    .Q(_y[13])
);

DFFPOSX1 _1884_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_34_),
    .Q(_y[14])
);

DFFPOSX1 _1885_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_35_),
    .Q(_y[15])
);

DFFPOSX1 _1886_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_36_),
    .Q(Yin3[0])
);

DFFPOSX1 _1887_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_37_),
    .Q(Yin3[1])
);

DFFPOSX1 _1888_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_38_),
    .Q(Yin3[2])
);

DFFPOSX1 _1889_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_39_),
    .Q(Yin3[3])
);

DFFPOSX1 _1890_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_40_),
    .Q(Yin2[0])
);

DFFPOSX1 _1891_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_41_),
    .Q(Yin2[1])
);

DFFPOSX1 _1892_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_42_),
    .Q(Yin2[2])
);

DFFPOSX1 _1893_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_43_),
    .Q(Yin2[3])
);

DFFPOSX1 _1894_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_44_),
    .Q(Yin1[0])
);

DFFPOSX1 _1895_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_45_),
    .Q(Yin1[1])
);

DFFPOSX1 _1896_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_46_),
    .Q(Yin1[2])
);

DFFPOSX1 _1897_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_47_),
    .Q(Yin1[3])
);

DFFPOSX1 _1898_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_48_),
    .Q(Yin0[0])
);

DFFPOSX1 _1899_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_49_),
    .Q(Yin0[1])
);

DFFPOSX1 _1900_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_50_),
    .Q(Yin0[2])
);

DFFPOSX1 _1901_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_51_),
    .Q(Yin0[3])
);

DFFPOSX1 _1902_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_52_),
    .Q(XinHL[0])
);

DFFPOSX1 _1903_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_53_),
    .Q(XinHL[1])
);

DFFPOSX1 _1904_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_54_),
    .Q(XinHL[2])
);

DFFPOSX1 _1905_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_55_),
    .Q(XinHL[3])
);

DFFPOSX1 _1906_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(Rdy),
    .Q(LoadCtl[0])
);

DFFPOSX1 _1907_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(LoadCtl_0_bF$buf4),
    .Q(LoadCtl[1])
);

DFFPOSX1 _1908_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(LoadCtl[1]),
    .Q(LoadCtl[2])
);

DFFPOSX1 _1909_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(LoadCtl[2]),
    .Q(LoadCtl[3])
);

DFFPOSX1 _1910_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(LoadCtl[3]),
    .Q(LoadCtl[4])
);

BUFX2 _1911_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf2),
    .Y(Vld)
);

BUFX2 _1912_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_920_[0]),
    .Y(Xout[0])
);

BUFX2 _1913_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_920_[1]),
    .Y(Xout[1])
);

BUFX2 _1914_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_920_[2]),
    .Y(Xout[2])
);

BUFX2 _1915_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_920_[3]),
    .Y(Xout[3])
);

BUFX2 _1916_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_921_[0]),
    .Y(Yout[0])
);

BUFX2 _1917_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_921_[1]),
    .Y(Yout[1])
);

BUFX2 _1918_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_921_[2]),
    .Y(Yout[2])
);

BUFX2 _1919_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_921_[3]),
    .Y(Yout[3])
);

NOR2X1 _922_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl[1]),
    .B(LoadCtl_0_bF$buf3),
    .Y(_104_)
);

INVX2 _923_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_104_),
    .Y(_105_)
);

INVX1 _924_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(y[8]),
    .Y(_106_)
);

NAND2X1 _925_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl[2]),
    .B(_106_),
    .Y(_107_)
);

OAI21X1 _926_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl[2]),
    .B(y[12]),
    .C(_107_),
    .Y(_108_)
);

INVX2 _927_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl[1]),
    .Y(_109_)
);

NOR2X1 _928_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf2),
    .B(_109_),
    .Y(_110_)
);

AOI22X1 _929_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf1),
    .B(y[0]),
    .C(_110_),
    .D(y[4]),
    .Y(_111_)
);

OAI21X1 _930_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_105_),
    .B(_108_),
    .C(_111_),
    .Y(_921_[0])
);

INVX1 _931_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(y[9]),
    .Y(_112_)
);

NAND2X1 _932_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl[2]),
    .B(_112_),
    .Y(_113_)
);

OAI21X1 _933_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl[2]),
    .B(y[13]),
    .C(_113_),
    .Y(_114_)
);

AOI22X1 _934_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf0),
    .B(y[1]),
    .C(_110_),
    .D(y[5]),
    .Y(_115_)
);

OAI21X1 _935_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_105_),
    .B(_114_),
    .C(_115_),
    .Y(_921_[1])
);

INVX1 _936_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(y[10]),
    .Y(_116_)
);

NAND2X1 _937_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl[2]),
    .B(_116_),
    .Y(_117_)
);

OAI21X1 _938_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl[2]),
    .B(y[14]),
    .C(_117_),
    .Y(_118_)
);

AOI22X1 _939_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf4),
    .B(y[2]),
    .C(_110_),
    .D(y[6]),
    .Y(_119_)
);

OAI21X1 _940_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_105_),
    .B(_118_),
    .C(_119_),
    .Y(_921_[2])
);

INVX1 _941_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(y[11]),
    .Y(_120_)
);

NAND2X1 _942_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl[2]),
    .B(_120_),
    .Y(_121_)
);

OAI21X1 _943_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl[2]),
    .B(y[15]),
    .C(_121_),
    .Y(_122_)
);

AOI22X1 _944_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf3),
    .B(y[3]),
    .C(_110_),
    .D(y[7]),
    .Y(_123_)
);

OAI21X1 _945_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_105_),
    .B(_122_),
    .C(_123_),
    .Y(_921_[3])
);

INVX1 _946_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[0]),
    .Y(_124_)
);

NAND2X1 _947_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf2),
    .B(XinHL[0]),
    .Y(_125_)
);

OAI21X1 _948_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf1),
    .B(_124_),
    .C(_125_),
    .Y(_920_[0])
);

INVX1 _949_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[1]),
    .Y(_126_)
);

NAND2X1 _950_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf0),
    .B(XinHL[1]),
    .Y(_127_)
);

OAI21X1 _951_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf4),
    .B(_126_),
    .C(_127_),
    .Y(_920_[1])
);

INVX2 _952_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[2]),
    .Y(_128_)
);

NAND2X1 _953_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf3),
    .B(XinHL[2]),
    .Y(_129_)
);

OAI21X1 _954_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf2),
    .B(_128_),
    .C(_129_),
    .Y(_920_[2])
);

INVX2 _955_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(XinH[3]),
    .Y(_130_)
);

NAND2X1 _956_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf1),
    .B(XinHL[3]),
    .Y(_131_)
);

OAI21X1 _957_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_0_bF$buf0),
    .B(_130_),
    .C(_131_),
    .Y(_920_[3])
);

NAND2X1 _958_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[0]),
    .B(_110_),
    .Y(_132_)
);

OAI21X1 _959_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_124_),
    .B(_110_),
    .C(_132_),
    .Y(_0_)
);

NAND2X1 _960_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[1]),
    .B(_110_),
    .Y(_133_)
);

OAI21X1 _961_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_126_),
    .B(_110_),
    .C(_133_),
    .Y(_1_)
);

NAND2X1 _962_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[2]),
    .B(_110_),
    .Y(_134_)
);

OAI21X1 _963_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_128_),
    .B(_110_),
    .C(_134_),
    .Y(_2_)
);

NAND2X1 _964_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Xin[3]),
    .B(_110_),
    .Y(_135_)
);

OAI21X1 _965_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_130_),
    .B(_110_),
    .C(_135_),
    .Y(_3_)
);

INVX1 _966_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(y[0]),
    .Y(_136_)
);

NAND2X1 _967_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_y[0]),
    .B(LoadCtl_4_bF$buf1),
    .Y(_137_)
);

OAI21X1 _968_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf0),
    .B(_136_),
    .C(_137_),
    .Y(_4_)
);

INVX1 _969_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(y[1]),
    .Y(_138_)
);

NAND2X1 _970_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf4),
    .B(_y[1]),
    .Y(_139_)
);

OAI21X1 _971_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf3),
    .B(_138_),
    .C(_139_),
    .Y(_5_)
);

INVX1 _972_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(y[2]),
    .Y(_140_)
);

NAND2X1 _973_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf2),
    .B(_y[2]),
    .Y(_141_)
);

OAI21X1 _974_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf1),
    .B(_140_),
    .C(_141_),
    .Y(_6_)
);

INVX1 _975_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(y[3]),
    .Y(_142_)
);

NAND2X1 _976_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf0),
    .B(_y[3]),
    .Y(_143_)
);

OAI21X1 _977_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf4),
    .B(_142_),
    .C(_143_),
    .Y(_7_)
);

INVX1 _978_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(y[4]),
    .Y(_144_)
);

NAND2X1 _979_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf3),
    .B(_y[4]),
    .Y(_145_)
);

OAI21X1 _980_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf2),
    .B(_144_),
    .C(_145_),
    .Y(_8_)
);

INVX1 _981_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(y[5]),
    .Y(_146_)
);

NAND2X1 _982_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf1),
    .B(_y[5]),
    .Y(_147_)
);

OAI21X1 _983_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf0),
    .B(_146_),
    .C(_147_),
    .Y(_9_)
);

INVX8 _984_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf4),
    .Y(_148_)
);

INVX1 _985_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_y[6]),
    .Y(_149_)
);

NAND2X1 _986_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(y[6]),
    .B(_148__bF$buf1),
    .Y(_150_)
);

OAI21X1 _987_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_148__bF$buf0),
    .B(_149_),
    .C(_150_),
    .Y(_10_)
);

INVX1 _988_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_y[7]),
    .Y(_151_)
);

NAND2X1 _989_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(y[7]),
    .B(_148__bF$buf4),
    .Y(_152_)
);

OAI21X1 _990_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_148__bF$buf3),
    .B(_151_),
    .C(_152_),
    .Y(_11_)
);

NAND2X1 _991_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf3),
    .B(_y[8]),
    .Y(_153_)
);

OAI21X1 _992_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf2),
    .B(_106_),
    .C(_153_),
    .Y(_12_)
);

NAND2X1 _993_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf1),
    .B(_y[9]),
    .Y(_154_)
);

OAI21X1 _994_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf0),
    .B(_112_),
    .C(_154_),
    .Y(_13_)
);

NAND2X1 _995_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf4),
    .B(_y[10]),
    .Y(_155_)
);

OAI21X1 _996_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf3),
    .B(_116_),
    .C(_155_),
    .Y(_14_)
);

NAND2X1 _997_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf2),
    .B(_y[11]),
    .Y(_156_)
);

OAI21X1 _998_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCtl_4_bF$buf1),
    .B(_120_),
    .C(_156_),
    .Y(_15_)
);

INVX1 _999_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(y[12]),
    .Y(_157_)
);

endmodule

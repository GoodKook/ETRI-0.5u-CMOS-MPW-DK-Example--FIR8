VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fir_pe
  CLASS BLOCK ;
  FOREIGN fir_pe ;
  ORIGIN 6.000 6.000 ;
  SIZE 1023.000 BY 990.000 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 975.300 1026.450 977.700 ;
        RECT 1017.450 899.700 1026.450 975.300 ;
        RECT 0.600 897.300 1026.450 899.700 ;
        RECT 1017.450 821.700 1026.450 897.300 ;
        RECT 0.600 819.300 1026.450 821.700 ;
        RECT 1017.450 743.700 1026.450 819.300 ;
        RECT 0.600 741.300 1026.450 743.700 ;
        RECT 1017.450 665.700 1026.450 741.300 ;
        RECT 0.600 663.300 1026.450 665.700 ;
        RECT 1017.450 587.700 1026.450 663.300 ;
        RECT 0.600 585.300 1026.450 587.700 ;
        RECT 1017.450 509.700 1026.450 585.300 ;
        RECT 0.600 507.300 1026.450 509.700 ;
        RECT 1017.450 431.700 1026.450 507.300 ;
        RECT 0.600 429.300 1026.450 431.700 ;
        RECT 1017.450 353.700 1026.450 429.300 ;
        RECT 0.600 351.300 1026.450 353.700 ;
        RECT 1017.450 275.700 1026.450 351.300 ;
        RECT 0.600 273.300 1026.450 275.700 ;
        RECT 1017.450 197.700 1026.450 273.300 ;
        RECT 0.600 195.300 1026.450 197.700 ;
        RECT 1017.450 119.700 1026.450 195.300 ;
        RECT 0.600 117.300 1026.450 119.700 ;
        RECT 1017.450 41.700 1026.450 117.300 ;
        RECT 0.600 39.300 1026.450 41.700 ;
        RECT 1017.450 0.300 1026.450 39.300 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -9.450 938.700 -0.450 977.700 ;
        RECT -9.450 936.300 1016.400 938.700 ;
        RECT -9.450 860.700 -0.450 936.300 ;
        RECT -9.450 858.300 1016.400 860.700 ;
        RECT -9.450 782.700 -0.450 858.300 ;
        RECT -9.450 780.300 1016.400 782.700 ;
        RECT -9.450 704.700 -0.450 780.300 ;
        RECT -9.450 702.300 1016.400 704.700 ;
        RECT -9.450 626.700 -0.450 702.300 ;
        RECT -9.450 624.300 1016.400 626.700 ;
        RECT -9.450 548.700 -0.450 624.300 ;
        RECT -9.450 546.300 1016.400 548.700 ;
        RECT -9.450 470.700 -0.450 546.300 ;
        RECT -9.450 468.300 1016.400 470.700 ;
        RECT -9.450 392.700 -0.450 468.300 ;
        RECT -9.450 390.300 1016.400 392.700 ;
        RECT -9.450 314.700 -0.450 390.300 ;
        RECT -9.450 312.300 1016.400 314.700 ;
        RECT -9.450 236.700 -0.450 312.300 ;
        RECT -9.450 234.300 1016.400 236.700 ;
        RECT -9.450 158.700 -0.450 234.300 ;
        RECT -9.450 156.300 1016.400 158.700 ;
        RECT -9.450 80.700 -0.450 156.300 ;
        RECT -9.450 78.300 1016.400 80.700 ;
        RECT -9.450 2.700 -0.450 78.300 ;
        RECT -9.450 0.300 1016.400 2.700 ;
    END
  END vdd
  PIN Cin[7]
    PORT
      LAYER metal1 ;
        RECT 391.950 963.450 394.050 964.050 ;
        RECT 397.950 963.450 400.050 964.050 ;
        RECT 391.950 962.550 400.050 963.450 ;
        RECT 391.950 961.950 394.050 962.550 ;
        RECT 397.950 961.950 400.050 962.550 ;
        RECT 391.950 951.450 394.050 952.050 ;
        RECT 400.950 951.450 403.050 952.050 ;
        RECT 391.950 950.550 403.050 951.450 ;
        RECT 391.950 949.950 394.050 950.550 ;
        RECT 400.950 949.950 403.050 950.550 ;
        RECT 472.950 642.450 475.050 643.050 ;
        RECT 490.950 642.450 493.050 642.750 ;
        RECT 472.950 641.550 493.050 642.450 ;
        RECT 472.950 640.950 475.050 641.550 ;
        RECT 490.950 640.650 493.050 641.550 ;
        RECT 627.000 495.450 631.050 496.050 ;
        RECT 626.550 493.950 631.050 495.450 ;
        RECT 626.550 490.050 627.450 493.950 ;
        RECT 626.550 488.550 631.050 490.050 ;
        RECT 627.000 487.950 631.050 488.550 ;
        RECT 643.950 450.450 648.000 451.050 ;
        RECT 643.950 448.950 648.450 450.450 ;
        RECT 647.550 444.450 648.450 448.950 ;
        RECT 652.950 444.450 655.050 445.050 ;
        RECT 647.550 443.550 655.050 444.450 ;
        RECT 652.950 442.950 655.050 443.550 ;
      LAYER via1 ;
        RECT 628.950 493.950 631.050 496.050 ;
        RECT 628.950 487.950 631.050 490.050 ;
      LAYER metal2 ;
        RECT 398.400 964.050 399.450 984.450 ;
        RECT 391.950 961.950 394.050 964.050 ;
        RECT 397.950 961.950 400.050 964.050 ;
        RECT 392.400 952.050 393.450 961.950 ;
        RECT 391.950 949.950 394.050 952.050 ;
        RECT 400.950 949.950 403.050 952.050 ;
        RECT 392.400 878.400 393.600 880.650 ;
        RECT 392.400 871.050 393.450 878.400 ;
        RECT 401.400 871.050 402.450 949.950 ;
        RECT 391.950 868.950 394.050 871.050 ;
        RECT 400.950 868.950 403.050 871.050 ;
        RECT 427.950 868.950 430.050 871.050 ;
        RECT 428.400 787.050 429.450 868.950 ;
        RECT 553.950 811.950 556.050 814.050 ;
        RECT 685.950 811.950 688.050 814.050 ;
        RECT 554.400 808.050 555.450 811.950 ;
        RECT 520.950 805.950 523.050 808.050 ;
        RECT 553.800 805.950 555.900 808.050 ;
        RECT 458.400 800.400 459.600 802.650 ;
        RECT 458.400 787.050 459.450 800.400 ;
        RECT 521.400 787.050 522.450 805.950 ;
        RECT 686.400 801.900 687.450 811.950 ;
        RECT 692.400 801.900 693.600 802.650 ;
        RECT 685.950 799.800 688.050 801.900 ;
        RECT 691.950 799.800 694.050 801.900 ;
        RECT 397.950 784.950 400.050 787.050 ;
        RECT 427.950 784.950 430.050 787.050 ;
        RECT 457.950 784.950 460.050 787.050 ;
        RECT 520.950 784.950 523.050 787.050 ;
        RECT 398.400 766.050 399.450 784.950 ;
        RECT 364.950 762.000 367.050 766.050 ;
        RECT 397.950 763.950 400.050 766.050 ;
        RECT 365.400 760.350 366.600 762.000 ;
        RECT 398.400 730.050 399.450 763.950 ;
        RECT 382.950 727.950 385.050 730.050 ;
        RECT 397.950 727.950 400.050 730.050 ;
        RECT 323.400 678.000 324.600 679.650 ;
        RECT 322.950 673.950 325.050 678.000 ;
        RECT 383.400 676.050 384.450 727.950 ;
        RECT 382.950 673.950 385.050 676.050 ;
        RECT 472.950 673.950 475.050 676.050 ;
        RECT 473.400 643.050 474.450 673.950 ;
        RECT 472.950 640.950 475.050 643.050 ;
        RECT 490.950 640.650 493.050 642.750 ;
        RECT 491.400 547.050 492.450 640.650 ;
        RECT 490.950 544.950 493.050 547.050 ;
        RECT 568.950 544.950 571.050 547.050 ;
        RECT 569.400 541.050 570.450 544.950 ;
        RECT 568.950 538.950 571.050 541.050 ;
        RECT 595.950 538.950 598.050 541.050 ;
        RECT 596.400 529.050 597.450 538.950 ;
        RECT 595.950 526.950 598.050 529.050 ;
        RECT 619.950 527.100 622.050 529.200 ;
        RECT 620.400 526.350 621.600 527.100 ;
        RECT 628.800 520.950 630.900 523.050 ;
        RECT 629.400 496.050 630.450 520.950 ;
        RECT 628.950 493.950 631.050 496.050 ;
        RECT 628.950 487.950 631.050 490.050 ;
        RECT 629.400 454.050 630.450 487.950 ;
        RECT 628.950 451.950 631.050 454.050 ;
        RECT 643.950 448.950 646.050 454.050 ;
        RECT 652.950 442.950 655.050 445.050 ;
        RECT 653.400 421.050 654.450 442.950 ;
        RECT 652.950 418.950 655.050 421.050 ;
        RECT 662.400 411.900 663.600 412.650 ;
        RECT 661.950 409.800 664.050 411.900 ;
      LAYER via2 ;
        RECT 364.950 763.950 367.050 766.050 ;
        RECT 643.950 451.950 646.050 454.050 ;
      LAYER metal3 ;
        RECT 391.950 870.600 394.050 871.050 ;
        RECT 400.950 870.600 403.050 871.050 ;
        RECT 427.950 870.600 430.050 871.050 ;
        RECT 391.950 869.400 430.050 870.600 ;
        RECT 391.950 868.950 394.050 869.400 ;
        RECT 400.950 868.950 403.050 869.400 ;
        RECT 427.950 868.950 430.050 869.400 ;
        RECT 553.950 813.600 556.050 814.050 ;
        RECT 685.950 813.600 688.050 814.050 ;
        RECT 553.950 812.400 688.050 813.600 ;
        RECT 553.950 811.950 556.050 812.400 ;
        RECT 685.950 811.950 688.050 812.400 ;
        RECT 520.950 807.600 523.050 808.050 ;
        RECT 553.800 807.600 555.900 808.050 ;
        RECT 520.950 806.400 555.900 807.600 ;
        RECT 520.950 805.950 523.050 806.400 ;
        RECT 553.800 805.950 555.900 806.400 ;
        RECT 685.950 801.450 688.050 801.900 ;
        RECT 691.950 801.450 694.050 801.900 ;
        RECT 685.950 800.250 694.050 801.450 ;
        RECT 685.950 799.800 688.050 800.250 ;
        RECT 691.950 799.800 694.050 800.250 ;
        RECT 397.950 786.600 400.050 787.050 ;
        RECT 427.950 786.600 430.050 787.050 ;
        RECT 457.950 786.600 460.050 787.050 ;
        RECT 520.950 786.600 523.050 787.050 ;
        RECT 397.950 785.400 523.050 786.600 ;
        RECT 397.950 784.950 400.050 785.400 ;
        RECT 427.950 784.950 430.050 785.400 ;
        RECT 457.950 784.950 460.050 785.400 ;
        RECT 520.950 784.950 523.050 785.400 ;
        RECT 364.950 765.600 367.050 766.050 ;
        RECT 397.950 765.600 400.050 766.050 ;
        RECT 364.950 764.400 400.050 765.600 ;
        RECT 364.950 763.950 367.050 764.400 ;
        RECT 397.950 763.950 400.050 764.400 ;
        RECT 382.950 729.600 385.050 730.050 ;
        RECT 397.950 729.600 400.050 730.050 ;
        RECT 382.950 728.400 400.050 729.600 ;
        RECT 382.950 727.950 385.050 728.400 ;
        RECT 397.950 727.950 400.050 728.400 ;
        RECT 322.950 675.600 325.050 676.050 ;
        RECT 382.950 675.600 385.050 676.050 ;
        RECT 472.950 675.600 475.050 676.050 ;
        RECT 322.950 674.400 475.050 675.600 ;
        RECT 322.950 673.950 325.050 674.400 ;
        RECT 382.950 673.950 385.050 674.400 ;
        RECT 472.950 673.950 475.050 674.400 ;
        RECT 490.950 546.600 493.050 547.050 ;
        RECT 568.950 546.600 571.050 547.050 ;
        RECT 490.950 545.400 571.050 546.600 ;
        RECT 490.950 544.950 493.050 545.400 ;
        RECT 568.950 544.950 571.050 545.400 ;
        RECT 568.950 540.600 571.050 541.050 ;
        RECT 595.950 540.600 598.050 541.050 ;
        RECT 568.950 539.400 598.050 540.600 ;
        RECT 568.950 538.950 571.050 539.400 ;
        RECT 595.950 538.950 598.050 539.400 ;
        RECT 595.950 525.600 598.050 529.050 ;
        RECT 619.950 527.100 622.050 529.200 ;
        RECT 620.400 525.600 621.600 527.100 ;
        RECT 595.950 525.000 627.600 525.600 ;
        RECT 596.400 524.400 627.600 525.000 ;
        RECT 626.400 523.050 627.600 524.400 ;
        RECT 626.400 521.400 630.900 523.050 ;
        RECT 627.000 520.950 630.900 521.400 ;
        RECT 628.950 453.600 631.050 454.050 ;
        RECT 643.950 453.600 646.050 454.050 ;
        RECT 628.950 452.400 646.050 453.600 ;
        RECT 628.950 451.950 631.050 452.400 ;
        RECT 643.950 451.950 646.050 452.400 ;
        RECT 652.950 420.600 657.000 421.050 ;
        RECT 652.950 418.950 657.600 420.600 ;
        RECT 656.400 411.600 657.600 418.950 ;
        RECT 661.950 411.600 664.050 411.900 ;
        RECT 656.400 410.400 664.050 411.600 ;
        RECT 661.950 409.800 664.050 410.400 ;
    END
  END Cin[7]
  PIN Cin[6]
    PORT
      LAYER metal1 ;
        RECT 343.950 810.450 346.050 811.050 ;
        RECT 352.950 810.450 355.050 811.050 ;
        RECT 343.950 809.550 355.050 810.450 ;
        RECT 343.950 808.950 346.050 809.550 ;
        RECT 352.950 808.950 355.050 809.550 ;
        RECT 751.950 732.450 754.050 733.050 ;
        RECT 757.950 732.450 760.050 733.050 ;
        RECT 751.950 731.550 760.050 732.450 ;
        RECT 751.950 730.950 754.050 731.550 ;
        RECT 757.950 730.950 760.050 731.550 ;
        RECT 772.950 657.450 775.050 658.050 ;
        RECT 767.550 656.550 775.050 657.450 ;
        RECT 767.550 651.450 768.450 656.550 ;
        RECT 772.950 655.950 775.050 656.550 ;
        RECT 772.950 651.450 775.050 652.050 ;
        RECT 767.550 650.550 775.050 651.450 ;
        RECT 772.950 649.950 775.050 650.550 ;
        RECT 781.950 609.450 784.050 610.050 ;
        RECT 787.950 609.450 790.050 610.050 ;
        RECT 781.950 608.550 790.050 609.450 ;
        RECT 781.950 607.950 784.050 608.550 ;
        RECT 787.950 607.950 790.050 608.550 ;
      LAYER metal2 ;
        RECT 449.400 979.050 450.450 984.450 ;
        RECT 448.950 976.950 451.050 979.050 ;
        RECT 463.950 976.950 466.050 979.050 ;
        RECT 373.950 889.950 376.050 892.050 ;
        RECT 374.400 859.050 375.450 889.950 ;
        RECT 464.400 889.200 465.450 976.950 ;
        RECT 439.950 885.000 442.050 889.050 ;
        RECT 463.950 887.100 466.050 889.200 ;
        RECT 475.950 886.950 478.050 889.050 ;
        RECT 440.400 883.350 441.600 885.000 ;
        RECT 476.400 871.050 477.450 886.950 ;
        RECT 658.950 883.950 661.050 886.050 ;
        RECT 685.950 884.100 688.050 886.200 ;
        RECT 694.950 884.100 697.050 886.200 ;
        RECT 475.950 868.950 478.050 871.050 ;
        RECT 568.950 868.950 571.050 871.050 ;
        RECT 343.950 856.950 346.050 859.050 ;
        RECT 373.950 856.950 376.050 859.050 ;
        RECT 344.400 841.200 345.450 856.950 ;
        RECT 569.400 850.050 570.450 868.950 ;
        RECT 659.400 856.050 660.450 883.950 ;
        RECT 686.400 883.350 687.600 884.100 ;
        RECT 695.400 865.050 696.450 884.100 ;
        RECT 694.950 862.950 697.050 865.050 ;
        RECT 724.950 862.950 727.050 865.050 ;
        RECT 628.950 853.950 631.050 856.050 ;
        RECT 658.950 853.950 661.050 856.050 ;
        RECT 629.400 850.050 630.450 853.950 ;
        RECT 568.950 847.950 571.050 850.050 ;
        RECT 628.950 847.950 631.050 850.050 ;
        RECT 337.950 838.950 340.050 841.050 ;
        RECT 343.950 839.100 346.050 841.200 ;
        RECT 629.400 840.600 630.450 847.950 ;
        RECT 338.400 817.050 339.450 838.950 ;
        RECT 344.400 838.350 345.600 839.100 ;
        RECT 629.400 838.350 630.600 840.600 ;
        RECT 337.950 814.950 340.050 817.050 ;
        RECT 343.950 814.950 346.050 817.050 ;
        RECT 344.400 811.050 345.450 814.950 ;
        RECT 725.400 814.050 726.450 862.950 ;
        RECT 715.950 811.950 718.050 814.050 ;
        RECT 724.950 811.950 727.050 814.050 ;
        RECT 748.950 811.950 751.050 814.050 ;
        RECT 343.950 808.950 346.050 811.050 ;
        RECT 352.950 808.950 355.050 811.050 ;
        RECT 344.400 807.600 345.450 808.950 ;
        RECT 344.400 805.350 345.600 807.600 ;
        RECT 353.400 790.050 354.450 808.950 ;
        RECT 716.400 807.600 717.450 811.950 ;
        RECT 716.400 805.350 717.600 807.600 ;
        RECT 749.400 807.450 750.450 811.950 ;
        RECT 749.400 806.400 753.450 807.450 ;
        RECT 331.950 787.950 334.050 790.050 ;
        RECT 352.950 787.950 355.050 790.050 ;
        RECT 332.400 763.200 333.450 787.950 ;
        RECT 316.950 761.100 319.050 763.200 ;
        RECT 317.400 760.350 318.600 761.100 ;
        RECT 322.950 760.950 325.050 763.050 ;
        RECT 331.950 761.100 334.050 763.200 ;
        RECT 323.400 732.450 324.450 760.950 ;
        RECT 752.400 733.050 753.450 806.400 ;
        RECT 320.400 731.400 324.450 732.450 ;
        RECT 320.400 729.600 321.450 731.400 ;
        RECT 751.950 730.950 754.050 733.050 ;
        RECT 757.950 730.950 760.050 733.050 ;
        RECT 320.400 727.350 321.600 729.600 ;
        RECT 758.400 708.450 759.450 730.950 ;
        RECT 755.400 707.400 759.450 708.450 ;
        RECT 755.400 664.050 756.450 707.400 ;
        RECT 754.950 661.950 757.050 664.050 ;
        RECT 772.950 661.950 775.050 664.050 ;
        RECT 773.400 658.050 774.450 661.950 ;
        RECT 772.950 655.950 775.050 658.050 ;
        RECT 772.950 649.950 775.050 652.050 ;
        RECT 773.400 637.050 774.450 649.950 ;
        RECT 772.950 634.950 775.050 637.050 ;
        RECT 781.950 634.950 784.050 637.050 ;
        RECT 782.400 610.050 783.450 634.950 ;
        RECT 781.950 606.000 784.050 610.050 ;
        RECT 787.950 607.950 790.050 610.050 ;
        RECT 782.400 604.350 783.600 606.000 ;
        RECT 788.400 598.050 789.450 607.950 ;
        RECT 775.950 595.950 778.050 598.050 ;
        RECT 787.950 595.950 790.050 598.050 ;
        RECT 776.400 550.050 777.450 595.950 ;
        RECT 715.950 547.950 718.050 550.050 ;
        RECT 775.950 547.950 778.050 550.050 ;
        RECT 716.400 496.200 717.450 547.950 ;
        RECT 634.950 494.100 637.050 496.200 ;
        RECT 715.950 494.100 718.050 496.200 ;
        RECT 724.950 494.100 727.050 496.200 ;
        RECT 635.400 493.350 636.600 494.100 ;
        RECT 619.950 487.950 622.050 490.050 ;
        RECT 620.400 427.050 621.450 487.950 ;
        RECT 716.400 427.050 717.450 494.100 ;
        RECT 725.400 493.350 726.600 494.100 ;
        RECT 763.950 449.100 766.050 451.200 ;
        RECT 775.950 449.100 778.050 451.200 ;
        RECT 764.400 427.050 765.450 449.100 ;
        RECT 776.400 448.350 777.600 449.100 ;
        RECT 619.950 424.950 622.050 427.050 ;
        RECT 685.950 424.950 688.050 427.050 ;
        RECT 715.950 424.950 718.050 427.050 ;
        RECT 763.950 424.950 766.050 427.050 ;
        RECT 686.400 417.600 687.450 424.950 ;
        RECT 764.400 417.600 765.450 424.950 ;
        RECT 686.400 415.350 687.600 417.600 ;
        RECT 764.400 415.350 765.600 417.600 ;
      LAYER via2 ;
        RECT 439.950 886.950 442.050 889.050 ;
      LAYER metal3 ;
        RECT 448.950 978.600 451.050 979.050 ;
        RECT 463.950 978.600 466.050 979.050 ;
        RECT 448.950 977.400 466.050 978.600 ;
        RECT 448.950 976.950 451.050 977.400 ;
        RECT 463.950 976.950 466.050 977.400 ;
        RECT 373.950 891.600 376.050 892.050 ;
        RECT 373.950 890.400 441.600 891.600 ;
        RECT 373.950 889.950 376.050 890.400 ;
        RECT 440.400 889.050 441.600 890.400 ;
        RECT 439.950 888.600 442.050 889.050 ;
        RECT 463.950 888.600 466.050 889.200 ;
        RECT 475.950 888.600 478.050 889.050 ;
        RECT 439.950 887.400 478.050 888.600 ;
        RECT 439.950 886.950 442.050 887.400 ;
        RECT 463.950 887.100 466.050 887.400 ;
        RECT 475.950 886.950 478.050 887.400 ;
        RECT 658.950 885.600 661.050 886.050 ;
        RECT 685.950 885.750 688.050 886.200 ;
        RECT 694.950 885.750 697.050 886.200 ;
        RECT 685.950 885.600 697.050 885.750 ;
        RECT 658.950 884.550 697.050 885.600 ;
        RECT 658.950 884.400 688.050 884.550 ;
        RECT 658.950 883.950 661.050 884.400 ;
        RECT 685.950 884.100 688.050 884.400 ;
        RECT 694.950 884.100 697.050 884.550 ;
        RECT 475.950 870.600 478.050 871.050 ;
        RECT 568.950 870.600 571.050 871.050 ;
        RECT 475.950 869.400 571.050 870.600 ;
        RECT 475.950 868.950 478.050 869.400 ;
        RECT 568.950 868.950 571.050 869.400 ;
        RECT 694.950 864.600 697.050 865.050 ;
        RECT 724.950 864.600 727.050 865.050 ;
        RECT 694.950 863.400 727.050 864.600 ;
        RECT 694.950 862.950 697.050 863.400 ;
        RECT 724.950 862.950 727.050 863.400 ;
        RECT 343.950 858.600 346.050 859.050 ;
        RECT 373.950 858.600 376.050 859.050 ;
        RECT 343.950 857.400 376.050 858.600 ;
        RECT 343.950 856.950 346.050 857.400 ;
        RECT 373.950 856.950 376.050 857.400 ;
        RECT 628.950 855.600 631.050 856.050 ;
        RECT 658.950 855.600 661.050 856.050 ;
        RECT 628.950 854.400 661.050 855.600 ;
        RECT 628.950 853.950 631.050 854.400 ;
        RECT 658.950 853.950 661.050 854.400 ;
        RECT 568.950 849.600 571.050 850.050 ;
        RECT 628.950 849.600 631.050 850.050 ;
        RECT 568.950 848.400 631.050 849.600 ;
        RECT 568.950 847.950 571.050 848.400 ;
        RECT 628.950 847.950 631.050 848.400 ;
        RECT 337.950 840.600 340.050 841.050 ;
        RECT 343.950 840.600 346.050 841.200 ;
        RECT 337.950 839.400 346.050 840.600 ;
        RECT 337.950 838.950 340.050 839.400 ;
        RECT 343.950 839.100 346.050 839.400 ;
        RECT 337.950 816.600 340.050 817.050 ;
        RECT 343.950 816.600 346.050 817.050 ;
        RECT 337.950 815.400 346.050 816.600 ;
        RECT 337.950 814.950 340.050 815.400 ;
        RECT 343.950 814.950 346.050 815.400 ;
        RECT 715.950 813.600 718.050 814.050 ;
        RECT 724.950 813.600 727.050 814.050 ;
        RECT 748.950 813.600 751.050 814.050 ;
        RECT 715.950 812.400 751.050 813.600 ;
        RECT 715.950 811.950 718.050 812.400 ;
        RECT 724.950 811.950 727.050 812.400 ;
        RECT 748.950 811.950 751.050 812.400 ;
        RECT 331.950 789.600 334.050 790.050 ;
        RECT 352.950 789.600 355.050 790.050 ;
        RECT 331.950 788.400 355.050 789.600 ;
        RECT 331.950 787.950 334.050 788.400 ;
        RECT 352.950 787.950 355.050 788.400 ;
        RECT 316.950 762.750 319.050 763.200 ;
        RECT 322.950 762.750 325.050 763.050 ;
        RECT 331.950 762.750 334.050 763.200 ;
        RECT 316.950 761.550 334.050 762.750 ;
        RECT 316.950 761.100 319.050 761.550 ;
        RECT 322.950 760.950 325.050 761.550 ;
        RECT 331.950 761.100 334.050 761.550 ;
        RECT 754.950 663.600 757.050 664.050 ;
        RECT 772.950 663.600 775.050 664.050 ;
        RECT 754.950 662.400 775.050 663.600 ;
        RECT 754.950 661.950 757.050 662.400 ;
        RECT 772.950 661.950 775.050 662.400 ;
        RECT 772.950 636.600 775.050 637.050 ;
        RECT 781.950 636.600 784.050 637.050 ;
        RECT 772.950 635.400 784.050 636.600 ;
        RECT 772.950 634.950 775.050 635.400 ;
        RECT 781.950 634.950 784.050 635.400 ;
        RECT 775.950 597.600 778.050 598.050 ;
        RECT 787.950 597.600 790.050 598.050 ;
        RECT 775.950 596.400 790.050 597.600 ;
        RECT 775.950 595.950 778.050 596.400 ;
        RECT 787.950 595.950 790.050 596.400 ;
        RECT 715.950 549.600 718.050 550.050 ;
        RECT 775.950 549.600 778.050 550.050 ;
        RECT 715.950 548.400 778.050 549.600 ;
        RECT 715.950 547.950 718.050 548.400 ;
        RECT 775.950 547.950 778.050 548.400 ;
        RECT 634.950 494.100 637.050 496.200 ;
        RECT 715.950 495.750 718.050 496.200 ;
        RECT 724.950 495.750 727.050 496.200 ;
        RECT 715.950 494.550 727.050 495.750 ;
        RECT 715.950 494.100 718.050 494.550 ;
        RECT 724.950 494.100 727.050 494.550 ;
        RECT 619.950 489.600 622.050 490.050 ;
        RECT 635.400 489.600 636.600 494.100 ;
        RECT 619.950 488.400 636.600 489.600 ;
        RECT 619.950 487.950 622.050 488.400 ;
        RECT 763.950 450.750 766.050 451.200 ;
        RECT 775.950 450.750 778.050 451.200 ;
        RECT 763.950 449.550 778.050 450.750 ;
        RECT 763.950 449.100 766.050 449.550 ;
        RECT 775.950 449.100 778.050 449.550 ;
        RECT 619.950 426.600 622.050 427.050 ;
        RECT 685.950 426.600 688.050 427.050 ;
        RECT 715.950 426.600 718.050 427.050 ;
        RECT 763.950 426.600 766.050 427.050 ;
        RECT 619.950 425.400 766.050 426.600 ;
        RECT 619.950 424.950 622.050 425.400 ;
        RECT 685.950 424.950 688.050 425.400 ;
        RECT 715.950 424.950 718.050 425.400 ;
        RECT 763.950 424.950 766.050 425.400 ;
    END
  END Cin[6]
  PIN Cin[5]
    PORT
      LAYER metal1 ;
        RECT 340.950 753.450 343.050 754.050 ;
        RECT 352.950 753.450 355.050 754.050 ;
        RECT 340.950 752.550 355.050 753.450 ;
        RECT 340.950 751.950 343.050 752.550 ;
        RECT 352.950 751.950 355.050 752.550 ;
        RECT 693.000 528.450 697.050 529.050 ;
        RECT 692.550 526.950 697.050 528.450 ;
        RECT 692.550 523.050 693.450 526.950 ;
        RECT 692.550 521.550 697.050 523.050 ;
        RECT 693.000 520.950 697.050 521.550 ;
        RECT 703.950 453.450 706.050 454.050 ;
        RECT 698.550 452.550 706.050 453.450 ;
        RECT 698.550 450.450 699.450 452.550 ;
        RECT 703.950 451.950 706.050 452.550 ;
        RECT 695.550 449.550 699.450 450.450 ;
        RECT 695.550 442.050 696.450 449.550 ;
        RECT 693.000 441.900 696.450 442.050 ;
        RECT 691.950 440.550 696.450 441.900 ;
        RECT 691.950 439.950 696.000 440.550 ;
        RECT 691.950 439.800 694.050 439.950 ;
      LAYER via1 ;
        RECT 694.950 526.950 697.050 529.050 ;
        RECT 694.950 520.950 697.050 523.050 ;
      LAYER metal2 ;
        RECT 425.400 979.050 426.450 984.450 ;
        RECT 418.950 976.950 421.050 979.050 ;
        RECT 424.950 976.950 427.050 979.050 ;
        RECT 419.400 886.050 420.450 976.950 ;
        RECT 418.950 883.950 421.050 886.050 ;
        RECT 424.950 884.100 427.050 886.200 ;
        RECT 433.950 884.100 436.050 886.200 ;
        RECT 425.400 877.050 426.450 884.100 ;
        RECT 434.400 883.350 435.600 884.100 ;
        RECT 424.950 874.950 427.050 877.050 ;
        RECT 430.950 874.650 433.050 876.750 ;
        RECT 431.400 841.200 432.450 874.650 ;
        RECT 430.950 839.100 433.050 841.200 ;
        RECT 436.950 839.100 439.050 841.200 ;
        RECT 431.400 811.050 432.450 839.100 ;
        RECT 437.400 838.350 438.600 839.100 ;
        RECT 337.950 807.000 340.050 811.050 ;
        RECT 358.950 808.950 361.050 811.050 ;
        RECT 430.950 808.950 433.050 811.050 ;
        RECT 338.400 805.350 339.600 807.000 ;
        RECT 359.400 796.050 360.450 808.950 ;
        RECT 721.950 806.100 724.050 808.200 ;
        RECT 722.400 805.350 723.600 806.100 ;
        RECT 709.950 799.950 712.050 802.050 ;
        RECT 358.950 793.950 361.050 796.050 ;
        RECT 370.950 793.950 373.050 796.050 ;
        RECT 341.400 756.000 342.600 757.650 ;
        RECT 340.950 751.950 343.050 756.000 ;
        RECT 352.950 748.950 355.050 754.050 ;
        RECT 371.400 751.050 372.450 793.950 ;
        RECT 710.400 784.050 711.450 799.950 ;
        RECT 685.950 781.950 688.050 784.050 ;
        RECT 709.950 781.950 712.050 784.050 ;
        RECT 370.950 748.950 373.050 751.050 ;
        RECT 341.400 722.400 342.600 724.650 ;
        RECT 341.400 715.050 342.450 722.400 ;
        RECT 353.400 715.050 354.450 748.950 ;
        RECT 686.400 721.050 687.450 781.950 ;
        RECT 685.950 718.950 688.050 721.050 ;
        RECT 700.950 718.950 703.050 721.050 ;
        RECT 340.950 712.950 343.050 715.050 ;
        RECT 352.950 712.950 355.050 715.050 ;
        RECT 553.950 712.950 556.050 715.050 ;
        RECT 554.400 664.050 555.450 712.950 ;
        RECT 701.400 664.050 702.450 718.950 ;
        RECT 553.950 661.950 556.050 664.050 ;
        RECT 577.950 661.800 580.050 663.900 ;
        RECT 700.950 661.950 703.050 664.050 ;
        RECT 578.400 625.050 579.450 661.800 ;
        RECT 667.950 658.950 670.050 661.050 ;
        RECT 668.400 651.600 669.450 658.950 ;
        RECT 668.400 649.350 669.600 651.600 ;
        RECT 701.400 643.050 702.450 661.950 ;
        RECT 710.400 645.000 711.600 646.650 ;
        RECT 700.950 640.950 703.050 643.050 ;
        RECT 709.950 640.950 712.050 645.000 ;
        RECT 701.400 625.050 702.450 640.950 ;
        RECT 577.950 622.950 580.050 625.050 ;
        RECT 700.950 622.950 703.050 625.050 ;
        RECT 701.400 598.050 702.450 622.950 ;
        RECT 700.950 595.950 703.050 598.050 ;
        RECT 706.950 595.950 709.050 598.050 ;
        RECT 707.400 559.050 708.450 595.950 ;
        RECT 694.950 556.950 697.050 559.050 ;
        RECT 706.950 556.950 709.050 559.050 ;
        RECT 695.400 529.050 696.450 556.950 ;
        RECT 694.950 526.950 697.050 529.050 ;
        RECT 694.950 520.950 697.050 523.050 ;
        RECT 695.400 502.050 696.450 520.950 ;
        RECT 694.950 499.950 697.050 502.050 ;
        RECT 706.950 496.950 709.050 499.050 ;
        RECT 707.400 477.450 708.450 496.950 ;
        RECT 704.400 476.400 708.450 477.450 ;
        RECT 704.400 454.050 705.450 476.400 ;
        RECT 703.950 451.950 706.050 454.050 ;
        RECT 691.950 439.800 694.050 441.900 ;
        RECT 692.400 418.200 693.450 439.800 ;
        RECT 691.950 416.100 694.050 418.200 ;
        RECT 712.950 416.100 715.050 418.200 ;
        RECT 736.950 416.100 739.050 418.200 ;
        RECT 692.400 415.350 693.600 416.100 ;
        RECT 713.400 415.350 714.600 416.100 ;
        RECT 737.400 415.350 738.600 416.100 ;
      LAYER via2 ;
        RECT 337.950 808.950 340.050 811.050 ;
      LAYER metal3 ;
        RECT 418.950 978.600 421.050 979.050 ;
        RECT 424.950 978.600 427.050 979.050 ;
        RECT 418.950 977.400 427.050 978.600 ;
        RECT 418.950 976.950 421.050 977.400 ;
        RECT 424.950 976.950 427.050 977.400 ;
        RECT 418.950 885.600 421.050 886.050 ;
        RECT 424.950 885.750 427.050 886.200 ;
        RECT 433.950 885.750 436.050 886.200 ;
        RECT 424.950 885.600 436.050 885.750 ;
        RECT 418.950 884.550 436.050 885.600 ;
        RECT 418.950 884.400 427.050 884.550 ;
        RECT 418.950 883.950 421.050 884.400 ;
        RECT 424.950 884.100 427.050 884.400 ;
        RECT 433.950 884.100 436.050 884.550 ;
        RECT 424.950 876.600 427.050 877.050 ;
        RECT 430.950 876.600 433.050 876.750 ;
        RECT 424.950 875.400 433.050 876.600 ;
        RECT 424.950 874.950 427.050 875.400 ;
        RECT 430.950 874.650 433.050 875.400 ;
        RECT 430.950 840.750 433.050 841.200 ;
        RECT 436.950 840.750 439.050 841.200 ;
        RECT 430.950 839.550 439.050 840.750 ;
        RECT 430.950 839.100 433.050 839.550 ;
        RECT 436.950 839.100 439.050 839.550 ;
        RECT 337.950 810.600 340.050 811.050 ;
        RECT 358.950 810.600 361.050 811.050 ;
        RECT 430.950 810.600 433.050 811.050 ;
        RECT 337.950 809.400 433.050 810.600 ;
        RECT 337.950 808.950 340.050 809.400 ;
        RECT 358.950 808.950 361.050 809.400 ;
        RECT 430.950 808.950 433.050 809.400 ;
        RECT 721.950 806.100 724.050 808.200 ;
        RECT 709.950 801.600 712.050 802.050 ;
        RECT 722.400 801.600 723.600 806.100 ;
        RECT 709.950 800.400 723.600 801.600 ;
        RECT 709.950 799.950 712.050 800.400 ;
        RECT 358.950 795.600 361.050 796.050 ;
        RECT 370.950 795.600 373.050 796.050 ;
        RECT 358.950 794.400 373.050 795.600 ;
        RECT 358.950 793.950 361.050 794.400 ;
        RECT 370.950 793.950 373.050 794.400 ;
        RECT 685.950 783.600 688.050 784.050 ;
        RECT 709.950 783.600 712.050 784.050 ;
        RECT 685.950 782.400 712.050 783.600 ;
        RECT 685.950 781.950 688.050 782.400 ;
        RECT 709.950 781.950 712.050 782.400 ;
        RECT 352.950 750.600 355.050 751.050 ;
        RECT 370.950 750.600 373.050 751.050 ;
        RECT 352.950 749.400 373.050 750.600 ;
        RECT 352.950 748.950 355.050 749.400 ;
        RECT 370.950 748.950 373.050 749.400 ;
        RECT 685.950 720.600 688.050 721.050 ;
        RECT 700.950 720.600 703.050 721.050 ;
        RECT 685.950 719.400 703.050 720.600 ;
        RECT 685.950 718.950 688.050 719.400 ;
        RECT 700.950 718.950 703.050 719.400 ;
        RECT 340.950 714.600 343.050 715.050 ;
        RECT 352.950 714.600 355.050 715.050 ;
        RECT 553.950 714.600 556.050 715.050 ;
        RECT 340.950 713.400 556.050 714.600 ;
        RECT 340.950 712.950 343.050 713.400 ;
        RECT 352.950 712.950 355.050 713.400 ;
        RECT 553.950 712.950 556.050 713.400 ;
        RECT 553.950 663.600 556.050 664.050 ;
        RECT 577.950 663.600 580.050 663.900 ;
        RECT 700.950 663.600 703.050 664.050 ;
        RECT 553.950 662.400 580.050 663.600 ;
        RECT 553.950 661.950 556.050 662.400 ;
        RECT 577.950 661.800 580.050 662.400 ;
        RECT 680.400 662.400 703.050 663.600 ;
        RECT 667.950 660.600 670.050 661.050 ;
        RECT 680.400 660.600 681.600 662.400 ;
        RECT 700.950 661.950 703.050 662.400 ;
        RECT 667.950 659.400 681.600 660.600 ;
        RECT 667.950 658.950 670.050 659.400 ;
        RECT 700.950 642.600 703.050 643.050 ;
        RECT 709.950 642.600 712.050 643.050 ;
        RECT 700.950 641.400 712.050 642.600 ;
        RECT 700.950 640.950 703.050 641.400 ;
        RECT 709.950 640.950 712.050 641.400 ;
        RECT 577.950 624.600 580.050 625.050 ;
        RECT 700.950 624.600 703.050 625.050 ;
        RECT 577.950 623.400 703.050 624.600 ;
        RECT 577.950 622.950 580.050 623.400 ;
        RECT 700.950 622.950 703.050 623.400 ;
        RECT 700.950 597.600 703.050 598.050 ;
        RECT 706.950 597.600 709.050 598.050 ;
        RECT 700.950 596.400 709.050 597.600 ;
        RECT 700.950 595.950 703.050 596.400 ;
        RECT 706.950 595.950 709.050 596.400 ;
        RECT 694.950 558.600 697.050 559.050 ;
        RECT 706.950 558.600 709.050 559.050 ;
        RECT 694.950 557.400 709.050 558.600 ;
        RECT 694.950 556.950 697.050 557.400 ;
        RECT 706.950 556.950 709.050 557.400 ;
        RECT 694.950 501.600 697.050 502.050 ;
        RECT 694.950 500.400 705.600 501.600 ;
        RECT 694.950 499.950 697.050 500.400 ;
        RECT 704.400 499.050 705.600 500.400 ;
        RECT 704.400 497.400 709.050 499.050 ;
        RECT 705.000 496.950 709.050 497.400 ;
        RECT 691.950 417.600 694.050 418.200 ;
        RECT 712.950 417.600 715.050 418.200 ;
        RECT 736.950 417.600 739.050 418.200 ;
        RECT 691.950 416.400 739.050 417.600 ;
        RECT 691.950 416.100 694.050 416.400 ;
        RECT 712.950 416.100 715.050 416.400 ;
        RECT 736.950 416.100 739.050 416.400 ;
    END
  END Cin[5]
  PIN Cin[4]
    PORT
      LAYER metal1 ;
        RECT 487.950 963.450 490.050 964.050 ;
        RECT 493.950 963.450 496.050 964.050 ;
        RECT 487.950 962.550 496.050 963.450 ;
        RECT 487.950 961.950 490.050 962.550 ;
        RECT 493.950 961.950 496.050 962.550 ;
        RECT 682.950 456.450 685.050 457.050 ;
        RECT 706.950 456.450 709.050 457.050 ;
        RECT 682.950 455.550 709.050 456.450 ;
        RECT 682.950 454.950 685.050 455.550 ;
        RECT 706.950 454.950 709.050 455.550 ;
        RECT 706.950 363.450 709.050 363.750 ;
        RECT 718.950 363.450 721.050 364.050 ;
        RECT 706.950 362.550 721.050 363.450 ;
        RECT 706.950 361.650 709.050 362.550 ;
        RECT 718.950 361.950 721.050 362.550 ;
        RECT 607.950 264.450 610.050 265.200 ;
        RECT 607.950 263.550 615.450 264.450 ;
        RECT 607.950 263.100 610.050 263.550 ;
        RECT 614.550 261.450 615.450 263.550 ;
        RECT 614.550 260.550 618.450 261.450 ;
        RECT 617.550 256.050 618.450 260.550 ;
        RECT 613.950 254.550 618.450 256.050 ;
        RECT 613.950 253.950 618.000 254.550 ;
      LAYER metal2 ;
        RECT 494.400 964.050 495.450 984.450 ;
        RECT 487.950 961.950 490.050 964.050 ;
        RECT 493.950 961.950 496.050 964.050 ;
        RECT 488.400 904.050 489.450 961.950 ;
        RECT 487.950 901.950 490.050 904.050 ;
        RECT 511.950 901.950 514.050 904.050 ;
        RECT 484.950 811.950 487.050 814.050 ;
        RECT 499.950 811.950 502.050 814.050 ;
        RECT 485.400 807.600 486.450 811.950 ;
        RECT 500.400 808.200 501.450 811.950 ;
        RECT 512.400 808.200 513.450 901.950 ;
        RECT 485.400 805.350 486.600 807.600 ;
        RECT 499.950 806.100 502.050 808.200 ;
        RECT 511.950 806.100 514.050 808.200 ;
        RECT 500.400 766.050 501.450 806.100 ;
        RECT 512.400 805.350 513.600 806.100 ;
        RECT 746.400 800.400 747.600 802.650 ;
        RECT 746.400 789.450 747.450 800.400 ;
        RECT 743.400 788.400 747.450 789.450 ;
        RECT 743.400 781.050 744.450 788.400 ;
        RECT 658.950 778.950 661.050 781.050 ;
        RECT 742.950 778.950 745.050 781.050 ;
        RECT 659.400 766.050 660.450 778.950 ;
        RECT 499.950 763.950 502.050 766.050 ;
        RECT 580.950 763.950 583.050 766.050 ;
        RECT 658.950 763.950 661.050 766.050 ;
        RECT 581.400 754.050 582.450 763.950 ;
        RECT 580.950 751.950 583.050 754.050 ;
        RECT 589.950 751.950 592.050 754.050 ;
        RECT 560.400 722.400 561.600 724.650 ;
        RECT 560.400 703.050 561.450 722.400 ;
        RECT 590.400 703.050 591.450 751.950 ;
        RECT 559.950 700.950 562.050 703.050 ;
        RECT 589.950 700.950 592.050 703.050 ;
        RECT 628.950 700.950 631.050 703.050 ;
        RECT 629.400 678.450 630.450 700.950 ;
        RECT 629.400 678.000 633.450 678.450 ;
        RECT 629.400 677.400 634.050 678.000 ;
        RECT 631.950 673.950 634.050 677.400 ;
        RECT 655.950 673.950 658.050 676.050 ;
        RECT 656.400 640.050 657.450 673.950 ;
        RECT 646.950 637.950 649.050 640.050 ;
        RECT 655.950 637.950 658.050 640.050 ;
        RECT 647.400 589.050 648.450 637.950 ;
        RECT 646.950 586.950 649.050 589.050 ;
        RECT 658.950 586.950 661.050 589.050 ;
        RECT 659.400 519.450 660.450 586.950 ;
        RECT 659.400 518.400 663.450 519.450 ;
        RECT 662.400 484.050 663.450 518.400 ;
        RECT 661.950 481.950 664.050 484.050 ;
        RECT 679.950 481.950 682.050 484.050 ;
        RECT 680.400 474.450 681.450 481.950 ;
        RECT 680.400 473.400 684.450 474.450 ;
        RECT 683.400 457.050 684.450 473.400 ;
        RECT 682.950 454.950 685.050 457.050 ;
        RECT 706.950 454.950 709.050 460.050 ;
        RECT 718.950 457.950 721.050 460.050 ;
        RECT 754.950 457.950 757.050 460.050 ;
        RECT 719.400 444.450 720.450 457.950 ;
        RECT 755.400 450.600 756.450 457.950 ;
        RECT 755.400 448.350 756.600 450.600 ;
        RECT 719.400 443.400 723.450 444.450 ;
        RECT 722.400 411.450 723.450 443.400 ;
        RECT 719.400 410.400 723.450 411.450 ;
        RECT 719.400 364.050 720.450 410.400 ;
        RECT 706.950 361.650 709.050 363.750 ;
        RECT 718.950 361.950 721.050 364.050 ;
        RECT 707.400 337.050 708.450 361.650 ;
        RECT 706.950 334.950 709.050 337.050 ;
        RECT 655.950 331.950 658.050 334.050 ;
        RECT 740.400 333.900 741.600 334.650 ;
        RECT 656.400 325.050 657.450 331.950 ;
        RECT 739.950 331.800 742.050 333.900 ;
        RECT 622.950 322.950 625.050 325.050 ;
        RECT 655.950 322.950 658.050 325.050 ;
        RECT 623.400 301.050 624.450 322.950 ;
        RECT 607.950 298.950 610.050 301.050 ;
        RECT 622.950 298.950 625.050 301.050 ;
        RECT 608.400 265.200 609.450 298.950 ;
        RECT 607.950 263.100 610.050 265.200 ;
        RECT 613.950 253.950 616.050 256.050 ;
        RECT 595.950 216.000 598.050 220.050 ;
        RECT 610.950 219.450 613.050 220.050 ;
        RECT 614.400 219.450 615.450 253.950 ;
        RECT 610.950 218.400 615.450 219.450 ;
        RECT 610.950 216.000 613.050 218.400 ;
        RECT 596.400 214.350 597.600 216.000 ;
        RECT 611.400 214.350 612.600 216.000 ;
      LAYER via2 ;
        RECT 706.950 457.950 709.050 460.050 ;
        RECT 595.950 217.950 598.050 220.050 ;
        RECT 610.950 217.950 613.050 220.050 ;
      LAYER metal3 ;
        RECT 487.950 903.600 490.050 904.050 ;
        RECT 511.950 903.600 514.050 904.050 ;
        RECT 487.950 902.400 514.050 903.600 ;
        RECT 487.950 901.950 490.050 902.400 ;
        RECT 511.950 901.950 514.050 902.400 ;
        RECT 484.950 813.600 487.050 814.050 ;
        RECT 499.950 813.600 502.050 814.050 ;
        RECT 484.950 812.400 502.050 813.600 ;
        RECT 484.950 811.950 487.050 812.400 ;
        RECT 499.950 811.950 502.050 812.400 ;
        RECT 499.950 807.750 502.050 808.200 ;
        RECT 511.950 807.750 514.050 808.200 ;
        RECT 499.950 806.550 514.050 807.750 ;
        RECT 499.950 806.100 502.050 806.550 ;
        RECT 511.950 806.100 514.050 806.550 ;
        RECT 658.950 780.600 661.050 781.050 ;
        RECT 742.950 780.600 745.050 781.050 ;
        RECT 658.950 779.400 745.050 780.600 ;
        RECT 658.950 778.950 661.050 779.400 ;
        RECT 742.950 778.950 745.050 779.400 ;
        RECT 499.950 765.600 502.050 766.050 ;
        RECT 580.950 765.600 583.050 766.050 ;
        RECT 658.950 765.600 661.050 766.050 ;
        RECT 499.950 764.400 661.050 765.600 ;
        RECT 499.950 763.950 502.050 764.400 ;
        RECT 580.950 763.950 583.050 764.400 ;
        RECT 658.950 763.950 661.050 764.400 ;
        RECT 580.950 753.600 583.050 754.050 ;
        RECT 589.950 753.600 592.050 754.050 ;
        RECT 580.950 752.400 592.050 753.600 ;
        RECT 580.950 751.950 583.050 752.400 ;
        RECT 589.950 751.950 592.050 752.400 ;
        RECT 559.950 702.600 562.050 703.050 ;
        RECT 589.950 702.600 592.050 703.050 ;
        RECT 628.950 702.600 631.050 703.050 ;
        RECT 559.950 701.400 631.050 702.600 ;
        RECT 559.950 700.950 562.050 701.400 ;
        RECT 589.950 700.950 592.050 701.400 ;
        RECT 628.950 700.950 631.050 701.400 ;
        RECT 631.950 675.600 634.050 676.050 ;
        RECT 655.950 675.600 658.050 676.050 ;
        RECT 631.950 674.400 658.050 675.600 ;
        RECT 631.950 673.950 634.050 674.400 ;
        RECT 655.950 673.950 658.050 674.400 ;
        RECT 646.950 639.600 649.050 640.050 ;
        RECT 655.950 639.600 658.050 640.050 ;
        RECT 646.950 638.400 658.050 639.600 ;
        RECT 646.950 637.950 649.050 638.400 ;
        RECT 655.950 637.950 658.050 638.400 ;
        RECT 646.950 588.600 649.050 589.050 ;
        RECT 658.950 588.600 661.050 589.050 ;
        RECT 646.950 587.400 661.050 588.600 ;
        RECT 646.950 586.950 649.050 587.400 ;
        RECT 658.950 586.950 661.050 587.400 ;
        RECT 661.950 483.600 664.050 484.050 ;
        RECT 679.950 483.600 682.050 484.050 ;
        RECT 661.950 482.400 682.050 483.600 ;
        RECT 661.950 481.950 664.050 482.400 ;
        RECT 679.950 481.950 682.050 482.400 ;
        RECT 706.950 459.600 709.050 460.050 ;
        RECT 718.950 459.600 721.050 460.050 ;
        RECT 754.950 459.600 757.050 460.050 ;
        RECT 706.950 458.400 757.050 459.600 ;
        RECT 706.950 457.950 709.050 458.400 ;
        RECT 718.950 457.950 721.050 458.400 ;
        RECT 754.950 457.950 757.050 458.400 ;
        RECT 706.950 336.600 709.050 337.050 ;
        RECT 686.400 335.400 738.600 336.600 ;
        RECT 655.950 333.600 658.050 334.050 ;
        RECT 686.400 333.600 687.600 335.400 ;
        RECT 706.950 334.950 709.050 335.400 ;
        RECT 655.950 332.400 687.600 333.600 ;
        RECT 737.400 333.600 738.600 335.400 ;
        RECT 739.950 333.600 742.050 333.900 ;
        RECT 737.400 332.400 742.050 333.600 ;
        RECT 655.950 331.950 658.050 332.400 ;
        RECT 739.950 331.800 742.050 332.400 ;
        RECT 622.950 324.600 625.050 325.050 ;
        RECT 655.950 324.600 658.050 325.050 ;
        RECT 622.950 323.400 658.050 324.600 ;
        RECT 622.950 322.950 625.050 323.400 ;
        RECT 655.950 322.950 658.050 323.400 ;
        RECT 607.950 300.600 610.050 301.050 ;
        RECT 622.950 300.600 625.050 301.050 ;
        RECT 607.950 299.400 625.050 300.600 ;
        RECT 607.950 298.950 610.050 299.400 ;
        RECT 622.950 298.950 625.050 299.400 ;
        RECT 595.950 219.600 598.050 220.050 ;
        RECT 610.950 219.600 613.050 220.050 ;
        RECT 595.950 218.400 613.050 219.600 ;
        RECT 595.950 217.950 598.050 218.400 ;
        RECT 610.950 217.950 613.050 218.400 ;
    END
  END Cin[4]
  PIN Cin[3]
    PORT
      LAYER metal1 ;
        RECT 640.950 720.450 643.050 721.050 ;
        RECT 652.950 720.450 655.050 721.050 ;
        RECT 640.950 719.550 655.050 720.450 ;
        RECT 640.950 718.950 643.050 719.550 ;
        RECT 652.950 718.950 655.050 719.550 ;
        RECT 598.950 606.450 603.000 607.050 ;
        RECT 598.950 604.950 603.450 606.450 ;
        RECT 602.550 601.050 603.450 604.950 ;
        RECT 598.950 599.550 603.450 601.050 ;
        RECT 598.950 598.950 603.000 599.550 ;
        RECT 679.950 375.450 682.050 376.050 ;
        RECT 674.550 374.550 682.050 375.450 ;
        RECT 674.550 372.450 675.450 374.550 ;
        RECT 679.950 373.950 682.050 374.550 ;
        RECT 671.550 371.550 675.450 372.450 ;
        RECT 671.550 367.050 672.450 371.550 ;
        RECT 671.550 365.550 676.050 367.050 ;
        RECT 672.000 364.950 676.050 365.550 ;
        RECT 673.950 339.450 676.050 343.050 ;
        RECT 673.950 339.000 678.450 339.450 ;
        RECT 674.550 338.550 678.450 339.000 ;
        RECT 677.550 334.050 678.450 338.550 ;
        RECT 673.950 332.550 678.450 334.050 ;
        RECT 673.950 331.950 678.000 332.550 ;
        RECT 391.950 129.450 394.050 130.050 ;
        RECT 400.950 129.450 403.050 130.050 ;
        RECT 391.950 128.550 403.050 129.450 ;
        RECT 391.950 127.950 394.050 128.550 ;
        RECT 400.950 127.950 403.050 128.550 ;
        RECT 685.950 36.450 688.050 37.050 ;
        RECT 694.950 36.450 697.050 37.050 ;
        RECT 685.950 35.550 697.050 36.450 ;
        RECT 685.950 34.950 688.050 35.550 ;
        RECT 694.950 34.950 697.050 35.550 ;
      LAYER via1 ;
        RECT 673.950 364.950 676.050 367.050 ;
        RECT 673.950 340.950 676.050 343.050 ;
      LAYER metal2 ;
        RECT 472.950 806.100 475.050 808.200 ;
        RECT 490.950 806.100 493.050 808.200 ;
        RECT 473.400 783.450 474.450 806.100 ;
        RECT 491.400 805.350 492.600 806.100 ;
        RECT 470.400 782.400 474.450 783.450 ;
        RECT 470.400 757.050 471.450 782.400 ;
        RECT 469.950 754.950 472.050 757.050 ;
        RECT 485.400 756.900 486.600 757.650 ;
        RECT 484.950 754.800 487.050 756.900 ;
        RECT 499.950 754.800 502.050 756.900 ;
        RECT 500.400 751.050 501.450 754.800 ;
        RECT 499.950 748.950 502.050 751.050 ;
        RECT 619.950 748.950 622.050 751.050 ;
        RECT 620.400 739.050 621.450 748.950 ;
        RECT 619.950 736.950 622.050 739.050 ;
        RECT 640.950 736.950 643.050 739.050 ;
        RECT 641.400 721.050 642.450 736.950 ;
        RECT 724.950 733.950 727.050 736.050 ;
        RECT 725.400 729.600 726.450 733.950 ;
        RECT 725.400 727.350 726.600 729.600 ;
        RECT 653.400 722.400 654.600 724.650 ;
        RECT 653.400 721.050 654.450 722.400 ;
        RECT 640.950 718.950 643.050 721.050 ;
        RECT 652.950 718.950 655.050 721.050 ;
        RECT 653.400 702.450 654.450 718.950 ;
        RECT 650.400 701.400 654.450 702.450 ;
        RECT 650.400 684.450 651.450 701.400 ;
        RECT 647.400 683.400 651.450 684.450 ;
        RECT 647.400 667.050 648.450 683.400 ;
        RECT 595.950 664.950 598.050 667.050 ;
        RECT 646.950 664.950 649.050 667.050 ;
        RECT 596.400 612.450 597.450 664.950 ;
        RECT 596.400 611.400 600.450 612.450 ;
        RECT 599.400 607.050 600.450 611.400 ;
        RECT 598.950 604.950 601.050 607.050 ;
        RECT 598.950 597.450 601.050 601.050 ;
        RECT 596.400 597.000 601.050 597.450 ;
        RECT 596.400 596.400 600.450 597.000 ;
        RECT 596.400 574.050 597.450 596.400 ;
        RECT 595.950 571.950 598.050 574.050 ;
        RECT 595.950 565.950 598.050 568.050 ;
        RECT 596.400 547.050 597.450 565.950 ;
        RECT 586.950 544.950 589.050 547.050 ;
        RECT 595.950 544.950 598.050 547.050 ;
        RECT 574.950 527.100 577.050 529.200 ;
        RECT 580.950 527.100 583.050 529.200 ;
        RECT 587.400 529.050 588.450 544.950 ;
        RECT 575.400 513.450 576.450 527.100 ;
        RECT 581.400 526.350 582.600 527.100 ;
        RECT 586.950 526.950 589.050 529.050 ;
        RECT 572.400 512.400 576.450 513.450 ;
        RECT 572.400 484.050 573.450 512.400 ;
        RECT 677.400 488.400 678.600 490.650 ;
        RECT 571.950 481.950 574.050 484.050 ;
        RECT 610.950 481.950 613.050 484.050 ;
        RECT 611.400 454.050 612.450 481.950 ;
        RECT 677.400 463.050 678.450 488.400 ;
        RECT 676.950 460.950 679.050 463.050 ;
        RECT 688.950 460.950 691.050 463.050 ;
        RECT 610.950 451.950 613.050 454.050 ;
        RECT 628.950 439.950 631.050 442.050 ;
        RECT 629.400 424.050 630.450 439.950 ;
        RECT 628.950 421.950 631.050 424.050 ;
        RECT 689.400 421.050 690.450 460.950 ;
        RECT 688.950 418.950 691.050 421.050 ;
        RECT 679.950 409.950 682.050 412.050 ;
        RECT 680.400 376.050 681.450 409.950 ;
        RECT 679.950 373.950 682.050 376.050 ;
        RECT 673.950 364.950 676.050 367.050 ;
        RECT 674.400 343.050 675.450 364.950 ;
        RECT 673.950 338.100 676.050 343.050 ;
        RECT 691.950 338.100 694.050 340.200 ;
        RECT 692.400 337.350 693.600 338.100 ;
        RECT 667.950 328.950 670.050 331.050 ;
        RECT 673.950 328.950 676.050 334.050 ;
        RECT 668.400 295.050 669.450 328.950 ;
        RECT 667.950 292.950 670.050 295.050 ;
        RECT 643.950 283.950 646.050 286.050 ;
        RECT 644.400 220.050 645.450 283.950 ;
        RECT 625.950 217.950 628.050 220.050 ;
        RECT 643.950 217.950 646.050 220.050 ;
        RECT 626.400 210.450 627.450 217.950 ;
        RECT 626.400 209.400 630.450 210.450 ;
        RECT 400.950 154.950 403.050 157.050 ;
        RECT 541.950 154.950 544.050 157.050 ;
        RECT 392.400 132.000 393.600 133.650 ;
        RECT 391.950 127.950 394.050 132.000 ;
        RECT 401.400 130.050 402.450 154.950 ;
        RECT 542.400 139.200 543.450 154.950 ;
        RECT 541.950 137.100 544.050 139.200 ;
        RECT 542.400 136.350 543.600 137.100 ;
        RECT 604.950 136.950 607.050 139.050 ;
        RECT 605.400 130.050 606.450 136.950 ;
        RECT 629.400 130.050 630.450 209.400 ;
        RECT 755.400 209.400 756.600 211.650 ;
        RECT 755.400 190.050 756.450 209.400 ;
        RECT 754.950 187.950 757.050 190.050 ;
        RECT 769.950 187.950 772.050 190.050 ;
        RECT 770.400 142.050 771.450 187.950 ;
        RECT 703.950 139.950 706.050 142.050 ;
        RECT 769.950 139.950 772.050 142.050 ;
        RECT 668.400 131.400 669.600 133.650 ;
        RECT 400.950 127.950 403.050 130.050 ;
        RECT 604.950 127.950 607.050 130.050 ;
        RECT 628.950 127.950 631.050 130.050 ;
        RECT 668.400 127.050 669.450 131.400 ;
        RECT 704.400 127.050 705.450 139.950 ;
        RECT 808.950 138.000 811.050 142.050 ;
        RECT 809.400 136.350 810.600 138.000 ;
        RECT 667.950 124.950 670.050 127.050 ;
        RECT 697.950 124.950 700.050 127.050 ;
        RECT 703.950 124.950 706.050 127.050 ;
        RECT 698.400 96.450 699.450 124.950 ;
        RECT 695.400 95.400 699.450 96.450 ;
        RECT 695.400 37.050 696.450 95.400 ;
        RECT 685.950 34.950 688.050 37.050 ;
        RECT 694.950 34.950 697.050 37.050 ;
        RECT 686.400 4.050 687.450 34.950 ;
        RECT 667.950 1.950 670.050 4.050 ;
        RECT 685.950 1.950 688.050 4.050 ;
        RECT 668.400 -3.600 669.450 1.950 ;
      LAYER via2 ;
        RECT 808.950 139.950 811.050 142.050 ;
      LAYER metal3 ;
        RECT 472.950 807.750 475.050 808.200 ;
        RECT 490.950 807.750 493.050 808.200 ;
        RECT 472.950 806.550 493.050 807.750 ;
        RECT 472.950 806.100 475.050 806.550 ;
        RECT 490.950 806.100 493.050 806.550 ;
        RECT 469.950 756.600 472.050 757.050 ;
        RECT 484.950 756.600 487.050 756.900 ;
        RECT 469.950 756.450 487.050 756.600 ;
        RECT 499.950 756.450 502.050 756.900 ;
        RECT 469.950 755.400 502.050 756.450 ;
        RECT 469.950 754.950 472.050 755.400 ;
        RECT 484.950 755.250 502.050 755.400 ;
        RECT 484.950 754.800 487.050 755.250 ;
        RECT 499.950 754.800 502.050 755.250 ;
        RECT 499.950 750.600 502.050 751.050 ;
        RECT 619.950 750.600 622.050 751.050 ;
        RECT 499.950 749.400 622.050 750.600 ;
        RECT 499.950 748.950 502.050 749.400 ;
        RECT 619.950 748.950 622.050 749.400 ;
        RECT 619.950 738.600 622.050 739.050 ;
        RECT 640.950 738.600 643.050 739.050 ;
        RECT 619.950 737.400 723.600 738.600 ;
        RECT 619.950 736.950 622.050 737.400 ;
        RECT 640.950 736.950 643.050 737.400 ;
        RECT 722.400 736.050 723.600 737.400 ;
        RECT 722.400 734.400 727.050 736.050 ;
        RECT 723.000 733.950 727.050 734.400 ;
        RECT 595.950 666.600 598.050 667.050 ;
        RECT 646.950 666.600 649.050 667.050 ;
        RECT 595.950 665.400 649.050 666.600 ;
        RECT 595.950 664.950 598.050 665.400 ;
        RECT 646.950 664.950 649.050 665.400 ;
        RECT 595.950 571.950 598.050 574.050 ;
        RECT 596.400 568.050 597.600 571.950 ;
        RECT 595.950 565.950 598.050 568.050 ;
        RECT 586.950 546.600 589.050 547.050 ;
        RECT 595.950 546.600 598.050 547.050 ;
        RECT 586.950 545.400 598.050 546.600 ;
        RECT 586.950 544.950 589.050 545.400 ;
        RECT 595.950 544.950 598.050 545.400 ;
        RECT 574.950 528.750 577.050 529.200 ;
        RECT 580.950 528.750 583.050 529.200 ;
        RECT 574.950 528.600 583.050 528.750 ;
        RECT 586.950 528.600 589.050 529.050 ;
        RECT 574.950 527.550 589.050 528.600 ;
        RECT 574.950 527.100 577.050 527.550 ;
        RECT 580.950 527.400 589.050 527.550 ;
        RECT 580.950 527.100 583.050 527.400 ;
        RECT 586.950 526.950 589.050 527.400 ;
        RECT 571.950 483.600 574.050 484.050 ;
        RECT 610.950 483.600 613.050 484.050 ;
        RECT 571.950 482.400 613.050 483.600 ;
        RECT 571.950 481.950 574.050 482.400 ;
        RECT 610.950 481.950 613.050 482.400 ;
        RECT 676.950 462.600 679.050 463.050 ;
        RECT 688.950 462.600 691.050 463.050 ;
        RECT 676.950 461.400 691.050 462.600 ;
        RECT 676.950 460.950 679.050 461.400 ;
        RECT 688.950 460.950 691.050 461.400 ;
        RECT 610.950 453.600 615.000 454.050 ;
        RECT 610.950 451.950 615.600 453.600 ;
        RECT 614.400 447.600 615.600 451.950 ;
        RECT 614.400 446.400 621.600 447.600 ;
        RECT 620.400 441.600 621.600 446.400 ;
        RECT 628.950 441.600 631.050 442.050 ;
        RECT 620.400 440.400 631.050 441.600 ;
        RECT 628.950 439.950 631.050 440.400 ;
        RECT 628.950 423.600 631.050 424.050 ;
        RECT 628.950 422.400 690.600 423.600 ;
        RECT 628.950 421.950 631.050 422.400 ;
        RECT 689.400 421.050 690.600 422.400 ;
        RECT 688.950 418.950 691.050 421.050 ;
        RECT 689.400 414.600 690.600 418.950 ;
        RECT 680.400 414.000 690.600 414.600 ;
        RECT 679.950 413.400 690.600 414.000 ;
        RECT 679.950 409.950 682.050 413.400 ;
        RECT 673.950 339.750 676.050 340.200 ;
        RECT 691.950 339.750 694.050 340.200 ;
        RECT 673.950 338.550 694.050 339.750 ;
        RECT 673.950 338.100 676.050 338.550 ;
        RECT 691.950 338.100 694.050 338.550 ;
        RECT 667.950 330.600 670.050 331.050 ;
        RECT 673.950 330.600 676.050 331.050 ;
        RECT 667.950 329.400 676.050 330.600 ;
        RECT 667.950 328.950 670.050 329.400 ;
        RECT 673.950 328.950 676.050 329.400 ;
        RECT 667.950 292.950 670.050 295.050 ;
        RECT 643.950 285.600 646.050 286.050 ;
        RECT 668.400 285.600 669.600 292.950 ;
        RECT 643.950 284.400 669.600 285.600 ;
        RECT 643.950 283.950 646.050 284.400 ;
        RECT 625.950 219.600 628.050 220.050 ;
        RECT 643.950 219.600 646.050 220.050 ;
        RECT 625.950 218.400 646.050 219.600 ;
        RECT 625.950 217.950 628.050 218.400 ;
        RECT 643.950 217.950 646.050 218.400 ;
        RECT 754.950 189.600 757.050 190.050 ;
        RECT 769.950 189.600 772.050 190.050 ;
        RECT 754.950 188.400 772.050 189.600 ;
        RECT 754.950 187.950 757.050 188.400 ;
        RECT 769.950 187.950 772.050 188.400 ;
        RECT 400.950 156.600 403.050 157.050 ;
        RECT 541.950 156.600 544.050 157.050 ;
        RECT 400.950 155.400 544.050 156.600 ;
        RECT 400.950 154.950 403.050 155.400 ;
        RECT 541.950 154.950 544.050 155.400 ;
        RECT 703.950 141.600 706.050 142.050 ;
        RECT 769.950 141.600 772.050 142.050 ;
        RECT 808.950 141.600 811.050 142.050 ;
        RECT 703.950 140.400 811.050 141.600 ;
        RECT 703.950 139.950 706.050 140.400 ;
        RECT 769.950 139.950 772.050 140.400 ;
        RECT 808.950 139.950 811.050 140.400 ;
        RECT 541.950 138.600 544.050 139.200 ;
        RECT 604.950 138.600 607.050 139.050 ;
        RECT 541.950 137.400 607.050 138.600 ;
        RECT 541.950 137.100 544.050 137.400 ;
        RECT 604.950 136.950 607.050 137.400 ;
        RECT 604.950 129.600 607.050 130.050 ;
        RECT 628.950 129.600 631.050 130.050 ;
        RECT 604.950 128.400 636.600 129.600 ;
        RECT 604.950 127.950 607.050 128.400 ;
        RECT 628.950 127.950 631.050 128.400 ;
        RECT 635.400 126.600 636.600 128.400 ;
        RECT 667.950 126.600 670.050 127.050 ;
        RECT 697.950 126.600 700.050 127.050 ;
        RECT 703.950 126.600 706.050 127.050 ;
        RECT 635.400 125.400 706.050 126.600 ;
        RECT 667.950 124.950 670.050 125.400 ;
        RECT 697.950 124.950 700.050 125.400 ;
        RECT 703.950 124.950 706.050 125.400 ;
        RECT 667.950 3.600 670.050 4.050 ;
        RECT 685.950 3.600 688.050 4.050 ;
        RECT 667.950 2.400 688.050 3.600 ;
        RECT 667.950 1.950 670.050 2.400 ;
        RECT 685.950 1.950 688.050 2.400 ;
    END
  END Cin[3]
  PIN Cin[2]
    PORT
      LAYER metal1 ;
        RECT 541.950 729.450 546.000 730.050 ;
        RECT 541.950 727.950 546.450 729.450 ;
        RECT 545.550 723.450 546.450 727.950 ;
        RECT 550.950 723.450 553.050 724.050 ;
        RECT 545.550 722.550 553.050 723.450 ;
        RECT 550.950 721.950 553.050 722.550 ;
        RECT 694.950 696.450 697.050 697.050 ;
        RECT 703.950 696.450 706.050 697.050 ;
        RECT 694.950 695.550 706.050 696.450 ;
        RECT 694.950 694.950 697.050 695.550 ;
        RECT 703.950 694.950 706.050 695.550 ;
        RECT 607.950 420.450 610.050 421.050 ;
        RECT 616.950 420.450 619.050 421.050 ;
        RECT 607.950 419.550 619.050 420.450 ;
        RECT 607.950 418.950 610.050 419.550 ;
        RECT 616.950 418.950 619.050 419.550 ;
        RECT 700.950 297.450 703.050 298.050 ;
        RECT 700.950 296.550 714.450 297.450 ;
        RECT 700.950 295.950 703.050 296.550 ;
        RECT 713.550 289.050 714.450 296.550 ;
        RECT 713.550 287.550 718.050 289.050 ;
        RECT 714.000 286.950 718.050 287.550 ;
        RECT 376.950 129.450 379.050 130.050 ;
        RECT 385.950 129.450 388.050 130.050 ;
        RECT 376.950 128.550 388.050 129.450 ;
        RECT 376.950 127.950 379.050 128.550 ;
        RECT 385.950 127.950 388.050 128.550 ;
      LAYER via1 ;
        RECT 715.950 286.950 718.050 289.050 ;
      LAYER metal2 ;
        RECT 716.400 755.400 717.600 757.650 ;
        RECT 716.400 748.050 717.450 755.400 ;
        RECT 679.950 745.950 682.050 748.050 ;
        RECT 715.950 745.950 718.050 748.050 ;
        RECT 484.950 733.950 487.050 736.050 ;
        RECT 541.950 733.950 544.050 736.050 ;
        RECT 485.400 729.600 486.450 733.950 ;
        RECT 542.400 730.050 543.450 733.950 ;
        RECT 680.400 730.200 681.450 745.950 ;
        RECT 485.400 727.350 486.600 729.600 ;
        RECT 541.950 727.950 544.050 730.050 ;
        RECT 664.950 728.100 667.050 730.200 ;
        RECT 679.950 728.100 682.050 730.200 ;
        RECT 550.950 721.950 553.050 724.050 ;
        RECT 551.400 697.050 552.450 721.950 ;
        RECT 665.400 714.450 666.450 728.100 ;
        RECT 680.400 727.350 681.600 728.100 ;
        RECT 662.400 713.400 666.450 714.450 ;
        RECT 698.400 722.400 699.600 724.650 ;
        RECT 662.400 697.050 663.450 713.400 ;
        RECT 698.400 712.050 699.450 722.400 ;
        RECT 697.950 709.950 700.050 712.050 ;
        RECT 703.950 709.950 706.050 712.050 ;
        RECT 704.400 697.050 705.450 709.950 ;
        RECT 550.950 694.950 553.050 697.050 ;
        RECT 661.950 694.950 664.050 697.050 ;
        RECT 694.950 694.950 697.050 697.050 ;
        RECT 703.950 694.950 706.050 697.050 ;
        RECT 662.400 691.050 663.450 694.950 ;
        RECT 695.400 691.050 696.450 694.950 ;
        RECT 661.950 688.950 664.050 691.050 ;
        RECT 694.950 688.950 697.050 691.050 ;
        RECT 695.400 681.450 696.450 688.950 ;
        RECT 695.400 680.400 699.450 681.450 ;
        RECT 698.400 580.050 699.450 680.400 ;
        RECT 655.950 577.950 658.050 580.050 ;
        RECT 697.950 577.950 700.050 580.050 ;
        RECT 656.400 568.050 657.450 577.950 ;
        RECT 655.950 565.950 658.050 568.050 ;
        RECT 664.950 565.950 667.050 568.050 ;
        RECT 665.400 517.050 666.450 565.950 ;
        RECT 664.950 514.950 667.050 517.050 ;
        RECT 685.950 514.950 688.050 517.050 ;
        RECT 686.400 481.050 687.450 514.950 ;
        RECT 655.950 478.950 658.050 481.050 ;
        RECT 685.950 478.950 688.050 481.050 ;
        RECT 656.400 451.200 657.450 478.950 ;
        RECT 646.950 449.100 649.050 451.200 ;
        RECT 655.950 449.100 658.050 451.200 ;
        RECT 635.400 444.900 636.600 445.650 ;
        RECT 647.400 445.050 648.450 449.100 ;
        RECT 656.400 448.350 657.600 449.100 ;
        RECT 634.950 442.800 637.050 444.900 ;
        RECT 646.950 442.950 649.050 445.050 ;
        RECT 635.400 433.050 636.450 442.800 ;
        RECT 616.950 430.950 619.050 433.050 ;
        RECT 634.950 430.950 637.050 433.050 ;
        RECT 617.400 421.050 618.450 430.950 ;
        RECT 607.950 418.950 610.050 421.050 ;
        RECT 616.950 418.950 619.050 421.050 ;
        RECT 608.400 403.050 609.450 418.950 ;
        RECT 586.950 400.950 589.050 403.050 ;
        RECT 607.950 400.950 610.050 403.050 ;
        RECT 587.400 372.600 588.450 400.950 ;
        RECT 608.400 391.050 609.450 400.950 ;
        RECT 607.950 388.950 610.050 391.050 ;
        RECT 646.950 388.950 649.050 391.050 ;
        RECT 587.400 370.350 588.600 372.600 ;
        RECT 647.400 349.050 648.450 388.950 ;
        RECT 688.950 352.950 691.050 355.050 ;
        RECT 694.950 352.950 697.050 355.050 ;
        RECT 689.400 349.050 690.450 352.950 ;
        RECT 646.950 346.950 649.050 349.050 ;
        RECT 688.950 346.950 691.050 349.050 ;
        RECT 695.400 343.050 696.450 352.950 ;
        RECT 694.950 340.950 697.050 343.050 ;
        RECT 700.950 340.950 703.050 343.050 ;
        RECT 701.400 298.050 702.450 340.950 ;
        RECT 700.950 295.950 703.050 298.050 ;
        RECT 781.950 293.100 784.050 295.200 ;
        RECT 782.400 292.350 783.600 293.100 ;
        RECT 751.950 289.800 754.050 291.900 ;
        RECT 715.950 286.950 718.050 289.050 ;
        RECT 716.400 283.050 717.450 286.950 ;
        RECT 752.400 283.050 753.450 289.800 ;
        RECT 715.950 280.950 718.050 283.050 ;
        RECT 721.950 280.950 724.050 283.050 ;
        RECT 733.950 280.950 736.050 283.050 ;
        RECT 751.950 280.950 754.050 283.050 ;
        RECT 722.400 226.050 723.450 280.950 ;
        RECT 734.400 261.600 735.450 280.950 ;
        RECT 734.400 259.350 735.600 261.600 ;
        RECT 700.950 223.950 703.050 226.050 ;
        RECT 721.950 223.950 724.050 226.050 ;
        RECT 701.400 205.050 702.450 223.950 ;
        RECT 667.950 202.950 670.050 205.050 ;
        RECT 700.950 202.950 703.050 205.050 ;
        RECT 625.950 190.950 628.050 193.050 ;
        RECT 649.950 190.950 652.050 193.050 ;
        RECT 364.950 142.950 367.050 145.050 ;
        RECT 376.950 142.950 379.050 145.050 ;
        RECT 365.400 138.600 366.450 142.950 ;
        RECT 365.400 136.350 366.600 138.600 ;
        RECT 377.400 130.050 378.450 142.950 ;
        RECT 626.400 142.050 627.450 190.950 ;
        RECT 650.400 187.050 651.450 190.950 ;
        RECT 668.400 187.050 669.450 202.950 ;
        RECT 649.950 184.950 652.050 187.050 ;
        RECT 667.950 184.950 670.050 187.050 ;
        RECT 668.400 183.600 669.450 184.950 ;
        RECT 668.400 181.350 669.600 183.600 ;
        RECT 625.950 139.950 628.050 142.050 ;
        RECT 386.400 132.000 387.600 133.650 ;
        RECT 376.950 127.950 379.050 130.050 ;
        RECT 385.950 129.450 388.050 132.000 ;
        RECT 385.950 129.000 390.450 129.450 ;
        RECT 385.950 128.400 391.050 129.000 ;
        RECT 385.950 127.950 388.050 128.400 ;
        RECT 388.950 124.950 391.050 128.400 ;
        RECT 394.950 124.950 397.050 127.050 ;
        RECT 395.400 73.050 396.450 124.950 ;
        RECT 370.950 70.950 373.050 73.050 ;
        RECT 394.950 70.950 397.050 73.050 ;
        RECT 371.400 60.450 372.450 70.950 ;
        RECT 371.400 59.400 375.450 60.450 ;
        RECT 374.400 31.050 375.450 59.400 ;
        RECT 373.950 28.950 376.050 31.050 ;
        RECT 382.950 28.950 385.050 31.050 ;
        RECT 383.400 -3.600 384.450 28.950 ;
      LAYER metal3 ;
        RECT 679.950 747.600 682.050 748.050 ;
        RECT 715.950 747.600 718.050 748.050 ;
        RECT 679.950 746.400 718.050 747.600 ;
        RECT 679.950 745.950 682.050 746.400 ;
        RECT 715.950 745.950 718.050 746.400 ;
        RECT 484.950 735.600 487.050 736.050 ;
        RECT 541.950 735.600 544.050 736.050 ;
        RECT 484.950 734.400 544.050 735.600 ;
        RECT 484.950 733.950 487.050 734.400 ;
        RECT 541.950 733.950 544.050 734.400 ;
        RECT 664.950 729.750 667.050 730.200 ;
        RECT 679.950 729.750 682.050 730.200 ;
        RECT 664.950 728.550 682.050 729.750 ;
        RECT 664.950 728.100 667.050 728.550 ;
        RECT 679.950 728.100 682.050 728.550 ;
        RECT 697.950 711.600 700.050 712.050 ;
        RECT 703.950 711.600 706.050 712.050 ;
        RECT 697.950 710.400 706.050 711.600 ;
        RECT 697.950 709.950 700.050 710.400 ;
        RECT 703.950 709.950 706.050 710.400 ;
        RECT 550.950 696.600 553.050 697.050 ;
        RECT 661.950 696.600 664.050 697.050 ;
        RECT 550.950 695.400 664.050 696.600 ;
        RECT 550.950 694.950 553.050 695.400 ;
        RECT 661.950 694.950 664.050 695.400 ;
        RECT 661.950 690.600 664.050 691.050 ;
        RECT 694.950 690.600 697.050 691.050 ;
        RECT 661.950 689.400 697.050 690.600 ;
        RECT 661.950 688.950 664.050 689.400 ;
        RECT 694.950 688.950 697.050 689.400 ;
        RECT 655.950 579.600 658.050 580.050 ;
        RECT 697.950 579.600 700.050 580.050 ;
        RECT 655.950 578.400 700.050 579.600 ;
        RECT 655.950 577.950 658.050 578.400 ;
        RECT 697.950 577.950 700.050 578.400 ;
        RECT 655.950 567.600 658.050 568.050 ;
        RECT 664.950 567.600 667.050 568.050 ;
        RECT 655.950 566.400 667.050 567.600 ;
        RECT 655.950 565.950 658.050 566.400 ;
        RECT 664.950 565.950 667.050 566.400 ;
        RECT 664.950 516.600 667.050 517.050 ;
        RECT 685.950 516.600 688.050 517.050 ;
        RECT 664.950 515.400 688.050 516.600 ;
        RECT 664.950 514.950 667.050 515.400 ;
        RECT 685.950 514.950 688.050 515.400 ;
        RECT 655.950 480.600 658.050 481.050 ;
        RECT 685.950 480.600 688.050 481.050 ;
        RECT 655.950 479.400 688.050 480.600 ;
        RECT 655.950 478.950 658.050 479.400 ;
        RECT 685.950 478.950 688.050 479.400 ;
        RECT 646.950 450.750 649.050 451.200 ;
        RECT 655.950 450.750 658.050 451.200 ;
        RECT 646.950 449.550 658.050 450.750 ;
        RECT 646.950 449.100 649.050 449.550 ;
        RECT 655.950 449.100 658.050 449.550 ;
        RECT 634.950 444.600 637.050 444.900 ;
        RECT 646.950 444.600 649.050 445.050 ;
        RECT 634.950 443.400 649.050 444.600 ;
        RECT 634.950 442.800 637.050 443.400 ;
        RECT 646.950 442.950 649.050 443.400 ;
        RECT 616.950 432.600 619.050 433.050 ;
        RECT 634.950 432.600 637.050 433.050 ;
        RECT 616.950 431.400 637.050 432.600 ;
        RECT 616.950 430.950 619.050 431.400 ;
        RECT 634.950 430.950 637.050 431.400 ;
        RECT 586.950 402.600 589.050 403.050 ;
        RECT 607.950 402.600 610.050 403.050 ;
        RECT 586.950 401.400 610.050 402.600 ;
        RECT 586.950 400.950 589.050 401.400 ;
        RECT 607.950 400.950 610.050 401.400 ;
        RECT 607.950 390.600 610.050 391.050 ;
        RECT 646.950 390.600 649.050 391.050 ;
        RECT 607.950 389.400 649.050 390.600 ;
        RECT 607.950 388.950 610.050 389.400 ;
        RECT 646.950 388.950 649.050 389.400 ;
        RECT 688.950 354.600 691.050 355.050 ;
        RECT 694.950 354.600 697.050 355.050 ;
        RECT 688.950 353.400 697.050 354.600 ;
        RECT 688.950 352.950 691.050 353.400 ;
        RECT 694.950 352.950 697.050 353.400 ;
        RECT 646.950 348.600 649.050 349.050 ;
        RECT 688.950 348.600 691.050 349.050 ;
        RECT 646.950 347.400 691.050 348.600 ;
        RECT 646.950 346.950 649.050 347.400 ;
        RECT 688.950 346.950 691.050 347.400 ;
        RECT 694.950 342.600 697.050 343.050 ;
        RECT 700.950 342.600 703.050 343.050 ;
        RECT 694.950 341.400 703.050 342.600 ;
        RECT 694.950 340.950 697.050 341.400 ;
        RECT 700.950 340.950 703.050 341.400 ;
        RECT 781.950 293.100 784.050 295.200 ;
        RECT 751.950 291.600 754.050 291.900 ;
        RECT 782.400 291.600 783.600 293.100 ;
        RECT 751.950 290.400 783.600 291.600 ;
        RECT 751.950 289.800 754.050 290.400 ;
        RECT 715.950 282.600 718.050 283.050 ;
        RECT 721.950 282.600 724.050 283.050 ;
        RECT 733.950 282.600 736.050 283.050 ;
        RECT 751.950 282.600 754.050 283.050 ;
        RECT 715.950 281.400 754.050 282.600 ;
        RECT 715.950 280.950 718.050 281.400 ;
        RECT 721.950 280.950 724.050 281.400 ;
        RECT 733.950 280.950 736.050 281.400 ;
        RECT 751.950 280.950 754.050 281.400 ;
        RECT 700.950 225.600 703.050 226.050 ;
        RECT 721.950 225.600 724.050 226.050 ;
        RECT 700.950 224.400 724.050 225.600 ;
        RECT 700.950 223.950 703.050 224.400 ;
        RECT 721.950 223.950 724.050 224.400 ;
        RECT 667.950 204.600 670.050 205.050 ;
        RECT 700.950 204.600 703.050 205.050 ;
        RECT 667.950 203.400 703.050 204.600 ;
        RECT 667.950 202.950 670.050 203.400 ;
        RECT 700.950 202.950 703.050 203.400 ;
        RECT 625.950 192.600 628.050 193.050 ;
        RECT 649.950 192.600 652.050 193.050 ;
        RECT 625.950 191.400 652.050 192.600 ;
        RECT 625.950 190.950 628.050 191.400 ;
        RECT 649.950 190.950 652.050 191.400 ;
        RECT 649.950 186.600 652.050 187.050 ;
        RECT 667.950 186.600 670.050 187.050 ;
        RECT 649.950 185.400 670.050 186.600 ;
        RECT 649.950 184.950 652.050 185.400 ;
        RECT 667.950 184.950 670.050 185.400 ;
        RECT 364.950 144.600 367.050 145.050 ;
        RECT 376.950 144.600 379.050 145.050 ;
        RECT 364.950 143.400 417.600 144.600 ;
        RECT 364.950 142.950 367.050 143.400 ;
        RECT 376.950 142.950 379.050 143.400 ;
        RECT 416.400 141.600 417.600 143.400 ;
        RECT 625.950 141.600 628.050 142.050 ;
        RECT 416.400 140.400 628.050 141.600 ;
        RECT 625.950 139.950 628.050 140.400 ;
        RECT 388.950 126.600 391.050 127.050 ;
        RECT 394.950 126.600 397.050 127.050 ;
        RECT 388.950 125.400 397.050 126.600 ;
        RECT 388.950 124.950 391.050 125.400 ;
        RECT 394.950 124.950 397.050 125.400 ;
        RECT 370.950 72.600 373.050 73.050 ;
        RECT 394.950 72.600 397.050 73.050 ;
        RECT 370.950 71.400 397.050 72.600 ;
        RECT 370.950 70.950 373.050 71.400 ;
        RECT 394.950 70.950 397.050 71.400 ;
        RECT 373.950 30.600 376.050 31.050 ;
        RECT 382.950 30.600 385.050 31.050 ;
        RECT 373.950 29.400 385.050 30.600 ;
        RECT 373.950 28.950 376.050 29.400 ;
        RECT 382.950 28.950 385.050 29.400 ;
    END
  END Cin[2]
  PIN Cin[1]
    PORT
      LAYER metal1 ;
        RECT 553.950 654.450 556.050 655.050 ;
        RECT 562.950 654.450 565.050 655.050 ;
        RECT 553.950 653.550 565.050 654.450 ;
        RECT 553.950 652.950 556.050 653.550 ;
        RECT 562.950 652.950 565.050 653.550 ;
        RECT 532.950 561.450 535.050 562.050 ;
        RECT 544.950 561.450 547.050 561.900 ;
        RECT 532.950 560.550 547.050 561.450 ;
        RECT 532.950 559.950 535.050 560.550 ;
        RECT 544.950 559.800 547.050 560.550 ;
      LAYER metal2 ;
        RECT 553.950 652.950 556.050 655.050 ;
        RECT 487.950 650.100 490.050 652.200 ;
        RECT 499.950 650.100 502.050 652.200 ;
        RECT 488.400 649.350 489.600 650.100 ;
        RECT 500.400 625.050 501.450 650.100 ;
        RECT 554.400 640.050 555.450 652.950 ;
        RECT 562.950 651.000 565.050 655.050 ;
        RECT 563.400 649.350 564.600 651.000 ;
        RECT 532.950 637.950 535.050 640.050 ;
        RECT 553.950 637.950 556.050 640.050 ;
        RECT 589.950 637.950 592.050 640.050 ;
        RECT 533.400 625.050 534.450 637.950 ;
        RECT 590.400 628.050 591.450 637.950 ;
        RECT 589.950 625.950 592.050 628.050 ;
        RECT 706.950 625.950 709.050 628.050 ;
        RECT 499.950 622.950 502.050 625.050 ;
        RECT 532.950 622.950 535.050 625.050 ;
        RECT 533.400 562.050 534.450 622.950 ;
        RECT 707.400 606.600 708.450 625.950 ;
        RECT 707.400 604.350 708.600 606.600 ;
        RECT 532.950 559.950 535.050 562.050 ;
        RECT 544.950 559.800 547.050 561.900 ;
        RECT 545.400 517.050 546.450 559.800 ;
        RECT 532.950 514.950 535.050 517.050 ;
        RECT 544.950 514.950 547.050 517.050 ;
        RECT 533.400 364.050 534.450 514.950 ;
        RECT 532.950 361.950 535.050 364.050 ;
        RECT 547.800 361.950 549.900 364.050 ;
        RECT 548.400 235.050 549.450 361.950 ;
        RECT 635.400 254.400 636.600 256.650 ;
        RECT 635.400 235.050 636.450 254.400 ;
        RECT 547.950 232.950 550.050 235.050 ;
        RECT 634.950 232.950 637.050 235.050 ;
        RECT 235.950 229.950 238.050 232.050 ;
        RECT 502.950 229.950 505.050 232.050 ;
        RECT 79.950 223.950 82.050 226.050 ;
        RECT 181.950 223.950 184.050 226.050 ;
        RECT 80.400 220.050 81.450 223.950 ;
        RECT 31.950 217.950 34.050 220.050 ;
        RECT 79.950 217.950 82.050 220.050 ;
        RECT 14.400 177.900 15.600 178.650 ;
        RECT 32.400 177.900 33.450 217.950 ;
        RECT 182.400 217.200 183.450 223.950 ;
        RECT 181.950 215.100 184.050 217.200 ;
        RECT 223.950 215.100 226.050 217.200 ;
        RECT 236.400 217.050 237.450 229.950 ;
        RECT 182.400 214.350 183.600 215.100 ;
        RECT 224.400 214.350 225.600 215.100 ;
        RECT 235.950 214.950 238.050 217.050 ;
        RECT 503.400 216.600 504.450 229.950 ;
        RECT 236.400 193.050 237.450 214.950 ;
        RECT 503.400 214.350 504.600 216.600 ;
        RECT 235.950 190.950 238.050 193.050 ;
        RECT 250.800 190.950 252.900 193.050 ;
        RECT 248.400 183.450 249.600 183.600 ;
        RECT 251.400 183.450 252.450 190.950 ;
        RECT 248.400 182.400 252.450 183.450 ;
        RECT 248.400 181.350 249.600 182.400 ;
        RECT 38.400 177.900 39.600 178.650 ;
        RECT 13.950 175.800 16.050 177.900 ;
        RECT 31.950 175.800 34.050 177.900 ;
        RECT 37.950 175.800 40.050 177.900 ;
      LAYER metal3 ;
        RECT 487.950 651.750 490.050 652.200 ;
        RECT 499.950 651.750 502.050 652.200 ;
        RECT 487.950 650.550 502.050 651.750 ;
        RECT 487.950 650.100 490.050 650.550 ;
        RECT 499.950 650.100 502.050 650.550 ;
        RECT 532.950 639.600 535.050 640.050 ;
        RECT 553.950 639.600 556.050 640.050 ;
        RECT 589.950 639.600 592.050 640.050 ;
        RECT 532.950 638.400 592.050 639.600 ;
        RECT 532.950 637.950 535.050 638.400 ;
        RECT 553.950 637.950 556.050 638.400 ;
        RECT 589.950 637.950 592.050 638.400 ;
        RECT 589.950 627.600 592.050 628.050 ;
        RECT 706.950 627.600 709.050 628.050 ;
        RECT 589.950 626.400 709.050 627.600 ;
        RECT 589.950 625.950 592.050 626.400 ;
        RECT 706.950 625.950 709.050 626.400 ;
        RECT 499.950 624.600 502.050 625.050 ;
        RECT 532.950 624.600 535.050 625.050 ;
        RECT 499.950 623.400 535.050 624.600 ;
        RECT 499.950 622.950 502.050 623.400 ;
        RECT 532.950 622.950 535.050 623.400 ;
        RECT 532.950 516.600 535.050 517.050 ;
        RECT 544.950 516.600 547.050 517.050 ;
        RECT 532.950 515.400 547.050 516.600 ;
        RECT 532.950 514.950 535.050 515.400 ;
        RECT 544.950 514.950 547.050 515.400 ;
        RECT 532.950 363.600 535.050 364.050 ;
        RECT 547.800 363.600 549.900 364.050 ;
        RECT 532.950 362.400 549.900 363.600 ;
        RECT 532.950 361.950 535.050 362.400 ;
        RECT 547.800 361.950 549.900 362.400 ;
        RECT 547.950 234.600 550.050 235.050 ;
        RECT 634.950 234.600 637.050 235.050 ;
        RECT 503.400 233.400 637.050 234.600 ;
        RECT 503.400 232.050 504.600 233.400 ;
        RECT 547.950 232.950 550.050 233.400 ;
        RECT 634.950 232.950 637.050 233.400 ;
        RECT 235.950 231.600 238.050 232.050 ;
        RECT 502.950 231.600 505.050 232.050 ;
        RECT 235.950 230.400 505.050 231.600 ;
        RECT 235.950 229.950 238.050 230.400 ;
        RECT 502.950 229.950 505.050 230.400 ;
        RECT 79.950 225.600 82.050 226.050 ;
        RECT 181.950 225.600 184.050 226.050 ;
        RECT 79.950 224.400 184.050 225.600 ;
        RECT 79.950 223.950 82.050 224.400 ;
        RECT 181.950 223.950 184.050 224.400 ;
        RECT 31.950 219.600 34.050 220.050 ;
        RECT 79.950 219.600 82.050 220.050 ;
        RECT 31.950 218.400 82.050 219.600 ;
        RECT 31.950 217.950 34.050 218.400 ;
        RECT 79.950 217.950 82.050 218.400 ;
        RECT 181.950 216.600 184.050 217.200 ;
        RECT 223.950 216.600 226.050 217.200 ;
        RECT 235.950 216.600 238.050 217.050 ;
        RECT 181.950 215.400 238.050 216.600 ;
        RECT 181.950 215.100 184.050 215.400 ;
        RECT 223.950 215.100 226.050 215.400 ;
        RECT 235.950 214.950 238.050 215.400 ;
        RECT 235.950 192.600 238.050 193.050 ;
        RECT 250.800 192.600 252.900 193.050 ;
        RECT 235.950 191.400 252.900 192.600 ;
        RECT 235.950 190.950 238.050 191.400 ;
        RECT 250.800 190.950 252.900 191.400 ;
        RECT 13.950 177.600 16.050 177.900 ;
        RECT 31.950 177.600 34.050 177.900 ;
        RECT -3.600 177.450 34.050 177.600 ;
        RECT 37.950 177.450 40.050 177.900 ;
        RECT -3.600 176.400 40.050 177.450 ;
        RECT 13.950 175.800 16.050 176.400 ;
        RECT 31.950 176.250 40.050 176.400 ;
        RECT 31.950 175.800 34.050 176.250 ;
        RECT 37.950 175.800 40.050 176.250 ;
    END
  END Cin[1]
  PIN Cin[0]
    PORT
      LAYER metal2 ;
        RECT 154.950 379.950 157.050 382.050 ;
        RECT 376.950 379.950 379.050 382.050 ;
        RECT 155.400 301.050 156.450 379.950 ;
        RECT 377.400 343.050 378.450 379.950 ;
        RECT 545.400 365.400 546.600 367.650 ;
        RECT 391.950 346.950 394.050 349.050 ;
        RECT 463.950 346.950 466.050 349.050 ;
        RECT 392.400 343.050 393.450 346.950 ;
        RECT 376.950 340.950 379.050 343.050 ;
        RECT 391.950 340.950 394.050 343.050 ;
        RECT 464.400 340.050 465.450 346.950 ;
        RECT 545.400 343.050 546.450 365.400 ;
        RECT 463.950 337.950 466.050 340.050 ;
        RECT 538.950 338.100 541.050 343.050 ;
        RECT 544.950 340.950 547.050 343.050 ;
        RECT 539.400 337.350 540.600 338.100 ;
        RECT 94.950 298.950 97.050 301.050 ;
        RECT 154.950 298.950 157.050 301.050 ;
        RECT 95.400 288.450 96.450 298.950 ;
        RECT 98.400 288.450 99.600 289.650 ;
        RECT 95.400 287.400 99.600 288.450 ;
        RECT 95.400 277.050 96.450 287.400 ;
        RECT 1.950 274.950 4.050 277.050 ;
        RECT 94.950 274.950 97.050 277.050 ;
        RECT 2.400 217.050 3.450 274.950 ;
        RECT 1.950 214.950 4.050 217.050 ;
        RECT 2.400 210.900 3.450 214.950 ;
        RECT 14.400 210.900 15.600 211.650 ;
        RECT 1.950 208.800 4.050 210.900 ;
        RECT 13.950 208.800 16.050 210.900 ;
      LAYER via2 ;
        RECT 538.950 340.950 541.050 343.050 ;
      LAYER metal3 ;
        RECT 154.950 381.600 157.050 382.050 ;
        RECT 376.950 381.600 379.050 382.050 ;
        RECT 154.950 380.400 379.050 381.600 ;
        RECT 154.950 379.950 157.050 380.400 ;
        RECT 376.950 379.950 379.050 380.400 ;
        RECT 391.950 348.600 394.050 349.050 ;
        RECT 463.950 348.600 466.050 349.050 ;
        RECT 391.950 347.400 466.050 348.600 ;
        RECT 391.950 346.950 394.050 347.400 ;
        RECT 463.950 346.950 466.050 347.400 ;
        RECT 376.950 342.600 379.050 343.050 ;
        RECT 391.950 342.600 394.050 343.050 ;
        RECT 376.950 341.400 394.050 342.600 ;
        RECT 376.950 340.950 379.050 341.400 ;
        RECT 391.950 340.950 394.050 341.400 ;
        RECT 538.950 342.600 541.050 343.050 ;
        RECT 544.950 342.600 547.050 343.050 ;
        RECT 538.950 341.400 547.050 342.600 ;
        RECT 538.950 340.950 541.050 341.400 ;
        RECT 544.950 340.950 547.050 341.400 ;
        RECT 463.950 339.600 466.050 340.050 ;
        RECT 538.950 339.600 541.050 340.200 ;
        RECT 463.950 338.400 541.050 339.600 ;
        RECT 463.950 337.950 466.050 338.400 ;
        RECT 538.950 338.100 541.050 338.400 ;
        RECT 94.950 300.600 97.050 301.050 ;
        RECT 154.950 300.600 157.050 301.050 ;
        RECT 94.950 299.400 157.050 300.600 ;
        RECT 94.950 298.950 97.050 299.400 ;
        RECT 154.950 298.950 157.050 299.400 ;
        RECT 1.950 276.600 4.050 277.050 ;
        RECT 94.950 276.600 97.050 277.050 ;
        RECT 1.950 275.400 97.050 276.600 ;
        RECT 1.950 274.950 4.050 275.400 ;
        RECT 94.950 274.950 97.050 275.400 ;
        RECT 1.950 216.600 4.050 217.050 ;
        RECT -3.600 215.400 4.050 216.600 ;
        RECT 1.950 214.950 4.050 215.400 ;
        RECT 1.950 210.450 4.050 210.900 ;
        RECT 13.950 210.450 16.050 210.900 ;
        RECT 1.950 209.250 16.050 210.450 ;
        RECT 1.950 208.800 4.050 209.250 ;
        RECT 13.950 208.800 16.050 209.250 ;
    END
  END Cin[0]
  PIN Rdy
    PORT
      LAYER metal2 ;
        RECT 14.400 411.900 15.600 412.650 ;
        RECT 13.950 409.800 16.050 411.900 ;
      LAYER metal3 ;
        RECT 13.950 411.600 16.050 411.900 ;
        RECT -3.600 410.400 16.050 411.600 ;
        RECT 13.950 409.800 16.050 410.400 ;
    END
  END Rdy
  PIN Vld
    PORT
      LAYER metal2 ;
        RECT 413.400 20.400 414.600 22.650 ;
        RECT 413.400 -2.550 414.450 20.400 ;
        RECT 413.400 -3.600 417.450 -2.550 ;
    END
  END Vld
  PIN Xin[3]
    PORT
      LAYER metal2 ;
        RECT 200.400 410.400 201.600 412.650 ;
        RECT 200.400 388.050 201.450 410.400 ;
        RECT 7.950 385.950 10.050 388.050 ;
        RECT 58.950 385.950 61.050 388.050 ;
        RECT 199.950 385.950 202.050 388.050 ;
        RECT 8.400 379.050 9.450 385.950 ;
        RECT 7.950 376.950 10.050 379.050 ;
        RECT 59.400 372.600 60.450 385.950 ;
        RECT 59.400 370.350 60.600 372.600 ;
      LAYER metal3 ;
        RECT 7.950 387.600 10.050 388.050 ;
        RECT 58.950 387.600 61.050 388.050 ;
        RECT 199.950 387.600 202.050 388.050 ;
        RECT 7.950 386.400 202.050 387.600 ;
        RECT 7.950 385.950 10.050 386.400 ;
        RECT 58.950 385.950 61.050 386.400 ;
        RECT 199.950 385.950 202.050 386.400 ;
        RECT 7.950 378.600 10.050 379.050 ;
        RECT -3.600 377.400 10.050 378.600 ;
        RECT -3.600 371.400 -2.400 377.400 ;
        RECT 7.950 376.950 10.050 377.400 ;
    END
  END Xin[3]
  PIN Xin[2]
    PORT
      LAYER metal2 ;
        RECT 455.400 254.400 456.600 256.650 ;
        RECT 455.400 241.050 456.450 254.400 ;
        RECT 454.950 238.950 457.050 241.050 ;
        RECT 463.950 238.950 466.050 241.050 ;
        RECT 449.400 176.400 450.600 178.650 ;
        RECT 449.400 172.050 450.450 176.400 ;
        RECT 464.400 172.050 465.450 238.950 ;
        RECT 448.950 171.450 451.050 172.050 ;
        RECT 448.950 170.400 453.450 171.450 ;
        RECT 448.950 169.950 451.050 170.400 ;
        RECT 452.400 27.450 453.450 170.400 ;
        RECT 463.950 169.950 466.050 172.050 ;
        RECT 449.400 26.400 453.450 27.450 ;
        RECT 449.400 -2.550 450.450 26.400 ;
        RECT 449.400 -3.600 453.450 -2.550 ;
      LAYER metal3 ;
        RECT 454.950 240.600 457.050 241.050 ;
        RECT 463.950 240.600 466.050 241.050 ;
        RECT 454.950 239.400 466.050 240.600 ;
        RECT 454.950 238.950 457.050 239.400 ;
        RECT 463.950 238.950 466.050 239.400 ;
        RECT 448.950 171.600 451.050 172.050 ;
        RECT 463.950 171.600 466.050 172.050 ;
        RECT 448.950 170.400 466.050 171.600 ;
        RECT 448.950 169.950 451.050 170.400 ;
        RECT 463.950 169.950 466.050 170.400 ;
    END
  END Xin[2]
  PIN Xin[1]
    PORT
      LAYER metal1 ;
        RECT 319.950 105.450 322.050 106.050 ;
        RECT 325.950 105.450 328.050 106.050 ;
        RECT 319.950 104.550 328.050 105.450 ;
        RECT 319.950 103.950 322.050 104.550 ;
        RECT 325.950 103.950 328.050 104.550 ;
      LAYER metal2 ;
        RECT 401.400 254.400 402.600 256.650 ;
        RECT 401.400 241.050 402.450 254.400 ;
        RECT 400.950 238.950 403.050 241.050 ;
        RECT 325.950 235.950 328.050 238.050 ;
        RECT 293.400 176.400 294.600 178.650 ;
        RECT 293.400 172.050 294.450 176.400 ;
        RECT 326.400 172.050 327.450 235.950 ;
        RECT 292.950 169.950 295.050 172.050 ;
        RECT 325.950 169.950 328.050 172.050 ;
        RECT 326.400 106.050 327.450 169.950 ;
        RECT 319.950 103.950 322.050 106.050 ;
        RECT 325.950 103.950 328.050 106.050 ;
        RECT 320.400 34.050 321.450 103.950 ;
        RECT 307.950 31.950 310.050 34.050 ;
        RECT 319.950 31.950 322.050 34.050 ;
        RECT 308.400 4.050 309.450 31.950 ;
        RECT 289.950 1.950 292.050 4.050 ;
        RECT 307.950 1.950 310.050 4.050 ;
        RECT 290.400 -3.600 291.450 1.950 ;
      LAYER metal3 ;
        RECT 400.950 240.600 403.050 241.050 ;
        RECT 347.400 239.400 403.050 240.600 ;
        RECT 325.950 237.600 328.050 238.050 ;
        RECT 347.400 237.600 348.600 239.400 ;
        RECT 400.950 238.950 403.050 239.400 ;
        RECT 325.950 236.400 348.600 237.600 ;
        RECT 325.950 235.950 328.050 236.400 ;
        RECT 292.950 171.600 295.050 172.050 ;
        RECT 325.950 171.600 328.050 172.050 ;
        RECT 292.950 170.400 328.050 171.600 ;
        RECT 292.950 169.950 295.050 170.400 ;
        RECT 325.950 169.950 328.050 170.400 ;
        RECT 307.950 33.600 310.050 34.050 ;
        RECT 319.950 33.600 322.050 34.050 ;
        RECT 307.950 32.400 322.050 33.600 ;
        RECT 307.950 31.950 310.050 32.400 ;
        RECT 319.950 31.950 322.050 32.400 ;
        RECT 289.950 3.600 292.050 4.050 ;
        RECT 307.950 3.600 310.050 4.050 ;
        RECT 289.950 2.400 310.050 3.600 ;
        RECT 289.950 1.950 292.050 2.400 ;
        RECT 307.950 1.950 310.050 2.400 ;
    END
  END Xin[1]
  PIN Xin[0]
    PORT
      LAYER metal2 ;
        RECT 185.400 332.400 186.600 334.650 ;
        RECT 185.400 313.050 186.450 332.400 ;
        RECT 184.950 310.950 187.050 313.050 ;
        RECT 10.950 307.950 13.050 310.050 ;
        RECT 11.400 295.050 12.450 307.950 ;
        RECT 185.400 295.200 186.450 310.950 ;
        RECT 10.950 292.950 13.050 295.050 ;
        RECT 169.950 293.100 172.050 295.200 ;
        RECT 184.950 293.100 187.050 295.200 ;
        RECT 170.400 292.350 171.600 293.100 ;
      LAYER metal3 ;
        RECT 184.950 312.600 187.050 313.050 ;
        RECT 29.400 311.400 187.050 312.600 ;
        RECT 10.950 309.600 13.050 310.050 ;
        RECT 29.400 309.600 30.600 311.400 ;
        RECT 184.950 310.950 187.050 311.400 ;
        RECT 10.950 308.400 30.600 309.600 ;
        RECT 10.950 307.950 13.050 308.400 ;
        RECT 10.950 294.600 13.050 295.050 ;
        RECT -3.600 293.400 13.050 294.600 ;
        RECT 10.950 292.950 13.050 293.400 ;
        RECT 169.950 294.750 172.050 295.200 ;
        RECT 184.950 294.750 187.050 295.200 ;
        RECT 169.950 293.550 187.050 294.750 ;
        RECT 169.950 293.100 172.050 293.550 ;
        RECT 184.950 293.100 187.050 293.550 ;
    END
  END Xin[0]
  PIN Xout[3]
    PORT
      LAYER metal2 ;
        RECT 13.950 527.100 16.050 529.200 ;
        RECT 14.400 526.350 15.600 527.100 ;
      LAYER metal3 ;
        RECT 13.950 528.600 16.050 529.200 ;
        RECT -3.600 527.400 16.050 528.600 ;
        RECT 13.950 527.100 16.050 527.400 ;
    END
  END Xout[3]
  PIN Xout[2]
    PORT
      LAYER metal2 ;
        RECT 16.950 450.000 19.050 454.050 ;
        RECT 17.400 448.350 18.600 450.000 ;
      LAYER via2 ;
        RECT 16.950 451.950 19.050 454.050 ;
      LAYER metal3 ;
        RECT -3.600 453.600 -2.400 456.600 ;
        RECT 16.950 453.600 19.050 454.050 ;
        RECT -3.600 452.400 19.050 453.600 ;
        RECT 16.950 451.950 19.050 452.400 ;
    END
  END Xout[2]
  PIN Xout[1]
    PORT
      LAYER metal2 ;
        RECT 374.400 20.400 375.600 22.650 ;
        RECT 374.400 -2.550 375.450 20.400 ;
        RECT 371.400 -3.600 375.450 -2.550 ;
    END
  END Xout[1]
  PIN Xout[0]
    PORT
      LAYER metal2 ;
        RECT 14.400 255.900 15.600 256.650 ;
        RECT 13.950 253.800 16.050 255.900 ;
      LAYER metal3 ;
        RECT 13.950 255.600 16.050 255.900 ;
        RECT -3.600 254.400 16.050 255.600 ;
        RECT 13.950 253.800 16.050 254.400 ;
    END
  END Xout[0]
  PIN Yin[3]
    PORT
      LAYER metal2 ;
        RECT 17.400 566.400 18.600 568.650 ;
        RECT 17.400 559.050 18.450 566.400 ;
        RECT 16.950 556.950 19.050 559.050 ;
        RECT 22.950 556.950 25.050 559.050 ;
        RECT 23.400 520.050 24.450 556.950 ;
        RECT 35.400 522.000 36.600 523.650 ;
        RECT 22.950 519.450 25.050 520.050 ;
        RECT 22.950 518.400 27.450 519.450 ;
        RECT 22.950 517.950 25.050 518.400 ;
        RECT 26.400 429.450 27.450 518.400 ;
        RECT 34.950 517.950 37.050 522.000 ;
        RECT 23.400 428.400 27.450 429.450 ;
        RECT 23.400 373.050 24.450 428.400 ;
        RECT 7.950 370.950 10.050 373.050 ;
        RECT 22.950 370.950 25.050 373.050 ;
        RECT 8.400 301.050 9.450 370.950 ;
        RECT 7.950 298.950 10.050 301.050 ;
        RECT 13.950 298.950 16.050 301.050 ;
        RECT 14.400 294.600 15.450 298.950 ;
        RECT 14.400 292.350 15.600 294.600 ;
      LAYER metal3 ;
        RECT 16.950 558.600 19.050 559.050 ;
        RECT 22.950 558.600 25.050 559.050 ;
        RECT 16.950 557.400 25.050 558.600 ;
        RECT 16.950 556.950 19.050 557.400 ;
        RECT 22.950 556.950 25.050 557.400 ;
        RECT 22.950 519.600 25.050 520.050 ;
        RECT 34.950 519.600 37.050 520.050 ;
        RECT 22.950 518.400 37.050 519.600 ;
        RECT 22.950 517.950 25.050 518.400 ;
        RECT 34.950 517.950 37.050 518.400 ;
        RECT 7.950 372.600 10.050 373.050 ;
        RECT 22.950 372.600 25.050 373.050 ;
        RECT 7.950 371.400 25.050 372.600 ;
        RECT 7.950 370.950 10.050 371.400 ;
        RECT 22.950 370.950 25.050 371.400 ;
        RECT 7.950 300.600 10.050 301.050 ;
        RECT 13.950 300.600 16.050 301.050 ;
        RECT -3.600 299.400 16.050 300.600 ;
        RECT 7.950 298.950 10.050 299.400 ;
        RECT 13.950 298.950 16.050 299.400 ;
    END
  END Yin[3]
  PIN Yin[2]
    PORT
      LAYER metal2 ;
        RECT 14.400 722.400 15.600 724.650 ;
        RECT 14.400 685.050 15.450 722.400 ;
        RECT 13.950 682.950 16.050 685.050 ;
        RECT 14.400 651.600 15.450 682.950 ;
        RECT 14.400 649.350 15.600 651.600 ;
      LAYER metal3 ;
        RECT 13.950 684.600 16.050 685.050 ;
        RECT -3.600 683.400 16.050 684.600 ;
        RECT 13.950 682.950 16.050 683.400 ;
    END
  END Yin[2]
  PIN Yin[1]
    PORT
      LAYER metal1 ;
        RECT 22.950 732.450 25.050 733.050 ;
        RECT 34.950 732.450 37.050 733.050 ;
        RECT 22.950 731.550 37.050 732.450 ;
        RECT 22.950 730.950 25.050 731.550 ;
        RECT 34.950 730.950 37.050 731.550 ;
      LAYER metal2 ;
        RECT 169.950 761.100 172.050 763.200 ;
        RECT 178.950 761.100 181.050 763.200 ;
        RECT 170.400 760.350 171.600 761.100 ;
        RECT 179.400 748.050 180.450 761.100 ;
        RECT 103.950 745.950 106.050 748.050 ;
        RECT 178.950 745.950 181.050 748.050 ;
        RECT 104.400 742.050 105.450 745.950 ;
        RECT 36.000 741.450 40.050 742.050 ;
        RECT 35.400 739.950 40.050 741.450 ;
        RECT 103.800 739.950 105.900 742.050 ;
        RECT 35.400 733.050 36.450 739.950 ;
        RECT 22.950 727.950 25.050 733.050 ;
        RECT 34.950 729.000 37.050 733.050 ;
        RECT 35.400 727.350 36.600 729.000 ;
      LAYER via2 ;
        RECT 37.950 739.950 40.050 742.050 ;
      LAYER metal3 ;
        RECT 169.950 762.750 172.050 763.200 ;
        RECT 178.950 762.750 181.050 763.200 ;
        RECT 169.950 761.550 181.050 762.750 ;
        RECT 169.950 761.100 172.050 761.550 ;
        RECT 178.950 761.100 181.050 761.550 ;
        RECT 103.950 747.600 106.050 748.050 ;
        RECT 178.950 747.600 181.050 748.050 ;
        RECT 103.950 746.400 181.050 747.600 ;
        RECT 103.950 745.950 106.050 746.400 ;
        RECT 178.950 745.950 181.050 746.400 ;
        RECT 37.950 741.600 40.050 742.050 ;
        RECT 103.800 741.600 105.900 742.050 ;
        RECT 37.950 740.400 105.900 741.600 ;
        RECT 37.950 739.950 40.050 740.400 ;
        RECT 103.800 739.950 105.900 740.400 ;
        RECT 22.950 729.600 25.050 730.050 ;
        RECT -3.600 728.400 25.050 729.600 ;
        RECT 22.950 727.950 25.050 728.400 ;
    END
  END Yin[1]
  PIN Yin[0]
    PORT
      LAYER metal2 ;
        RECT 17.400 365.400 18.600 367.650 ;
        RECT 17.400 346.050 18.450 365.400 ;
        RECT 4.950 343.950 7.050 346.050 ;
        RECT 16.950 343.950 19.050 346.050 ;
        RECT 5.400 334.050 6.450 343.950 ;
        RECT 4.950 331.950 7.050 334.050 ;
        RECT 14.400 333.000 15.600 334.650 ;
        RECT 13.950 328.950 16.050 333.000 ;
      LAYER metal3 ;
        RECT 4.950 345.600 7.050 346.050 ;
        RECT 16.950 345.600 19.050 346.050 ;
        RECT 4.950 344.400 19.050 345.600 ;
        RECT 4.950 343.950 7.050 344.400 ;
        RECT 16.950 343.950 19.050 344.400 ;
        RECT 4.950 333.600 7.050 334.050 ;
        RECT -3.600 332.400 7.050 333.600 ;
        RECT 4.950 331.950 7.050 332.400 ;
        RECT 5.400 330.600 6.600 331.950 ;
        RECT 13.950 330.600 16.050 331.050 ;
        RECT 5.400 329.400 16.050 330.600 ;
        RECT 13.950 328.950 16.050 329.400 ;
    END
  END Yin[0]
  PIN Yout[3]
    PORT
      LAYER metal2 ;
        RECT 14.400 489.900 15.600 490.650 ;
        RECT 13.950 487.800 16.050 489.900 ;
      LAYER metal3 ;
        RECT 13.950 489.600 16.050 489.900 ;
        RECT -3.600 488.400 16.050 489.600 ;
        RECT 13.950 487.800 16.050 488.400 ;
    END
  END Yout[3]
  PIN Yout[2]
    PORT
      LAYER metal2 ;
        RECT 37.950 449.100 40.050 451.200 ;
        RECT 38.400 448.350 39.600 449.100 ;
      LAYER metal3 ;
        RECT 37.950 450.600 40.050 451.200 ;
        RECT -3.600 449.400 40.050 450.600 ;
        RECT 37.950 449.100 40.050 449.400 ;
    END
  END Yout[2]
  PIN Yout[1]
    PORT
      LAYER metal2 ;
        RECT 370.950 214.950 373.050 217.050 ;
        RECT 379.950 215.100 382.050 217.200 ;
        RECT 371.400 141.450 372.450 214.950 ;
        RECT 380.400 214.350 381.600 215.100 ;
        RECT 371.400 140.400 375.450 141.450 ;
        RECT 374.400 64.050 375.450 140.400 ;
        RECT 373.950 61.950 376.050 64.050 ;
        RECT 379.950 61.950 382.050 64.050 ;
        RECT 380.400 4.050 381.450 61.950 ;
        RECT 364.950 1.950 367.050 4.050 ;
        RECT 379.950 1.950 382.050 4.050 ;
        RECT 365.400 -3.600 366.450 1.950 ;
      LAYER metal3 ;
        RECT 370.950 216.600 373.050 217.050 ;
        RECT 379.950 216.600 382.050 217.200 ;
        RECT 370.950 215.400 382.050 216.600 ;
        RECT 370.950 214.950 373.050 215.400 ;
        RECT 379.950 215.100 382.050 215.400 ;
        RECT 373.950 63.600 376.050 64.050 ;
        RECT 379.950 63.600 382.050 64.050 ;
        RECT 373.950 62.400 382.050 63.600 ;
        RECT 373.950 61.950 376.050 62.400 ;
        RECT 379.950 61.950 382.050 62.400 ;
        RECT 364.950 3.600 367.050 4.050 ;
        RECT 379.950 3.600 382.050 4.050 ;
        RECT 364.950 2.400 382.050 3.600 ;
        RECT 364.950 1.950 367.050 2.400 ;
        RECT 379.950 1.950 382.050 2.400 ;
    END
  END Yout[1]
  PIN Yout[0]
    PORT
      LAYER metal2 ;
        RECT 389.400 20.400 390.600 22.650 ;
        RECT 389.400 -2.550 390.450 20.400 ;
        RECT 389.400 -3.600 393.450 -2.550 ;
    END
  END Yout[0]
  PIN clk
    PORT
      LAYER metal2 ;
        RECT 182.400 606.450 183.600 606.600 ;
        RECT 179.400 605.400 183.600 606.450 ;
        RECT 179.400 580.050 180.450 605.400 ;
        RECT 182.400 604.350 183.600 605.400 ;
        RECT 85.950 577.950 88.050 580.050 ;
        RECT 178.950 577.950 181.050 580.050 ;
        RECT 62.400 566.400 63.600 568.650 ;
        RECT 62.400 553.050 63.450 566.400 ;
        RECT 86.400 553.050 87.450 577.950 ;
        RECT 28.950 550.950 31.050 553.050 ;
        RECT 61.950 550.950 64.050 553.050 ;
        RECT 85.950 550.950 88.050 553.050 ;
        RECT 29.400 496.050 30.450 550.950 ;
        RECT 313.950 527.100 316.050 529.200 ;
        RECT 319.950 527.100 322.050 529.200 ;
        RECT 28.950 493.950 31.050 496.050 ;
        RECT 40.950 493.950 43.050 496.050 ;
        RECT 38.400 489.450 39.600 490.650 ;
        RECT 41.400 489.450 42.450 493.950 ;
        RECT 38.400 488.400 42.450 489.450 ;
        RECT 38.400 469.050 39.450 488.400 ;
        RECT 37.950 466.950 40.050 469.050 ;
        RECT 163.950 466.950 166.050 469.050 ;
        RECT 164.400 463.050 165.450 466.950 ;
        RECT 314.400 463.050 315.450 527.100 ;
        RECT 320.400 526.350 321.600 527.100 ;
        RECT 163.950 460.950 166.050 463.050 ;
        RECT 313.950 460.950 316.050 463.050 ;
        RECT 164.400 385.050 165.450 460.950 ;
        RECT 413.400 410.400 414.600 412.650 ;
        RECT 413.400 385.050 414.450 410.400 ;
        RECT 163.950 382.950 166.050 385.050 ;
        RECT 265.950 382.950 268.050 385.050 ;
        RECT 412.950 382.950 415.050 385.050 ;
        RECT 164.400 372.600 165.450 382.950 ;
        RECT 266.400 372.600 267.450 382.950 ;
        RECT 164.400 370.350 165.600 372.600 ;
        RECT 266.400 370.350 267.600 372.600 ;
      LAYER metal3 ;
        RECT 85.950 579.600 88.050 580.050 ;
        RECT 178.950 579.600 181.050 580.050 ;
        RECT 85.950 578.400 181.050 579.600 ;
        RECT 85.950 577.950 88.050 578.400 ;
        RECT 178.950 577.950 181.050 578.400 ;
        RECT 28.950 552.600 31.050 553.050 ;
        RECT 61.950 552.600 64.050 553.050 ;
        RECT 85.950 552.600 88.050 553.050 ;
        RECT 28.950 551.400 88.050 552.600 ;
        RECT 28.950 550.950 31.050 551.400 ;
        RECT 61.950 550.950 64.050 551.400 ;
        RECT 85.950 550.950 88.050 551.400 ;
        RECT 313.950 528.750 316.050 529.200 ;
        RECT 319.950 528.750 322.050 529.200 ;
        RECT 313.950 527.550 322.050 528.750 ;
        RECT 313.950 527.100 316.050 527.550 ;
        RECT 319.950 527.100 322.050 527.550 ;
        RECT 28.950 495.600 31.050 496.050 ;
        RECT 40.950 495.600 43.050 496.050 ;
        RECT -3.600 494.400 43.050 495.600 ;
        RECT 28.950 493.950 31.050 494.400 ;
        RECT 40.950 493.950 43.050 494.400 ;
        RECT 37.950 468.600 40.050 469.050 ;
        RECT 163.950 468.600 166.050 469.050 ;
        RECT 37.950 467.400 166.050 468.600 ;
        RECT 37.950 466.950 40.050 467.400 ;
        RECT 163.950 466.950 166.050 467.400 ;
        RECT 163.950 462.600 166.050 463.050 ;
        RECT 313.950 462.600 316.050 463.050 ;
        RECT 163.950 461.400 316.050 462.600 ;
        RECT 163.950 460.950 166.050 461.400 ;
        RECT 313.950 460.950 316.050 461.400 ;
        RECT 163.950 384.600 166.050 385.050 ;
        RECT 265.950 384.600 268.050 385.050 ;
        RECT 412.950 384.600 415.050 385.050 ;
        RECT 163.950 383.400 415.050 384.600 ;
        RECT 163.950 382.950 166.050 383.400 ;
        RECT 265.950 382.950 268.050 383.400 ;
        RECT 412.950 382.950 415.050 383.400 ;
    END
  END clk
  OBS
      LAYER metal1 ;
        RECT 14.100 974.400 15.300 975.000 ;
        RECT 14.100 971.400 15.900 974.400 ;
        RECT 17.100 971.400 18.900 974.400 ;
        RECT 17.400 967.200 18.300 971.400 ;
        RECT 20.100 969.000 21.900 975.000 ;
        RECT 23.100 968.400 24.900 974.400 ;
        RECT 38.400 968.400 40.200 975.000 ;
        RECT 17.400 966.300 22.800 967.200 ;
        RECT 20.700 965.400 22.800 966.300 ;
        RECT 14.400 961.050 16.200 962.850 ;
        RECT 14.100 958.950 16.200 961.050 ;
        RECT 17.400 958.950 19.500 961.050 ;
        RECT 18.000 957.150 19.800 958.950 ;
        RECT 20.700 954.900 21.600 965.400 ;
        RECT 24.000 961.050 24.900 968.400 ;
        RECT 43.500 967.200 45.300 974.400 ;
        RECT 62.400 968.400 64.200 975.000 ;
        RECT 67.500 967.200 69.300 974.400 ;
        RECT 41.100 966.300 45.300 967.200 ;
        RECT 65.100 966.300 69.300 967.200 ;
        RECT 38.250 961.050 40.050 962.850 ;
        RECT 41.100 961.050 42.300 966.300 ;
        RECT 44.100 961.050 45.900 962.850 ;
        RECT 62.250 961.050 64.050 962.850 ;
        RECT 65.100 961.050 66.300 966.300 ;
        RECT 83.100 965.400 84.900 975.000 ;
        RECT 89.700 966.000 91.500 974.400 ;
        RECT 110.100 971.400 111.900 975.000 ;
        RECT 113.100 971.400 114.900 974.400 ;
        RECT 89.700 964.800 93.000 966.000 ;
        RECT 68.100 961.050 69.900 962.850 ;
        RECT 83.100 961.050 84.900 962.850 ;
        RECT 89.100 961.050 90.900 962.850 ;
        RECT 92.100 961.050 93.000 964.800 ;
        RECT 113.100 961.050 114.300 971.400 ;
        RECT 128.100 969.300 129.900 974.400 ;
        RECT 131.100 970.200 132.900 975.000 ;
        RECT 134.100 969.300 135.900 974.400 ;
        RECT 128.100 967.950 135.900 969.300 ;
        RECT 137.100 968.400 138.900 974.400 ;
        RECT 152.100 971.400 153.900 974.400 ;
        RECT 155.100 971.400 156.900 975.000 ;
        RECT 137.100 966.300 138.300 968.400 ;
        RECT 134.700 965.400 138.300 966.300 ;
        RECT 131.100 961.050 132.900 962.850 ;
        RECT 134.700 961.050 135.900 965.400 ;
        RECT 137.100 961.050 138.900 962.850 ;
        RECT 152.700 961.050 153.900 971.400 ;
        RECT 170.400 968.400 172.200 975.000 ;
        RECT 175.500 967.200 177.300 974.400 ;
        RECT 191.100 971.400 192.900 975.000 ;
        RECT 194.100 971.400 195.900 974.400 ;
        RECT 173.100 966.300 177.300 967.200 ;
        RECT 170.250 961.050 172.050 962.850 ;
        RECT 173.100 961.050 174.300 966.300 ;
        RECT 176.100 961.050 177.900 962.850 ;
        RECT 194.100 961.050 195.300 971.400 ;
        RECT 211.500 966.000 213.300 974.400 ;
        RECT 210.000 964.800 213.300 966.000 ;
        RECT 218.100 965.400 219.900 975.000 ;
        RECT 238.500 966.000 240.300 974.400 ;
        RECT 237.000 964.800 240.300 966.000 ;
        RECT 245.100 965.400 246.900 975.000 ;
        RECT 262.500 966.000 264.300 974.400 ;
        RECT 261.000 964.800 264.300 966.000 ;
        RECT 269.100 965.400 270.900 975.000 ;
        RECT 285.000 968.400 286.800 975.000 ;
        RECT 289.500 969.600 291.300 974.400 ;
        RECT 292.500 971.400 294.300 975.000 ;
        RECT 289.500 968.400 294.600 969.600 ;
        RECT 312.000 968.400 313.800 975.000 ;
        RECT 316.500 969.600 318.300 974.400 ;
        RECT 319.500 971.400 321.300 975.000 ;
        RECT 316.500 968.400 321.600 969.600 ;
        RECT 210.000 961.050 210.900 964.800 ;
        RECT 220.950 963.450 223.050 964.050 ;
        RECT 229.950 963.450 232.050 964.050 ;
        RECT 212.100 961.050 213.900 962.850 ;
        RECT 218.100 961.050 219.900 962.850 ;
        RECT 220.950 962.550 232.050 963.450 ;
        RECT 220.950 961.950 223.050 962.550 ;
        RECT 229.950 961.950 232.050 962.550 ;
        RECT 237.000 961.050 237.900 964.800 ;
        RECT 239.100 961.050 240.900 962.850 ;
        RECT 245.100 961.050 246.900 962.850 ;
        RECT 261.000 961.050 261.900 964.800 ;
        RECT 263.100 961.050 264.900 962.850 ;
        RECT 269.100 961.050 270.900 962.850 ;
        RECT 284.100 961.050 285.900 962.850 ;
        RECT 290.250 961.050 292.050 962.850 ;
        RECT 293.700 961.050 294.600 968.400 ;
        RECT 311.100 961.050 312.900 962.850 ;
        RECT 317.250 961.050 319.050 962.850 ;
        RECT 320.700 961.050 321.600 968.400 ;
        RECT 335.100 969.300 336.900 974.400 ;
        RECT 338.100 970.200 339.900 975.000 ;
        RECT 341.100 969.300 342.900 974.400 ;
        RECT 335.100 967.950 342.900 969.300 ;
        RECT 344.100 968.400 345.900 974.400 ;
        RECT 359.100 971.400 360.900 975.000 ;
        RECT 362.100 971.400 363.900 974.400 ;
        RECT 344.100 966.300 345.300 968.400 ;
        RECT 341.700 965.400 345.300 966.300 ;
        RECT 338.100 961.050 339.900 962.850 ;
        RECT 341.700 961.050 342.900 965.400 ;
        RECT 344.100 961.050 345.900 962.850 ;
        RECT 362.100 961.050 363.300 971.400 ;
        RECT 377.700 967.200 379.500 974.400 ;
        RECT 382.800 968.400 384.600 975.000 ;
        RECT 377.700 966.300 381.900 967.200 ;
        RECT 377.100 961.050 378.900 962.850 ;
        RECT 380.700 961.050 381.900 966.300 ;
        RECT 401.100 965.400 402.900 975.000 ;
        RECT 407.700 966.000 409.500 974.400 ;
        RECT 407.700 964.800 411.000 966.000 ;
        RECT 425.100 965.400 426.900 975.000 ;
        RECT 431.700 966.000 433.500 974.400 ;
        RECT 452.700 967.200 454.500 974.400 ;
        RECT 457.800 968.400 459.600 975.000 ;
        RECT 452.700 966.300 456.900 967.200 ;
        RECT 431.700 964.800 435.000 966.000 ;
        RECT 382.950 961.050 384.750 962.850 ;
        RECT 401.100 961.050 402.900 962.850 ;
        RECT 407.100 961.050 408.900 962.850 ;
        RECT 410.100 961.050 411.000 964.800 ;
        RECT 425.100 961.050 426.900 962.850 ;
        RECT 431.100 961.050 432.900 962.850 ;
        RECT 434.100 961.050 435.000 964.800 ;
        RECT 452.100 961.050 453.900 962.850 ;
        RECT 455.700 961.050 456.900 966.300 ;
        RECT 475.500 966.000 477.300 974.400 ;
        RECT 474.000 964.800 477.300 966.000 ;
        RECT 482.100 965.400 483.900 975.000 ;
        RECT 498.000 968.400 499.800 975.000 ;
        RECT 502.500 969.600 504.300 974.400 ;
        RECT 505.500 971.400 507.300 975.000 ;
        RECT 502.500 968.400 507.600 969.600 ;
        RECT 457.950 961.050 459.750 962.850 ;
        RECT 474.000 961.050 474.900 964.800 ;
        RECT 476.100 961.050 477.900 962.850 ;
        RECT 482.100 961.050 483.900 962.850 ;
        RECT 497.100 961.050 498.900 962.850 ;
        RECT 503.250 961.050 505.050 962.850 ;
        RECT 506.700 961.050 507.600 968.400 ;
        RECT 521.100 969.300 522.900 974.400 ;
        RECT 524.100 970.200 525.900 975.000 ;
        RECT 527.100 969.300 528.900 974.400 ;
        RECT 521.100 967.950 528.900 969.300 ;
        RECT 530.100 968.400 531.900 974.400 ;
        RECT 548.700 971.400 550.500 975.000 ;
        RECT 551.700 969.600 553.500 974.400 ;
        RECT 548.400 968.400 553.500 969.600 ;
        RECT 556.200 968.400 558.000 975.000 ;
        RECT 572.100 971.400 573.900 974.400 ;
        RECT 575.100 971.400 576.900 975.000 ;
        RECT 530.100 966.300 531.300 968.400 ;
        RECT 527.700 965.400 531.300 966.300 ;
        RECT 524.100 961.050 525.900 962.850 ;
        RECT 527.700 961.050 528.900 965.400 ;
        RECT 535.950 963.450 538.050 964.050 ;
        RECT 544.950 963.450 547.050 964.050 ;
        RECT 530.100 961.050 531.900 962.850 ;
        RECT 535.950 962.550 547.050 963.450 ;
        RECT 535.950 961.950 538.050 962.550 ;
        RECT 544.950 961.950 547.050 962.550 ;
        RECT 548.400 961.050 549.300 968.400 ;
        RECT 550.950 961.050 552.750 962.850 ;
        RECT 557.100 961.050 558.900 962.850 ;
        RECT 572.700 961.050 573.900 971.400 ;
        RECT 593.100 965.400 594.900 975.000 ;
        RECT 599.700 966.000 601.500 974.400 ;
        RECT 619.500 966.000 621.300 974.400 ;
        RECT 599.700 964.800 603.000 966.000 ;
        RECT 593.100 961.050 594.900 962.850 ;
        RECT 599.100 961.050 600.900 962.850 ;
        RECT 602.100 961.050 603.000 964.800 ;
        RECT 618.000 964.800 621.300 966.000 ;
        RECT 626.100 965.400 627.900 975.000 ;
        RECT 641.400 968.400 643.200 975.000 ;
        RECT 646.500 967.200 648.300 974.400 ;
        RECT 662.100 968.400 663.900 974.400 ;
        RECT 644.100 966.300 648.300 967.200 ;
        RECT 662.700 966.300 663.900 968.400 ;
        RECT 665.100 969.300 666.900 974.400 ;
        RECT 668.100 970.200 669.900 975.000 ;
        RECT 671.100 969.300 672.900 974.400 ;
        RECT 686.100 971.400 687.900 975.000 ;
        RECT 689.100 971.400 690.900 974.400 ;
        RECT 692.100 971.400 693.900 975.000 ;
        RECT 665.100 967.950 672.900 969.300 ;
        RECT 618.000 961.050 618.900 964.800 ;
        RECT 620.100 961.050 621.900 962.850 ;
        RECT 626.100 961.050 627.900 962.850 ;
        RECT 641.250 961.050 643.050 962.850 ;
        RECT 644.100 961.050 645.300 966.300 ;
        RECT 662.700 965.400 666.300 966.300 ;
        RECT 647.100 961.050 648.900 962.850 ;
        RECT 662.100 961.050 663.900 962.850 ;
        RECT 665.100 961.050 666.300 965.400 ;
        RECT 668.100 961.050 669.900 962.850 ;
        RECT 689.700 961.050 690.600 971.400 ;
        RECT 707.700 967.200 709.500 974.400 ;
        RECT 712.800 968.400 714.600 975.000 ;
        RECT 731.400 968.400 733.200 975.000 ;
        RECT 736.500 967.200 738.300 974.400 ;
        RECT 707.700 966.300 711.900 967.200 ;
        RECT 707.100 961.050 708.900 962.850 ;
        RECT 710.700 961.050 711.900 966.300 ;
        RECT 712.950 966.450 715.050 967.050 ;
        RECT 730.950 966.450 733.050 967.050 ;
        RECT 712.950 965.550 733.050 966.450 ;
        RECT 712.950 964.950 715.050 965.550 ;
        RECT 730.950 964.950 733.050 965.550 ;
        RECT 734.100 966.300 738.300 967.200 ;
        RECT 712.950 961.050 714.750 962.850 ;
        RECT 731.250 961.050 733.050 962.850 ;
        RECT 734.100 961.050 735.300 966.300 ;
        RECT 755.100 965.400 756.900 975.000 ;
        RECT 761.700 966.000 763.500 974.400 ;
        RECT 779.100 968.400 780.900 974.400 ;
        RECT 779.700 966.300 780.900 968.400 ;
        RECT 782.100 969.300 783.900 974.400 ;
        RECT 785.100 970.200 786.900 975.000 ;
        RECT 788.100 969.300 789.900 974.400 ;
        RECT 803.700 971.400 805.500 975.000 ;
        RECT 806.700 969.600 808.500 974.400 ;
        RECT 782.100 967.950 789.900 969.300 ;
        RECT 803.400 968.400 808.500 969.600 ;
        RECT 811.200 968.400 813.000 975.000 ;
        RECT 827.100 971.400 828.900 974.400 ;
        RECT 830.100 971.400 831.900 975.000 ;
        RECT 761.700 964.800 765.000 966.000 ;
        RECT 779.700 965.400 783.300 966.300 ;
        RECT 737.100 961.050 738.900 962.850 ;
        RECT 755.100 961.050 756.900 962.850 ;
        RECT 761.100 961.050 762.900 962.850 ;
        RECT 764.100 961.050 765.000 964.800 ;
        RECT 779.100 961.050 780.900 962.850 ;
        RECT 782.100 961.050 783.300 965.400 ;
        RECT 785.100 961.050 786.900 962.850 ;
        RECT 803.400 961.050 804.300 968.400 ;
        RECT 808.950 966.450 811.050 967.050 ;
        RECT 823.950 966.450 826.050 967.200 ;
        RECT 808.950 965.550 826.050 966.450 ;
        RECT 808.950 964.950 811.050 965.550 ;
        RECT 823.950 965.100 826.050 965.550 ;
        RECT 805.950 961.050 807.750 962.850 ;
        RECT 812.100 961.050 813.900 962.850 ;
        RECT 827.700 961.050 828.900 971.400 ;
        RECT 829.950 966.450 832.050 967.200 ;
        RECT 844.950 966.450 847.050 967.050 ;
        RECT 829.950 965.550 847.050 966.450 ;
        RECT 829.950 965.100 832.050 965.550 ;
        RECT 844.950 964.950 847.050 965.550 ;
        RECT 848.100 965.400 849.900 975.000 ;
        RECT 854.700 966.000 856.500 974.400 ;
        RECT 874.500 966.000 876.300 974.400 ;
        RECT 854.700 964.800 858.000 966.000 ;
        RECT 848.100 961.050 849.900 962.850 ;
        RECT 854.100 961.050 855.900 962.850 ;
        RECT 857.100 961.050 858.000 964.800 ;
        RECT 873.000 964.800 876.300 966.000 ;
        RECT 881.100 965.400 882.900 975.000 ;
        RECT 883.950 969.450 886.050 970.050 ;
        RECT 889.950 969.450 892.050 970.050 ;
        RECT 883.950 968.550 892.050 969.450 ;
        RECT 883.950 967.950 886.050 968.550 ;
        RECT 889.950 967.950 892.050 968.550 ;
        RECT 896.100 965.400 897.900 975.000 ;
        RECT 902.700 966.000 904.500 974.400 ;
        RECT 920.700 971.400 922.500 975.000 ;
        RECT 923.700 969.600 925.500 974.400 ;
        RECT 920.400 968.400 925.500 969.600 ;
        RECT 928.200 968.400 930.000 975.000 ;
        RECT 902.700 964.800 906.000 966.000 ;
        RECT 873.000 961.050 873.900 964.800 ;
        RECT 875.100 961.050 876.900 962.850 ;
        RECT 881.100 961.050 882.900 962.850 ;
        RECT 896.100 961.050 897.900 962.850 ;
        RECT 902.100 961.050 903.900 962.850 ;
        RECT 905.100 961.050 906.000 964.800 ;
        RECT 920.400 961.050 921.300 968.400 ;
        RECT 925.950 966.450 928.050 967.050 ;
        RECT 943.950 966.450 946.050 967.050 ;
        RECT 925.950 965.550 946.050 966.450 ;
        RECT 925.950 964.950 928.050 965.550 ;
        RECT 943.950 964.950 946.050 965.550 ;
        RECT 947.100 965.400 948.900 975.000 ;
        RECT 953.700 966.000 955.500 974.400 ;
        RECT 953.700 964.800 957.000 966.000 ;
        RECT 971.100 965.400 972.900 975.000 ;
        RECT 977.700 966.000 979.500 974.400 ;
        RECT 1000.500 966.000 1002.300 974.400 ;
        RECT 977.700 964.800 981.000 966.000 ;
        RECT 922.950 961.050 924.750 962.850 ;
        RECT 929.100 961.050 930.900 962.850 ;
        RECT 947.100 961.050 948.900 962.850 ;
        RECT 953.100 961.050 954.900 962.850 ;
        RECT 956.100 961.050 957.000 964.800 ;
        RECT 971.100 961.050 972.900 962.850 ;
        RECT 977.100 961.050 978.900 962.850 ;
        RECT 980.100 961.050 981.000 964.800 ;
        RECT 999.000 964.800 1002.300 966.000 ;
        RECT 1007.100 965.400 1008.900 975.000 ;
        RECT 999.000 961.050 999.900 964.800 ;
        RECT 1001.100 961.050 1002.900 962.850 ;
        RECT 1007.100 961.050 1008.900 962.850 ;
        RECT 22.800 958.950 24.900 961.050 ;
        RECT 37.950 958.950 40.050 961.050 ;
        RECT 40.950 958.950 43.050 961.050 ;
        RECT 43.950 958.950 46.050 961.050 ;
        RECT 61.950 958.950 64.050 961.050 ;
        RECT 64.950 958.950 67.050 961.050 ;
        RECT 67.950 958.950 70.050 961.050 ;
        RECT 82.950 958.950 85.050 961.050 ;
        RECT 85.950 958.950 88.050 961.050 ;
        RECT 88.950 958.950 91.050 961.050 ;
        RECT 91.950 958.950 94.050 961.050 ;
        RECT 109.950 958.950 112.050 961.050 ;
        RECT 112.950 958.950 115.050 961.050 ;
        RECT 127.950 958.950 130.050 961.050 ;
        RECT 130.950 958.950 133.050 961.050 ;
        RECT 133.950 958.950 136.050 961.050 ;
        RECT 136.950 958.950 139.050 961.050 ;
        RECT 151.950 958.950 154.050 961.050 ;
        RECT 154.950 958.950 157.050 961.050 ;
        RECT 169.950 958.950 172.050 961.050 ;
        RECT 172.950 958.950 175.050 961.050 ;
        RECT 175.950 958.950 178.050 961.050 ;
        RECT 190.950 958.950 193.050 961.050 ;
        RECT 193.950 958.950 196.050 961.050 ;
        RECT 208.950 958.950 211.050 961.050 ;
        RECT 211.950 958.950 214.050 961.050 ;
        RECT 214.950 958.950 217.050 961.050 ;
        RECT 217.950 958.950 220.050 961.050 ;
        RECT 235.950 958.950 238.050 961.050 ;
        RECT 238.950 958.950 241.050 961.050 ;
        RECT 241.950 958.950 244.050 961.050 ;
        RECT 244.950 958.950 247.050 961.050 ;
        RECT 259.950 958.950 262.050 961.050 ;
        RECT 262.950 958.950 265.050 961.050 ;
        RECT 265.950 958.950 268.050 961.050 ;
        RECT 268.950 958.950 271.050 961.050 ;
        RECT 283.950 958.950 286.050 961.050 ;
        RECT 286.950 958.950 289.050 961.050 ;
        RECT 289.950 958.950 292.050 961.050 ;
        RECT 292.950 958.950 295.050 961.050 ;
        RECT 310.950 958.950 313.050 961.050 ;
        RECT 313.950 958.950 316.050 961.050 ;
        RECT 316.950 958.950 319.050 961.050 ;
        RECT 319.950 958.950 322.050 961.050 ;
        RECT 334.950 958.950 337.050 961.050 ;
        RECT 337.950 958.950 340.050 961.050 ;
        RECT 340.950 958.950 343.050 961.050 ;
        RECT 343.950 958.950 346.050 961.050 ;
        RECT 358.950 958.950 361.050 961.050 ;
        RECT 361.950 958.950 364.050 961.050 ;
        RECT 376.950 958.950 379.050 961.050 ;
        RECT 379.950 958.950 382.050 961.050 ;
        RECT 382.950 958.950 385.050 961.050 ;
        RECT 400.950 958.950 403.050 961.050 ;
        RECT 403.950 958.950 406.050 961.050 ;
        RECT 406.950 958.950 409.050 961.050 ;
        RECT 409.950 958.950 412.050 961.050 ;
        RECT 424.950 958.950 427.050 961.050 ;
        RECT 427.950 958.950 430.050 961.050 ;
        RECT 430.950 958.950 433.050 961.050 ;
        RECT 433.950 958.950 436.050 961.050 ;
        RECT 451.950 958.950 454.050 961.050 ;
        RECT 454.950 958.950 457.050 961.050 ;
        RECT 457.950 958.950 460.050 961.050 ;
        RECT 472.950 958.950 475.050 961.050 ;
        RECT 475.950 958.950 478.050 961.050 ;
        RECT 478.950 958.950 481.050 961.050 ;
        RECT 481.950 958.950 484.050 961.050 ;
        RECT 496.950 958.950 499.050 961.050 ;
        RECT 499.950 958.950 502.050 961.050 ;
        RECT 502.950 958.950 505.050 961.050 ;
        RECT 505.950 958.950 508.050 961.050 ;
        RECT 520.950 958.950 523.050 961.050 ;
        RECT 523.950 958.950 526.050 961.050 ;
        RECT 526.950 958.950 529.050 961.050 ;
        RECT 529.950 958.950 532.050 961.050 ;
        RECT 547.950 958.950 550.050 961.050 ;
        RECT 550.950 958.950 553.050 961.050 ;
        RECT 553.950 958.950 556.050 961.050 ;
        RECT 556.950 958.950 559.050 961.050 ;
        RECT 571.950 958.950 574.050 961.050 ;
        RECT 574.950 958.950 577.050 961.050 ;
        RECT 592.950 958.950 595.050 961.050 ;
        RECT 595.950 958.950 598.050 961.050 ;
        RECT 598.950 958.950 601.050 961.050 ;
        RECT 601.950 958.950 604.050 961.050 ;
        RECT 616.950 958.950 619.050 961.050 ;
        RECT 619.950 958.950 622.050 961.050 ;
        RECT 622.950 958.950 625.050 961.050 ;
        RECT 625.950 958.950 628.050 961.050 ;
        RECT 640.950 958.950 643.050 961.050 ;
        RECT 643.950 958.950 646.050 961.050 ;
        RECT 646.950 958.950 649.050 961.050 ;
        RECT 661.950 958.950 664.050 961.050 ;
        RECT 664.950 958.950 667.050 961.050 ;
        RECT 667.950 958.950 670.050 961.050 ;
        RECT 670.950 958.950 673.050 961.050 ;
        RECT 685.950 958.950 688.050 961.050 ;
        RECT 688.950 958.950 691.050 961.050 ;
        RECT 691.950 958.950 694.050 961.050 ;
        RECT 706.950 958.950 709.050 961.050 ;
        RECT 709.950 958.950 712.050 961.050 ;
        RECT 712.950 958.950 715.050 961.050 ;
        RECT 730.950 958.950 733.050 961.050 ;
        RECT 733.950 958.950 736.050 961.050 ;
        RECT 736.950 958.950 739.050 961.050 ;
        RECT 754.950 958.950 757.050 961.050 ;
        RECT 757.950 958.950 760.050 961.050 ;
        RECT 760.950 958.950 763.050 961.050 ;
        RECT 763.950 958.950 766.050 961.050 ;
        RECT 778.950 958.950 781.050 961.050 ;
        RECT 781.950 958.950 784.050 961.050 ;
        RECT 784.950 958.950 787.050 961.050 ;
        RECT 787.950 958.950 790.050 961.050 ;
        RECT 802.950 958.950 805.050 961.050 ;
        RECT 805.950 958.950 808.050 961.050 ;
        RECT 808.950 958.950 811.050 961.050 ;
        RECT 811.950 958.950 814.050 961.050 ;
        RECT 826.950 958.950 829.050 961.050 ;
        RECT 829.950 958.950 832.050 961.050 ;
        RECT 847.950 958.950 850.050 961.050 ;
        RECT 850.950 958.950 853.050 961.050 ;
        RECT 853.950 958.950 856.050 961.050 ;
        RECT 856.950 958.950 859.050 961.050 ;
        RECT 871.950 958.950 874.050 961.050 ;
        RECT 874.950 958.950 877.050 961.050 ;
        RECT 877.950 958.950 880.050 961.050 ;
        RECT 880.950 958.950 883.050 961.050 ;
        RECT 895.950 958.950 898.050 961.050 ;
        RECT 898.950 958.950 901.050 961.050 ;
        RECT 901.950 958.950 904.050 961.050 ;
        RECT 904.950 958.950 907.050 961.050 ;
        RECT 919.950 958.950 922.050 961.050 ;
        RECT 922.950 958.950 925.050 961.050 ;
        RECT 925.950 958.950 928.050 961.050 ;
        RECT 928.950 958.950 931.050 961.050 ;
        RECT 946.950 958.950 949.050 961.050 ;
        RECT 949.950 958.950 952.050 961.050 ;
        RECT 952.950 958.950 955.050 961.050 ;
        RECT 955.950 958.950 958.050 961.050 ;
        RECT 970.950 958.950 973.050 961.050 ;
        RECT 973.950 958.950 976.050 961.050 ;
        RECT 976.950 958.950 979.050 961.050 ;
        RECT 979.950 958.950 982.050 961.050 ;
        RECT 997.950 958.950 1000.050 961.050 ;
        RECT 1000.950 958.950 1003.050 961.050 ;
        RECT 1003.950 958.950 1006.050 961.050 ;
        RECT 1006.950 958.950 1009.050 961.050 ;
        RECT 20.100 954.300 21.900 954.900 ;
        RECT 14.100 953.100 21.900 954.300 ;
        RECT 14.100 951.600 15.300 953.100 ;
        RECT 22.800 951.600 24.000 958.950 ;
        RECT 14.100 939.600 15.900 951.600 ;
        RECT 18.600 939.000 20.400 951.600 ;
        RECT 21.600 950.100 24.000 951.600 ;
        RECT 21.600 939.600 23.400 950.100 ;
        RECT 41.100 945.600 42.300 958.950 ;
        RECT 65.100 945.600 66.300 958.950 ;
        RECT 86.100 957.150 87.900 958.950 ;
        RECT 92.100 946.800 93.000 958.950 ;
        RECT 110.100 957.150 111.900 958.950 ;
        RECT 86.400 945.900 93.000 946.800 ;
        RECT 86.400 945.600 87.900 945.900 ;
        RECT 38.100 939.000 39.900 945.600 ;
        RECT 41.100 939.600 42.900 945.600 ;
        RECT 44.100 939.000 45.900 945.600 ;
        RECT 62.100 939.000 63.900 945.600 ;
        RECT 65.100 939.600 66.900 945.600 ;
        RECT 68.100 939.000 69.900 945.600 ;
        RECT 83.100 939.000 84.900 945.600 ;
        RECT 86.100 939.600 87.900 945.600 ;
        RECT 92.100 945.600 93.000 945.900 ;
        RECT 113.100 945.600 114.300 958.950 ;
        RECT 128.100 957.150 129.900 958.950 ;
        RECT 134.700 951.600 135.900 958.950 ;
        RECT 89.100 939.000 90.900 945.000 ;
        RECT 92.100 939.600 93.900 945.600 ;
        RECT 110.100 939.000 111.900 945.600 ;
        RECT 113.100 939.600 114.900 945.600 ;
        RECT 128.400 939.000 130.200 951.600 ;
        RECT 133.500 950.100 135.900 951.600 ;
        RECT 133.500 939.600 135.300 950.100 ;
        RECT 136.200 947.100 138.000 948.900 ;
        RECT 152.700 945.600 153.900 958.950 ;
        RECT 155.100 957.150 156.900 958.950 ;
        RECT 173.100 945.600 174.300 958.950 ;
        RECT 191.100 957.150 192.900 958.950 ;
        RECT 194.100 945.600 195.300 958.950 ;
        RECT 210.000 946.800 210.900 958.950 ;
        RECT 215.100 957.150 216.900 958.950 ;
        RECT 237.000 946.800 237.900 958.950 ;
        RECT 242.100 957.150 243.900 958.950 ;
        RECT 261.000 946.800 261.900 958.950 ;
        RECT 266.100 957.150 267.900 958.950 ;
        RECT 287.250 957.150 289.050 958.950 ;
        RECT 262.950 954.450 265.050 955.050 ;
        RECT 283.950 954.450 286.050 955.050 ;
        RECT 262.950 953.550 286.050 954.450 ;
        RECT 262.950 952.950 265.050 953.550 ;
        RECT 283.950 952.950 286.050 953.550 ;
        RECT 293.700 951.600 294.600 958.950 ;
        RECT 314.250 957.150 316.050 958.950 ;
        RECT 295.950 954.450 298.050 955.050 ;
        RECT 316.950 954.450 319.050 954.750 ;
        RECT 295.950 953.550 319.050 954.450 ;
        RECT 295.950 952.950 298.050 953.550 ;
        RECT 316.950 952.650 319.050 953.550 ;
        RECT 320.700 951.600 321.600 958.950 ;
        RECT 335.100 957.150 336.900 958.950 ;
        RECT 322.950 954.450 325.050 954.750 ;
        RECT 337.950 954.450 340.050 954.750 ;
        RECT 322.950 953.550 340.050 954.450 ;
        RECT 322.950 952.650 325.050 953.550 ;
        RECT 337.950 952.650 340.050 953.550 ;
        RECT 341.700 951.600 342.900 958.950 ;
        RECT 359.100 957.150 360.900 958.950 ;
        RECT 284.100 950.700 291.900 951.600 ;
        RECT 210.000 945.900 216.600 946.800 ;
        RECT 210.000 945.600 210.900 945.900 ;
        RECT 136.500 939.000 138.300 945.600 ;
        RECT 152.100 939.600 153.900 945.600 ;
        RECT 155.100 939.000 156.900 945.600 ;
        RECT 170.100 939.000 171.900 945.600 ;
        RECT 173.100 939.600 174.900 945.600 ;
        RECT 176.100 939.000 177.900 945.600 ;
        RECT 191.100 939.000 192.900 945.600 ;
        RECT 194.100 939.600 195.900 945.600 ;
        RECT 209.100 939.600 210.900 945.600 ;
        RECT 215.100 945.600 216.600 945.900 ;
        RECT 237.000 945.900 243.600 946.800 ;
        RECT 237.000 945.600 237.900 945.900 ;
        RECT 212.100 939.000 213.900 945.000 ;
        RECT 215.100 939.600 216.900 945.600 ;
        RECT 218.100 939.000 219.900 945.600 ;
        RECT 236.100 939.600 237.900 945.600 ;
        RECT 242.100 945.600 243.600 945.900 ;
        RECT 261.000 945.900 267.600 946.800 ;
        RECT 261.000 945.600 261.900 945.900 ;
        RECT 239.100 939.000 240.900 945.000 ;
        RECT 242.100 939.600 243.900 945.600 ;
        RECT 245.100 939.000 246.900 945.600 ;
        RECT 260.100 939.600 261.900 945.600 ;
        RECT 266.100 945.600 267.600 945.900 ;
        RECT 263.100 939.000 264.900 945.000 ;
        RECT 266.100 939.600 267.900 945.600 ;
        RECT 269.100 939.000 270.900 945.600 ;
        RECT 284.100 939.600 285.900 950.700 ;
        RECT 287.100 939.000 288.900 949.800 ;
        RECT 290.100 939.600 291.900 950.700 ;
        RECT 293.100 939.600 294.900 951.600 ;
        RECT 311.100 950.700 318.900 951.600 ;
        RECT 311.100 939.600 312.900 950.700 ;
        RECT 314.100 939.000 315.900 949.800 ;
        RECT 317.100 939.600 318.900 950.700 ;
        RECT 320.100 939.600 321.900 951.600 ;
        RECT 335.400 939.000 337.200 951.600 ;
        RECT 340.500 950.100 342.900 951.600 ;
        RECT 340.500 939.600 342.300 950.100 ;
        RECT 343.200 947.100 345.000 948.900 ;
        RECT 362.100 945.600 363.300 958.950 ;
        RECT 380.700 945.600 381.900 958.950 ;
        RECT 404.100 957.150 405.900 958.950 ;
        RECT 410.100 946.800 411.000 958.950 ;
        RECT 428.100 957.150 429.900 958.950 ;
        RECT 434.100 946.800 435.000 958.950 ;
        RECT 404.400 945.900 411.000 946.800 ;
        RECT 404.400 945.600 405.900 945.900 ;
        RECT 343.500 939.000 345.300 945.600 ;
        RECT 359.100 939.000 360.900 945.600 ;
        RECT 362.100 939.600 363.900 945.600 ;
        RECT 377.100 939.000 378.900 945.600 ;
        RECT 380.100 939.600 381.900 945.600 ;
        RECT 383.100 939.000 384.900 945.600 ;
        RECT 401.100 939.000 402.900 945.600 ;
        RECT 404.100 939.600 405.900 945.600 ;
        RECT 410.100 945.600 411.000 945.900 ;
        RECT 428.400 945.900 435.000 946.800 ;
        RECT 428.400 945.600 429.900 945.900 ;
        RECT 407.100 939.000 408.900 945.000 ;
        RECT 410.100 939.600 411.900 945.600 ;
        RECT 425.100 939.000 426.900 945.600 ;
        RECT 428.100 939.600 429.900 945.600 ;
        RECT 434.100 945.600 435.000 945.900 ;
        RECT 455.700 945.600 456.900 958.950 ;
        RECT 474.000 946.800 474.900 958.950 ;
        RECT 479.100 957.150 480.900 958.950 ;
        RECT 500.250 957.150 502.050 958.950 ;
        RECT 475.950 954.450 478.050 955.050 ;
        RECT 496.950 954.450 499.050 955.050 ;
        RECT 475.950 953.550 499.050 954.450 ;
        RECT 475.950 952.950 478.050 953.550 ;
        RECT 496.950 952.950 499.050 953.550 ;
        RECT 506.700 951.600 507.600 958.950 ;
        RECT 521.100 957.150 522.900 958.950 ;
        RECT 527.700 951.600 528.900 958.950 ;
        RECT 548.400 951.600 549.300 958.950 ;
        RECT 553.950 957.150 555.750 958.950 ;
        RECT 497.100 950.700 504.900 951.600 ;
        RECT 474.000 945.900 480.600 946.800 ;
        RECT 474.000 945.600 474.900 945.900 ;
        RECT 431.100 939.000 432.900 945.000 ;
        RECT 434.100 939.600 435.900 945.600 ;
        RECT 452.100 939.000 453.900 945.600 ;
        RECT 455.100 939.600 456.900 945.600 ;
        RECT 458.100 939.000 459.900 945.600 ;
        RECT 473.100 939.600 474.900 945.600 ;
        RECT 479.100 945.600 480.600 945.900 ;
        RECT 476.100 939.000 477.900 945.000 ;
        RECT 479.100 939.600 480.900 945.600 ;
        RECT 482.100 939.000 483.900 945.600 ;
        RECT 497.100 939.600 498.900 950.700 ;
        RECT 500.100 939.000 501.900 949.800 ;
        RECT 503.100 939.600 504.900 950.700 ;
        RECT 506.100 939.600 507.900 951.600 ;
        RECT 521.400 939.000 523.200 951.600 ;
        RECT 526.500 950.100 528.900 951.600 ;
        RECT 526.500 939.600 528.300 950.100 ;
        RECT 529.200 947.100 531.000 948.900 ;
        RECT 529.500 939.000 531.300 945.600 ;
        RECT 548.100 939.600 549.900 951.600 ;
        RECT 551.100 950.700 558.900 951.600 ;
        RECT 551.100 939.600 552.900 950.700 ;
        RECT 554.100 939.000 555.900 949.800 ;
        RECT 557.100 939.600 558.900 950.700 ;
        RECT 572.700 945.600 573.900 958.950 ;
        RECT 575.100 957.150 576.900 958.950 ;
        RECT 596.100 957.150 597.900 958.950 ;
        RECT 574.950 954.450 577.050 955.050 ;
        RECT 592.950 954.450 595.050 955.050 ;
        RECT 574.950 953.550 595.050 954.450 ;
        RECT 574.950 952.950 577.050 953.550 ;
        RECT 592.950 952.950 595.050 953.550 ;
        RECT 602.100 946.800 603.000 958.950 ;
        RECT 596.400 945.900 603.000 946.800 ;
        RECT 596.400 945.600 597.900 945.900 ;
        RECT 572.100 939.600 573.900 945.600 ;
        RECT 575.100 939.000 576.900 945.600 ;
        RECT 593.100 939.000 594.900 945.600 ;
        RECT 596.100 939.600 597.900 945.600 ;
        RECT 602.100 945.600 603.000 945.900 ;
        RECT 618.000 946.800 618.900 958.950 ;
        RECT 623.100 957.150 624.900 958.950 ;
        RECT 618.000 945.900 624.600 946.800 ;
        RECT 618.000 945.600 618.900 945.900 ;
        RECT 599.100 939.000 600.900 945.000 ;
        RECT 602.100 939.600 603.900 945.600 ;
        RECT 617.100 939.600 618.900 945.600 ;
        RECT 623.100 945.600 624.600 945.900 ;
        RECT 644.100 945.600 645.300 958.950 ;
        RECT 665.100 951.600 666.300 958.950 ;
        RECT 671.100 957.150 672.900 958.950 ;
        RECT 686.100 957.150 687.900 958.950 ;
        RECT 689.700 951.600 690.600 958.950 ;
        RECT 691.950 957.150 693.750 958.950 ;
        RECT 665.100 950.100 667.500 951.600 ;
        RECT 663.000 947.100 664.800 948.900 ;
        RECT 620.100 939.000 621.900 945.000 ;
        RECT 623.100 939.600 624.900 945.600 ;
        RECT 626.100 939.000 627.900 945.600 ;
        RECT 641.100 939.000 642.900 945.600 ;
        RECT 644.100 939.600 645.900 945.600 ;
        RECT 647.100 939.000 648.900 945.600 ;
        RECT 662.700 939.000 664.500 945.600 ;
        RECT 665.700 939.600 667.500 950.100 ;
        RECT 670.800 939.000 672.600 951.600 ;
        RECT 687.000 950.400 690.600 951.600 ;
        RECT 687.000 939.600 688.800 950.400 ;
        RECT 692.100 939.000 693.900 951.600 ;
        RECT 710.700 945.600 711.900 958.950 ;
        RECT 734.100 945.600 735.300 958.950 ;
        RECT 758.100 957.150 759.900 958.950 ;
        RECT 751.950 954.450 754.050 955.050 ;
        RECT 760.950 954.450 763.050 955.050 ;
        RECT 751.950 953.550 763.050 954.450 ;
        RECT 751.950 952.950 754.050 953.550 ;
        RECT 760.950 952.950 763.050 953.550 ;
        RECT 764.100 946.800 765.000 958.950 ;
        RECT 782.100 951.600 783.300 958.950 ;
        RECT 788.100 957.150 789.900 958.950 ;
        RECT 803.400 951.600 804.300 958.950 ;
        RECT 808.950 957.150 810.750 958.950 ;
        RECT 782.100 950.100 784.500 951.600 ;
        RECT 780.000 947.100 781.800 948.900 ;
        RECT 758.400 945.900 765.000 946.800 ;
        RECT 758.400 945.600 759.900 945.900 ;
        RECT 707.100 939.000 708.900 945.600 ;
        RECT 710.100 939.600 711.900 945.600 ;
        RECT 713.100 939.000 714.900 945.600 ;
        RECT 731.100 939.000 732.900 945.600 ;
        RECT 734.100 939.600 735.900 945.600 ;
        RECT 737.100 939.000 738.900 945.600 ;
        RECT 755.100 939.000 756.900 945.600 ;
        RECT 758.100 939.600 759.900 945.600 ;
        RECT 764.100 945.600 765.000 945.900 ;
        RECT 761.100 939.000 762.900 945.000 ;
        RECT 764.100 939.600 765.900 945.600 ;
        RECT 779.700 939.000 781.500 945.600 ;
        RECT 782.700 939.600 784.500 950.100 ;
        RECT 787.800 939.000 789.600 951.600 ;
        RECT 803.100 939.600 804.900 951.600 ;
        RECT 806.100 950.700 813.900 951.600 ;
        RECT 806.100 939.600 807.900 950.700 ;
        RECT 809.100 939.000 810.900 949.800 ;
        RECT 812.100 939.600 813.900 950.700 ;
        RECT 827.700 945.600 828.900 958.950 ;
        RECT 830.100 957.150 831.900 958.950 ;
        RECT 851.100 957.150 852.900 958.950 ;
        RECT 844.950 954.450 847.050 955.050 ;
        RECT 853.950 954.450 856.050 954.750 ;
        RECT 844.950 953.550 856.050 954.450 ;
        RECT 844.950 952.950 847.050 953.550 ;
        RECT 853.950 952.650 856.050 953.550 ;
        RECT 857.100 946.800 858.000 958.950 ;
        RECT 859.950 954.450 862.050 955.050 ;
        RECT 865.950 954.450 868.050 955.050 ;
        RECT 859.950 953.550 868.050 954.450 ;
        RECT 859.950 952.950 862.050 953.550 ;
        RECT 865.950 952.950 868.050 953.550 ;
        RECT 851.400 945.900 858.000 946.800 ;
        RECT 851.400 945.600 852.900 945.900 ;
        RECT 827.100 939.600 828.900 945.600 ;
        RECT 830.100 939.000 831.900 945.600 ;
        RECT 848.100 939.000 849.900 945.600 ;
        RECT 851.100 939.600 852.900 945.600 ;
        RECT 857.100 945.600 858.000 945.900 ;
        RECT 873.000 946.800 873.900 958.950 ;
        RECT 878.100 957.150 879.900 958.950 ;
        RECT 899.100 957.150 900.900 958.950 ;
        RECT 874.950 954.450 877.050 955.050 ;
        RECT 886.950 954.450 889.050 954.900 ;
        RECT 874.950 953.550 889.050 954.450 ;
        RECT 874.950 952.950 877.050 953.550 ;
        RECT 886.950 952.800 889.050 953.550 ;
        RECT 905.100 946.800 906.000 958.950 ;
        RECT 920.400 951.600 921.300 958.950 ;
        RECT 925.950 957.150 927.750 958.950 ;
        RECT 950.100 957.150 951.900 958.950 ;
        RECT 934.950 954.450 937.050 955.050 ;
        RECT 952.950 954.450 955.050 955.050 ;
        RECT 934.950 953.550 955.050 954.450 ;
        RECT 934.950 952.950 937.050 953.550 ;
        RECT 952.950 952.950 955.050 953.550 ;
        RECT 873.000 945.900 879.600 946.800 ;
        RECT 873.000 945.600 873.900 945.900 ;
        RECT 854.100 939.000 855.900 945.000 ;
        RECT 857.100 939.600 858.900 945.600 ;
        RECT 872.100 939.600 873.900 945.600 ;
        RECT 878.100 945.600 879.600 945.900 ;
        RECT 899.400 945.900 906.000 946.800 ;
        RECT 899.400 945.600 900.900 945.900 ;
        RECT 875.100 939.000 876.900 945.000 ;
        RECT 878.100 939.600 879.900 945.600 ;
        RECT 881.100 939.000 882.900 945.600 ;
        RECT 896.100 939.000 897.900 945.600 ;
        RECT 899.100 939.600 900.900 945.600 ;
        RECT 905.100 945.600 906.000 945.900 ;
        RECT 902.100 939.000 903.900 945.000 ;
        RECT 905.100 939.600 906.900 945.600 ;
        RECT 920.100 939.600 921.900 951.600 ;
        RECT 923.100 950.700 930.900 951.600 ;
        RECT 923.100 939.600 924.900 950.700 ;
        RECT 926.100 939.000 927.900 949.800 ;
        RECT 929.100 939.600 930.900 950.700 ;
        RECT 956.100 946.800 957.000 958.950 ;
        RECT 974.100 957.150 975.900 958.950 ;
        RECT 980.100 946.800 981.000 958.950 ;
        RECT 950.400 945.900 957.000 946.800 ;
        RECT 950.400 945.600 951.900 945.900 ;
        RECT 947.100 939.000 948.900 945.600 ;
        RECT 950.100 939.600 951.900 945.600 ;
        RECT 956.100 945.600 957.000 945.900 ;
        RECT 974.400 945.900 981.000 946.800 ;
        RECT 974.400 945.600 975.900 945.900 ;
        RECT 953.100 939.000 954.900 945.000 ;
        RECT 956.100 939.600 957.900 945.600 ;
        RECT 971.100 939.000 972.900 945.600 ;
        RECT 974.100 939.600 975.900 945.600 ;
        RECT 980.100 945.600 981.000 945.900 ;
        RECT 999.000 946.800 999.900 958.950 ;
        RECT 1004.100 957.150 1005.900 958.950 ;
        RECT 999.000 945.900 1005.600 946.800 ;
        RECT 999.000 945.600 999.900 945.900 ;
        RECT 977.100 939.000 978.900 945.000 ;
        RECT 980.100 939.600 981.900 945.600 ;
        RECT 998.100 939.600 999.900 945.600 ;
        RECT 1004.100 945.600 1005.600 945.900 ;
        RECT 1001.100 939.000 1002.900 945.000 ;
        RECT 1004.100 939.600 1005.900 945.600 ;
        RECT 1007.100 939.000 1008.900 945.600 ;
        RECT 17.400 923.400 19.200 936.000 ;
        RECT 22.500 924.900 24.300 935.400 ;
        RECT 25.500 929.400 27.300 936.000 ;
        RECT 44.100 929.400 45.900 936.000 ;
        RECT 47.100 929.400 48.900 935.400 ;
        RECT 50.100 930.000 51.900 936.000 ;
        RECT 47.400 929.100 48.900 929.400 ;
        RECT 53.100 929.400 54.900 935.400 ;
        RECT 68.100 929.400 69.900 936.000 ;
        RECT 71.100 929.400 72.900 935.400 ;
        RECT 74.100 929.400 75.900 936.000 ;
        RECT 89.100 929.400 90.900 935.400 ;
        RECT 92.100 929.400 93.900 936.000 ;
        RECT 110.100 929.400 111.900 936.000 ;
        RECT 113.100 929.400 114.900 935.400 ;
        RECT 116.100 930.000 117.900 936.000 ;
        RECT 53.100 929.100 54.000 929.400 ;
        RECT 47.400 928.200 54.000 929.100 ;
        RECT 25.200 926.100 27.000 927.900 ;
        RECT 22.500 923.400 24.900 924.900 ;
        RECT 17.100 916.050 18.900 917.850 ;
        RECT 23.700 916.050 24.900 923.400 ;
        RECT 47.100 916.050 48.900 917.850 ;
        RECT 53.100 916.050 54.000 928.200 ;
        RECT 71.100 916.050 72.300 929.400 ;
        RECT 89.700 916.050 90.900 929.400 ;
        RECT 113.400 929.100 114.900 929.400 ;
        RECT 119.100 929.400 120.900 935.400 ;
        RECT 119.100 929.100 120.000 929.400 ;
        RECT 113.400 928.200 120.000 929.100 ;
        RECT 92.100 916.050 93.900 917.850 ;
        RECT 113.100 916.050 114.900 917.850 ;
        RECT 119.100 916.050 120.000 928.200 ;
        RECT 134.100 924.300 135.900 935.400 ;
        RECT 137.100 925.200 138.900 936.000 ;
        RECT 140.100 924.300 141.900 935.400 ;
        RECT 134.100 923.400 141.900 924.300 ;
        RECT 143.100 923.400 144.900 935.400 ;
        RECT 158.100 929.400 159.900 936.000 ;
        RECT 161.100 929.400 162.900 935.400 ;
        RECT 164.100 929.400 165.900 936.000 ;
        RECT 179.100 929.400 180.900 936.000 ;
        RECT 182.100 929.400 183.900 935.400 ;
        RECT 185.100 930.000 186.900 936.000 ;
        RECT 137.250 916.050 139.050 917.850 ;
        RECT 143.700 916.050 144.600 923.400 ;
        RECT 161.700 916.050 162.900 929.400 ;
        RECT 182.400 929.100 183.900 929.400 ;
        RECT 188.100 929.400 189.900 935.400 ;
        RECT 188.100 929.100 189.000 929.400 ;
        RECT 182.400 928.200 189.000 929.100 ;
        RECT 182.100 916.050 183.900 917.850 ;
        RECT 188.100 916.050 189.000 928.200 ;
        RECT 203.400 923.400 205.200 936.000 ;
        RECT 208.500 924.900 210.300 935.400 ;
        RECT 211.500 929.400 213.300 936.000 ;
        RECT 211.200 926.100 213.000 927.900 ;
        RECT 208.500 923.400 210.900 924.900 ;
        RECT 227.400 923.400 229.200 936.000 ;
        RECT 232.500 924.900 234.300 935.400 ;
        RECT 235.500 929.400 237.300 936.000 ;
        RECT 251.100 929.400 252.900 935.400 ;
        RECT 254.100 929.400 255.900 936.000 ;
        RECT 272.100 929.400 273.900 935.400 ;
        RECT 275.100 930.000 276.900 936.000 ;
        RECT 235.200 926.100 237.000 927.900 ;
        RECT 241.950 925.950 247.050 928.050 ;
        RECT 232.500 923.400 234.900 924.900 ;
        RECT 203.100 916.050 204.900 917.850 ;
        RECT 209.700 916.050 210.900 923.400 ;
        RECT 227.100 916.050 228.900 917.850 ;
        RECT 233.700 916.050 234.900 923.400 ;
        RECT 235.950 924.450 238.050 925.050 ;
        RECT 247.950 924.450 250.050 924.900 ;
        RECT 235.950 923.550 250.050 924.450 ;
        RECT 235.950 922.950 238.050 923.550 ;
        RECT 247.950 922.800 250.050 923.550 ;
        RECT 251.700 916.050 252.900 929.400 ;
        RECT 273.000 929.100 273.900 929.400 ;
        RECT 278.100 929.400 279.900 935.400 ;
        RECT 281.100 929.400 282.900 936.000 ;
        RECT 296.100 929.400 297.900 935.400 ;
        RECT 299.100 930.000 300.900 936.000 ;
        RECT 278.100 929.100 279.600 929.400 ;
        RECT 273.000 928.200 279.600 929.100 ;
        RECT 297.000 929.100 297.900 929.400 ;
        RECT 302.100 929.400 303.900 935.400 ;
        RECT 305.100 929.400 306.900 936.000 ;
        RECT 320.100 929.400 321.900 936.000 ;
        RECT 323.100 929.400 324.900 935.400 ;
        RECT 326.100 929.400 327.900 936.000 ;
        RECT 344.100 929.400 345.900 935.400 ;
        RECT 347.100 929.400 348.900 936.000 ;
        RECT 362.700 929.400 364.500 936.000 ;
        RECT 302.100 929.100 303.600 929.400 ;
        RECT 297.000 928.200 303.600 929.100 ;
        RECT 254.100 916.050 255.900 917.850 ;
        RECT 273.000 916.050 273.900 928.200 ;
        RECT 278.100 916.050 279.900 917.850 ;
        RECT 297.000 916.050 297.900 928.200 ;
        RECT 302.100 916.050 303.900 917.850 ;
        RECT 323.700 916.050 324.900 929.400 ;
        RECT 344.700 916.050 345.900 929.400 ;
        RECT 363.000 926.100 364.800 927.900 ;
        RECT 365.700 924.900 367.500 935.400 ;
        RECT 365.100 923.400 367.500 924.900 ;
        RECT 370.800 923.400 372.600 936.000 ;
        RECT 386.700 929.400 388.500 936.000 ;
        RECT 387.000 926.100 388.800 927.900 ;
        RECT 389.700 924.900 391.500 935.400 ;
        RECT 389.100 923.400 391.500 924.900 ;
        RECT 394.800 923.400 396.600 936.000 ;
        RECT 410.100 929.400 411.900 936.000 ;
        RECT 413.100 929.400 414.900 935.400 ;
        RECT 428.100 929.400 429.900 936.000 ;
        RECT 431.100 929.400 432.900 935.400 ;
        RECT 347.100 916.050 348.900 917.850 ;
        RECT 365.100 916.050 366.300 923.400 ;
        RECT 371.100 916.050 372.900 917.850 ;
        RECT 389.100 916.050 390.300 923.400 ;
        RECT 395.100 916.050 396.900 917.850 ;
        RECT 410.100 916.050 411.900 917.850 ;
        RECT 413.100 916.050 414.300 929.400 ;
        RECT 428.100 916.050 429.900 917.850 ;
        RECT 431.100 916.050 432.300 929.400 ;
        RECT 446.100 924.300 447.900 935.400 ;
        RECT 449.100 925.200 450.900 936.000 ;
        RECT 452.100 924.300 453.900 935.400 ;
        RECT 446.100 923.400 453.900 924.300 ;
        RECT 455.100 923.400 456.900 935.400 ;
        RECT 473.100 929.400 474.900 936.000 ;
        RECT 476.100 929.400 477.900 935.400 ;
        RECT 479.100 930.000 480.900 936.000 ;
        RECT 476.400 929.100 477.900 929.400 ;
        RECT 482.100 929.400 483.900 935.400 ;
        RECT 497.700 929.400 499.500 936.000 ;
        RECT 482.100 929.100 483.000 929.400 ;
        RECT 476.400 928.200 483.000 929.100 ;
        RECT 449.250 916.050 451.050 917.850 ;
        RECT 455.700 916.050 456.600 923.400 ;
        RECT 460.950 921.450 463.050 922.050 ;
        RECT 475.950 921.450 478.050 925.050 ;
        RECT 460.950 921.000 478.050 921.450 ;
        RECT 460.950 920.550 477.450 921.000 ;
        RECT 460.950 919.950 463.050 920.550 ;
        RECT 476.100 916.050 477.900 917.850 ;
        RECT 482.100 916.050 483.000 928.200 ;
        RECT 498.000 926.100 499.800 927.900 ;
        RECT 500.700 924.900 502.500 935.400 ;
        RECT 500.100 923.400 502.500 924.900 ;
        RECT 505.800 923.400 507.600 936.000 ;
        RECT 524.100 929.400 525.900 935.400 ;
        RECT 527.100 929.400 528.900 936.000 ;
        RECT 500.100 916.050 501.300 923.400 ;
        RECT 506.100 916.050 507.900 917.850 ;
        RECT 524.700 916.050 525.900 929.400 ;
        RECT 542.100 923.400 543.900 935.400 ;
        RECT 545.100 924.300 546.900 935.400 ;
        RECT 548.100 925.200 549.900 936.000 ;
        RECT 551.100 924.300 552.900 935.400 ;
        RECT 569.100 929.400 570.900 936.000 ;
        RECT 572.100 929.400 573.900 935.400 ;
        RECT 575.100 929.400 576.900 936.000 ;
        RECT 590.100 929.400 591.900 935.400 ;
        RECT 593.100 930.000 594.900 936.000 ;
        RECT 562.950 927.450 565.050 928.050 ;
        RECT 568.950 927.450 571.050 928.050 ;
        RECT 562.950 926.550 571.050 927.450 ;
        RECT 562.950 925.950 565.050 926.550 ;
        RECT 568.950 925.950 571.050 926.550 ;
        RECT 545.100 923.400 552.900 924.300 ;
        RECT 527.100 916.050 528.900 917.850 ;
        RECT 542.400 916.050 543.300 923.400 ;
        RECT 564.000 918.450 568.050 919.050 ;
        RECT 547.950 916.050 549.750 917.850 ;
        RECT 563.550 916.950 568.050 918.450 ;
        RECT 16.950 913.950 19.050 916.050 ;
        RECT 19.950 913.950 22.050 916.050 ;
        RECT 22.950 913.950 25.050 916.050 ;
        RECT 25.950 913.950 28.050 916.050 ;
        RECT 43.950 913.950 46.050 916.050 ;
        RECT 46.950 913.950 49.050 916.050 ;
        RECT 49.950 913.950 52.050 916.050 ;
        RECT 52.950 913.950 55.050 916.050 ;
        RECT 67.950 913.950 70.050 916.050 ;
        RECT 70.950 913.950 73.050 916.050 ;
        RECT 73.950 913.950 76.050 916.050 ;
        RECT 88.950 913.950 91.050 916.050 ;
        RECT 91.950 913.950 94.050 916.050 ;
        RECT 109.950 913.950 112.050 916.050 ;
        RECT 112.950 913.950 115.050 916.050 ;
        RECT 115.950 913.950 118.050 916.050 ;
        RECT 118.950 913.950 121.050 916.050 ;
        RECT 133.950 913.950 136.050 916.050 ;
        RECT 136.950 913.950 139.050 916.050 ;
        RECT 139.950 913.950 142.050 916.050 ;
        RECT 142.950 913.950 145.050 916.050 ;
        RECT 157.950 913.950 160.050 916.050 ;
        RECT 160.950 913.950 163.050 916.050 ;
        RECT 163.950 913.950 166.050 916.050 ;
        RECT 178.950 913.950 181.050 916.050 ;
        RECT 181.950 913.950 184.050 916.050 ;
        RECT 184.950 913.950 187.050 916.050 ;
        RECT 187.950 913.950 190.050 916.050 ;
        RECT 202.950 913.950 205.050 916.050 ;
        RECT 205.950 913.950 208.050 916.050 ;
        RECT 208.950 913.950 211.050 916.050 ;
        RECT 211.950 913.950 214.050 916.050 ;
        RECT 226.950 913.950 229.050 916.050 ;
        RECT 229.950 913.950 232.050 916.050 ;
        RECT 232.950 913.950 235.050 916.050 ;
        RECT 235.950 913.950 238.050 916.050 ;
        RECT 250.950 913.950 253.050 916.050 ;
        RECT 253.950 913.950 256.050 916.050 ;
        RECT 271.950 913.950 274.050 916.050 ;
        RECT 274.950 913.950 277.050 916.050 ;
        RECT 277.950 913.950 280.050 916.050 ;
        RECT 280.950 913.950 283.050 916.050 ;
        RECT 295.950 913.950 298.050 916.050 ;
        RECT 298.950 913.950 301.050 916.050 ;
        RECT 301.950 913.950 304.050 916.050 ;
        RECT 304.950 913.950 307.050 916.050 ;
        RECT 319.950 913.950 322.050 916.050 ;
        RECT 322.950 913.950 325.050 916.050 ;
        RECT 325.950 913.950 328.050 916.050 ;
        RECT 343.950 913.950 346.050 916.050 ;
        RECT 346.950 913.950 349.050 916.050 ;
        RECT 361.950 913.950 364.050 916.050 ;
        RECT 364.950 913.950 367.050 916.050 ;
        RECT 367.950 913.950 370.050 916.050 ;
        RECT 370.950 913.950 373.050 916.050 ;
        RECT 385.950 913.950 388.050 916.050 ;
        RECT 388.950 913.950 391.050 916.050 ;
        RECT 391.950 913.950 394.050 916.050 ;
        RECT 394.950 913.950 397.050 916.050 ;
        RECT 409.950 913.950 412.050 916.050 ;
        RECT 412.950 913.950 415.050 916.050 ;
        RECT 427.950 913.950 430.050 916.050 ;
        RECT 430.950 913.950 433.050 916.050 ;
        RECT 445.950 913.950 448.050 916.050 ;
        RECT 448.950 913.950 451.050 916.050 ;
        RECT 451.950 913.950 454.050 916.050 ;
        RECT 454.950 913.950 457.050 916.050 ;
        RECT 472.950 913.950 475.050 916.050 ;
        RECT 475.950 913.950 478.050 916.050 ;
        RECT 478.950 913.950 481.050 916.050 ;
        RECT 481.950 913.950 484.050 916.050 ;
        RECT 496.950 913.950 499.050 916.050 ;
        RECT 499.950 913.950 502.050 916.050 ;
        RECT 502.950 913.950 505.050 916.050 ;
        RECT 505.950 913.950 508.050 916.050 ;
        RECT 523.950 913.950 526.050 916.050 ;
        RECT 526.950 913.950 529.050 916.050 ;
        RECT 541.950 913.950 544.050 916.050 ;
        RECT 544.950 913.950 547.050 916.050 ;
        RECT 547.950 913.950 550.050 916.050 ;
        RECT 550.950 913.950 553.050 916.050 ;
        RECT 20.100 912.150 21.900 913.950 ;
        RECT 23.700 909.600 24.900 913.950 ;
        RECT 26.100 912.150 27.900 913.950 ;
        RECT 44.100 912.150 45.900 913.950 ;
        RECT 50.100 912.150 51.900 913.950 ;
        RECT 53.100 910.200 54.000 913.950 ;
        RECT 68.250 912.150 70.050 913.950 ;
        RECT 23.700 908.700 27.300 909.600 ;
        RECT 17.100 905.700 24.900 907.050 ;
        RECT 17.100 900.600 18.900 905.700 ;
        RECT 20.100 900.000 21.900 904.800 ;
        RECT 23.100 900.600 24.900 905.700 ;
        RECT 26.100 906.600 27.300 908.700 ;
        RECT 26.100 900.600 27.900 906.600 ;
        RECT 44.100 900.000 45.900 909.600 ;
        RECT 50.700 909.000 54.000 910.200 ;
        RECT 50.700 900.600 52.500 909.000 ;
        RECT 71.100 908.700 72.300 913.950 ;
        RECT 74.100 912.150 75.900 913.950 ;
        RECT 71.100 907.800 75.300 908.700 ;
        RECT 68.400 900.000 70.200 906.600 ;
        RECT 73.500 900.600 75.300 907.800 ;
        RECT 89.700 903.600 90.900 913.950 ;
        RECT 110.100 912.150 111.900 913.950 ;
        RECT 116.100 912.150 117.900 913.950 ;
        RECT 119.100 910.200 120.000 913.950 ;
        RECT 134.100 912.150 135.900 913.950 ;
        RECT 140.250 912.150 142.050 913.950 ;
        RECT 89.100 900.600 90.900 903.600 ;
        RECT 92.100 900.000 93.900 903.600 ;
        RECT 110.100 900.000 111.900 909.600 ;
        RECT 116.700 909.000 120.000 910.200 ;
        RECT 121.950 909.450 124.050 910.050 ;
        RECT 139.950 909.450 142.050 910.050 ;
        RECT 116.700 900.600 118.500 909.000 ;
        RECT 121.950 908.550 142.050 909.450 ;
        RECT 121.950 907.950 124.050 908.550 ;
        RECT 139.950 907.950 142.050 908.550 ;
        RECT 143.700 906.600 144.600 913.950 ;
        RECT 158.100 912.150 159.900 913.950 ;
        RECT 161.700 908.700 162.900 913.950 ;
        RECT 163.950 912.150 165.750 913.950 ;
        RECT 179.100 912.150 180.900 913.950 ;
        RECT 185.100 912.150 186.900 913.950 ;
        RECT 188.100 910.200 189.000 913.950 ;
        RECT 206.100 912.150 207.900 913.950 ;
        RECT 135.000 900.000 136.800 906.600 ;
        RECT 139.500 905.400 144.600 906.600 ;
        RECT 158.700 907.800 162.900 908.700 ;
        RECT 139.500 900.600 141.300 905.400 ;
        RECT 142.500 900.000 144.300 903.600 ;
        RECT 158.700 900.600 160.500 907.800 ;
        RECT 163.800 900.000 165.600 906.600 ;
        RECT 179.100 900.000 180.900 909.600 ;
        RECT 185.700 909.000 189.000 910.200 ;
        RECT 209.700 909.600 210.900 913.950 ;
        RECT 212.100 912.150 213.900 913.950 ;
        RECT 230.100 912.150 231.900 913.950 ;
        RECT 233.700 909.600 234.900 913.950 ;
        RECT 236.100 912.150 237.900 913.950 ;
        RECT 185.700 900.600 187.500 909.000 ;
        RECT 209.700 908.700 213.300 909.600 ;
        RECT 233.700 908.700 237.300 909.600 ;
        RECT 203.100 905.700 210.900 907.050 ;
        RECT 203.100 900.600 204.900 905.700 ;
        RECT 206.100 900.000 207.900 904.800 ;
        RECT 209.100 900.600 210.900 905.700 ;
        RECT 212.100 906.600 213.300 908.700 ;
        RECT 212.100 900.600 213.900 906.600 ;
        RECT 227.100 905.700 234.900 907.050 ;
        RECT 227.100 900.600 228.900 905.700 ;
        RECT 230.100 900.000 231.900 904.800 ;
        RECT 233.100 900.600 234.900 905.700 ;
        RECT 236.100 906.600 237.300 908.700 ;
        RECT 236.100 900.600 237.900 906.600 ;
        RECT 251.700 903.600 252.900 913.950 ;
        RECT 273.000 910.200 273.900 913.950 ;
        RECT 275.100 912.150 276.900 913.950 ;
        RECT 281.100 912.150 282.900 913.950 ;
        RECT 297.000 910.200 297.900 913.950 ;
        RECT 299.100 912.150 300.900 913.950 ;
        RECT 305.100 912.150 306.900 913.950 ;
        RECT 320.100 912.150 321.900 913.950 ;
        RECT 273.000 909.000 276.300 910.200 ;
        RECT 251.100 900.600 252.900 903.600 ;
        RECT 254.100 900.000 255.900 903.600 ;
        RECT 274.500 900.600 276.300 909.000 ;
        RECT 281.100 900.000 282.900 909.600 ;
        RECT 297.000 909.000 300.300 910.200 ;
        RECT 298.500 900.600 300.300 909.000 ;
        RECT 305.100 900.000 306.900 909.600 ;
        RECT 323.700 908.700 324.900 913.950 ;
        RECT 325.950 912.150 327.750 913.950 ;
        RECT 320.700 907.800 324.900 908.700 ;
        RECT 320.700 900.600 322.500 907.800 ;
        RECT 325.800 900.000 327.600 906.600 ;
        RECT 344.700 903.600 345.900 913.950 ;
        RECT 362.100 912.150 363.900 913.950 ;
        RECT 365.100 909.600 366.300 913.950 ;
        RECT 368.100 912.150 369.900 913.950 ;
        RECT 386.100 912.150 387.900 913.950 ;
        RECT 389.100 909.600 390.300 913.950 ;
        RECT 392.100 912.150 393.900 913.950 ;
        RECT 362.700 908.700 366.300 909.600 ;
        RECT 386.700 908.700 390.300 909.600 ;
        RECT 362.700 906.600 363.900 908.700 ;
        RECT 344.100 900.600 345.900 903.600 ;
        RECT 347.100 900.000 348.900 903.600 ;
        RECT 362.100 900.600 363.900 906.600 ;
        RECT 365.100 905.700 372.900 907.050 ;
        RECT 386.700 906.600 387.900 908.700 ;
        RECT 365.100 900.600 366.900 905.700 ;
        RECT 368.100 900.000 369.900 904.800 ;
        RECT 371.100 900.600 372.900 905.700 ;
        RECT 386.100 900.600 387.900 906.600 ;
        RECT 389.100 905.700 396.900 907.050 ;
        RECT 389.100 900.600 390.900 905.700 ;
        RECT 392.100 900.000 393.900 904.800 ;
        RECT 395.100 900.600 396.900 905.700 ;
        RECT 413.100 903.600 414.300 913.950 ;
        RECT 431.100 903.600 432.300 913.950 ;
        RECT 446.100 912.150 447.900 913.950 ;
        RECT 452.250 912.150 454.050 913.950 ;
        RECT 455.700 906.600 456.600 913.950 ;
        RECT 473.100 912.150 474.900 913.950 ;
        RECT 479.100 912.150 480.900 913.950 ;
        RECT 482.100 910.200 483.000 913.950 ;
        RECT 497.100 912.150 498.900 913.950 ;
        RECT 410.100 900.000 411.900 903.600 ;
        RECT 413.100 900.600 414.900 903.600 ;
        RECT 428.100 900.000 429.900 903.600 ;
        RECT 431.100 900.600 432.900 903.600 ;
        RECT 447.000 900.000 448.800 906.600 ;
        RECT 451.500 905.400 456.600 906.600 ;
        RECT 451.500 900.600 453.300 905.400 ;
        RECT 454.500 900.000 456.300 903.600 ;
        RECT 473.100 900.000 474.900 909.600 ;
        RECT 479.700 909.000 483.000 910.200 ;
        RECT 500.100 909.600 501.300 913.950 ;
        RECT 503.100 912.150 504.900 913.950 ;
        RECT 479.700 900.600 481.500 909.000 ;
        RECT 497.700 908.700 501.300 909.600 ;
        RECT 497.700 906.600 498.900 908.700 ;
        RECT 497.100 900.600 498.900 906.600 ;
        RECT 500.100 905.700 507.900 907.050 ;
        RECT 500.100 900.600 501.900 905.700 ;
        RECT 503.100 900.000 504.900 904.800 ;
        RECT 506.100 900.600 507.900 905.700 ;
        RECT 524.700 903.600 525.900 913.950 ;
        RECT 542.400 906.600 543.300 913.950 ;
        RECT 544.950 912.150 546.750 913.950 ;
        RECT 551.100 912.150 552.900 913.950 ;
        RECT 553.950 912.450 556.050 913.050 ;
        RECT 563.550 912.450 564.450 916.950 ;
        RECT 572.100 916.050 573.300 929.400 ;
        RECT 591.000 929.100 591.900 929.400 ;
        RECT 596.100 929.400 597.900 935.400 ;
        RECT 599.100 929.400 600.900 936.000 ;
        RECT 596.100 929.100 597.600 929.400 ;
        RECT 591.000 928.200 597.600 929.100 ;
        RECT 591.000 916.050 591.900 928.200 ;
        RECT 614.100 923.400 615.900 935.400 ;
        RECT 617.100 924.000 618.900 936.000 ;
        RECT 620.100 929.400 621.900 935.400 ;
        RECT 623.100 929.400 624.900 936.000 ;
        RECT 596.100 916.050 597.900 917.850 ;
        RECT 614.700 916.050 615.600 923.400 ;
        RECT 618.000 916.050 619.800 917.850 ;
        RECT 568.950 913.950 571.050 916.050 ;
        RECT 571.950 913.950 574.050 916.050 ;
        RECT 574.950 913.950 577.050 916.050 ;
        RECT 589.950 913.950 592.050 916.050 ;
        RECT 592.950 913.950 595.050 916.050 ;
        RECT 595.950 913.950 598.050 916.050 ;
        RECT 598.950 913.950 601.050 916.050 ;
        RECT 614.100 913.950 616.200 916.050 ;
        RECT 617.400 913.950 619.500 916.050 ;
        RECT 553.950 911.550 564.450 912.450 ;
        RECT 569.250 912.150 571.050 913.950 ;
        RECT 553.950 910.950 556.050 911.550 ;
        RECT 572.100 908.700 573.300 913.950 ;
        RECT 575.100 912.150 576.900 913.950 ;
        RECT 591.000 910.200 591.900 913.950 ;
        RECT 593.100 912.150 594.900 913.950 ;
        RECT 599.100 912.150 600.900 913.950 ;
        RECT 591.000 909.000 594.300 910.200 ;
        RECT 572.100 907.800 576.300 908.700 ;
        RECT 542.400 905.400 547.500 906.600 ;
        RECT 524.100 900.600 525.900 903.600 ;
        RECT 527.100 900.000 528.900 903.600 ;
        RECT 542.700 900.000 544.500 903.600 ;
        RECT 545.700 900.600 547.500 905.400 ;
        RECT 550.200 900.000 552.000 906.600 ;
        RECT 569.400 900.000 571.200 906.600 ;
        RECT 574.500 900.600 576.300 907.800 ;
        RECT 592.500 900.600 594.300 909.000 ;
        RECT 599.100 900.000 600.900 909.600 ;
        RECT 614.700 906.600 615.600 913.950 ;
        RECT 621.000 909.300 621.900 929.400 ;
        RECT 641.100 924.300 642.900 935.400 ;
        RECT 644.100 925.200 645.900 936.000 ;
        RECT 647.100 924.300 648.900 935.400 ;
        RECT 641.100 923.400 648.900 924.300 ;
        RECT 650.100 923.400 651.900 935.400 ;
        RECT 665.100 923.400 666.900 935.400 ;
        RECT 668.100 924.300 669.900 935.400 ;
        RECT 671.100 925.200 672.900 936.000 ;
        RECT 674.100 924.300 675.900 935.400 ;
        RECT 692.100 929.400 693.900 935.400 ;
        RECT 695.100 929.400 696.900 936.000 ;
        RECT 668.100 923.400 675.900 924.300 ;
        RECT 644.250 916.050 646.050 917.850 ;
        RECT 650.700 916.050 651.600 923.400 ;
        RECT 665.400 916.050 666.300 923.400 ;
        RECT 670.950 916.050 672.750 917.850 ;
        RECT 692.700 916.050 693.900 929.400 ;
        RECT 710.400 923.400 712.200 936.000 ;
        RECT 715.500 924.900 717.300 935.400 ;
        RECT 718.500 929.400 720.300 936.000 ;
        RECT 718.200 926.100 720.000 927.900 ;
        RECT 715.500 923.400 717.900 924.900 ;
        RECT 734.400 923.400 736.200 936.000 ;
        RECT 739.500 924.900 741.300 935.400 ;
        RECT 742.500 929.400 744.300 936.000 ;
        RECT 758.100 929.400 759.900 935.400 ;
        RECT 761.100 929.400 762.900 936.000 ;
        RECT 742.200 926.100 744.000 927.900 ;
        RECT 739.500 923.400 741.900 924.900 ;
        RECT 695.100 916.050 696.900 917.850 ;
        RECT 710.100 916.050 711.900 917.850 ;
        RECT 716.700 916.050 717.900 923.400 ;
        RECT 718.950 921.450 721.050 922.050 ;
        RECT 733.950 921.450 736.050 922.050 ;
        RECT 718.950 920.550 736.050 921.450 ;
        RECT 718.950 919.950 721.050 920.550 ;
        RECT 733.950 919.950 736.050 920.550 ;
        RECT 734.100 916.050 735.900 917.850 ;
        RECT 740.700 916.050 741.900 923.400 ;
        RECT 758.700 916.050 759.900 929.400 ;
        RECT 776.100 924.300 777.900 935.400 ;
        RECT 779.100 925.200 780.900 936.000 ;
        RECT 782.100 924.300 783.900 935.400 ;
        RECT 776.100 923.400 783.900 924.300 ;
        RECT 785.100 923.400 786.900 935.400 ;
        RECT 803.400 923.400 805.200 936.000 ;
        RECT 808.500 924.900 810.300 935.400 ;
        RECT 811.500 929.400 813.300 936.000 ;
        RECT 830.100 929.400 831.900 936.000 ;
        RECT 833.100 929.400 834.900 935.400 ;
        RECT 836.100 929.400 837.900 936.000 ;
        RECT 851.100 929.400 852.900 936.000 ;
        RECT 854.100 929.400 855.900 935.400 ;
        RECT 857.100 929.400 858.900 936.000 ;
        RECT 811.200 926.100 813.000 927.900 ;
        RECT 808.500 923.400 810.900 924.900 ;
        RECT 761.100 916.050 762.900 917.850 ;
        RECT 779.250 916.050 781.050 917.850 ;
        RECT 785.700 916.050 786.600 923.400 ;
        RECT 803.100 916.050 804.900 917.850 ;
        RECT 809.700 916.050 810.900 923.400 ;
        RECT 833.100 916.050 834.300 929.400 ;
        RECT 854.100 916.050 855.300 929.400 ;
        RECT 872.400 923.400 874.200 936.000 ;
        RECT 877.500 924.900 879.300 935.400 ;
        RECT 880.500 929.400 882.300 936.000 ;
        RECT 880.200 926.100 882.000 927.900 ;
        RECT 877.500 923.400 879.900 924.900 ;
        RECT 896.100 923.400 897.900 935.400 ;
        RECT 899.100 924.300 900.900 935.400 ;
        RECT 902.100 925.200 903.900 936.000 ;
        RECT 905.100 924.300 906.900 935.400 ;
        RECT 923.100 929.400 924.900 936.000 ;
        RECT 926.100 929.400 927.900 935.400 ;
        RECT 899.100 923.400 906.900 924.300 ;
        RECT 862.950 921.450 865.050 922.050 ;
        RECT 874.950 921.450 877.050 922.050 ;
        RECT 862.950 920.550 877.050 921.450 ;
        RECT 862.950 919.950 865.050 920.550 ;
        RECT 874.950 919.950 877.050 920.550 ;
        RECT 872.100 916.050 873.900 917.850 ;
        RECT 878.700 916.050 879.900 923.400 ;
        RECT 896.400 916.050 897.300 923.400 ;
        RECT 904.950 921.450 907.050 922.050 ;
        RECT 922.950 921.450 925.050 922.200 ;
        RECT 904.950 920.550 925.050 921.450 ;
        RECT 904.950 919.950 907.050 920.550 ;
        RECT 922.950 920.100 925.050 920.550 ;
        RECT 901.950 916.050 903.750 917.850 ;
        RECT 622.800 913.950 624.900 916.050 ;
        RECT 640.950 913.950 643.050 916.050 ;
        RECT 643.950 913.950 646.050 916.050 ;
        RECT 646.950 913.950 649.050 916.050 ;
        RECT 649.950 913.950 652.050 916.050 ;
        RECT 664.950 913.950 667.050 916.050 ;
        RECT 667.950 913.950 670.050 916.050 ;
        RECT 670.950 913.950 673.050 916.050 ;
        RECT 673.950 913.950 676.050 916.050 ;
        RECT 691.950 913.950 694.050 916.050 ;
        RECT 694.950 913.950 697.050 916.050 ;
        RECT 709.950 913.950 712.050 916.050 ;
        RECT 712.950 913.950 715.050 916.050 ;
        RECT 715.950 913.950 718.050 916.050 ;
        RECT 718.950 913.950 721.050 916.050 ;
        RECT 733.950 913.950 736.050 916.050 ;
        RECT 736.950 913.950 739.050 916.050 ;
        RECT 739.950 913.950 742.050 916.050 ;
        RECT 742.950 913.950 745.050 916.050 ;
        RECT 757.950 913.950 760.050 916.050 ;
        RECT 760.950 913.950 763.050 916.050 ;
        RECT 775.950 913.950 778.050 916.050 ;
        RECT 778.950 913.950 781.050 916.050 ;
        RECT 781.950 913.950 784.050 916.050 ;
        RECT 784.950 913.950 787.050 916.050 ;
        RECT 802.950 913.950 805.050 916.050 ;
        RECT 805.950 913.950 808.050 916.050 ;
        RECT 808.950 913.950 811.050 916.050 ;
        RECT 811.950 913.950 814.050 916.050 ;
        RECT 829.950 913.950 832.050 916.050 ;
        RECT 832.950 913.950 835.050 916.050 ;
        RECT 835.950 913.950 838.050 916.050 ;
        RECT 850.950 913.950 853.050 916.050 ;
        RECT 853.950 913.950 856.050 916.050 ;
        RECT 856.950 913.950 859.050 916.050 ;
        RECT 871.950 913.950 874.050 916.050 ;
        RECT 874.950 913.950 877.050 916.050 ;
        RECT 877.950 913.950 880.050 916.050 ;
        RECT 880.950 913.950 883.050 916.050 ;
        RECT 895.950 913.950 898.050 916.050 ;
        RECT 898.950 913.950 901.050 916.050 ;
        RECT 901.950 913.950 904.050 916.050 ;
        RECT 904.950 913.950 907.050 916.050 ;
        RECT 923.100 913.950 925.200 916.050 ;
        RECT 622.950 912.150 624.750 913.950 ;
        RECT 641.100 912.150 642.900 913.950 ;
        RECT 647.250 912.150 649.050 913.950 ;
        RECT 616.500 908.400 624.900 909.300 ;
        RECT 616.500 907.500 618.300 908.400 ;
        RECT 614.700 904.800 617.400 906.600 ;
        RECT 615.600 900.600 617.400 904.800 ;
        RECT 618.600 900.000 620.400 906.600 ;
        RECT 623.100 900.600 624.900 908.400 ;
        RECT 650.700 906.600 651.600 913.950 ;
        RECT 642.000 900.000 643.800 906.600 ;
        RECT 646.500 905.400 651.600 906.600 ;
        RECT 665.400 906.600 666.300 913.950 ;
        RECT 667.950 912.150 669.750 913.950 ;
        RECT 674.100 912.150 675.900 913.950 ;
        RECT 665.400 905.400 670.500 906.600 ;
        RECT 646.500 900.600 648.300 905.400 ;
        RECT 649.500 900.000 651.300 903.600 ;
        RECT 665.700 900.000 667.500 903.600 ;
        RECT 668.700 900.600 670.500 905.400 ;
        RECT 673.200 900.000 675.000 906.600 ;
        RECT 692.700 903.600 693.900 913.950 ;
        RECT 713.100 912.150 714.900 913.950 ;
        RECT 716.700 909.600 717.900 913.950 ;
        RECT 719.100 912.150 720.900 913.950 ;
        RECT 737.100 912.150 738.900 913.950 ;
        RECT 740.700 909.600 741.900 913.950 ;
        RECT 743.100 912.150 744.900 913.950 ;
        RECT 716.700 908.700 720.300 909.600 ;
        RECT 740.700 908.700 744.300 909.600 ;
        RECT 710.100 905.700 717.900 907.050 ;
        RECT 692.100 900.600 693.900 903.600 ;
        RECT 695.100 900.000 696.900 903.600 ;
        RECT 710.100 900.600 711.900 905.700 ;
        RECT 713.100 900.000 714.900 904.800 ;
        RECT 716.100 900.600 717.900 905.700 ;
        RECT 719.100 906.600 720.300 908.700 ;
        RECT 719.100 900.600 720.900 906.600 ;
        RECT 734.100 905.700 741.900 907.050 ;
        RECT 734.100 900.600 735.900 905.700 ;
        RECT 737.100 900.000 738.900 904.800 ;
        RECT 740.100 900.600 741.900 905.700 ;
        RECT 743.100 906.600 744.300 908.700 ;
        RECT 743.100 900.600 744.900 906.600 ;
        RECT 758.700 903.600 759.900 913.950 ;
        RECT 776.100 912.150 777.900 913.950 ;
        RECT 782.250 912.150 784.050 913.950 ;
        RECT 785.700 906.600 786.600 913.950 ;
        RECT 806.100 912.150 807.900 913.950 ;
        RECT 809.700 909.600 810.900 913.950 ;
        RECT 812.100 912.150 813.900 913.950 ;
        RECT 830.250 912.150 832.050 913.950 ;
        RECT 809.700 908.700 813.300 909.600 ;
        RECT 758.100 900.600 759.900 903.600 ;
        RECT 761.100 900.000 762.900 903.600 ;
        RECT 777.000 900.000 778.800 906.600 ;
        RECT 781.500 905.400 786.600 906.600 ;
        RECT 803.100 905.700 810.900 907.050 ;
        RECT 781.500 900.600 783.300 905.400 ;
        RECT 784.500 900.000 786.300 903.600 ;
        RECT 803.100 900.600 804.900 905.700 ;
        RECT 806.100 900.000 807.900 904.800 ;
        RECT 809.100 900.600 810.900 905.700 ;
        RECT 812.100 906.600 813.300 908.700 ;
        RECT 833.100 908.700 834.300 913.950 ;
        RECT 836.100 912.150 837.900 913.950 ;
        RECT 851.250 912.150 853.050 913.950 ;
        RECT 854.100 908.700 855.300 913.950 ;
        RECT 857.100 912.150 858.900 913.950 ;
        RECT 875.100 912.150 876.900 913.950 ;
        RECT 878.700 909.600 879.900 913.950 ;
        RECT 881.100 912.150 882.900 913.950 ;
        RECT 878.700 908.700 882.300 909.600 ;
        RECT 833.100 907.800 837.300 908.700 ;
        RECT 854.100 907.800 858.300 908.700 ;
        RECT 812.100 900.600 813.900 906.600 ;
        RECT 830.400 900.000 832.200 906.600 ;
        RECT 835.500 900.600 837.300 907.800 ;
        RECT 851.400 900.000 853.200 906.600 ;
        RECT 856.500 900.600 858.300 907.800 ;
        RECT 872.100 905.700 879.900 907.050 ;
        RECT 872.100 900.600 873.900 905.700 ;
        RECT 875.100 900.000 876.900 904.800 ;
        RECT 878.100 900.600 879.900 905.700 ;
        RECT 881.100 906.600 882.300 908.700 ;
        RECT 896.400 906.600 897.300 913.950 ;
        RECT 898.950 912.150 900.750 913.950 ;
        RECT 905.100 912.150 906.900 913.950 ;
        RECT 923.250 912.150 925.050 913.950 ;
        RECT 926.100 909.300 927.000 929.400 ;
        RECT 929.100 924.000 930.900 936.000 ;
        RECT 932.100 923.400 933.900 935.400 ;
        RECT 950.100 929.400 951.900 936.000 ;
        RECT 953.100 929.400 954.900 935.400 ;
        RECT 956.100 930.000 957.900 936.000 ;
        RECT 953.400 929.100 954.900 929.400 ;
        RECT 959.100 929.400 960.900 935.400 ;
        RECT 959.100 929.100 960.000 929.400 ;
        RECT 953.400 928.200 960.000 929.100 ;
        RECT 928.200 916.050 930.000 917.850 ;
        RECT 932.400 916.050 933.300 923.400 ;
        RECT 934.950 921.450 937.050 922.050 ;
        RECT 955.950 921.450 958.050 922.050 ;
        RECT 934.950 920.550 958.050 921.450 ;
        RECT 934.950 919.950 937.050 920.550 ;
        RECT 955.950 919.950 958.050 920.550 ;
        RECT 953.100 916.050 954.900 917.850 ;
        RECT 959.100 916.050 960.000 928.200 ;
        RECT 974.400 923.400 976.200 936.000 ;
        RECT 979.500 924.900 981.300 935.400 ;
        RECT 982.500 929.400 984.300 936.000 ;
        RECT 982.200 926.100 984.000 927.900 ;
        RECT 979.500 923.400 981.900 924.900 ;
        RECT 1001.100 924.300 1002.900 935.400 ;
        RECT 1004.100 925.200 1005.900 936.000 ;
        RECT 1007.100 924.300 1008.900 935.400 ;
        RECT 1001.100 923.400 1008.900 924.300 ;
        RECT 1010.100 923.400 1011.900 935.400 ;
        RECT 974.100 916.050 975.900 917.850 ;
        RECT 980.700 916.050 981.900 923.400 ;
        RECT 982.950 921.450 985.050 922.050 ;
        RECT 991.950 921.450 994.050 922.050 ;
        RECT 1006.950 921.450 1009.050 922.050 ;
        RECT 982.950 920.550 994.050 921.450 ;
        RECT 982.950 919.950 985.050 920.550 ;
        RECT 991.950 919.950 994.050 920.550 ;
        RECT 998.550 920.550 1009.050 921.450 ;
        RECT 988.950 918.450 991.050 919.050 ;
        RECT 998.550 918.450 999.450 920.550 ;
        RECT 1006.950 919.950 1009.050 920.550 ;
        RECT 988.950 917.550 999.450 918.450 ;
        RECT 988.950 916.950 991.050 917.550 ;
        RECT 1004.250 916.050 1006.050 917.850 ;
        RECT 1010.700 916.050 1011.600 923.400 ;
        RECT 928.500 913.950 930.600 916.050 ;
        RECT 931.800 913.950 933.900 916.050 ;
        RECT 949.950 913.950 952.050 916.050 ;
        RECT 952.950 913.950 955.050 916.050 ;
        RECT 955.950 913.950 958.050 916.050 ;
        RECT 958.950 913.950 961.050 916.050 ;
        RECT 973.950 913.950 976.050 916.050 ;
        RECT 976.950 913.950 979.050 916.050 ;
        RECT 979.950 913.950 982.050 916.050 ;
        RECT 982.950 913.950 985.050 916.050 ;
        RECT 1000.950 913.950 1003.050 916.050 ;
        RECT 1003.950 913.950 1006.050 916.050 ;
        RECT 1006.950 913.950 1009.050 916.050 ;
        RECT 1009.950 913.950 1012.050 916.050 ;
        RECT 923.100 908.400 931.500 909.300 ;
        RECT 881.100 900.600 882.900 906.600 ;
        RECT 896.400 905.400 901.500 906.600 ;
        RECT 896.700 900.000 898.500 903.600 ;
        RECT 899.700 900.600 901.500 905.400 ;
        RECT 904.200 900.000 906.000 906.600 ;
        RECT 923.100 900.600 924.900 908.400 ;
        RECT 929.700 907.500 931.500 908.400 ;
        RECT 932.400 906.600 933.300 913.950 ;
        RECT 950.100 912.150 951.900 913.950 ;
        RECT 956.100 912.150 957.900 913.950 ;
        RECT 959.100 910.200 960.000 913.950 ;
        RECT 977.100 912.150 978.900 913.950 ;
        RECT 927.600 900.000 929.400 906.600 ;
        RECT 930.600 904.800 933.300 906.600 ;
        RECT 930.600 900.600 932.400 904.800 ;
        RECT 950.100 900.000 951.900 909.600 ;
        RECT 956.700 909.000 960.000 910.200 ;
        RECT 980.700 909.600 981.900 913.950 ;
        RECT 983.100 912.150 984.900 913.950 ;
        RECT 1001.100 912.150 1002.900 913.950 ;
        RECT 1007.250 912.150 1009.050 913.950 ;
        RECT 956.700 900.600 958.500 909.000 ;
        RECT 980.700 908.700 984.300 909.600 ;
        RECT 974.100 905.700 981.900 907.050 ;
        RECT 974.100 900.600 975.900 905.700 ;
        RECT 977.100 900.000 978.900 904.800 ;
        RECT 980.100 900.600 981.900 905.700 ;
        RECT 983.100 906.600 984.300 908.700 ;
        RECT 1010.700 906.600 1011.600 913.950 ;
        RECT 983.100 900.600 984.900 906.600 ;
        RECT 1002.000 900.000 1003.800 906.600 ;
        RECT 1006.500 905.400 1011.600 906.600 ;
        RECT 1006.500 900.600 1008.300 905.400 ;
        RECT 1009.500 900.000 1011.300 903.600 ;
        RECT 17.100 890.400 18.900 896.400 ;
        RECT 20.100 891.000 21.900 897.000 ;
        RECT 26.700 896.400 27.900 897.000 ;
        RECT 23.100 893.400 24.900 896.400 ;
        RECT 26.100 893.400 27.900 896.400 ;
        RECT 17.100 883.050 18.000 890.400 ;
        RECT 23.700 889.200 24.600 893.400 ;
        RECT 41.400 890.400 43.200 897.000 ;
        RECT 46.500 889.200 48.300 896.400 ;
        RECT 62.400 890.400 64.200 897.000 ;
        RECT 67.500 889.200 69.300 896.400 ;
        RECT 83.100 890.400 84.900 896.400 ;
        RECT 19.200 888.300 24.600 889.200 ;
        RECT 44.100 888.300 48.300 889.200 ;
        RECT 65.100 888.300 69.300 889.200 ;
        RECT 83.700 888.300 84.900 890.400 ;
        RECT 86.100 891.300 87.900 896.400 ;
        RECT 89.100 892.200 90.900 897.000 ;
        RECT 92.100 891.300 93.900 896.400 ;
        RECT 107.100 893.400 108.900 897.000 ;
        RECT 110.100 893.400 111.900 896.400 ;
        RECT 86.100 889.950 93.900 891.300 ;
        RECT 19.200 887.400 21.300 888.300 ;
        RECT 17.100 880.950 19.200 883.050 ;
        RECT 18.000 873.600 19.200 880.950 ;
        RECT 20.400 876.900 21.300 887.400 ;
        RECT 25.800 883.050 27.600 884.850 ;
        RECT 41.250 883.050 43.050 884.850 ;
        RECT 44.100 883.050 45.300 888.300 ;
        RECT 47.100 883.050 48.900 884.850 ;
        RECT 62.250 883.050 64.050 884.850 ;
        RECT 65.100 883.050 66.300 888.300 ;
        RECT 83.700 887.400 87.300 888.300 ;
        RECT 68.100 883.050 69.900 884.850 ;
        RECT 83.100 883.050 84.900 884.850 ;
        RECT 86.100 883.050 87.300 887.400 ;
        RECT 89.100 883.050 90.900 884.850 ;
        RECT 110.100 883.050 111.300 893.400 ;
        RECT 127.500 888.000 129.300 896.400 ;
        RECT 126.000 886.800 129.300 888.000 ;
        RECT 134.100 887.400 135.900 897.000 ;
        RECT 152.100 890.400 153.900 896.400 ;
        RECT 155.100 891.000 156.900 897.000 ;
        RECT 161.700 896.400 162.900 897.000 ;
        RECT 158.100 893.400 159.900 896.400 ;
        RECT 161.100 893.400 162.900 896.400 ;
        RECT 179.100 893.400 180.900 897.000 ;
        RECT 182.100 893.400 183.900 896.400 ;
        RECT 185.100 893.400 186.900 897.000 ;
        RECT 126.000 883.050 126.900 886.800 ;
        RECT 128.100 883.050 129.900 884.850 ;
        RECT 134.100 883.050 135.900 884.850 ;
        RECT 152.100 883.050 153.000 890.400 ;
        RECT 158.700 889.200 159.600 893.400 ;
        RECT 154.200 888.300 159.600 889.200 ;
        RECT 154.200 887.400 156.300 888.300 ;
        RECT 22.500 880.950 24.600 883.050 ;
        RECT 25.800 880.950 27.900 883.050 ;
        RECT 40.950 880.950 43.050 883.050 ;
        RECT 43.950 880.950 46.050 883.050 ;
        RECT 46.950 880.950 49.050 883.050 ;
        RECT 61.950 880.950 64.050 883.050 ;
        RECT 64.950 880.950 67.050 883.050 ;
        RECT 67.950 880.950 70.050 883.050 ;
        RECT 82.950 880.950 85.050 883.050 ;
        RECT 85.950 880.950 88.050 883.050 ;
        RECT 88.950 880.950 91.050 883.050 ;
        RECT 91.950 880.950 94.050 883.050 ;
        RECT 106.950 880.950 109.050 883.050 ;
        RECT 109.950 880.950 112.050 883.050 ;
        RECT 124.950 880.950 127.050 883.050 ;
        RECT 127.950 880.950 130.050 883.050 ;
        RECT 130.950 880.950 133.050 883.050 ;
        RECT 133.950 880.950 136.050 883.050 ;
        RECT 152.100 880.950 154.200 883.050 ;
        RECT 22.200 879.150 24.000 880.950 ;
        RECT 20.100 876.300 21.900 876.900 ;
        RECT 20.100 875.100 27.900 876.300 ;
        RECT 26.700 873.600 27.900 875.100 ;
        RECT 18.000 872.100 20.400 873.600 ;
        RECT 18.600 861.600 20.400 872.100 ;
        RECT 21.600 861.000 23.400 873.600 ;
        RECT 26.100 861.600 27.900 873.600 ;
        RECT 44.100 867.600 45.300 880.950 ;
        RECT 65.100 867.600 66.300 880.950 ;
        RECT 86.100 873.600 87.300 880.950 ;
        RECT 92.100 879.150 93.900 880.950 ;
        RECT 107.100 879.150 108.900 880.950 ;
        RECT 86.100 872.100 88.500 873.600 ;
        RECT 84.000 869.100 85.800 870.900 ;
        RECT 41.100 861.000 42.900 867.600 ;
        RECT 44.100 861.600 45.900 867.600 ;
        RECT 47.100 861.000 48.900 867.600 ;
        RECT 62.100 861.000 63.900 867.600 ;
        RECT 65.100 861.600 66.900 867.600 ;
        RECT 68.100 861.000 69.900 867.600 ;
        RECT 83.700 861.000 85.500 867.600 ;
        RECT 86.700 861.600 88.500 872.100 ;
        RECT 91.800 861.000 93.600 873.600 ;
        RECT 110.100 867.600 111.300 880.950 ;
        RECT 126.000 868.800 126.900 880.950 ;
        RECT 131.100 879.150 132.900 880.950 ;
        RECT 153.000 873.600 154.200 880.950 ;
        RECT 155.400 876.900 156.300 887.400 ;
        RECT 160.800 883.050 162.600 884.850 ;
        RECT 182.700 883.050 183.600 893.400 ;
        RECT 200.100 890.400 201.900 896.400 ;
        RECT 200.700 888.300 201.900 890.400 ;
        RECT 203.100 891.300 204.900 896.400 ;
        RECT 206.100 892.200 207.900 897.000 ;
        RECT 209.100 891.300 210.900 896.400 ;
        RECT 235.200 893.400 237.900 896.400 ;
        RECT 239.100 893.400 240.900 897.000 ;
        RECT 242.100 893.400 243.900 896.400 ;
        RECT 245.100 893.400 247.200 897.000 ;
        RECT 235.200 892.500 236.100 893.400 ;
        RECT 242.400 892.500 243.300 893.400 ;
        RECT 203.100 889.950 210.900 891.300 ;
        RECT 214.950 891.450 217.050 892.050 ;
        RECT 220.950 891.450 223.050 892.050 ;
        RECT 214.950 890.550 223.050 891.450 ;
        RECT 214.950 889.950 217.050 890.550 ;
        RECT 220.950 889.950 223.050 890.550 ;
        RECT 230.700 891.600 243.300 892.500 ;
        RECT 200.700 887.400 204.300 888.300 ;
        RECT 200.100 883.050 201.900 884.850 ;
        RECT 203.100 883.050 204.300 887.400 ;
        RECT 211.950 885.450 214.050 886.050 ;
        RECT 220.950 885.450 223.050 885.900 ;
        RECT 206.100 883.050 207.900 884.850 ;
        RECT 211.950 884.550 223.050 885.450 ;
        RECT 211.950 883.950 214.050 884.550 ;
        RECT 220.950 883.800 223.050 884.550 ;
        RECT 230.700 883.050 231.900 891.600 ;
        RECT 263.100 891.300 264.900 896.400 ;
        RECT 266.100 892.200 267.900 897.000 ;
        RECT 269.100 891.300 270.900 896.400 ;
        RECT 263.100 889.950 270.900 891.300 ;
        RECT 272.100 890.400 273.900 896.400 ;
        RECT 287.700 893.400 289.500 897.000 ;
        RECT 290.700 891.600 292.500 896.400 ;
        RECT 287.400 890.400 292.500 891.600 ;
        RECT 295.200 890.400 297.000 897.000 ;
        RECT 232.950 888.450 235.050 889.050 ;
        RECT 256.950 888.450 259.050 889.050 ;
        RECT 232.950 887.550 259.050 888.450 ;
        RECT 272.100 888.300 273.300 890.400 ;
        RECT 232.950 886.950 235.050 887.550 ;
        RECT 256.950 886.950 259.050 887.550 ;
        RECT 269.700 887.400 273.300 888.300 ;
        RECT 239.250 883.050 241.050 884.850 ;
        RECT 266.100 883.050 267.900 884.850 ;
        RECT 269.700 883.050 270.900 887.400 ;
        RECT 272.100 883.050 273.900 884.850 ;
        RECT 287.400 883.050 288.300 890.400 ;
        RECT 316.500 888.000 318.300 896.400 ;
        RECT 315.000 886.800 318.300 888.000 ;
        RECT 323.100 887.400 324.900 897.000 ;
        RECT 341.100 891.300 342.900 896.400 ;
        RECT 344.100 892.200 345.900 897.000 ;
        RECT 347.100 891.300 348.900 896.400 ;
        RECT 341.100 889.950 348.900 891.300 ;
        RECT 350.100 890.400 351.900 896.400 ;
        RECT 365.100 893.400 366.900 896.400 ;
        RECT 368.100 893.400 369.900 897.000 ;
        RECT 350.100 888.300 351.300 890.400 ;
        RECT 347.700 887.400 351.300 888.300 ;
        RECT 289.950 883.050 291.750 884.850 ;
        RECT 296.100 883.050 297.900 884.850 ;
        RECT 315.000 883.050 315.900 886.800 ;
        RECT 317.100 883.050 318.900 884.850 ;
        RECT 323.100 883.050 324.900 884.850 ;
        RECT 344.100 883.050 345.900 884.850 ;
        RECT 347.700 883.050 348.900 887.400 ;
        RECT 350.100 883.050 351.900 884.850 ;
        RECT 365.700 883.050 366.900 893.400 ;
        RECT 386.400 890.400 388.200 897.000 ;
        RECT 391.500 889.200 393.300 896.400 ;
        RECT 389.100 888.300 393.300 889.200 ;
        RECT 407.700 889.200 409.500 896.400 ;
        RECT 412.800 890.400 414.600 897.000 ;
        RECT 433.500 890.400 435.300 897.000 ;
        RECT 438.000 890.400 439.800 896.400 ;
        RECT 442.500 890.400 444.300 897.000 ;
        RECT 458.100 891.300 459.900 896.400 ;
        RECT 461.100 892.200 462.900 897.000 ;
        RECT 464.100 891.300 465.900 896.400 ;
        RECT 407.700 888.300 411.900 889.200 ;
        RECT 386.250 883.050 388.050 884.850 ;
        RECT 389.100 883.050 390.300 888.300 ;
        RECT 392.100 883.050 393.900 884.850 ;
        RECT 407.100 883.050 408.900 884.850 ;
        RECT 410.700 883.050 411.900 888.300 ;
        RECT 412.950 883.050 414.750 884.850 ;
        RECT 431.100 883.050 432.900 884.850 ;
        RECT 437.700 883.050 438.900 890.400 ;
        RECT 458.100 889.950 465.900 891.300 ;
        RECT 467.100 890.400 468.900 896.400 ;
        RECT 487.800 893.400 489.900 897.000 ;
        RECT 491.100 893.400 492.900 896.400 ;
        RECT 494.100 893.400 495.900 897.000 ;
        RECT 497.100 893.400 499.800 896.400 ;
        RECT 491.700 892.500 492.600 893.400 ;
        RECT 498.900 892.500 499.800 893.400 ;
        RECT 478.950 891.450 481.050 892.050 ;
        RECT 487.950 891.450 490.050 892.050 ;
        RECT 491.700 891.600 504.300 892.500 ;
        RECT 478.950 890.550 490.050 891.450 ;
        RECT 467.100 888.300 468.300 890.400 ;
        RECT 478.950 889.950 481.050 890.550 ;
        RECT 487.950 889.950 490.050 890.550 ;
        RECT 464.700 887.400 468.300 888.300 ;
        RECT 472.950 888.450 475.050 889.050 ;
        RECT 496.950 888.450 499.050 889.050 ;
        RECT 472.950 887.550 499.050 888.450 ;
        RECT 442.950 883.050 444.750 884.850 ;
        RECT 461.100 883.050 462.900 884.850 ;
        RECT 464.700 883.050 465.900 887.400 ;
        RECT 472.950 886.950 475.050 887.550 ;
        RECT 496.950 886.950 499.050 887.550 ;
        RECT 467.100 883.050 468.900 884.850 ;
        RECT 493.950 883.050 495.750 884.850 ;
        RECT 503.100 883.050 504.300 891.600 ;
        RECT 521.400 890.400 523.200 897.000 ;
        RECT 526.500 889.200 528.300 896.400 ;
        RECT 524.100 888.300 528.300 889.200 ;
        RECT 521.250 883.050 523.050 884.850 ;
        RECT 524.100 883.050 525.300 888.300 ;
        RECT 545.100 887.400 546.900 897.000 ;
        RECT 551.700 888.000 553.500 896.400 ;
        RECT 569.100 890.400 570.900 896.400 ;
        RECT 569.700 888.300 570.900 890.400 ;
        RECT 572.100 891.300 573.900 896.400 ;
        RECT 575.100 892.200 576.900 897.000 ;
        RECT 578.100 891.300 579.900 896.400 ;
        RECT 572.100 889.950 579.900 891.300 ;
        RECT 580.950 891.450 583.050 892.050 ;
        RECT 589.950 891.450 592.050 895.050 ;
        RECT 580.950 891.000 592.050 891.450 ;
        RECT 593.100 891.300 594.900 896.400 ;
        RECT 596.100 892.200 597.900 897.000 ;
        RECT 599.100 891.300 600.900 896.400 ;
        RECT 580.950 890.550 591.450 891.000 ;
        RECT 580.950 889.950 583.050 890.550 ;
        RECT 593.100 889.950 600.900 891.300 ;
        RECT 602.100 890.400 603.900 896.400 ;
        RECT 602.100 888.300 603.300 890.400 ;
        RECT 551.700 886.800 555.000 888.000 ;
        RECT 569.700 887.400 573.300 888.300 ;
        RECT 527.100 883.050 528.900 884.850 ;
        RECT 545.100 883.050 546.900 884.850 ;
        RECT 551.100 883.050 552.900 884.850 ;
        RECT 554.100 883.050 555.000 886.800 ;
        RECT 569.100 883.050 570.900 884.850 ;
        RECT 572.100 883.050 573.300 887.400 ;
        RECT 599.700 887.400 603.300 888.300 ;
        RECT 617.100 887.400 618.900 897.000 ;
        RECT 623.700 888.000 625.500 896.400 ;
        RECT 643.500 888.000 645.300 896.400 ;
        RECT 575.100 883.050 576.900 884.850 ;
        RECT 596.100 883.050 597.900 884.850 ;
        RECT 599.700 883.050 600.900 887.400 ;
        RECT 623.700 886.800 627.000 888.000 ;
        RECT 602.100 883.050 603.900 884.850 ;
        RECT 617.100 883.050 618.900 884.850 ;
        RECT 623.100 883.050 624.900 884.850 ;
        RECT 626.100 883.050 627.000 886.800 ;
        RECT 642.000 886.800 645.300 888.000 ;
        RECT 650.100 887.400 651.900 897.000 ;
        RECT 665.100 893.400 666.900 897.000 ;
        RECT 668.100 893.400 669.900 896.400 ;
        RECT 642.000 883.050 642.900 886.800 ;
        RECT 644.100 883.050 645.900 884.850 ;
        RECT 650.100 883.050 651.900 884.850 ;
        RECT 668.100 883.050 669.300 893.400 ;
        RECT 684.600 892.200 686.400 896.400 ;
        RECT 683.700 890.400 686.400 892.200 ;
        RECT 687.600 890.400 689.400 897.000 ;
        RECT 683.700 883.050 684.600 890.400 ;
        RECT 685.500 888.600 687.300 889.500 ;
        RECT 692.100 888.600 693.900 896.400 ;
        RECT 710.100 890.400 711.900 896.400 ;
        RECT 685.500 887.700 693.900 888.600 ;
        RECT 710.700 888.300 711.900 890.400 ;
        RECT 713.100 891.300 714.900 896.400 ;
        RECT 716.100 892.200 717.900 897.000 ;
        RECT 719.100 891.300 720.900 896.400 ;
        RECT 734.100 893.400 735.900 897.000 ;
        RECT 737.100 893.400 738.900 896.400 ;
        RECT 713.100 889.950 720.900 891.300 ;
        RECT 157.500 880.950 159.600 883.050 ;
        RECT 160.800 880.950 162.900 883.050 ;
        RECT 178.950 880.950 181.050 883.050 ;
        RECT 181.950 880.950 184.050 883.050 ;
        RECT 184.950 880.950 187.050 883.050 ;
        RECT 199.950 880.950 202.050 883.050 ;
        RECT 202.950 880.950 205.050 883.050 ;
        RECT 205.950 880.950 208.050 883.050 ;
        RECT 208.950 880.950 211.050 883.050 ;
        RECT 230.400 880.950 232.500 883.050 ;
        RECT 235.950 880.950 238.050 883.050 ;
        RECT 238.950 880.950 241.050 883.050 ;
        RECT 245.100 880.950 247.200 883.050 ;
        RECT 262.950 880.950 265.050 883.050 ;
        RECT 265.950 880.950 268.050 883.050 ;
        RECT 268.950 880.950 271.050 883.050 ;
        RECT 271.950 880.950 274.050 883.050 ;
        RECT 286.950 880.950 289.050 883.050 ;
        RECT 289.950 880.950 292.050 883.050 ;
        RECT 292.950 880.950 295.050 883.050 ;
        RECT 295.950 880.950 298.050 883.050 ;
        RECT 313.950 880.950 316.050 883.050 ;
        RECT 316.950 880.950 319.050 883.050 ;
        RECT 319.950 880.950 322.050 883.050 ;
        RECT 322.950 880.950 325.050 883.050 ;
        RECT 340.950 880.950 343.050 883.050 ;
        RECT 343.950 880.950 346.050 883.050 ;
        RECT 346.950 880.950 349.050 883.050 ;
        RECT 349.950 880.950 352.050 883.050 ;
        RECT 364.950 880.950 367.050 883.050 ;
        RECT 367.950 880.950 370.050 883.050 ;
        RECT 385.950 880.950 388.050 883.050 ;
        RECT 388.950 880.950 391.050 883.050 ;
        RECT 391.950 880.950 394.050 883.050 ;
        RECT 406.950 880.950 409.050 883.050 ;
        RECT 409.950 880.950 412.050 883.050 ;
        RECT 412.950 880.950 415.050 883.050 ;
        RECT 430.950 880.950 433.050 883.050 ;
        RECT 433.950 880.950 436.050 883.050 ;
        RECT 436.950 880.950 439.050 883.050 ;
        RECT 439.950 880.950 442.050 883.050 ;
        RECT 442.950 880.950 445.050 883.050 ;
        RECT 457.950 880.950 460.050 883.050 ;
        RECT 460.950 880.950 463.050 883.050 ;
        RECT 463.950 880.950 466.050 883.050 ;
        RECT 466.950 880.950 469.050 883.050 ;
        RECT 487.800 880.950 489.900 883.050 ;
        RECT 493.950 880.950 496.050 883.050 ;
        RECT 496.950 880.950 499.050 883.050 ;
        RECT 502.500 880.950 504.600 883.050 ;
        RECT 520.950 880.950 523.050 883.050 ;
        RECT 523.950 880.950 526.050 883.050 ;
        RECT 526.950 880.950 529.050 883.050 ;
        RECT 544.950 880.950 547.050 883.050 ;
        RECT 547.950 880.950 550.050 883.050 ;
        RECT 550.950 880.950 553.050 883.050 ;
        RECT 553.950 880.950 556.050 883.050 ;
        RECT 568.950 880.950 571.050 883.050 ;
        RECT 571.950 880.950 574.050 883.050 ;
        RECT 574.950 880.950 577.050 883.050 ;
        RECT 577.950 880.950 580.050 883.050 ;
        RECT 592.950 880.950 595.050 883.050 ;
        RECT 595.950 880.950 598.050 883.050 ;
        RECT 598.950 880.950 601.050 883.050 ;
        RECT 601.950 880.950 604.050 883.050 ;
        RECT 616.950 880.950 619.050 883.050 ;
        RECT 619.950 880.950 622.050 883.050 ;
        RECT 622.950 880.950 625.050 883.050 ;
        RECT 625.950 880.950 628.050 883.050 ;
        RECT 640.950 880.950 643.050 883.050 ;
        RECT 643.950 880.950 646.050 883.050 ;
        RECT 646.950 880.950 649.050 883.050 ;
        RECT 649.950 880.950 652.050 883.050 ;
        RECT 664.950 880.950 667.050 883.050 ;
        RECT 667.950 880.950 670.050 883.050 ;
        RECT 683.100 880.950 685.200 883.050 ;
        RECT 686.400 880.950 688.500 883.050 ;
        RECT 157.200 879.150 159.000 880.950 ;
        RECT 179.100 879.150 180.900 880.950 ;
        RECT 155.100 876.300 156.900 876.900 ;
        RECT 155.100 875.100 162.900 876.300 ;
        RECT 161.700 873.600 162.900 875.100 ;
        RECT 182.700 873.600 183.600 880.950 ;
        RECT 184.950 879.150 186.750 880.950 ;
        RECT 203.100 873.600 204.300 880.950 ;
        RECT 209.100 879.150 210.900 880.950 ;
        RECT 153.000 872.100 155.400 873.600 ;
        RECT 126.000 867.900 132.600 868.800 ;
        RECT 126.000 867.600 126.900 867.900 ;
        RECT 107.100 861.000 108.900 867.600 ;
        RECT 110.100 861.600 111.900 867.600 ;
        RECT 125.100 861.600 126.900 867.600 ;
        RECT 131.100 867.600 132.600 867.900 ;
        RECT 128.100 861.000 129.900 867.000 ;
        RECT 131.100 861.600 132.900 867.600 ;
        RECT 134.100 861.000 135.900 867.600 ;
        RECT 153.600 861.600 155.400 872.100 ;
        RECT 156.600 861.000 158.400 873.600 ;
        RECT 161.100 861.600 162.900 873.600 ;
        RECT 180.000 872.400 183.600 873.600 ;
        RECT 180.000 861.600 181.800 872.400 ;
        RECT 185.100 861.000 186.900 873.600 ;
        RECT 203.100 872.100 205.500 873.600 ;
        RECT 201.000 869.100 202.800 870.900 ;
        RECT 200.700 861.000 202.500 867.600 ;
        RECT 203.700 861.600 205.500 872.100 ;
        RECT 208.800 861.000 210.600 873.600 ;
        RECT 227.100 862.500 228.900 871.800 ;
        RECT 230.700 871.200 231.900 880.950 ;
        RECT 235.950 879.150 237.750 880.950 ;
        RECT 245.100 879.150 246.900 880.950 ;
        RECT 263.100 879.150 264.900 880.950 ;
        RECT 238.950 876.450 241.050 877.050 ;
        RECT 265.950 876.450 268.050 877.050 ;
        RECT 238.950 875.550 268.050 876.450 ;
        RECT 238.950 874.950 241.050 875.550 ;
        RECT 265.950 874.950 268.050 875.550 ;
        RECT 269.700 873.600 270.900 880.950 ;
        RECT 287.400 873.600 288.300 880.950 ;
        RECT 292.950 879.150 294.750 880.950 ;
        RECT 289.950 876.450 292.050 877.050 ;
        RECT 301.950 876.450 304.050 877.050 ;
        RECT 289.950 875.550 304.050 876.450 ;
        RECT 289.950 874.950 292.050 875.550 ;
        RECT 301.950 874.950 304.050 875.550 ;
        RECT 230.100 863.400 231.900 871.200 ;
        RECT 233.100 871.200 240.900 872.100 ;
        RECT 233.100 862.500 234.900 871.200 ;
        RECT 227.100 861.600 234.900 862.500 ;
        RECT 236.100 862.500 237.900 870.300 ;
        RECT 239.100 863.400 240.900 871.200 ;
        RECT 242.100 871.500 249.900 872.400 ;
        RECT 242.100 862.500 243.900 871.500 ;
        RECT 236.100 861.600 243.900 862.500 ;
        RECT 245.100 861.000 246.900 870.600 ;
        RECT 248.100 861.600 249.900 871.500 ;
        RECT 263.400 861.000 265.200 873.600 ;
        RECT 268.500 872.100 270.900 873.600 ;
        RECT 268.500 861.600 270.300 872.100 ;
        RECT 271.200 869.100 273.000 870.900 ;
        RECT 271.500 861.000 273.300 867.600 ;
        RECT 287.100 861.600 288.900 873.600 ;
        RECT 290.100 872.700 297.900 873.600 ;
        RECT 290.100 861.600 291.900 872.700 ;
        RECT 293.100 861.000 294.900 871.800 ;
        RECT 296.100 861.600 297.900 872.700 ;
        RECT 315.000 868.800 315.900 880.950 ;
        RECT 320.100 879.150 321.900 880.950 ;
        RECT 341.100 879.150 342.900 880.950 ;
        RECT 347.700 873.600 348.900 880.950 ;
        RECT 315.000 867.900 321.600 868.800 ;
        RECT 315.000 867.600 315.900 867.900 ;
        RECT 314.100 861.600 315.900 867.600 ;
        RECT 320.100 867.600 321.600 867.900 ;
        RECT 317.100 861.000 318.900 867.000 ;
        RECT 320.100 861.600 321.900 867.600 ;
        RECT 323.100 861.000 324.900 867.600 ;
        RECT 341.400 861.000 343.200 873.600 ;
        RECT 346.500 872.100 348.900 873.600 ;
        RECT 346.500 861.600 348.300 872.100 ;
        RECT 349.200 869.100 351.000 870.900 ;
        RECT 365.700 867.600 366.900 880.950 ;
        RECT 368.100 879.150 369.900 880.950 ;
        RECT 389.100 867.600 390.300 880.950 ;
        RECT 410.700 867.600 411.900 880.950 ;
        RECT 434.100 879.150 435.900 880.950 ;
        RECT 438.000 875.400 438.900 880.950 ;
        RECT 439.950 879.150 441.750 880.950 ;
        RECT 458.100 879.150 459.900 880.950 ;
        RECT 434.100 874.500 438.900 875.400 ;
        RECT 442.950 876.450 445.050 877.050 ;
        RECT 451.950 876.450 454.050 877.050 ;
        RECT 442.950 875.550 454.050 876.450 ;
        RECT 442.950 874.950 445.050 875.550 ;
        RECT 451.950 874.950 454.050 875.550 ;
        RECT 349.500 861.000 351.300 867.600 ;
        RECT 365.100 861.600 366.900 867.600 ;
        RECT 368.100 861.000 369.900 867.600 ;
        RECT 386.100 861.000 387.900 867.600 ;
        RECT 389.100 861.600 390.900 867.600 ;
        RECT 392.100 861.000 393.900 867.600 ;
        RECT 407.100 861.000 408.900 867.600 ;
        RECT 410.100 861.600 411.900 867.600 ;
        RECT 413.100 861.000 414.900 867.600 ;
        RECT 431.100 862.500 432.900 873.600 ;
        RECT 434.100 863.400 435.900 874.500 ;
        RECT 464.700 873.600 465.900 880.950 ;
        RECT 488.100 879.150 489.900 880.950 ;
        RECT 497.250 879.150 499.050 880.950 ;
        RECT 437.100 872.400 444.900 873.300 ;
        RECT 437.100 862.500 438.900 872.400 ;
        RECT 431.100 861.600 438.900 862.500 ;
        RECT 440.100 861.000 441.900 871.500 ;
        RECT 443.100 861.600 444.900 872.400 ;
        RECT 458.400 861.000 460.200 873.600 ;
        RECT 463.500 872.100 465.900 873.600 ;
        RECT 463.500 861.600 465.300 872.100 ;
        RECT 485.100 871.500 492.900 872.400 ;
        RECT 466.200 869.100 468.000 870.900 ;
        RECT 466.500 861.000 468.300 867.600 ;
        RECT 485.100 861.600 486.900 871.500 ;
        RECT 488.100 861.000 489.900 870.600 ;
        RECT 491.100 862.500 492.900 871.500 ;
        RECT 494.100 871.200 501.900 872.100 ;
        RECT 494.100 863.400 495.900 871.200 ;
        RECT 497.100 862.500 498.900 870.300 ;
        RECT 491.100 861.600 498.900 862.500 ;
        RECT 500.100 862.500 501.900 871.200 ;
        RECT 503.100 871.200 504.300 880.950 ;
        RECT 508.950 876.450 511.050 877.050 ;
        RECT 520.950 876.450 523.050 877.050 ;
        RECT 508.950 875.550 523.050 876.450 ;
        RECT 508.950 874.950 511.050 875.550 ;
        RECT 520.950 874.950 523.050 875.550 ;
        RECT 503.100 863.400 504.900 871.200 ;
        RECT 506.100 862.500 507.900 871.800 ;
        RECT 524.100 867.600 525.300 880.950 ;
        RECT 548.100 879.150 549.900 880.950 ;
        RECT 538.950 876.450 541.050 877.050 ;
        RECT 544.950 876.450 547.050 877.050 ;
        RECT 538.950 875.550 547.050 876.450 ;
        RECT 538.950 874.950 541.050 875.550 ;
        RECT 544.950 874.950 547.050 875.550 ;
        RECT 554.100 868.800 555.000 880.950 ;
        RECT 572.100 873.600 573.300 880.950 ;
        RECT 578.100 879.150 579.900 880.950 ;
        RECT 593.100 879.150 594.900 880.950 ;
        RECT 599.700 873.600 600.900 880.950 ;
        RECT 620.100 879.150 621.900 880.950 ;
        RECT 601.950 876.450 604.050 877.050 ;
        RECT 622.950 876.450 625.050 877.050 ;
        RECT 601.950 875.550 625.050 876.450 ;
        RECT 601.950 874.950 604.050 875.550 ;
        RECT 622.950 874.950 625.050 875.550 ;
        RECT 572.100 872.100 574.500 873.600 ;
        RECT 570.000 869.100 571.800 870.900 ;
        RECT 548.400 867.900 555.000 868.800 ;
        RECT 548.400 867.600 549.900 867.900 ;
        RECT 500.100 861.600 507.900 862.500 ;
        RECT 521.100 861.000 522.900 867.600 ;
        RECT 524.100 861.600 525.900 867.600 ;
        RECT 527.100 861.000 528.900 867.600 ;
        RECT 545.100 861.000 546.900 867.600 ;
        RECT 548.100 861.600 549.900 867.600 ;
        RECT 554.100 867.600 555.000 867.900 ;
        RECT 551.100 861.000 552.900 867.000 ;
        RECT 554.100 861.600 555.900 867.600 ;
        RECT 569.700 861.000 571.500 867.600 ;
        RECT 572.700 861.600 574.500 872.100 ;
        RECT 577.800 861.000 579.600 873.600 ;
        RECT 593.400 861.000 595.200 873.600 ;
        RECT 598.500 872.100 600.900 873.600 ;
        RECT 598.500 861.600 600.300 872.100 ;
        RECT 601.200 869.100 603.000 870.900 ;
        RECT 626.100 868.800 627.000 880.950 ;
        RECT 620.400 867.900 627.000 868.800 ;
        RECT 620.400 867.600 621.900 867.900 ;
        RECT 601.500 861.000 603.300 867.600 ;
        RECT 617.100 861.000 618.900 867.600 ;
        RECT 620.100 861.600 621.900 867.600 ;
        RECT 626.100 867.600 627.000 867.900 ;
        RECT 642.000 868.800 642.900 880.950 ;
        RECT 647.100 879.150 648.900 880.950 ;
        RECT 665.100 879.150 666.900 880.950 ;
        RECT 642.000 867.900 648.600 868.800 ;
        RECT 642.000 867.600 642.900 867.900 ;
        RECT 623.100 861.000 624.900 867.000 ;
        RECT 626.100 861.600 627.900 867.600 ;
        RECT 641.100 861.600 642.900 867.600 ;
        RECT 647.100 867.600 648.600 867.900 ;
        RECT 668.100 867.600 669.300 880.950 ;
        RECT 683.700 873.600 684.600 880.950 ;
        RECT 687.000 879.150 688.800 880.950 ;
        RECT 644.100 861.000 645.900 867.000 ;
        RECT 647.100 861.600 648.900 867.600 ;
        RECT 650.100 861.000 651.900 867.600 ;
        RECT 665.100 861.000 666.900 867.600 ;
        RECT 668.100 861.600 669.900 867.600 ;
        RECT 683.100 861.600 684.900 873.600 ;
        RECT 686.100 861.000 687.900 873.000 ;
        RECT 690.000 867.600 690.900 887.700 ;
        RECT 710.700 887.400 714.300 888.300 ;
        RECT 691.950 883.050 693.750 884.850 ;
        RECT 710.100 883.050 711.900 884.850 ;
        RECT 713.100 883.050 714.300 887.400 ;
        RECT 716.100 883.050 717.900 884.850 ;
        RECT 737.100 883.050 738.300 893.400 ;
        RECT 755.100 887.400 756.900 897.000 ;
        RECT 761.700 888.000 763.500 896.400 ;
        RECT 780.000 890.400 781.800 897.000 ;
        RECT 784.500 891.600 786.300 896.400 ;
        RECT 787.500 893.400 789.300 897.000 ;
        RECT 784.500 890.400 789.600 891.600 ;
        RECT 761.700 886.800 765.000 888.000 ;
        RECT 755.100 883.050 756.900 884.850 ;
        RECT 761.100 883.050 762.900 884.850 ;
        RECT 764.100 883.050 765.000 886.800 ;
        RECT 779.100 883.050 780.900 884.850 ;
        RECT 785.250 883.050 787.050 884.850 ;
        RECT 788.700 883.050 789.600 890.400 ;
        RECT 803.100 887.400 804.900 897.000 ;
        RECT 809.700 888.000 811.500 896.400 ;
        RECT 809.700 886.800 813.000 888.000 ;
        RECT 830.100 887.400 831.900 897.000 ;
        RECT 836.700 888.000 838.500 896.400 ;
        RECT 854.100 890.400 855.900 896.400 ;
        RECT 854.700 888.300 855.900 890.400 ;
        RECT 857.100 891.300 858.900 896.400 ;
        RECT 860.100 892.200 861.900 897.000 ;
        RECT 863.100 891.300 864.900 896.400 ;
        RECT 878.100 893.400 879.900 897.000 ;
        RECT 881.100 893.400 882.900 896.400 ;
        RECT 884.100 893.400 885.900 897.000 ;
        RECT 857.100 889.950 864.900 891.300 ;
        RECT 836.700 886.800 840.000 888.000 ;
        RECT 854.700 887.400 858.300 888.300 ;
        RECT 803.100 883.050 804.900 884.850 ;
        RECT 809.100 883.050 810.900 884.850 ;
        RECT 812.100 883.050 813.000 886.800 ;
        RECT 830.100 883.050 831.900 884.850 ;
        RECT 836.100 883.050 837.900 884.850 ;
        RECT 839.100 883.050 840.000 886.800 ;
        RECT 854.100 883.050 855.900 884.850 ;
        RECT 857.100 883.050 858.300 887.400 ;
        RECT 860.100 883.050 861.900 884.850 ;
        RECT 881.700 883.050 882.600 893.400 ;
        RECT 899.700 889.200 901.500 896.400 ;
        RECT 904.800 890.400 906.600 897.000 ;
        RECT 920.700 890.400 922.500 897.000 ;
        RECT 925.200 890.400 927.000 896.400 ;
        RECT 929.700 890.400 931.500 897.000 ;
        RECT 899.700 888.300 903.900 889.200 ;
        RECT 899.100 883.050 900.900 884.850 ;
        RECT 902.700 883.050 903.900 888.300 ;
        RECT 904.950 883.050 906.750 884.850 ;
        RECT 920.250 883.050 922.050 884.850 ;
        RECT 926.100 883.050 927.300 890.400 ;
        RECT 949.500 888.000 951.300 896.400 ;
        RECT 948.000 886.800 951.300 888.000 ;
        RECT 956.100 887.400 957.900 897.000 ;
        RECT 972.000 890.400 973.800 897.000 ;
        RECT 976.500 891.600 978.300 896.400 ;
        RECT 979.500 893.400 981.300 897.000 ;
        RECT 976.500 890.400 981.600 891.600 ;
        RECT 958.950 888.450 961.050 889.050 ;
        RECT 973.950 888.450 976.050 889.050 ;
        RECT 958.950 887.550 976.050 888.450 ;
        RECT 958.950 886.950 961.050 887.550 ;
        RECT 973.950 886.950 976.050 887.550 ;
        RECT 932.100 883.050 933.900 884.850 ;
        RECT 948.000 883.050 948.900 886.800 ;
        RECT 950.100 883.050 951.900 884.850 ;
        RECT 956.100 883.050 957.900 884.850 ;
        RECT 971.100 883.050 972.900 884.850 ;
        RECT 977.250 883.050 979.050 884.850 ;
        RECT 980.700 883.050 981.600 890.400 ;
        RECT 995.100 887.400 996.900 897.000 ;
        RECT 1001.700 888.000 1003.500 896.400 ;
        RECT 1001.700 886.800 1005.000 888.000 ;
        RECT 995.100 883.050 996.900 884.850 ;
        RECT 1001.100 883.050 1002.900 884.850 ;
        RECT 1004.100 883.050 1005.000 886.800 ;
        RECT 691.800 880.950 693.900 883.050 ;
        RECT 709.950 880.950 712.050 883.050 ;
        RECT 712.950 880.950 715.050 883.050 ;
        RECT 715.950 880.950 718.050 883.050 ;
        RECT 718.950 880.950 721.050 883.050 ;
        RECT 733.950 880.950 736.050 883.050 ;
        RECT 736.950 880.950 739.050 883.050 ;
        RECT 754.950 880.950 757.050 883.050 ;
        RECT 757.950 880.950 760.050 883.050 ;
        RECT 760.950 880.950 763.050 883.050 ;
        RECT 763.950 880.950 766.050 883.050 ;
        RECT 778.950 880.950 781.050 883.050 ;
        RECT 781.950 880.950 784.050 883.050 ;
        RECT 784.950 880.950 787.050 883.050 ;
        RECT 787.950 880.950 790.050 883.050 ;
        RECT 802.950 880.950 805.050 883.050 ;
        RECT 805.950 880.950 808.050 883.050 ;
        RECT 808.950 880.950 811.050 883.050 ;
        RECT 811.950 880.950 814.050 883.050 ;
        RECT 829.950 880.950 832.050 883.050 ;
        RECT 832.950 880.950 835.050 883.050 ;
        RECT 835.950 880.950 838.050 883.050 ;
        RECT 838.950 880.950 841.050 883.050 ;
        RECT 853.950 880.950 856.050 883.050 ;
        RECT 856.950 880.950 859.050 883.050 ;
        RECT 859.950 880.950 862.050 883.050 ;
        RECT 862.950 880.950 865.050 883.050 ;
        RECT 877.950 880.950 880.050 883.050 ;
        RECT 880.950 880.950 883.050 883.050 ;
        RECT 883.950 880.950 886.050 883.050 ;
        RECT 898.950 880.950 901.050 883.050 ;
        RECT 901.950 880.950 904.050 883.050 ;
        RECT 904.950 880.950 907.050 883.050 ;
        RECT 919.950 880.950 922.050 883.050 ;
        RECT 922.950 880.950 925.050 883.050 ;
        RECT 925.950 880.950 928.050 883.050 ;
        RECT 928.950 880.950 931.050 883.050 ;
        RECT 931.950 880.950 934.050 883.050 ;
        RECT 946.950 880.950 949.050 883.050 ;
        RECT 949.950 880.950 952.050 883.050 ;
        RECT 952.950 880.950 955.050 883.050 ;
        RECT 955.950 880.950 958.050 883.050 ;
        RECT 970.950 880.950 973.050 883.050 ;
        RECT 973.950 880.950 976.050 883.050 ;
        RECT 976.950 880.950 979.050 883.050 ;
        RECT 979.950 880.950 982.050 883.050 ;
        RECT 994.950 880.950 997.050 883.050 ;
        RECT 997.950 880.950 1000.050 883.050 ;
        RECT 1000.950 880.950 1003.050 883.050 ;
        RECT 1003.950 880.950 1006.050 883.050 ;
        RECT 713.100 873.600 714.300 880.950 ;
        RECT 719.100 879.150 720.900 880.950 ;
        RECT 734.100 879.150 735.900 880.950 ;
        RECT 713.100 872.100 715.500 873.600 ;
        RECT 711.000 869.100 712.800 870.900 ;
        RECT 689.100 861.600 690.900 867.600 ;
        RECT 692.100 861.000 693.900 867.600 ;
        RECT 710.700 861.000 712.500 867.600 ;
        RECT 713.700 861.600 715.500 872.100 ;
        RECT 718.800 861.000 720.600 873.600 ;
        RECT 737.100 867.600 738.300 880.950 ;
        RECT 758.100 879.150 759.900 880.950 ;
        RECT 764.100 868.800 765.000 880.950 ;
        RECT 782.250 879.150 784.050 880.950 ;
        RECT 788.700 873.600 789.600 880.950 ;
        RECT 806.100 879.150 807.900 880.950 ;
        RECT 799.950 876.450 802.050 877.050 ;
        RECT 808.950 876.450 811.050 877.050 ;
        RECT 799.950 875.550 811.050 876.450 ;
        RECT 799.950 874.950 802.050 875.550 ;
        RECT 808.950 874.950 811.050 875.550 ;
        RECT 758.400 867.900 765.000 868.800 ;
        RECT 758.400 867.600 759.900 867.900 ;
        RECT 734.100 861.000 735.900 867.600 ;
        RECT 737.100 861.600 738.900 867.600 ;
        RECT 755.100 861.000 756.900 867.600 ;
        RECT 758.100 861.600 759.900 867.600 ;
        RECT 764.100 867.600 765.000 867.900 ;
        RECT 779.100 872.700 786.900 873.600 ;
        RECT 761.100 861.000 762.900 867.000 ;
        RECT 764.100 861.600 765.900 867.600 ;
        RECT 779.100 861.600 780.900 872.700 ;
        RECT 782.100 861.000 783.900 871.800 ;
        RECT 785.100 861.600 786.900 872.700 ;
        RECT 788.100 861.600 789.900 873.600 ;
        RECT 812.100 868.800 813.000 880.950 ;
        RECT 833.100 879.150 834.900 880.950 ;
        RECT 839.100 868.800 840.000 880.950 ;
        RECT 857.100 873.600 858.300 880.950 ;
        RECT 863.100 879.150 864.900 880.950 ;
        RECT 878.100 879.150 879.900 880.950 ;
        RECT 881.700 873.600 882.600 880.950 ;
        RECT 883.950 879.150 885.750 880.950 ;
        RECT 857.100 872.100 859.500 873.600 ;
        RECT 855.000 869.100 856.800 870.900 ;
        RECT 806.400 867.900 813.000 868.800 ;
        RECT 806.400 867.600 807.900 867.900 ;
        RECT 803.100 861.000 804.900 867.600 ;
        RECT 806.100 861.600 807.900 867.600 ;
        RECT 812.100 867.600 813.000 867.900 ;
        RECT 833.400 867.900 840.000 868.800 ;
        RECT 833.400 867.600 834.900 867.900 ;
        RECT 809.100 861.000 810.900 867.000 ;
        RECT 812.100 861.600 813.900 867.600 ;
        RECT 830.100 861.000 831.900 867.600 ;
        RECT 833.100 861.600 834.900 867.600 ;
        RECT 839.100 867.600 840.000 867.900 ;
        RECT 836.100 861.000 837.900 867.000 ;
        RECT 839.100 861.600 840.900 867.600 ;
        RECT 854.700 861.000 856.500 867.600 ;
        RECT 857.700 861.600 859.500 872.100 ;
        RECT 862.800 861.000 864.600 873.600 ;
        RECT 879.000 872.400 882.600 873.600 ;
        RECT 879.000 861.600 880.800 872.400 ;
        RECT 884.100 861.000 885.900 873.600 ;
        RECT 902.700 867.600 903.900 880.950 ;
        RECT 923.250 879.150 925.050 880.950 ;
        RECT 926.100 875.400 927.000 880.950 ;
        RECT 929.100 879.150 930.900 880.950 ;
        RECT 926.100 874.500 930.900 875.400 ;
        RECT 920.100 872.400 927.900 873.300 ;
        RECT 904.950 870.450 907.050 871.050 ;
        RECT 913.950 870.450 916.050 871.050 ;
        RECT 904.950 869.550 916.050 870.450 ;
        RECT 904.950 868.950 907.050 869.550 ;
        RECT 913.950 868.950 916.050 869.550 ;
        RECT 899.100 861.000 900.900 867.600 ;
        RECT 902.100 861.600 903.900 867.600 ;
        RECT 905.100 861.000 906.900 867.600 ;
        RECT 920.100 861.600 921.900 872.400 ;
        RECT 923.100 861.000 924.900 871.500 ;
        RECT 926.100 862.500 927.900 872.400 ;
        RECT 929.100 863.400 930.900 874.500 ;
        RECT 932.100 862.500 933.900 873.600 ;
        RECT 948.000 868.800 948.900 880.950 ;
        RECT 953.100 879.150 954.900 880.950 ;
        RECT 974.250 879.150 976.050 880.950 ;
        RECT 980.700 873.600 981.600 880.950 ;
        RECT 998.100 879.150 999.900 880.950 ;
        RECT 971.100 872.700 978.900 873.600 ;
        RECT 948.000 867.900 954.600 868.800 ;
        RECT 948.000 867.600 948.900 867.900 ;
        RECT 926.100 861.600 933.900 862.500 ;
        RECT 947.100 861.600 948.900 867.600 ;
        RECT 953.100 867.600 954.600 867.900 ;
        RECT 950.100 861.000 951.900 867.000 ;
        RECT 953.100 861.600 954.900 867.600 ;
        RECT 956.100 861.000 957.900 867.600 ;
        RECT 971.100 861.600 972.900 872.700 ;
        RECT 974.100 861.000 975.900 871.800 ;
        RECT 977.100 861.600 978.900 872.700 ;
        RECT 980.100 861.600 981.900 873.600 ;
        RECT 1004.100 868.800 1005.000 880.950 ;
        RECT 998.400 867.900 1005.000 868.800 ;
        RECT 998.400 867.600 999.900 867.900 ;
        RECT 995.100 861.000 996.900 867.600 ;
        RECT 998.100 861.600 999.900 867.600 ;
        RECT 1004.100 867.600 1005.000 867.900 ;
        RECT 1001.100 861.000 1002.900 867.000 ;
        RECT 1004.100 861.600 1005.900 867.600 ;
        RECT 17.100 846.600 18.900 857.400 ;
        RECT 20.100 847.500 21.900 858.000 ;
        RECT 17.100 845.400 21.900 846.600 ;
        RECT 19.800 844.500 21.900 845.400 ;
        RECT 24.600 845.400 26.400 857.400 ;
        RECT 29.100 847.500 30.900 858.000 ;
        RECT 32.100 846.300 33.900 857.400 ;
        RECT 47.100 851.400 48.900 858.000 ;
        RECT 50.100 851.400 51.900 857.400 ;
        RECT 53.100 851.400 54.900 858.000 ;
        RECT 29.400 845.400 33.900 846.300 ;
        RECT 24.600 844.050 25.800 845.400 ;
        RECT 24.300 843.000 25.800 844.050 ;
        RECT 29.400 843.300 31.500 845.400 ;
        RECT 24.300 841.050 25.200 843.000 ;
        RECT 17.400 838.050 19.200 839.850 ;
        RECT 23.100 838.950 25.200 841.050 ;
        RECT 26.100 841.500 28.200 841.800 ;
        RECT 26.100 839.700 30.000 841.500 ;
        RECT 17.100 835.950 19.200 838.050 ;
        RECT 23.700 838.800 25.200 838.950 ;
        RECT 23.700 837.900 26.100 838.800 ;
        RECT 21.900 835.200 23.700 837.000 ;
        RECT 21.900 833.100 24.000 835.200 ;
        RECT 24.900 832.200 26.100 837.900 ;
        RECT 27.000 838.050 28.800 838.500 ;
        RECT 50.100 838.050 51.300 851.400 ;
        RECT 68.100 846.300 69.900 857.400 ;
        RECT 71.100 847.200 72.900 858.000 ;
        RECT 74.100 846.300 75.900 857.400 ;
        RECT 68.100 845.400 75.900 846.300 ;
        RECT 77.100 845.400 78.900 857.400 ;
        RECT 92.100 851.400 93.900 858.000 ;
        RECT 95.100 851.400 96.900 857.400 ;
        RECT 98.100 852.000 99.900 858.000 ;
        RECT 95.400 851.100 96.900 851.400 ;
        RECT 101.100 851.400 102.900 857.400 ;
        RECT 116.100 851.400 117.900 857.400 ;
        RECT 119.100 851.400 120.900 858.000 ;
        RECT 101.100 851.100 102.000 851.400 ;
        RECT 95.400 850.200 102.000 851.100 ;
        RECT 71.250 838.050 73.050 839.850 ;
        RECT 77.700 838.050 78.600 845.400 ;
        RECT 95.100 838.050 96.900 839.850 ;
        RECT 101.100 838.050 102.000 850.200 ;
        RECT 116.700 838.050 117.900 851.400 ;
        RECT 134.400 845.400 136.200 858.000 ;
        RECT 139.500 846.900 141.300 857.400 ;
        RECT 142.500 851.400 144.300 858.000 ;
        RECT 161.100 851.400 162.900 857.400 ;
        RECT 164.100 851.400 165.900 858.000 ;
        RECT 142.200 848.100 144.000 849.900 ;
        RECT 139.500 845.400 141.900 846.900 ;
        RECT 119.100 838.050 120.900 839.850 ;
        RECT 134.100 838.050 135.900 839.850 ;
        RECT 140.700 838.050 141.900 845.400 ;
        RECT 161.700 838.050 162.900 851.400 ;
        RECT 168.150 847.200 169.950 857.400 ;
        RECT 167.550 845.400 169.950 847.200 ;
        RECT 171.150 845.400 172.950 858.000 ;
        RECT 176.550 848.400 178.350 857.400 ;
        RECT 181.350 851.400 183.150 858.000 ;
        RECT 184.350 850.500 186.150 857.400 ;
        RECT 187.350 851.400 189.150 858.000 ;
        RECT 191.850 851.400 193.650 857.400 ;
        RECT 180.450 849.450 187.050 850.500 ;
        RECT 180.450 848.700 182.250 849.450 ;
        RECT 185.250 848.700 187.050 849.450 ;
        RECT 191.550 849.300 193.650 851.400 ;
        RECT 176.250 847.500 178.350 848.400 ;
        RECT 188.850 847.800 190.650 848.400 ;
        RECT 176.250 846.300 184.050 847.500 ;
        RECT 182.250 845.700 184.050 846.300 ;
        RECT 184.950 846.900 190.650 847.800 ;
        RECT 167.550 844.500 168.450 845.400 ;
        RECT 184.950 844.800 185.850 846.900 ;
        RECT 188.850 846.600 190.650 846.900 ;
        RECT 191.550 846.600 194.550 848.400 ;
        RECT 191.550 845.700 192.750 846.600 ;
        RECT 177.450 844.500 185.850 844.800 ;
        RECT 167.550 843.900 185.850 844.500 ;
        RECT 187.950 844.800 192.750 845.700 ;
        RECT 196.650 845.400 198.450 858.000 ;
        RECT 199.650 845.400 201.450 857.400 ;
        RECT 218.100 851.400 219.900 858.000 ;
        RECT 221.100 851.400 222.900 857.400 ;
        RECT 239.100 851.400 240.900 858.000 ;
        RECT 242.100 851.400 243.900 857.400 ;
        RECT 245.100 851.400 246.900 858.000 ;
        RECT 263.100 851.400 264.900 858.000 ;
        RECT 266.100 851.400 267.900 857.400 ;
        RECT 281.100 851.400 282.900 858.000 ;
        RECT 284.100 851.400 285.900 857.400 ;
        RECT 287.100 851.400 288.900 858.000 ;
        RECT 305.100 851.400 306.900 857.400 ;
        RECT 308.100 851.400 309.900 858.000 ;
        RECT 167.550 843.300 179.250 843.900 ;
        RECT 164.100 838.050 165.900 839.850 ;
        RECT 27.000 836.700 33.900 838.050 ;
        RECT 31.800 835.950 33.900 836.700 ;
        RECT 46.950 835.950 49.050 838.050 ;
        RECT 49.950 835.950 52.050 838.050 ;
        RECT 52.950 835.950 55.050 838.050 ;
        RECT 67.950 835.950 70.050 838.050 ;
        RECT 70.950 835.950 73.050 838.050 ;
        RECT 73.950 835.950 76.050 838.050 ;
        RECT 76.950 835.950 79.050 838.050 ;
        RECT 91.950 835.950 94.050 838.050 ;
        RECT 94.950 835.950 97.050 838.050 ;
        RECT 97.950 835.950 100.050 838.050 ;
        RECT 100.950 835.950 103.050 838.050 ;
        RECT 115.950 835.950 118.050 838.050 ;
        RECT 118.950 835.950 121.050 838.050 ;
        RECT 133.950 835.950 136.050 838.050 ;
        RECT 136.950 835.950 139.050 838.050 ;
        RECT 139.950 835.950 142.050 838.050 ;
        RECT 142.950 835.950 145.050 838.050 ;
        RECT 160.950 835.950 163.050 838.050 ;
        RECT 163.950 835.950 166.050 838.050 ;
        RECT 19.800 829.500 21.900 830.700 ;
        RECT 23.100 830.100 26.100 832.200 ;
        RECT 27.000 833.400 28.800 835.200 ;
        RECT 31.800 834.150 33.600 835.950 ;
        RECT 47.250 834.150 49.050 835.950 ;
        RECT 27.000 831.300 29.100 833.400 ;
        RECT 27.000 830.400 33.300 831.300 ;
        RECT 17.100 828.600 21.900 829.500 ;
        RECT 24.900 828.600 26.100 830.100 ;
        RECT 32.100 828.600 33.300 830.400 ;
        RECT 50.100 830.700 51.300 835.950 ;
        RECT 53.100 834.150 54.900 835.950 ;
        RECT 68.100 834.150 69.900 835.950 ;
        RECT 74.250 834.150 76.050 835.950 ;
        RECT 50.100 829.800 54.300 830.700 ;
        RECT 17.100 822.600 18.900 828.600 ;
        RECT 20.100 822.000 21.900 827.700 ;
        RECT 24.600 822.600 26.400 828.600 ;
        RECT 29.100 822.000 30.900 827.700 ;
        RECT 32.100 822.600 33.900 828.600 ;
        RECT 47.400 822.000 49.200 828.600 ;
        RECT 52.500 822.600 54.300 829.800 ;
        RECT 77.700 828.600 78.600 835.950 ;
        RECT 92.100 834.150 93.900 835.950 ;
        RECT 98.100 834.150 99.900 835.950 ;
        RECT 101.100 832.200 102.000 835.950 ;
        RECT 69.000 822.000 70.800 828.600 ;
        RECT 73.500 827.400 78.600 828.600 ;
        RECT 73.500 822.600 75.300 827.400 ;
        RECT 76.500 822.000 78.300 825.600 ;
        RECT 92.100 822.000 93.900 831.600 ;
        RECT 98.700 831.000 102.000 832.200 ;
        RECT 98.700 822.600 100.500 831.000 ;
        RECT 116.700 825.600 117.900 835.950 ;
        RECT 137.100 834.150 138.900 835.950 ;
        RECT 140.700 831.600 141.900 835.950 ;
        RECT 143.100 834.150 144.900 835.950 ;
        RECT 140.700 830.700 144.300 831.600 ;
        RECT 134.100 827.700 141.900 829.050 ;
        RECT 116.100 822.600 117.900 825.600 ;
        RECT 119.100 822.000 120.900 825.600 ;
        RECT 134.100 822.600 135.900 827.700 ;
        RECT 137.100 822.000 138.900 826.800 ;
        RECT 140.100 822.600 141.900 827.700 ;
        RECT 143.100 828.600 144.300 830.700 ;
        RECT 143.100 822.600 144.900 828.600 ;
        RECT 161.700 825.600 162.900 835.950 ;
        RECT 167.550 828.600 168.450 843.300 ;
        RECT 177.450 843.000 179.250 843.300 ;
        RECT 169.950 835.950 172.050 838.050 ;
        RECT 179.100 836.400 181.200 838.050 ;
        RECT 169.950 833.400 171.750 835.950 ;
        RECT 173.100 835.200 181.200 836.400 ;
        RECT 173.100 834.600 174.900 835.200 ;
        RECT 176.100 833.400 177.900 834.000 ;
        RECT 169.950 832.200 177.900 833.400 ;
        RECT 187.950 832.200 188.850 844.800 ;
        RECT 191.550 842.100 193.650 842.700 ;
        RECT 197.550 842.100 199.350 842.550 ;
        RECT 191.550 840.900 199.350 842.100 ;
        RECT 191.550 840.600 193.650 840.900 ;
        RECT 197.550 840.750 199.350 840.900 ;
        RECT 200.250 838.050 201.450 845.400 ;
        RECT 218.100 838.050 219.900 839.850 ;
        RECT 221.100 838.050 222.300 851.400 ;
        RECT 242.100 838.050 243.300 851.400 ;
        RECT 263.100 838.050 264.900 839.850 ;
        RECT 266.100 838.050 267.300 851.400 ;
        RECT 284.100 838.050 285.300 851.400 ;
        RECT 305.700 838.050 306.900 851.400 ;
        RECT 323.100 845.400 324.900 858.000 ;
        RECT 328.200 846.600 330.000 857.400 ;
        RECT 344.100 851.400 345.900 858.000 ;
        RECT 347.100 851.400 348.900 857.400 ;
        RECT 350.100 851.400 351.900 858.000 ;
        RECT 365.700 851.400 367.500 858.000 ;
        RECT 326.400 845.400 330.000 846.600 ;
        RECT 308.100 838.050 309.900 839.850 ;
        RECT 323.250 838.050 325.050 839.850 ;
        RECT 326.400 838.050 327.300 845.400 ;
        RECT 329.100 838.050 330.900 839.850 ;
        RECT 347.700 838.050 348.900 851.400 ;
        RECT 366.000 848.100 367.800 849.900 ;
        RECT 368.700 846.900 370.500 857.400 ;
        RECT 368.100 845.400 370.500 846.900 ;
        RECT 373.800 845.400 375.600 858.000 ;
        RECT 389.100 845.400 390.900 857.400 ;
        RECT 392.100 846.300 393.900 857.400 ;
        RECT 395.100 847.200 396.900 858.000 ;
        RECT 398.100 846.300 399.900 857.400 ;
        RECT 392.100 845.400 399.900 846.300 ;
        RECT 413.100 845.400 414.900 857.400 ;
        RECT 416.100 846.000 417.900 858.000 ;
        RECT 419.100 851.400 420.900 857.400 ;
        RECT 422.100 851.400 423.900 858.000 ;
        RECT 437.100 851.400 438.900 858.000 ;
        RECT 440.100 851.400 441.900 857.400 ;
        RECT 443.100 851.400 444.900 858.000 ;
        RECT 368.100 838.050 369.300 845.400 ;
        RECT 374.100 838.050 375.900 839.850 ;
        RECT 389.400 838.050 390.300 845.400 ;
        RECT 394.950 838.050 396.750 839.850 ;
        RECT 413.700 838.050 414.600 845.400 ;
        RECT 417.000 838.050 418.800 839.850 ;
        RECT 196.950 837.750 201.450 838.050 ;
        RECT 195.150 835.950 201.450 837.750 ;
        RECT 217.950 835.950 220.050 838.050 ;
        RECT 220.950 835.950 223.050 838.050 ;
        RECT 238.950 835.950 241.050 838.050 ;
        RECT 241.950 835.950 244.050 838.050 ;
        RECT 244.950 835.950 247.050 838.050 ;
        RECT 262.950 835.950 265.050 838.050 ;
        RECT 265.950 835.950 268.050 838.050 ;
        RECT 280.950 835.950 283.050 838.050 ;
        RECT 283.950 835.950 286.050 838.050 ;
        RECT 286.950 835.950 289.050 838.050 ;
        RECT 304.950 835.950 307.050 838.050 ;
        RECT 307.950 835.950 310.050 838.050 ;
        RECT 322.950 835.950 325.050 838.050 ;
        RECT 325.950 835.950 328.050 838.050 ;
        RECT 328.950 835.950 331.050 838.050 ;
        RECT 343.950 835.950 346.050 838.050 ;
        RECT 346.950 835.950 349.050 838.050 ;
        RECT 349.950 835.950 352.050 838.050 ;
        RECT 364.950 835.950 367.050 838.050 ;
        RECT 367.950 835.950 370.050 838.050 ;
        RECT 370.950 835.950 373.050 838.050 ;
        RECT 373.950 835.950 376.050 838.050 ;
        RECT 388.950 835.950 391.050 838.050 ;
        RECT 391.950 835.950 394.050 838.050 ;
        RECT 394.950 835.950 397.050 838.050 ;
        RECT 397.950 835.950 400.050 838.050 ;
        RECT 413.100 835.950 415.200 838.050 ;
        RECT 416.400 835.950 418.500 838.050 ;
        RECT 176.850 831.000 188.850 832.200 ;
        RECT 176.850 829.200 177.900 831.000 ;
        RECT 187.050 830.400 188.850 831.000 ;
        RECT 167.550 826.800 169.950 828.600 ;
        RECT 161.100 822.600 162.900 825.600 ;
        RECT 164.100 822.000 165.900 825.600 ;
        RECT 168.150 822.600 169.950 826.800 ;
        RECT 171.150 822.000 172.950 828.600 ;
        RECT 173.850 826.200 175.950 827.700 ;
        RECT 176.850 827.400 178.650 829.200 ;
        RECT 200.250 828.600 201.450 835.950 ;
        RECT 179.850 827.550 181.650 828.300 ;
        RECT 179.850 826.500 184.800 827.550 ;
        RECT 173.850 825.600 177.750 826.200 ;
        RECT 183.750 825.600 184.800 826.500 ;
        RECT 191.250 825.600 193.650 827.700 ;
        RECT 174.150 824.700 177.750 825.600 ;
        RECT 175.950 822.600 177.750 824.700 ;
        RECT 180.450 822.000 182.250 825.600 ;
        RECT 183.750 822.600 185.550 825.600 ;
        RECT 186.750 822.000 188.550 825.600 ;
        RECT 191.250 822.600 193.050 825.600 ;
        RECT 196.350 822.000 198.150 828.600 ;
        RECT 199.650 822.600 201.450 828.600 ;
        RECT 221.100 825.600 222.300 835.950 ;
        RECT 239.250 834.150 241.050 835.950 ;
        RECT 242.100 830.700 243.300 835.950 ;
        RECT 245.100 834.150 246.900 835.950 ;
        RECT 242.100 829.800 246.300 830.700 ;
        RECT 218.100 822.000 219.900 825.600 ;
        RECT 221.100 822.600 222.900 825.600 ;
        RECT 239.400 822.000 241.200 828.600 ;
        RECT 244.500 822.600 246.300 829.800 ;
        RECT 266.100 825.600 267.300 835.950 ;
        RECT 281.250 834.150 283.050 835.950 ;
        RECT 284.100 830.700 285.300 835.950 ;
        RECT 287.100 834.150 288.900 835.950 ;
        RECT 284.100 829.800 288.300 830.700 ;
        RECT 263.100 822.000 264.900 825.600 ;
        RECT 266.100 822.600 267.900 825.600 ;
        RECT 281.400 822.000 283.200 828.600 ;
        RECT 286.500 822.600 288.300 829.800 ;
        RECT 305.700 825.600 306.900 835.950 ;
        RECT 326.400 825.600 327.300 835.950 ;
        RECT 344.100 834.150 345.900 835.950 ;
        RECT 347.700 830.700 348.900 835.950 ;
        RECT 349.950 834.150 351.750 835.950 ;
        RECT 365.100 834.150 366.900 835.950 ;
        RECT 368.100 831.600 369.300 835.950 ;
        RECT 371.100 834.150 372.900 835.950 ;
        RECT 344.700 829.800 348.900 830.700 ;
        RECT 365.700 830.700 369.300 831.600 ;
        RECT 305.100 822.600 306.900 825.600 ;
        RECT 308.100 822.000 309.900 825.600 ;
        RECT 323.100 822.000 324.900 825.600 ;
        RECT 326.100 822.600 327.900 825.600 ;
        RECT 329.100 822.000 330.900 825.600 ;
        RECT 344.700 822.600 346.500 829.800 ;
        RECT 365.700 828.600 366.900 830.700 ;
        RECT 349.800 822.000 351.600 828.600 ;
        RECT 365.100 822.600 366.900 828.600 ;
        RECT 368.100 827.700 375.900 829.050 ;
        RECT 368.100 822.600 369.900 827.700 ;
        RECT 371.100 822.000 372.900 826.800 ;
        RECT 374.100 822.600 375.900 827.700 ;
        RECT 389.400 828.600 390.300 835.950 ;
        RECT 391.950 834.150 393.750 835.950 ;
        RECT 398.100 834.150 399.900 835.950 ;
        RECT 413.700 828.600 414.600 835.950 ;
        RECT 420.000 831.300 420.900 851.400 ;
        RECT 440.700 838.050 441.900 851.400 ;
        RECT 459.000 846.600 460.800 857.400 ;
        RECT 459.000 845.400 462.600 846.600 ;
        RECT 464.100 845.400 465.900 858.000 ;
        RECT 479.100 851.400 480.900 858.000 ;
        RECT 482.100 851.400 483.900 857.400 ;
        RECT 485.100 851.400 486.900 858.000 ;
        RECT 500.100 851.400 501.900 858.000 ;
        RECT 503.100 851.400 504.900 857.400 ;
        RECT 458.100 838.050 459.900 839.850 ;
        RECT 461.700 838.050 462.600 845.400 ;
        RECT 463.950 838.050 465.750 839.850 ;
        RECT 482.100 838.050 483.300 851.400 ;
        RECT 421.800 835.950 423.900 838.050 ;
        RECT 436.950 835.950 439.050 838.050 ;
        RECT 439.950 835.950 442.050 838.050 ;
        RECT 442.950 835.950 445.050 838.050 ;
        RECT 457.950 835.950 460.050 838.050 ;
        RECT 460.950 835.950 463.050 838.050 ;
        RECT 463.950 835.950 466.050 838.050 ;
        RECT 478.950 835.950 481.050 838.050 ;
        RECT 481.950 835.950 484.050 838.050 ;
        RECT 484.950 835.950 487.050 838.050 ;
        RECT 500.100 835.950 502.200 838.050 ;
        RECT 421.950 834.150 423.750 835.950 ;
        RECT 437.100 834.150 438.900 835.950 ;
        RECT 415.500 830.400 423.900 831.300 ;
        RECT 440.700 830.700 441.900 835.950 ;
        RECT 442.950 834.150 444.750 835.950 ;
        RECT 415.500 829.500 417.300 830.400 ;
        RECT 389.400 827.400 394.500 828.600 ;
        RECT 389.700 822.000 391.500 825.600 ;
        RECT 392.700 822.600 394.500 827.400 ;
        RECT 397.200 822.000 399.000 828.600 ;
        RECT 413.700 826.800 416.400 828.600 ;
        RECT 414.600 822.600 416.400 826.800 ;
        RECT 417.600 822.000 419.400 828.600 ;
        RECT 422.100 822.600 423.900 830.400 ;
        RECT 437.700 829.800 441.900 830.700 ;
        RECT 437.700 822.600 439.500 829.800 ;
        RECT 442.800 822.000 444.600 828.600 ;
        RECT 461.700 825.600 462.600 835.950 ;
        RECT 479.250 834.150 481.050 835.950 ;
        RECT 482.100 830.700 483.300 835.950 ;
        RECT 485.100 834.150 486.900 835.950 ;
        RECT 500.250 834.150 502.050 835.950 ;
        RECT 503.100 831.300 504.000 851.400 ;
        RECT 506.100 846.000 507.900 858.000 ;
        RECT 509.100 845.400 510.900 857.400 ;
        RECT 524.100 851.400 525.900 858.000 ;
        RECT 527.100 851.400 528.900 857.400 ;
        RECT 530.100 851.400 531.900 858.000 ;
        RECT 548.100 851.400 549.900 857.400 ;
        RECT 551.100 852.000 552.900 858.000 ;
        RECT 505.200 838.050 507.000 839.850 ;
        RECT 509.400 838.050 510.300 845.400 ;
        RECT 527.100 838.050 528.300 851.400 ;
        RECT 549.000 851.100 549.900 851.400 ;
        RECT 554.100 851.400 555.900 857.400 ;
        RECT 557.100 851.400 558.900 858.000 ;
        RECT 575.100 851.400 576.900 858.000 ;
        RECT 578.100 851.400 579.900 857.400 ;
        RECT 581.100 852.000 582.900 858.000 ;
        RECT 554.100 851.100 555.600 851.400 ;
        RECT 549.000 850.200 555.600 851.100 ;
        RECT 578.400 851.100 579.900 851.400 ;
        RECT 584.100 851.400 585.900 857.400 ;
        RECT 599.100 851.400 600.900 858.000 ;
        RECT 602.100 851.400 603.900 857.400 ;
        RECT 605.100 851.400 606.900 858.000 ;
        RECT 623.100 851.400 624.900 858.000 ;
        RECT 626.100 851.400 627.900 857.400 ;
        RECT 629.100 851.400 630.900 858.000 ;
        RECT 647.100 851.400 648.900 858.000 ;
        RECT 650.100 851.400 651.900 857.400 ;
        RECT 665.100 851.400 666.900 858.000 ;
        RECT 668.100 851.400 669.900 857.400 ;
        RECT 671.100 851.400 672.900 858.000 ;
        RECT 689.100 851.400 690.900 858.000 ;
        RECT 692.100 851.400 693.900 857.400 ;
        RECT 695.100 851.400 696.900 858.000 ;
        RECT 710.100 851.400 711.900 858.000 ;
        RECT 713.100 851.400 714.900 857.400 ;
        RECT 716.100 851.400 717.900 858.000 ;
        RECT 584.100 851.100 585.000 851.400 ;
        RECT 578.400 850.200 585.000 851.100 ;
        RECT 549.000 838.050 549.900 850.200 ;
        RECT 554.100 838.050 555.900 839.850 ;
        RECT 578.100 838.050 579.900 839.850 ;
        RECT 584.100 838.050 585.000 850.200 ;
        RECT 602.100 838.050 603.300 851.400 ;
        RECT 626.100 838.050 627.300 851.400 ;
        RECT 647.100 838.050 648.900 839.850 ;
        RECT 650.100 838.050 651.300 851.400 ;
        RECT 668.100 838.050 669.300 851.400 ;
        RECT 692.100 838.050 693.300 851.400 ;
        RECT 694.950 843.450 697.050 844.200 ;
        RECT 703.950 843.450 706.050 844.050 ;
        RECT 694.950 842.550 706.050 843.450 ;
        RECT 694.950 842.100 697.050 842.550 ;
        RECT 703.950 841.950 706.050 842.550 ;
        RECT 713.100 838.050 714.300 851.400 ;
        RECT 731.100 845.400 732.900 858.000 ;
        RECT 736.200 846.600 738.000 857.400 ;
        RECT 734.400 845.400 738.000 846.600 ;
        RECT 752.400 845.400 754.200 858.000 ;
        RECT 757.500 846.900 759.300 857.400 ;
        RECT 760.500 851.400 762.300 858.000 ;
        RECT 760.200 848.100 762.000 849.900 ;
        RECT 779.100 847.500 780.900 857.400 ;
        RECT 782.100 848.400 783.900 858.000 ;
        RECT 785.100 856.500 792.900 857.400 ;
        RECT 785.100 847.500 786.900 856.500 ;
        RECT 757.500 845.400 759.900 846.900 ;
        RECT 779.100 846.600 786.900 847.500 ;
        RECT 788.100 847.800 789.900 855.600 ;
        RECT 791.100 848.700 792.900 856.500 ;
        RECT 794.100 856.500 801.900 857.400 ;
        RECT 794.100 847.800 795.900 856.500 ;
        RECT 788.100 846.900 795.900 847.800 ;
        RECT 797.100 847.800 798.900 855.600 ;
        RECT 731.250 838.050 733.050 839.850 ;
        RECT 734.400 838.050 735.300 845.400 ;
        RECT 737.100 838.050 738.900 839.850 ;
        RECT 752.100 838.050 753.900 839.850 ;
        RECT 758.700 838.050 759.900 845.400 ;
        RECT 782.100 838.050 783.900 839.850 ;
        RECT 791.250 838.050 793.050 839.850 ;
        RECT 797.100 838.050 798.300 847.800 ;
        RECT 800.100 847.200 801.900 856.500 ;
        RECT 815.400 845.400 817.200 858.000 ;
        RECT 820.500 846.900 822.300 857.400 ;
        RECT 823.500 851.400 825.300 858.000 ;
        RECT 842.100 851.400 843.900 858.000 ;
        RECT 845.100 851.400 846.900 857.400 ;
        RECT 848.100 852.000 849.900 858.000 ;
        RECT 845.400 851.100 846.900 851.400 ;
        RECT 851.100 851.400 852.900 857.400 ;
        RECT 851.100 851.100 852.000 851.400 ;
        RECT 845.400 850.200 852.000 851.100 ;
        RECT 823.200 848.100 825.000 849.900 ;
        RECT 820.500 845.400 822.900 846.900 ;
        RECT 815.100 838.050 816.900 839.850 ;
        RECT 821.700 838.050 822.900 845.400 ;
        RECT 845.100 838.050 846.900 839.850 ;
        RECT 851.100 838.050 852.000 850.200 ;
        RECT 866.100 845.400 867.900 857.400 ;
        RECT 869.100 846.300 870.900 857.400 ;
        RECT 872.100 847.200 873.900 858.000 ;
        RECT 875.100 846.300 876.900 857.400 ;
        RECT 890.100 851.400 891.900 858.000 ;
        RECT 893.100 851.400 894.900 857.400 ;
        RECT 896.100 852.000 897.900 858.000 ;
        RECT 893.400 851.100 894.900 851.400 ;
        RECT 899.100 851.400 900.900 857.400 ;
        RECT 899.100 851.100 900.000 851.400 ;
        RECT 893.400 850.200 900.000 851.100 ;
        RECT 869.100 845.400 876.900 846.300 ;
        RECT 866.400 838.050 867.300 845.400 ;
        RECT 868.950 843.450 871.050 844.050 ;
        RECT 895.950 843.450 898.050 844.050 ;
        RECT 868.950 842.550 898.050 843.450 ;
        RECT 868.950 841.950 871.050 842.550 ;
        RECT 895.950 841.950 898.050 842.550 ;
        RECT 885.000 840.450 889.050 841.050 ;
        RECT 871.950 838.050 873.750 839.850 ;
        RECT 884.550 838.950 889.050 840.450 ;
        RECT 505.500 835.950 507.600 838.050 ;
        RECT 508.800 835.950 510.900 838.050 ;
        RECT 523.950 835.950 526.050 838.050 ;
        RECT 526.950 835.950 529.050 838.050 ;
        RECT 529.950 835.950 532.050 838.050 ;
        RECT 547.950 835.950 550.050 838.050 ;
        RECT 550.950 835.950 553.050 838.050 ;
        RECT 553.950 835.950 556.050 838.050 ;
        RECT 556.950 835.950 559.050 838.050 ;
        RECT 574.950 835.950 577.050 838.050 ;
        RECT 577.950 835.950 580.050 838.050 ;
        RECT 580.950 835.950 583.050 838.050 ;
        RECT 583.950 835.950 586.050 838.050 ;
        RECT 598.950 835.950 601.050 838.050 ;
        RECT 601.950 835.950 604.050 838.050 ;
        RECT 604.950 835.950 607.050 838.050 ;
        RECT 622.950 835.950 625.050 838.050 ;
        RECT 625.950 835.950 628.050 838.050 ;
        RECT 628.950 835.950 631.050 838.050 ;
        RECT 646.950 835.950 649.050 838.050 ;
        RECT 649.950 835.950 652.050 838.050 ;
        RECT 664.950 835.950 667.050 838.050 ;
        RECT 667.950 835.950 670.050 838.050 ;
        RECT 670.950 835.950 673.050 838.050 ;
        RECT 688.950 835.950 691.050 838.050 ;
        RECT 691.950 835.950 694.050 838.050 ;
        RECT 694.950 835.950 697.050 838.050 ;
        RECT 709.950 835.950 712.050 838.050 ;
        RECT 712.950 835.950 715.050 838.050 ;
        RECT 715.950 835.950 718.050 838.050 ;
        RECT 730.950 835.950 733.050 838.050 ;
        RECT 733.950 835.950 736.050 838.050 ;
        RECT 736.950 835.950 739.050 838.050 ;
        RECT 751.950 835.950 754.050 838.050 ;
        RECT 754.950 835.950 757.050 838.050 ;
        RECT 757.950 835.950 760.050 838.050 ;
        RECT 760.950 835.950 763.050 838.050 ;
        RECT 781.800 835.950 783.900 838.050 ;
        RECT 787.950 835.950 790.050 838.050 ;
        RECT 790.950 835.950 793.050 838.050 ;
        RECT 796.500 835.950 798.600 838.050 ;
        RECT 814.950 835.950 817.050 838.050 ;
        RECT 817.950 835.950 820.050 838.050 ;
        RECT 820.950 835.950 823.050 838.050 ;
        RECT 823.950 835.950 826.050 838.050 ;
        RECT 841.950 835.950 844.050 838.050 ;
        RECT 844.950 835.950 847.050 838.050 ;
        RECT 847.950 835.950 850.050 838.050 ;
        RECT 850.950 835.950 853.050 838.050 ;
        RECT 865.950 835.950 868.050 838.050 ;
        RECT 868.950 835.950 871.050 838.050 ;
        RECT 871.950 835.950 874.050 838.050 ;
        RECT 874.950 835.950 877.050 838.050 ;
        RECT 482.100 829.800 486.300 830.700 ;
        RECT 458.100 822.000 459.900 825.600 ;
        RECT 461.100 822.600 462.900 825.600 ;
        RECT 464.100 822.000 465.900 825.600 ;
        RECT 479.400 822.000 481.200 828.600 ;
        RECT 484.500 822.600 486.300 829.800 ;
        RECT 500.100 830.400 508.500 831.300 ;
        RECT 500.100 822.600 501.900 830.400 ;
        RECT 506.700 829.500 508.500 830.400 ;
        RECT 509.400 828.600 510.300 835.950 ;
        RECT 524.250 834.150 526.050 835.950 ;
        RECT 527.100 830.700 528.300 835.950 ;
        RECT 530.100 834.150 531.900 835.950 ;
        RECT 549.000 832.200 549.900 835.950 ;
        RECT 551.100 834.150 552.900 835.950 ;
        RECT 557.100 834.150 558.900 835.950 ;
        RECT 575.100 834.150 576.900 835.950 ;
        RECT 581.100 834.150 582.900 835.950 ;
        RECT 584.100 832.200 585.000 835.950 ;
        RECT 586.950 834.450 589.050 835.050 ;
        RECT 592.950 834.450 595.050 835.050 ;
        RECT 586.950 833.550 595.050 834.450 ;
        RECT 599.250 834.150 601.050 835.950 ;
        RECT 586.950 832.950 589.050 833.550 ;
        RECT 592.950 832.950 595.050 833.550 ;
        RECT 549.000 831.000 552.300 832.200 ;
        RECT 527.100 829.800 531.300 830.700 ;
        RECT 504.600 822.000 506.400 828.600 ;
        RECT 507.600 826.800 510.300 828.600 ;
        RECT 507.600 822.600 509.400 826.800 ;
        RECT 524.400 822.000 526.200 828.600 ;
        RECT 529.500 822.600 531.300 829.800 ;
        RECT 550.500 822.600 552.300 831.000 ;
        RECT 557.100 822.000 558.900 831.600 ;
        RECT 575.100 822.000 576.900 831.600 ;
        RECT 581.700 831.000 585.000 832.200 ;
        RECT 581.700 822.600 583.500 831.000 ;
        RECT 602.100 830.700 603.300 835.950 ;
        RECT 605.100 834.150 606.900 835.950 ;
        RECT 623.250 834.150 625.050 835.950 ;
        RECT 626.100 830.700 627.300 835.950 ;
        RECT 629.100 834.150 630.900 835.950 ;
        RECT 602.100 829.800 606.300 830.700 ;
        RECT 626.100 829.800 630.300 830.700 ;
        RECT 599.400 822.000 601.200 828.600 ;
        RECT 604.500 822.600 606.300 829.800 ;
        RECT 623.400 822.000 625.200 828.600 ;
        RECT 628.500 822.600 630.300 829.800 ;
        RECT 650.100 825.600 651.300 835.950 ;
        RECT 665.250 834.150 667.050 835.950 ;
        RECT 668.100 830.700 669.300 835.950 ;
        RECT 671.100 834.150 672.900 835.950 ;
        RECT 689.250 834.150 691.050 835.950 ;
        RECT 692.100 830.700 693.300 835.950 ;
        RECT 695.100 834.150 696.900 835.950 ;
        RECT 710.250 834.150 712.050 835.950 ;
        RECT 713.100 830.700 714.300 835.950 ;
        RECT 716.100 834.150 717.900 835.950 ;
        RECT 668.100 829.800 672.300 830.700 ;
        RECT 692.100 829.800 696.300 830.700 ;
        RECT 713.100 829.800 717.300 830.700 ;
        RECT 647.100 822.000 648.900 825.600 ;
        RECT 650.100 822.600 651.900 825.600 ;
        RECT 665.400 822.000 667.200 828.600 ;
        RECT 670.500 822.600 672.300 829.800 ;
        RECT 689.400 822.000 691.200 828.600 ;
        RECT 694.500 822.600 696.300 829.800 ;
        RECT 710.400 822.000 712.200 828.600 ;
        RECT 715.500 822.600 717.300 829.800 ;
        RECT 734.400 825.600 735.300 835.950 ;
        RECT 755.100 834.150 756.900 835.950 ;
        RECT 758.700 831.600 759.900 835.950 ;
        RECT 761.100 834.150 762.900 835.950 ;
        RECT 787.950 834.150 789.750 835.950 ;
        RECT 758.700 830.700 762.300 831.600 ;
        RECT 752.100 827.700 759.900 829.050 ;
        RECT 731.100 822.000 732.900 825.600 ;
        RECT 734.100 822.600 735.900 825.600 ;
        RECT 737.100 822.000 738.900 825.600 ;
        RECT 752.100 822.600 753.900 827.700 ;
        RECT 755.100 822.000 756.900 826.800 ;
        RECT 758.100 822.600 759.900 827.700 ;
        RECT 761.100 828.600 762.300 830.700 ;
        RECT 772.950 831.450 775.050 832.050 ;
        RECT 790.950 831.450 793.050 832.050 ;
        RECT 772.950 830.550 793.050 831.450 ;
        RECT 772.950 829.950 775.050 830.550 ;
        RECT 790.950 829.950 793.050 830.550 ;
        RECT 761.100 822.600 762.900 828.600 ;
        RECT 766.950 828.450 769.050 829.050 ;
        RECT 781.950 828.450 784.050 829.050 ;
        RECT 766.950 827.550 784.050 828.450 ;
        RECT 766.950 826.950 769.050 827.550 ;
        RECT 781.950 826.950 784.050 827.550 ;
        RECT 797.100 827.400 798.300 835.950 ;
        RECT 818.100 834.150 819.900 835.950 ;
        RECT 821.700 831.600 822.900 835.950 ;
        RECT 824.100 834.150 825.900 835.950 ;
        RECT 842.100 834.150 843.900 835.950 ;
        RECT 848.100 834.150 849.900 835.950 ;
        RECT 851.100 832.200 852.000 835.950 ;
        RECT 821.700 830.700 825.300 831.600 ;
        RECT 785.700 826.500 798.300 827.400 ;
        RECT 815.100 827.700 822.900 829.050 ;
        RECT 785.700 825.600 786.600 826.500 ;
        RECT 792.900 825.600 793.800 826.500 ;
        RECT 781.800 822.000 783.900 825.600 ;
        RECT 785.100 822.600 786.900 825.600 ;
        RECT 788.100 822.000 789.900 825.600 ;
        RECT 791.100 822.600 793.800 825.600 ;
        RECT 815.100 822.600 816.900 827.700 ;
        RECT 818.100 822.000 819.900 826.800 ;
        RECT 821.100 822.600 822.900 827.700 ;
        RECT 824.100 828.600 825.300 830.700 ;
        RECT 824.100 822.600 825.900 828.600 ;
        RECT 842.100 822.000 843.900 831.600 ;
        RECT 848.700 831.000 852.000 832.200 ;
        RECT 848.700 822.600 850.500 831.000 ;
        RECT 866.400 828.600 867.300 835.950 ;
        RECT 868.950 834.150 870.750 835.950 ;
        RECT 875.100 834.150 876.900 835.950 ;
        RECT 877.950 834.450 880.050 835.050 ;
        RECT 884.550 834.450 885.450 838.950 ;
        RECT 893.100 838.050 894.900 839.850 ;
        RECT 899.100 838.050 900.000 850.200 ;
        RECT 914.400 845.400 916.200 858.000 ;
        RECT 919.500 846.900 921.300 857.400 ;
        RECT 922.500 851.400 924.300 858.000 ;
        RECT 922.200 848.100 924.000 849.900 ;
        RECT 938.100 847.500 939.900 857.400 ;
        RECT 941.100 848.400 942.900 858.000 ;
        RECT 944.100 856.500 951.900 857.400 ;
        RECT 944.100 847.500 945.900 856.500 ;
        RECT 919.500 845.400 921.900 846.900 ;
        RECT 938.100 846.600 945.900 847.500 ;
        RECT 947.100 847.800 948.900 855.600 ;
        RECT 950.100 848.700 951.900 856.500 ;
        RECT 953.100 856.500 960.900 857.400 ;
        RECT 953.100 847.800 954.900 856.500 ;
        RECT 947.100 846.900 954.900 847.800 ;
        RECT 956.100 847.800 957.900 855.600 ;
        RECT 901.950 840.450 906.000 841.050 ;
        RECT 901.950 838.950 906.450 840.450 ;
        RECT 889.950 835.950 892.050 838.050 ;
        RECT 892.950 835.950 895.050 838.050 ;
        RECT 895.950 835.950 898.050 838.050 ;
        RECT 898.950 835.950 901.050 838.050 ;
        RECT 877.950 833.550 885.450 834.450 ;
        RECT 890.100 834.150 891.900 835.950 ;
        RECT 896.100 834.150 897.900 835.950 ;
        RECT 877.950 832.950 880.050 833.550 ;
        RECT 899.100 832.200 900.000 835.950 ;
        RECT 905.550 835.050 906.450 838.950 ;
        RECT 914.100 838.050 915.900 839.850 ;
        RECT 920.700 838.050 921.900 845.400 ;
        RECT 940.950 843.450 943.050 844.050 ;
        RECT 952.950 843.450 955.050 844.050 ;
        RECT 940.950 842.550 955.050 843.450 ;
        RECT 940.950 841.950 943.050 842.550 ;
        RECT 952.950 841.950 955.050 842.550 ;
        RECT 925.950 840.450 928.050 841.050 ;
        RECT 934.950 840.450 937.050 841.050 ;
        RECT 925.950 839.550 937.050 840.450 ;
        RECT 925.950 838.950 928.050 839.550 ;
        RECT 934.950 838.950 937.050 839.550 ;
        RECT 941.100 838.050 942.900 839.850 ;
        RECT 950.250 838.050 952.050 839.850 ;
        RECT 956.100 838.050 957.300 847.800 ;
        RECT 959.100 847.200 960.900 856.500 ;
        RECT 977.100 845.400 978.900 857.400 ;
        RECT 980.100 846.300 981.900 857.400 ;
        RECT 983.100 847.200 984.900 858.000 ;
        RECT 986.100 846.300 987.900 857.400 ;
        RECT 1004.100 851.400 1005.900 857.400 ;
        RECT 1007.100 851.400 1008.900 858.000 ;
        RECT 980.100 845.400 987.900 846.300 ;
        RECT 977.400 838.050 978.300 845.400 ;
        RECT 979.950 843.450 982.050 844.200 ;
        RECT 985.950 843.450 988.050 844.050 ;
        RECT 979.950 842.550 988.050 843.450 ;
        RECT 979.950 842.100 982.050 842.550 ;
        RECT 985.950 841.950 988.050 842.550 ;
        RECT 988.950 840.450 993.000 841.050 ;
        RECT 982.950 838.050 984.750 839.850 ;
        RECT 988.950 838.950 993.450 840.450 ;
        RECT 913.950 835.950 916.050 838.050 ;
        RECT 916.950 835.950 919.050 838.050 ;
        RECT 919.950 835.950 922.050 838.050 ;
        RECT 922.950 835.950 925.050 838.050 ;
        RECT 940.800 835.950 942.900 838.050 ;
        RECT 946.950 835.950 949.050 838.050 ;
        RECT 949.950 835.950 952.050 838.050 ;
        RECT 955.500 835.950 957.600 838.050 ;
        RECT 958.950 837.450 961.050 838.050 ;
        RECT 958.950 836.550 972.450 837.450 ;
        RECT 958.950 835.950 961.050 836.550 ;
        RECT 901.950 833.550 906.450 835.050 ;
        RECT 917.100 834.150 918.900 835.950 ;
        RECT 901.950 832.950 906.000 833.550 ;
        RECT 866.400 827.400 871.500 828.600 ;
        RECT 866.700 822.000 868.500 825.600 ;
        RECT 869.700 822.600 871.500 827.400 ;
        RECT 874.200 822.000 876.000 828.600 ;
        RECT 890.100 822.000 891.900 831.600 ;
        RECT 896.700 831.000 900.000 832.200 ;
        RECT 920.700 831.600 921.900 835.950 ;
        RECT 923.100 834.150 924.900 835.950 ;
        RECT 946.950 834.150 948.750 835.950 ;
        RECT 896.700 822.600 898.500 831.000 ;
        RECT 920.700 830.700 924.300 831.600 ;
        RECT 914.100 827.700 921.900 829.050 ;
        RECT 914.100 822.600 915.900 827.700 ;
        RECT 917.100 822.000 918.900 826.800 ;
        RECT 920.100 822.600 921.900 827.700 ;
        RECT 923.100 828.600 924.300 830.700 ;
        RECT 923.100 822.600 924.900 828.600 ;
        RECT 956.100 827.400 957.300 835.950 ;
        RECT 971.550 835.050 972.450 836.550 ;
        RECT 976.950 835.950 979.050 838.050 ;
        RECT 979.950 835.950 982.050 838.050 ;
        RECT 982.950 835.950 985.050 838.050 ;
        RECT 985.950 835.950 988.050 838.050 ;
        RECT 971.550 833.550 976.050 835.050 ;
        RECT 972.000 832.950 976.050 833.550 ;
        RECT 977.400 828.600 978.300 835.950 ;
        RECT 979.950 834.150 981.750 835.950 ;
        RECT 986.100 834.150 987.900 835.950 ;
        RECT 979.950 831.450 982.050 832.050 ;
        RECT 992.550 831.450 993.450 838.950 ;
        RECT 1004.700 838.050 1005.900 851.400 ;
        RECT 1007.100 838.050 1008.900 839.850 ;
        RECT 1003.950 835.950 1006.050 838.050 ;
        RECT 1006.950 835.950 1009.050 838.050 ;
        RECT 979.950 830.550 993.450 831.450 ;
        RECT 979.950 829.950 982.050 830.550 ;
        RECT 977.400 827.400 982.500 828.600 ;
        RECT 944.700 826.500 957.300 827.400 ;
        RECT 944.700 825.600 945.600 826.500 ;
        RECT 951.900 825.600 952.800 826.500 ;
        RECT 940.800 822.000 942.900 825.600 ;
        RECT 944.100 822.600 945.900 825.600 ;
        RECT 947.100 822.000 948.900 825.600 ;
        RECT 950.100 822.600 952.800 825.600 ;
        RECT 977.700 822.000 979.500 825.600 ;
        RECT 980.700 822.600 982.500 827.400 ;
        RECT 985.200 822.000 987.000 828.600 ;
        RECT 1004.700 825.600 1005.900 835.950 ;
        RECT 1004.100 822.600 1005.900 825.600 ;
        RECT 1007.100 822.000 1008.900 825.600 ;
        RECT 14.100 815.400 15.900 818.400 ;
        RECT 17.100 815.400 18.900 819.000 ;
        RECT 14.700 805.050 15.900 815.400 ;
        RECT 20.550 812.400 22.350 818.400 ;
        RECT 23.850 812.400 25.650 819.000 ;
        RECT 28.950 815.400 30.750 818.400 ;
        RECT 33.450 815.400 35.250 819.000 ;
        RECT 36.450 815.400 38.250 818.400 ;
        RECT 39.750 815.400 41.550 819.000 ;
        RECT 44.250 816.300 46.050 818.400 ;
        RECT 44.250 815.400 47.850 816.300 ;
        RECT 28.350 813.300 30.750 815.400 ;
        RECT 37.200 814.500 38.250 815.400 ;
        RECT 44.250 814.800 48.150 815.400 ;
        RECT 37.200 813.450 42.150 814.500 ;
        RECT 40.350 812.700 42.150 813.450 ;
        RECT 20.550 805.050 21.750 812.400 ;
        RECT 43.350 811.800 45.150 813.600 ;
        RECT 46.050 813.300 48.150 814.800 ;
        RECT 49.050 812.400 50.850 819.000 ;
        RECT 52.050 814.200 53.850 818.400 ;
        RECT 71.100 815.400 72.900 818.400 ;
        RECT 74.100 815.400 75.900 819.000 ;
        RECT 52.050 812.400 54.450 814.200 ;
        RECT 33.150 810.000 34.950 810.600 ;
        RECT 44.100 810.000 45.150 811.800 ;
        RECT 33.150 808.800 45.150 810.000 ;
        RECT 13.950 802.950 16.050 805.050 ;
        RECT 16.950 802.950 19.050 805.050 ;
        RECT 20.550 803.250 26.850 805.050 ;
        RECT 20.550 802.950 25.050 803.250 ;
        RECT 14.700 789.600 15.900 802.950 ;
        RECT 17.100 801.150 18.900 802.950 ;
        RECT 20.550 795.600 21.750 802.950 ;
        RECT 22.650 800.100 24.450 800.250 ;
        RECT 28.350 800.100 30.450 800.400 ;
        RECT 22.650 798.900 30.450 800.100 ;
        RECT 22.650 798.450 24.450 798.900 ;
        RECT 28.350 798.300 30.450 798.900 ;
        RECT 33.150 796.200 34.050 808.800 ;
        RECT 44.100 807.600 52.050 808.800 ;
        RECT 44.100 807.000 45.900 807.600 ;
        RECT 47.100 805.800 48.900 806.400 ;
        RECT 40.800 804.600 48.900 805.800 ;
        RECT 50.250 805.050 52.050 807.600 ;
        RECT 40.800 802.950 42.900 804.600 ;
        RECT 49.950 802.950 52.050 805.050 ;
        RECT 42.750 797.700 44.550 798.000 ;
        RECT 53.550 797.700 54.450 812.400 ;
        RECT 71.700 805.050 72.900 815.400 ;
        RECT 89.100 809.400 90.900 819.000 ;
        RECT 95.700 810.000 97.500 818.400 ;
        RECT 117.000 812.400 118.800 819.000 ;
        RECT 121.500 813.600 123.300 818.400 ;
        RECT 124.500 815.400 126.300 819.000 ;
        RECT 121.500 812.400 126.600 813.600 ;
        RECT 95.700 808.800 99.000 810.000 ;
        RECT 89.100 805.050 90.900 806.850 ;
        RECT 95.100 805.050 96.900 806.850 ;
        RECT 98.100 805.050 99.000 808.800 ;
        RECT 116.100 805.050 117.900 806.850 ;
        RECT 122.250 805.050 124.050 806.850 ;
        RECT 125.700 805.050 126.600 812.400 ;
        RECT 140.700 811.200 142.500 818.400 ;
        RECT 145.800 812.400 147.600 819.000 ;
        RECT 161.100 812.400 162.900 818.400 ;
        RECT 140.700 810.300 144.900 811.200 ;
        RECT 140.100 805.050 141.900 806.850 ;
        RECT 143.700 805.050 144.900 810.300 ;
        RECT 161.700 810.300 162.900 812.400 ;
        RECT 164.100 813.300 165.900 818.400 ;
        RECT 167.100 814.200 168.900 819.000 ;
        RECT 170.100 813.300 171.900 818.400 ;
        RECT 164.100 811.950 171.900 813.300 ;
        RECT 188.100 812.400 189.900 818.400 ;
        RECT 188.700 810.300 189.900 812.400 ;
        RECT 191.100 813.300 192.900 818.400 ;
        RECT 194.100 814.200 195.900 819.000 ;
        RECT 197.100 813.300 198.900 818.400 ;
        RECT 201.150 814.200 202.950 818.400 ;
        RECT 191.100 811.950 198.900 813.300 ;
        RECT 200.550 812.400 202.950 814.200 ;
        RECT 204.150 812.400 205.950 819.000 ;
        RECT 208.950 816.300 210.750 818.400 ;
        RECT 207.150 815.400 210.750 816.300 ;
        RECT 213.450 815.400 215.250 819.000 ;
        RECT 216.750 815.400 218.550 818.400 ;
        RECT 219.750 815.400 221.550 819.000 ;
        RECT 224.250 815.400 226.050 818.400 ;
        RECT 206.850 814.800 210.750 815.400 ;
        RECT 206.850 813.300 208.950 814.800 ;
        RECT 216.750 814.500 217.800 815.400 ;
        RECT 161.700 809.400 165.300 810.300 ;
        RECT 188.700 809.400 192.300 810.300 ;
        RECT 145.950 805.050 147.750 806.850 ;
        RECT 161.100 805.050 162.900 806.850 ;
        RECT 164.100 805.050 165.300 809.400 ;
        RECT 167.100 805.050 168.900 806.850 ;
        RECT 188.100 805.050 189.900 806.850 ;
        RECT 191.100 805.050 192.300 809.400 ;
        RECT 194.100 805.050 195.900 806.850 ;
        RECT 70.950 802.950 73.050 805.050 ;
        RECT 73.950 802.950 76.050 805.050 ;
        RECT 88.950 802.950 91.050 805.050 ;
        RECT 91.950 802.950 94.050 805.050 ;
        RECT 94.950 802.950 97.050 805.050 ;
        RECT 97.950 802.950 100.050 805.050 ;
        RECT 115.950 802.950 118.050 805.050 ;
        RECT 118.950 802.950 121.050 805.050 ;
        RECT 121.950 802.950 124.050 805.050 ;
        RECT 124.950 802.950 127.050 805.050 ;
        RECT 139.950 802.950 142.050 805.050 ;
        RECT 142.950 802.950 145.050 805.050 ;
        RECT 145.950 802.950 148.050 805.050 ;
        RECT 160.950 802.950 163.050 805.050 ;
        RECT 163.950 802.950 166.050 805.050 ;
        RECT 166.950 802.950 169.050 805.050 ;
        RECT 169.950 802.950 172.050 805.050 ;
        RECT 187.950 802.950 190.050 805.050 ;
        RECT 190.950 802.950 193.050 805.050 ;
        RECT 193.950 802.950 196.050 805.050 ;
        RECT 196.950 802.950 199.050 805.050 ;
        RECT 42.750 797.100 54.450 797.700 ;
        RECT 14.100 783.600 15.900 789.600 ;
        RECT 17.100 783.000 18.900 789.600 ;
        RECT 20.550 783.600 22.350 795.600 ;
        RECT 23.550 783.000 25.350 795.600 ;
        RECT 29.250 795.300 34.050 796.200 ;
        RECT 36.150 796.500 54.450 797.100 ;
        RECT 36.150 796.200 44.550 796.500 ;
        RECT 29.250 794.400 30.450 795.300 ;
        RECT 27.450 792.600 30.450 794.400 ;
        RECT 31.350 794.100 33.150 794.400 ;
        RECT 36.150 794.100 37.050 796.200 ;
        RECT 53.550 795.600 54.450 796.500 ;
        RECT 31.350 793.200 37.050 794.100 ;
        RECT 37.950 794.700 39.750 795.300 ;
        RECT 37.950 793.500 45.750 794.700 ;
        RECT 31.350 792.600 33.150 793.200 ;
        RECT 43.650 792.600 45.750 793.500 ;
        RECT 28.350 789.600 30.450 791.700 ;
        RECT 34.950 791.550 36.750 792.300 ;
        RECT 39.750 791.550 41.550 792.300 ;
        RECT 34.950 790.500 41.550 791.550 ;
        RECT 28.350 783.600 30.150 789.600 ;
        RECT 32.850 783.000 34.650 789.600 ;
        RECT 35.850 783.600 37.650 790.500 ;
        RECT 38.850 783.000 40.650 789.600 ;
        RECT 43.650 783.600 45.450 792.600 ;
        RECT 49.050 783.000 50.850 795.600 ;
        RECT 52.050 793.800 54.450 795.600 ;
        RECT 52.050 783.600 53.850 793.800 ;
        RECT 71.700 789.600 72.900 802.950 ;
        RECT 74.100 801.150 75.900 802.950 ;
        RECT 92.100 801.150 93.900 802.950 ;
        RECT 73.950 798.450 76.050 799.050 ;
        RECT 94.950 798.450 97.050 799.050 ;
        RECT 73.950 797.550 97.050 798.450 ;
        RECT 73.950 796.950 76.050 797.550 ;
        RECT 94.950 796.950 97.050 797.550 ;
        RECT 98.100 790.800 99.000 802.950 ;
        RECT 119.250 801.150 121.050 802.950 ;
        RECT 125.700 795.600 126.600 802.950 ;
        RECT 92.400 789.900 99.000 790.800 ;
        RECT 92.400 789.600 93.900 789.900 ;
        RECT 71.100 783.600 72.900 789.600 ;
        RECT 74.100 783.000 75.900 789.600 ;
        RECT 89.100 783.000 90.900 789.600 ;
        RECT 92.100 783.600 93.900 789.600 ;
        RECT 98.100 789.600 99.000 789.900 ;
        RECT 116.100 794.700 123.900 795.600 ;
        RECT 95.100 783.000 96.900 789.000 ;
        RECT 98.100 783.600 99.900 789.600 ;
        RECT 116.100 783.600 117.900 794.700 ;
        RECT 119.100 783.000 120.900 793.800 ;
        RECT 122.100 783.600 123.900 794.700 ;
        RECT 125.100 783.600 126.900 795.600 ;
        RECT 143.700 789.600 144.900 802.950 ;
        RECT 164.100 795.600 165.300 802.950 ;
        RECT 170.100 801.150 171.900 802.950 ;
        RECT 191.100 795.600 192.300 802.950 ;
        RECT 197.100 801.150 198.900 802.950 ;
        RECT 200.550 797.700 201.450 812.400 ;
        RECT 209.850 811.800 211.650 813.600 ;
        RECT 212.850 813.450 217.800 814.500 ;
        RECT 212.850 812.700 214.650 813.450 ;
        RECT 224.250 813.300 226.650 815.400 ;
        RECT 229.350 812.400 231.150 819.000 ;
        RECT 232.650 812.400 234.450 818.400 ;
        RECT 209.850 810.000 210.900 811.800 ;
        RECT 220.050 810.000 221.850 810.600 ;
        RECT 209.850 808.800 221.850 810.000 ;
        RECT 202.950 807.600 210.900 808.800 ;
        RECT 202.950 805.050 204.750 807.600 ;
        RECT 209.100 807.000 210.900 807.600 ;
        RECT 206.100 805.800 207.900 806.400 ;
        RECT 202.950 802.950 205.050 805.050 ;
        RECT 206.100 804.600 214.200 805.800 ;
        RECT 212.100 802.950 214.200 804.600 ;
        RECT 210.450 797.700 212.250 798.000 ;
        RECT 200.550 797.100 212.250 797.700 ;
        RECT 200.550 796.500 218.850 797.100 ;
        RECT 200.550 795.600 201.450 796.500 ;
        RECT 210.450 796.200 218.850 796.500 ;
        RECT 164.100 794.100 166.500 795.600 ;
        RECT 162.000 791.100 163.800 792.900 ;
        RECT 140.100 783.000 141.900 789.600 ;
        RECT 143.100 783.600 144.900 789.600 ;
        RECT 146.100 783.000 147.900 789.600 ;
        RECT 161.700 783.000 163.500 789.600 ;
        RECT 164.700 783.600 166.500 794.100 ;
        RECT 169.800 783.000 171.600 795.600 ;
        RECT 191.100 794.100 193.500 795.600 ;
        RECT 189.000 791.100 190.800 792.900 ;
        RECT 188.700 783.000 190.500 789.600 ;
        RECT 191.700 783.600 193.500 794.100 ;
        RECT 196.800 783.000 198.600 795.600 ;
        RECT 200.550 793.800 202.950 795.600 ;
        RECT 201.150 783.600 202.950 793.800 ;
        RECT 204.150 783.000 205.950 795.600 ;
        RECT 215.250 794.700 217.050 795.300 ;
        RECT 209.250 793.500 217.050 794.700 ;
        RECT 217.950 794.100 218.850 796.200 ;
        RECT 220.950 796.200 221.850 808.800 ;
        RECT 233.250 805.050 234.450 812.400 ;
        RECT 248.100 813.300 249.900 818.400 ;
        RECT 251.100 814.200 252.900 819.000 ;
        RECT 254.100 813.300 255.900 818.400 ;
        RECT 248.100 811.950 255.900 813.300 ;
        RECT 257.100 812.400 258.900 818.400 ;
        RECT 272.100 812.400 273.900 818.400 ;
        RECT 275.100 813.300 276.900 819.000 ;
        RECT 279.300 813.000 281.100 818.400 ;
        RECT 283.800 813.300 285.600 819.000 ;
        RECT 257.100 810.300 258.300 812.400 ;
        RECT 254.700 809.400 258.300 810.300 ;
        RECT 272.100 811.500 273.600 812.400 ;
        RECT 272.100 810.000 276.600 811.500 ;
        RECT 274.500 809.400 276.600 810.000 ;
        RECT 280.200 810.900 281.100 813.000 ;
        RECT 287.100 812.400 288.900 818.400 ;
        RECT 305.100 812.400 306.900 818.400 ;
        RECT 308.100 813.300 309.900 819.000 ;
        RECT 312.600 812.400 314.400 818.400 ;
        RECT 317.100 813.300 318.900 819.000 ;
        RECT 320.100 812.400 321.900 818.400 ;
        RECT 322.950 816.450 325.050 817.050 ;
        RECT 331.950 816.450 334.050 817.050 ;
        RECT 322.950 815.550 334.050 816.450 ;
        RECT 322.950 814.950 325.050 815.550 ;
        RECT 331.950 814.950 334.050 815.550 ;
        RECT 337.500 812.400 339.300 819.000 ;
        RECT 342.000 812.400 343.800 818.400 ;
        RECT 346.500 812.400 348.300 819.000 ;
        RECT 365.400 812.400 367.200 819.000 ;
        RECT 284.400 811.500 288.900 812.400 ;
        RECT 251.100 805.050 252.900 806.850 ;
        RECT 254.700 805.050 255.900 809.400 ;
        RECT 277.500 807.900 279.300 809.700 ;
        RECT 280.200 808.800 283.200 810.900 ;
        RECT 284.400 809.100 286.500 811.500 ;
        RECT 305.700 810.600 306.900 812.400 ;
        RECT 312.900 810.900 314.100 812.400 ;
        RECT 317.100 811.500 321.900 812.400 ;
        RECT 305.700 809.700 312.000 810.600 ;
        RECT 276.900 807.000 279.000 807.900 ;
        RECT 257.100 805.050 258.900 806.850 ;
        RECT 272.400 805.800 279.000 807.000 ;
        RECT 272.400 805.200 274.200 805.800 ;
        RECT 228.150 803.250 234.450 805.050 ;
        RECT 229.950 802.950 234.450 803.250 ;
        RECT 247.950 802.950 250.050 805.050 ;
        RECT 250.950 802.950 253.050 805.050 ;
        RECT 253.950 802.950 256.050 805.050 ;
        RECT 256.950 802.950 259.050 805.050 ;
        RECT 272.100 802.950 274.200 805.200 ;
        RECT 224.550 800.100 226.650 800.400 ;
        RECT 230.550 800.100 232.350 800.250 ;
        RECT 224.550 798.900 232.350 800.100 ;
        RECT 224.550 798.300 226.650 798.900 ;
        RECT 230.550 798.450 232.350 798.900 ;
        RECT 220.950 795.300 225.750 796.200 ;
        RECT 233.250 795.600 234.450 802.950 ;
        RECT 248.100 801.150 249.900 802.950 ;
        RECT 254.700 795.600 255.900 802.950 ;
        RECT 276.900 802.800 279.000 804.900 ;
        RECT 276.900 801.000 278.700 802.800 ;
        RECT 280.200 802.050 281.100 808.800 ;
        RECT 309.900 807.600 312.000 809.700 ;
        RECT 282.000 804.900 284.100 807.000 ;
        RECT 305.400 805.050 307.200 806.850 ;
        RECT 310.200 805.800 312.000 807.600 ;
        RECT 312.900 808.800 315.900 810.900 ;
        RECT 317.100 810.300 319.200 811.500 ;
        RECT 282.000 803.100 283.800 804.900 ;
        RECT 286.800 802.950 288.900 805.050 ;
        RECT 305.100 804.300 307.200 805.050 ;
        RECT 305.100 802.950 312.000 804.300 ;
        RECT 280.200 800.700 283.200 802.050 ;
        RECT 286.800 801.150 288.600 802.950 ;
        RECT 310.200 802.500 312.000 802.950 ;
        RECT 312.900 803.100 314.100 808.800 ;
        RECT 315.000 805.800 317.100 807.900 ;
        RECT 315.300 804.000 317.100 805.800 ;
        RECT 335.100 805.050 336.900 806.850 ;
        RECT 341.700 805.050 342.900 812.400 ;
        RECT 370.500 811.200 372.300 818.400 ;
        RECT 389.100 815.400 390.900 818.400 ;
        RECT 392.100 815.400 393.900 819.000 ;
        RECT 368.100 810.300 372.300 811.200 ;
        RECT 360.000 807.450 364.050 808.050 ;
        RECT 346.950 805.050 348.750 806.850 ;
        RECT 359.550 805.950 364.050 807.450 ;
        RECT 312.900 802.200 315.300 803.100 ;
        RECT 313.800 802.050 315.300 802.200 ;
        RECT 319.800 802.950 321.900 805.050 ;
        RECT 334.950 802.950 337.050 805.050 ;
        RECT 337.950 802.950 340.050 805.050 ;
        RECT 340.950 802.950 343.050 805.050 ;
        RECT 343.950 802.950 346.050 805.050 ;
        RECT 346.950 802.950 349.050 805.050 ;
        RECT 281.100 799.950 283.200 800.700 ;
        RECT 278.400 797.700 280.200 799.500 ;
        RECT 274.800 796.800 280.200 797.700 ;
        RECT 274.800 795.900 276.900 796.800 ;
        RECT 224.550 794.400 225.750 795.300 ;
        RECT 221.850 794.100 223.650 794.400 ;
        RECT 209.250 792.600 211.350 793.500 ;
        RECT 217.950 793.200 223.650 794.100 ;
        RECT 221.850 792.600 223.650 793.200 ;
        RECT 224.550 792.600 227.550 794.400 ;
        RECT 209.550 783.600 211.350 792.600 ;
        RECT 213.450 791.550 215.250 792.300 ;
        RECT 218.250 791.550 220.050 792.300 ;
        RECT 213.450 790.500 220.050 791.550 ;
        RECT 214.350 783.000 216.150 789.600 ;
        RECT 217.350 783.600 219.150 790.500 ;
        RECT 224.550 789.600 226.650 791.700 ;
        RECT 220.350 783.000 222.150 789.600 ;
        RECT 224.850 783.600 226.650 789.600 ;
        RECT 229.650 783.000 231.450 795.600 ;
        RECT 232.650 783.600 234.450 795.600 ;
        RECT 248.400 783.000 250.200 795.600 ;
        RECT 253.500 794.100 255.900 795.600 ;
        RECT 272.100 794.700 276.900 795.900 ;
        RECT 281.700 795.600 282.900 799.950 ;
        RECT 309.000 799.500 312.900 801.300 ;
        RECT 310.800 799.200 312.900 799.500 ;
        RECT 313.800 799.950 315.900 802.050 ;
        RECT 319.800 801.150 321.600 802.950 ;
        RECT 338.100 801.150 339.900 802.950 ;
        RECT 313.800 798.000 314.700 799.950 ;
        RECT 279.600 794.700 282.900 795.600 ;
        RECT 283.800 795.600 285.900 796.500 ;
        RECT 307.500 795.600 309.600 797.700 ;
        RECT 313.200 796.950 314.700 798.000 ;
        RECT 328.950 798.450 331.050 798.900 ;
        RECT 334.950 798.450 337.050 799.050 ;
        RECT 328.950 797.550 337.050 798.450 ;
        RECT 313.200 795.600 314.400 796.950 ;
        RECT 328.950 796.800 331.050 797.550 ;
        RECT 334.950 796.950 337.050 797.550 ;
        RECT 342.000 797.400 342.900 802.950 ;
        RECT 343.950 801.150 345.750 802.950 ;
        RECT 349.950 801.450 352.050 802.050 ;
        RECT 359.550 801.450 360.450 805.950 ;
        RECT 365.250 805.050 367.050 806.850 ;
        RECT 368.100 805.050 369.300 810.300 ;
        RECT 371.100 805.050 372.900 806.850 ;
        RECT 389.700 805.050 390.900 815.400 ;
        RECT 407.100 809.400 408.900 819.000 ;
        RECT 413.700 810.000 415.500 818.400 ;
        RECT 434.100 810.600 435.900 818.400 ;
        RECT 438.600 812.400 440.400 819.000 ;
        RECT 441.600 814.200 443.400 818.400 ;
        RECT 441.600 812.400 444.300 814.200 ;
        RECT 440.700 810.600 442.500 811.500 ;
        RECT 413.700 808.800 417.000 810.000 ;
        RECT 434.100 809.700 442.500 810.600 ;
        RECT 407.100 805.050 408.900 806.850 ;
        RECT 413.100 805.050 414.900 806.850 ;
        RECT 416.100 805.050 417.000 808.800 ;
        RECT 434.250 805.050 436.050 806.850 ;
        RECT 364.950 802.950 367.050 805.050 ;
        RECT 367.950 802.950 370.050 805.050 ;
        RECT 370.950 802.950 373.050 805.050 ;
        RECT 388.950 802.950 391.050 805.050 ;
        RECT 391.950 802.950 394.050 805.050 ;
        RECT 406.950 802.950 409.050 805.050 ;
        RECT 409.950 802.950 412.050 805.050 ;
        RECT 412.950 802.950 415.050 805.050 ;
        RECT 415.950 802.950 418.050 805.050 ;
        RECT 434.100 802.950 436.200 805.050 ;
        RECT 349.950 800.550 360.450 801.450 ;
        RECT 349.950 799.950 352.050 800.550 ;
        RECT 338.100 796.500 342.900 797.400 ;
        RECT 253.500 783.600 255.300 794.100 ;
        RECT 256.200 791.100 258.000 792.900 ;
        RECT 256.500 783.000 258.300 789.600 ;
        RECT 272.100 783.600 273.900 794.700 ;
        RECT 275.100 783.000 276.900 793.500 ;
        RECT 279.600 783.600 281.400 794.700 ;
        RECT 283.800 794.400 288.900 795.600 ;
        RECT 283.800 783.000 285.900 793.500 ;
        RECT 287.100 783.600 288.900 794.400 ;
        RECT 305.100 794.700 309.600 795.600 ;
        RECT 305.100 783.600 306.900 794.700 ;
        RECT 308.100 783.000 309.900 793.500 ;
        RECT 312.600 783.600 314.400 795.600 ;
        RECT 317.100 795.600 319.200 796.500 ;
        RECT 317.100 794.400 321.900 795.600 ;
        RECT 317.100 783.000 318.900 793.500 ;
        RECT 320.100 783.600 321.900 794.400 ;
        RECT 335.100 784.500 336.900 795.600 ;
        RECT 338.100 785.400 339.900 796.500 ;
        RECT 341.100 794.400 348.900 795.300 ;
        RECT 341.100 784.500 342.900 794.400 ;
        RECT 335.100 783.600 342.900 784.500 ;
        RECT 344.100 783.000 345.900 793.500 ;
        RECT 347.100 783.600 348.900 794.400 ;
        RECT 368.100 789.600 369.300 802.950 ;
        RECT 389.700 789.600 390.900 802.950 ;
        RECT 392.100 801.150 393.900 802.950 ;
        RECT 410.100 801.150 411.900 802.950 ;
        RECT 416.100 790.800 417.000 802.950 ;
        RECT 410.400 789.900 417.000 790.800 ;
        RECT 410.400 789.600 411.900 789.900 ;
        RECT 365.100 783.000 366.900 789.600 ;
        RECT 368.100 783.600 369.900 789.600 ;
        RECT 371.100 783.000 372.900 789.600 ;
        RECT 389.100 783.600 390.900 789.600 ;
        RECT 392.100 783.000 393.900 789.600 ;
        RECT 407.100 783.000 408.900 789.600 ;
        RECT 410.100 783.600 411.900 789.600 ;
        RECT 416.100 789.600 417.000 789.900 ;
        RECT 437.100 789.600 438.000 809.700 ;
        RECT 443.400 805.050 444.300 812.400 ;
        RECT 458.700 811.200 460.500 818.400 ;
        RECT 463.800 812.400 465.600 819.000 ;
        RECT 482.700 812.400 484.500 819.000 ;
        RECT 487.200 812.400 489.000 818.400 ;
        RECT 491.700 812.400 493.500 819.000 ;
        RECT 510.600 814.200 512.400 818.400 ;
        RECT 509.700 812.400 512.400 814.200 ;
        RECT 513.600 812.400 515.400 819.000 ;
        RECT 458.700 810.300 462.900 811.200 ;
        RECT 458.100 805.050 459.900 806.850 ;
        RECT 461.700 805.050 462.900 810.300 ;
        RECT 463.950 805.050 465.750 806.850 ;
        RECT 482.250 805.050 484.050 806.850 ;
        RECT 488.100 805.050 489.300 812.400 ;
        RECT 494.100 805.050 495.900 806.850 ;
        RECT 509.700 805.050 510.600 812.400 ;
        RECT 511.500 810.600 513.300 811.500 ;
        RECT 518.100 810.600 519.900 818.400 ;
        RECT 533.100 813.300 534.900 818.400 ;
        RECT 536.100 814.200 537.900 819.000 ;
        RECT 539.100 813.300 540.900 818.400 ;
        RECT 533.100 811.950 540.900 813.300 ;
        RECT 542.100 812.400 543.900 818.400 ;
        RECT 557.100 815.400 558.900 819.000 ;
        RECT 560.100 815.400 561.900 818.400 ;
        RECT 511.500 809.700 519.900 810.600 ;
        RECT 542.100 810.300 543.300 812.400 ;
        RECT 439.500 802.950 441.600 805.050 ;
        RECT 442.800 802.950 444.900 805.050 ;
        RECT 457.950 802.950 460.050 805.050 ;
        RECT 460.950 802.950 463.050 805.050 ;
        RECT 463.950 802.950 466.050 805.050 ;
        RECT 481.950 802.950 484.050 805.050 ;
        RECT 484.950 802.950 487.050 805.050 ;
        RECT 487.950 802.950 490.050 805.050 ;
        RECT 490.950 802.950 493.050 805.050 ;
        RECT 493.950 802.950 496.050 805.050 ;
        RECT 509.100 802.950 511.200 805.050 ;
        RECT 512.400 802.950 514.500 805.050 ;
        RECT 439.200 801.150 441.000 802.950 ;
        RECT 443.400 795.600 444.300 802.950 ;
        RECT 413.100 783.000 414.900 789.000 ;
        RECT 416.100 783.600 417.900 789.600 ;
        RECT 434.100 783.000 435.900 789.600 ;
        RECT 437.100 783.600 438.900 789.600 ;
        RECT 440.100 783.000 441.900 795.000 ;
        RECT 443.100 783.600 444.900 795.600 ;
        RECT 461.700 789.600 462.900 802.950 ;
        RECT 485.250 801.150 487.050 802.950 ;
        RECT 488.100 797.400 489.000 802.950 ;
        RECT 491.100 801.150 492.900 802.950 ;
        RECT 488.100 796.500 492.900 797.400 ;
        RECT 482.100 794.400 489.900 795.300 ;
        RECT 458.100 783.000 459.900 789.600 ;
        RECT 461.100 783.600 462.900 789.600 ;
        RECT 464.100 783.000 465.900 789.600 ;
        RECT 482.100 783.600 483.900 794.400 ;
        RECT 485.100 783.000 486.900 793.500 ;
        RECT 488.100 784.500 489.900 794.400 ;
        RECT 491.100 785.400 492.900 796.500 ;
        RECT 509.700 795.600 510.600 802.950 ;
        RECT 513.000 801.150 514.800 802.950 ;
        RECT 494.100 784.500 495.900 795.600 ;
        RECT 488.100 783.600 495.900 784.500 ;
        RECT 509.100 783.600 510.900 795.600 ;
        RECT 512.100 783.000 513.900 795.000 ;
        RECT 516.000 789.600 516.900 809.700 ;
        RECT 539.700 809.400 543.300 810.300 ;
        RECT 528.000 807.450 532.050 808.050 ;
        RECT 517.950 805.050 519.750 806.850 ;
        RECT 527.550 805.950 532.050 807.450 ;
        RECT 517.800 802.950 519.900 805.050 ;
        RECT 527.550 802.050 528.450 805.950 ;
        RECT 536.100 805.050 537.900 806.850 ;
        RECT 539.700 805.050 540.900 809.400 ;
        RECT 542.100 805.050 543.900 806.850 ;
        RECT 560.100 805.050 561.300 815.400 ;
        RECT 578.400 812.400 580.200 819.000 ;
        RECT 583.500 811.200 585.300 818.400 ;
        RECT 599.100 815.400 600.900 818.400 ;
        RECT 602.100 815.400 603.900 819.000 ;
        RECT 581.100 810.300 585.300 811.200 ;
        RECT 578.250 805.050 580.050 806.850 ;
        RECT 581.100 805.050 582.300 810.300 ;
        RECT 584.100 805.050 585.900 806.850 ;
        RECT 599.700 805.050 600.900 815.400 ;
        RECT 617.100 812.400 618.900 818.400 ;
        RECT 620.100 813.300 621.900 819.000 ;
        RECT 624.300 813.000 626.100 818.400 ;
        RECT 628.800 813.300 630.600 819.000 ;
        RECT 617.100 811.500 618.600 812.400 ;
        RECT 617.100 810.000 621.600 811.500 ;
        RECT 619.500 809.400 621.600 810.000 ;
        RECT 625.200 810.900 626.100 813.000 ;
        RECT 632.100 812.400 633.900 818.400 ;
        RECT 629.400 811.500 633.900 812.400 ;
        RECT 622.500 807.900 624.300 809.700 ;
        RECT 625.200 808.800 628.200 810.900 ;
        RECT 629.400 809.100 631.500 811.500 ;
        RECT 647.100 809.400 648.900 819.000 ;
        RECT 653.700 810.000 655.500 818.400 ;
        RECT 671.700 811.200 673.500 818.400 ;
        RECT 676.800 812.400 678.600 819.000 ;
        RECT 692.700 811.200 694.500 818.400 ;
        RECT 697.800 812.400 699.600 819.000 ;
        RECT 715.500 812.400 717.300 819.000 ;
        RECT 720.000 812.400 721.800 818.400 ;
        RECT 724.500 812.400 726.300 819.000 ;
        RECT 740.400 812.400 742.200 819.000 ;
        RECT 671.700 810.300 675.900 811.200 ;
        RECT 692.700 810.300 696.900 811.200 ;
        RECT 653.700 808.800 657.000 810.000 ;
        RECT 621.900 807.000 624.000 807.900 ;
        RECT 617.400 805.800 624.000 807.000 ;
        RECT 617.400 805.200 619.200 805.800 ;
        RECT 532.950 802.950 535.050 805.050 ;
        RECT 535.950 802.950 538.050 805.050 ;
        RECT 538.950 802.950 541.050 805.050 ;
        RECT 541.950 802.950 544.050 805.050 ;
        RECT 556.950 802.950 559.050 805.050 ;
        RECT 559.950 802.950 562.050 805.050 ;
        RECT 577.950 802.950 580.050 805.050 ;
        RECT 580.950 802.950 583.050 805.050 ;
        RECT 583.950 802.950 586.050 805.050 ;
        RECT 598.950 802.950 601.050 805.050 ;
        RECT 601.950 802.950 604.050 805.050 ;
        RECT 617.100 802.950 619.200 805.200 ;
        RECT 527.550 800.550 532.050 802.050 ;
        RECT 533.100 801.150 534.900 802.950 ;
        RECT 528.000 799.950 532.050 800.550 ;
        RECT 539.700 795.600 540.900 802.950 ;
        RECT 544.950 801.450 547.050 802.050 ;
        RECT 550.950 801.450 553.050 802.050 ;
        RECT 544.950 800.550 553.050 801.450 ;
        RECT 557.100 801.150 558.900 802.950 ;
        RECT 544.950 799.950 547.050 800.550 ;
        RECT 550.950 799.950 553.050 800.550 ;
        RECT 515.100 783.600 516.900 789.600 ;
        RECT 518.100 783.000 519.900 789.600 ;
        RECT 533.400 783.000 535.200 795.600 ;
        RECT 538.500 794.100 540.900 795.600 ;
        RECT 538.500 783.600 540.300 794.100 ;
        RECT 541.200 791.100 543.000 792.900 ;
        RECT 560.100 789.600 561.300 802.950 ;
        RECT 581.100 789.600 582.300 802.950 ;
        RECT 599.700 789.600 600.900 802.950 ;
        RECT 602.100 801.150 603.900 802.950 ;
        RECT 621.900 802.800 624.000 804.900 ;
        RECT 621.900 801.000 623.700 802.800 ;
        RECT 625.200 802.050 626.100 808.800 ;
        RECT 627.000 804.900 629.100 807.000 ;
        RECT 647.100 805.050 648.900 806.850 ;
        RECT 653.100 805.050 654.900 806.850 ;
        RECT 656.100 805.050 657.000 808.800 ;
        RECT 671.100 805.050 672.900 806.850 ;
        RECT 674.700 805.050 675.900 810.300 ;
        RECT 676.950 805.050 678.750 806.850 ;
        RECT 692.100 805.050 693.900 806.850 ;
        RECT 695.700 805.050 696.900 810.300 ;
        RECT 697.950 805.050 699.750 806.850 ;
        RECT 713.100 805.050 714.900 806.850 ;
        RECT 719.700 805.050 720.900 812.400 ;
        RECT 745.500 811.200 747.300 818.400 ;
        RECT 761.700 812.400 763.500 819.000 ;
        RECT 766.200 812.400 768.000 818.400 ;
        RECT 770.700 812.400 772.500 819.000 ;
        RECT 788.100 815.400 789.900 819.000 ;
        RECT 791.100 815.400 792.900 818.400 ;
        RECT 743.100 810.300 747.300 811.200 ;
        RECT 724.950 805.050 726.750 806.850 ;
        RECT 740.250 805.050 742.050 806.850 ;
        RECT 743.100 805.050 744.300 810.300 ;
        RECT 746.100 805.050 747.900 806.850 ;
        RECT 761.250 805.050 763.050 806.850 ;
        RECT 767.100 805.050 768.300 812.400 ;
        RECT 773.100 805.050 774.900 806.850 ;
        RECT 791.100 805.050 792.300 815.400 ;
        RECT 806.100 812.400 807.900 818.400 ;
        RECT 806.700 810.300 807.900 812.400 ;
        RECT 809.100 813.300 810.900 818.400 ;
        RECT 812.100 814.200 813.900 819.000 ;
        RECT 815.100 813.300 816.900 818.400 ;
        RECT 809.100 811.950 816.900 813.300 ;
        RECT 806.700 809.400 810.300 810.300 ;
        RECT 830.100 809.400 831.900 819.000 ;
        RECT 836.700 810.000 838.500 818.400 ;
        RECT 857.400 812.400 859.200 819.000 ;
        RECT 862.500 811.200 864.300 818.400 ;
        RECT 860.100 810.300 864.300 811.200 ;
        RECT 806.100 805.050 807.900 806.850 ;
        RECT 809.100 805.050 810.300 809.400 ;
        RECT 836.700 808.800 840.000 810.000 ;
        RECT 812.100 805.050 813.900 806.850 ;
        RECT 830.100 805.050 831.900 806.850 ;
        RECT 836.100 805.050 837.900 806.850 ;
        RECT 839.100 805.050 840.000 808.800 ;
        RECT 857.250 805.050 859.050 806.850 ;
        RECT 860.100 805.050 861.300 810.300 ;
        RECT 878.100 809.400 879.900 819.000 ;
        RECT 884.700 810.000 886.500 818.400 ;
        RECT 903.000 812.400 904.800 819.000 ;
        RECT 907.500 813.600 909.300 818.400 ;
        RECT 910.500 815.400 912.300 819.000 ;
        RECT 907.500 812.400 912.600 813.600 ;
        RECT 926.100 812.400 927.900 818.400 ;
        RECT 884.700 808.800 888.000 810.000 ;
        RECT 873.000 807.450 877.050 808.050 ;
        RECT 863.100 805.050 864.900 806.850 ;
        RECT 872.550 805.950 877.050 807.450 ;
        RECT 627.000 803.100 628.800 804.900 ;
        RECT 631.800 802.950 633.900 805.050 ;
        RECT 646.950 802.950 649.050 805.050 ;
        RECT 649.950 802.950 652.050 805.050 ;
        RECT 652.950 802.950 655.050 805.050 ;
        RECT 655.950 802.950 658.050 805.050 ;
        RECT 670.950 802.950 673.050 805.050 ;
        RECT 673.950 802.950 676.050 805.050 ;
        RECT 676.950 802.950 679.050 805.050 ;
        RECT 691.950 802.950 694.050 805.050 ;
        RECT 694.950 802.950 697.050 805.050 ;
        RECT 697.950 802.950 700.050 805.050 ;
        RECT 712.950 802.950 715.050 805.050 ;
        RECT 715.950 802.950 718.050 805.050 ;
        RECT 718.950 802.950 721.050 805.050 ;
        RECT 721.950 802.950 724.050 805.050 ;
        RECT 724.950 802.950 727.050 805.050 ;
        RECT 739.950 802.950 742.050 805.050 ;
        RECT 742.950 802.950 745.050 805.050 ;
        RECT 745.950 802.950 748.050 805.050 ;
        RECT 760.950 802.950 763.050 805.050 ;
        RECT 763.950 802.950 766.050 805.050 ;
        RECT 766.950 802.950 769.050 805.050 ;
        RECT 769.950 802.950 772.050 805.050 ;
        RECT 772.950 802.950 775.050 805.050 ;
        RECT 787.950 802.950 790.050 805.050 ;
        RECT 790.950 802.950 793.050 805.050 ;
        RECT 805.950 802.950 808.050 805.050 ;
        RECT 808.950 802.950 811.050 805.050 ;
        RECT 811.950 802.950 814.050 805.050 ;
        RECT 814.950 802.950 817.050 805.050 ;
        RECT 829.950 802.950 832.050 805.050 ;
        RECT 832.950 802.950 835.050 805.050 ;
        RECT 835.950 802.950 838.050 805.050 ;
        RECT 838.950 802.950 841.050 805.050 ;
        RECT 856.950 802.950 859.050 805.050 ;
        RECT 859.950 802.950 862.050 805.050 ;
        RECT 862.950 802.950 865.050 805.050 ;
        RECT 625.200 800.700 628.200 802.050 ;
        RECT 631.800 801.150 633.600 802.950 ;
        RECT 650.100 801.150 651.900 802.950 ;
        RECT 626.100 799.950 628.200 800.700 ;
        RECT 623.400 797.700 625.200 799.500 ;
        RECT 619.800 796.800 625.200 797.700 ;
        RECT 619.800 795.900 621.900 796.800 ;
        RECT 617.100 794.700 621.900 795.900 ;
        RECT 626.700 795.600 627.900 799.950 ;
        RECT 624.600 794.700 627.900 795.600 ;
        RECT 628.800 795.600 630.900 796.500 ;
        RECT 541.500 783.000 543.300 789.600 ;
        RECT 557.100 783.000 558.900 789.600 ;
        RECT 560.100 783.600 561.900 789.600 ;
        RECT 578.100 783.000 579.900 789.600 ;
        RECT 581.100 783.600 582.900 789.600 ;
        RECT 584.100 783.000 585.900 789.600 ;
        RECT 599.100 783.600 600.900 789.600 ;
        RECT 602.100 783.000 603.900 789.600 ;
        RECT 617.100 783.600 618.900 794.700 ;
        RECT 620.100 783.000 621.900 793.500 ;
        RECT 624.600 783.600 626.400 794.700 ;
        RECT 628.800 794.400 633.900 795.600 ;
        RECT 628.800 783.000 630.900 793.500 ;
        RECT 632.100 783.600 633.900 794.400 ;
        RECT 656.100 790.800 657.000 802.950 ;
        RECT 650.400 789.900 657.000 790.800 ;
        RECT 650.400 789.600 651.900 789.900 ;
        RECT 647.100 783.000 648.900 789.600 ;
        RECT 650.100 783.600 651.900 789.600 ;
        RECT 656.100 789.600 657.000 789.900 ;
        RECT 674.700 789.600 675.900 802.950 ;
        RECT 695.700 789.600 696.900 802.950 ;
        RECT 716.100 801.150 717.900 802.950 ;
        RECT 700.950 798.450 703.050 799.050 ;
        RECT 712.950 798.450 715.050 799.050 ;
        RECT 700.950 797.550 715.050 798.450 ;
        RECT 700.950 796.950 703.050 797.550 ;
        RECT 712.950 796.950 715.050 797.550 ;
        RECT 720.000 797.400 720.900 802.950 ;
        RECT 721.950 801.150 723.750 802.950 ;
        RECT 716.100 796.500 720.900 797.400 ;
        RECT 721.950 798.450 724.050 799.050 ;
        RECT 733.950 798.450 736.050 799.050 ;
        RECT 721.950 797.550 736.050 798.450 ;
        RECT 721.950 796.950 724.050 797.550 ;
        RECT 733.950 796.950 736.050 797.550 ;
        RECT 653.100 783.000 654.900 789.000 ;
        RECT 656.100 783.600 657.900 789.600 ;
        RECT 671.100 783.000 672.900 789.600 ;
        RECT 674.100 783.600 675.900 789.600 ;
        RECT 677.100 783.000 678.900 789.600 ;
        RECT 692.100 783.000 693.900 789.600 ;
        RECT 695.100 783.600 696.900 789.600 ;
        RECT 698.100 783.000 699.900 789.600 ;
        RECT 713.100 784.500 714.900 795.600 ;
        RECT 716.100 785.400 717.900 796.500 ;
        RECT 719.100 794.400 726.900 795.300 ;
        RECT 719.100 784.500 720.900 794.400 ;
        RECT 713.100 783.600 720.900 784.500 ;
        RECT 722.100 783.000 723.900 793.500 ;
        RECT 725.100 783.600 726.900 794.400 ;
        RECT 743.100 789.600 744.300 802.950 ;
        RECT 764.250 801.150 766.050 802.950 ;
        RECT 767.100 797.400 768.000 802.950 ;
        RECT 770.100 801.150 771.900 802.950 ;
        RECT 788.100 801.150 789.900 802.950 ;
        RECT 767.100 796.500 771.900 797.400 ;
        RECT 761.100 794.400 768.900 795.300 ;
        RECT 740.100 783.000 741.900 789.600 ;
        RECT 743.100 783.600 744.900 789.600 ;
        RECT 746.100 783.000 747.900 789.600 ;
        RECT 761.100 783.600 762.900 794.400 ;
        RECT 764.100 783.000 765.900 793.500 ;
        RECT 767.100 784.500 768.900 794.400 ;
        RECT 770.100 785.400 771.900 796.500 ;
        RECT 773.100 784.500 774.900 795.600 ;
        RECT 791.100 789.600 792.300 802.950 ;
        RECT 809.100 795.600 810.300 802.950 ;
        RECT 815.100 801.150 816.900 802.950 ;
        RECT 833.100 801.150 834.900 802.950 ;
        RECT 809.100 794.100 811.500 795.600 ;
        RECT 807.000 791.100 808.800 792.900 ;
        RECT 767.100 783.600 774.900 784.500 ;
        RECT 788.100 783.000 789.900 789.600 ;
        RECT 791.100 783.600 792.900 789.600 ;
        RECT 806.700 783.000 808.500 789.600 ;
        RECT 809.700 783.600 811.500 794.100 ;
        RECT 814.800 783.000 816.600 795.600 ;
        RECT 839.100 790.800 840.000 802.950 ;
        RECT 833.400 789.900 840.000 790.800 ;
        RECT 833.400 789.600 834.900 789.900 ;
        RECT 830.100 783.000 831.900 789.600 ;
        RECT 833.100 783.600 834.900 789.600 ;
        RECT 839.100 789.600 840.000 789.900 ;
        RECT 860.100 789.600 861.300 802.950 ;
        RECT 872.550 802.050 873.450 805.950 ;
        RECT 878.100 805.050 879.900 806.850 ;
        RECT 884.100 805.050 885.900 806.850 ;
        RECT 887.100 805.050 888.000 808.800 ;
        RECT 902.100 805.050 903.900 806.850 ;
        RECT 908.250 805.050 910.050 806.850 ;
        RECT 911.700 805.050 912.600 812.400 ;
        RECT 926.700 810.300 927.900 812.400 ;
        RECT 929.100 813.300 930.900 818.400 ;
        RECT 932.100 814.200 933.900 819.000 ;
        RECT 935.100 813.300 936.900 818.400 ;
        RECT 950.100 815.400 951.900 819.000 ;
        RECT 953.100 815.400 954.900 818.400 ;
        RECT 968.700 815.400 970.500 819.000 ;
        RECT 929.100 811.950 936.900 813.300 ;
        RECT 926.700 809.400 930.300 810.300 ;
        RECT 926.100 805.050 927.900 806.850 ;
        RECT 929.100 805.050 930.300 809.400 ;
        RECT 946.950 807.450 949.050 808.050 ;
        RECT 932.100 805.050 933.900 806.850 ;
        RECT 941.550 806.550 949.050 807.450 ;
        RECT 877.950 802.950 880.050 805.050 ;
        RECT 880.950 802.950 883.050 805.050 ;
        RECT 883.950 802.950 886.050 805.050 ;
        RECT 886.950 802.950 889.050 805.050 ;
        RECT 901.950 802.950 904.050 805.050 ;
        RECT 904.950 802.950 907.050 805.050 ;
        RECT 907.950 802.950 910.050 805.050 ;
        RECT 910.950 802.950 913.050 805.050 ;
        RECT 925.950 802.950 928.050 805.050 ;
        RECT 928.950 802.950 931.050 805.050 ;
        RECT 931.950 802.950 934.050 805.050 ;
        RECT 934.950 802.950 937.050 805.050 ;
        RECT 872.550 800.550 877.050 802.050 ;
        RECT 881.100 801.150 882.900 802.950 ;
        RECT 873.000 799.950 877.050 800.550 ;
        RECT 887.100 790.800 888.000 802.950 ;
        RECT 905.250 801.150 907.050 802.950 ;
        RECT 911.700 795.600 912.600 802.950 ;
        RECT 929.100 795.600 930.300 802.950 ;
        RECT 935.100 801.150 936.900 802.950 ;
        RECT 941.550 802.050 942.450 806.550 ;
        RECT 946.950 805.950 949.050 806.550 ;
        RECT 953.100 805.050 954.300 815.400 ;
        RECT 971.700 813.600 973.500 818.400 ;
        RECT 968.400 812.400 973.500 813.600 ;
        RECT 976.200 812.400 978.000 819.000 ;
        RECT 995.700 815.400 997.500 819.000 ;
        RECT 998.700 813.600 1000.500 818.400 ;
        RECT 995.400 812.400 1000.500 813.600 ;
        RECT 1003.200 812.400 1005.000 819.000 ;
        RECT 955.950 807.450 958.050 811.050 ;
        RECT 955.950 807.000 960.450 807.450 ;
        RECT 956.550 806.550 960.450 807.000 ;
        RECT 949.950 802.950 952.050 805.050 ;
        RECT 952.950 802.950 955.050 805.050 ;
        RECT 937.950 800.550 942.450 802.050 ;
        RECT 950.100 801.150 951.900 802.950 ;
        RECT 937.950 799.950 942.000 800.550 ;
        RECT 881.400 789.900 888.000 790.800 ;
        RECT 881.400 789.600 882.900 789.900 ;
        RECT 836.100 783.000 837.900 789.000 ;
        RECT 839.100 783.600 840.900 789.600 ;
        RECT 857.100 783.000 858.900 789.600 ;
        RECT 860.100 783.600 861.900 789.600 ;
        RECT 863.100 783.000 864.900 789.600 ;
        RECT 878.100 783.000 879.900 789.600 ;
        RECT 881.100 783.600 882.900 789.600 ;
        RECT 887.100 789.600 888.000 789.900 ;
        RECT 902.100 794.700 909.900 795.600 ;
        RECT 884.100 783.000 885.900 789.000 ;
        RECT 887.100 783.600 888.900 789.600 ;
        RECT 902.100 783.600 903.900 794.700 ;
        RECT 905.100 783.000 906.900 793.800 ;
        RECT 908.100 783.600 909.900 794.700 ;
        RECT 911.100 783.600 912.900 795.600 ;
        RECT 929.100 794.100 931.500 795.600 ;
        RECT 927.000 791.100 928.800 792.900 ;
        RECT 926.700 783.000 928.500 789.600 ;
        RECT 929.700 783.600 931.500 794.100 ;
        RECT 934.800 783.000 936.600 795.600 ;
        RECT 953.100 789.600 954.300 802.950 ;
        RECT 959.550 802.050 960.450 806.550 ;
        RECT 968.400 805.050 969.300 812.400 ;
        RECT 970.950 810.450 973.050 811.050 ;
        RECT 982.950 810.450 985.050 811.050 ;
        RECT 970.950 809.550 985.050 810.450 ;
        RECT 970.950 808.950 973.050 809.550 ;
        RECT 982.950 808.950 985.050 809.550 ;
        RECT 990.000 807.450 994.050 808.050 ;
        RECT 970.950 805.050 972.750 806.850 ;
        RECT 977.100 805.050 978.900 806.850 ;
        RECT 989.550 805.950 994.050 807.450 ;
        RECT 967.950 802.950 970.050 805.050 ;
        RECT 970.950 802.950 973.050 805.050 ;
        RECT 973.950 802.950 976.050 805.050 ;
        RECT 976.950 802.950 979.050 805.050 ;
        RECT 955.950 800.550 960.450 802.050 ;
        RECT 955.950 799.950 960.000 800.550 ;
        RECT 968.400 795.600 969.300 802.950 ;
        RECT 973.950 801.150 975.750 802.950 ;
        RECT 979.950 798.450 982.050 799.050 ;
        RECT 989.550 798.450 990.450 805.950 ;
        RECT 995.400 805.050 996.300 812.400 ;
        RECT 997.950 805.050 999.750 806.850 ;
        RECT 1004.100 805.050 1005.900 806.850 ;
        RECT 994.950 802.950 997.050 805.050 ;
        RECT 997.950 802.950 1000.050 805.050 ;
        RECT 1000.950 802.950 1003.050 805.050 ;
        RECT 1003.950 802.950 1006.050 805.050 ;
        RECT 979.950 797.550 990.450 798.450 ;
        RECT 979.950 796.950 982.050 797.550 ;
        RECT 995.400 795.600 996.300 802.950 ;
        RECT 1000.950 801.150 1002.750 802.950 ;
        RECT 950.100 783.000 951.900 789.600 ;
        RECT 953.100 783.600 954.900 789.600 ;
        RECT 968.100 783.600 969.900 795.600 ;
        RECT 971.100 794.700 978.900 795.600 ;
        RECT 971.100 783.600 972.900 794.700 ;
        RECT 974.100 783.000 975.900 793.800 ;
        RECT 977.100 783.600 978.900 794.700 ;
        RECT 995.100 783.600 996.900 795.600 ;
        RECT 998.100 794.700 1005.900 795.600 ;
        RECT 998.100 783.600 999.900 794.700 ;
        RECT 1001.100 783.000 1002.900 793.800 ;
        RECT 1004.100 783.600 1005.900 794.700 ;
        RECT 1006.950 792.450 1009.050 793.050 ;
        RECT 1012.950 792.450 1015.050 793.050 ;
        RECT 1006.950 791.550 1015.050 792.450 ;
        RECT 1006.950 790.950 1009.050 791.550 ;
        RECT 1012.950 790.950 1015.050 791.550 ;
        RECT 14.400 767.400 16.200 780.000 ;
        RECT 19.500 768.900 21.300 779.400 ;
        RECT 22.500 773.400 24.300 780.000 ;
        RECT 41.100 773.400 42.900 780.000 ;
        RECT 44.100 773.400 45.900 779.400 ;
        RECT 59.100 773.400 60.900 780.000 ;
        RECT 62.100 773.400 63.900 779.400 ;
        RECT 65.100 773.400 66.900 780.000 ;
        RECT 22.200 770.100 24.000 771.900 ;
        RECT 19.500 767.400 21.900 768.900 ;
        RECT 7.950 765.450 10.050 766.050 ;
        RECT 16.950 765.450 19.050 766.050 ;
        RECT 7.950 764.550 19.050 765.450 ;
        RECT 7.950 763.950 10.050 764.550 ;
        RECT 16.950 763.950 19.050 764.550 ;
        RECT 14.100 760.050 15.900 761.850 ;
        RECT 20.700 760.050 21.900 767.400 ;
        RECT 41.100 760.050 42.900 761.850 ;
        RECT 44.100 760.050 45.300 773.400 ;
        RECT 62.100 760.050 63.300 773.400 ;
        RECT 80.100 768.600 81.900 779.400 ;
        RECT 83.100 769.500 85.200 780.000 ;
        RECT 80.100 767.400 85.200 768.600 ;
        RECT 87.600 768.300 89.400 779.400 ;
        RECT 92.100 769.500 93.900 780.000 ;
        RECT 95.100 768.300 96.900 779.400 ;
        RECT 83.100 766.500 85.200 767.400 ;
        RECT 86.100 767.400 89.400 768.300 ;
        RECT 86.100 763.050 87.300 767.400 ;
        RECT 92.100 767.100 96.900 768.300 ;
        RECT 113.100 767.400 114.900 779.400 ;
        RECT 117.600 767.400 119.400 780.000 ;
        RECT 120.600 768.900 122.400 779.400 ;
        RECT 140.700 773.400 142.500 780.000 ;
        RECT 141.000 770.100 142.800 771.900 ;
        RECT 143.700 768.900 145.500 779.400 ;
        RECT 120.600 767.400 123.000 768.900 ;
        RECT 92.100 766.200 94.200 767.100 ;
        RECT 88.800 765.300 94.200 766.200 ;
        RECT 113.100 765.900 114.300 767.400 ;
        RECT 88.800 763.500 90.600 765.300 ;
        RECT 113.100 764.700 120.900 765.900 ;
        RECT 119.100 764.100 120.900 764.700 ;
        RECT 85.800 762.300 87.900 763.050 ;
        RECT 80.400 760.050 82.200 761.850 ;
        RECT 85.800 760.950 88.800 762.300 ;
        RECT 13.950 757.950 16.050 760.050 ;
        RECT 16.950 757.950 19.050 760.050 ;
        RECT 19.950 757.950 22.050 760.050 ;
        RECT 22.950 757.950 25.050 760.050 ;
        RECT 40.950 757.950 43.050 760.050 ;
        RECT 43.950 757.950 46.050 760.050 ;
        RECT 58.950 757.950 61.050 760.050 ;
        RECT 61.950 757.950 64.050 760.050 ;
        RECT 64.950 757.950 67.050 760.050 ;
        RECT 80.100 757.950 82.200 760.050 ;
        RECT 85.200 758.100 87.000 759.900 ;
        RECT 17.100 756.150 18.900 757.950 ;
        RECT 20.700 753.600 21.900 757.950 ;
        RECT 23.100 756.150 24.900 757.950 ;
        RECT 20.700 752.700 24.300 753.600 ;
        RECT 14.100 749.700 21.900 751.050 ;
        RECT 14.100 744.600 15.900 749.700 ;
        RECT 17.100 744.000 18.900 748.800 ;
        RECT 20.100 744.600 21.900 749.700 ;
        RECT 23.100 750.600 24.300 752.700 ;
        RECT 23.100 744.600 24.900 750.600 ;
        RECT 25.950 750.450 28.050 751.050 ;
        RECT 40.950 750.450 43.050 751.050 ;
        RECT 25.950 749.550 43.050 750.450 ;
        RECT 25.950 748.950 28.050 749.550 ;
        RECT 40.950 748.950 43.050 749.550 ;
        RECT 44.100 747.600 45.300 757.950 ;
        RECT 59.250 756.150 61.050 757.950 ;
        RECT 62.100 752.700 63.300 757.950 ;
        RECT 65.100 756.150 66.900 757.950 ;
        RECT 84.900 756.000 87.000 758.100 ;
        RECT 87.900 754.200 88.800 760.950 ;
        RECT 90.300 760.200 92.100 762.000 ;
        RECT 90.000 758.100 92.100 760.200 ;
        RECT 117.000 760.050 118.800 761.850 ;
        RECT 94.800 757.800 96.900 760.050 ;
        RECT 113.100 757.950 115.200 760.050 ;
        RECT 116.400 757.950 118.500 760.050 ;
        RECT 94.800 757.200 96.600 757.800 ;
        RECT 90.000 756.000 96.600 757.200 ;
        RECT 113.400 756.150 115.200 757.950 ;
        RECT 90.000 755.100 92.100 756.000 ;
        RECT 62.100 751.800 66.300 752.700 ;
        RECT 41.100 744.000 42.900 747.600 ;
        RECT 44.100 744.600 45.900 747.600 ;
        RECT 59.400 744.000 61.200 750.600 ;
        RECT 64.500 744.600 66.300 751.800 ;
        RECT 82.500 751.500 84.600 753.900 ;
        RECT 85.800 752.100 88.800 754.200 ;
        RECT 89.700 753.300 91.500 755.100 ;
        RECT 119.700 753.600 120.600 764.100 ;
        RECT 121.800 760.050 123.000 767.400 ;
        RECT 143.100 767.400 145.500 768.900 ;
        RECT 148.800 767.400 150.600 780.000 ;
        RECT 164.100 773.400 165.900 780.000 ;
        RECT 167.100 773.400 168.900 779.400 ;
        RECT 170.100 773.400 171.900 780.000 ;
        RECT 185.100 773.400 186.900 780.000 ;
        RECT 188.100 773.400 189.900 779.400 ;
        RECT 191.100 773.400 192.900 780.000 ;
        RECT 143.100 760.050 144.300 767.400 ;
        RECT 149.100 760.050 150.900 761.850 ;
        RECT 167.700 760.050 168.900 773.400 ;
        RECT 188.700 760.050 189.900 773.400 ;
        RECT 209.100 768.600 210.900 779.400 ;
        RECT 212.100 769.500 213.900 780.000 ;
        RECT 209.100 767.400 213.900 768.600 ;
        RECT 211.800 766.500 213.900 767.400 ;
        RECT 216.600 767.400 218.400 779.400 ;
        RECT 221.100 769.500 222.900 780.000 ;
        RECT 224.100 768.300 225.900 779.400 ;
        RECT 221.400 767.400 225.900 768.300 ;
        RECT 239.100 767.400 240.900 780.000 ;
        RECT 244.200 768.600 246.000 779.400 ;
        RECT 242.400 767.400 246.000 768.600 ;
        RECT 260.100 767.400 261.900 780.000 ;
        RECT 265.200 768.600 267.000 779.400 ;
        RECT 263.400 767.400 267.000 768.600 ;
        RECT 285.600 767.400 287.400 780.000 ;
        RECT 290.100 767.400 293.400 779.400 ;
        RECT 296.100 767.400 297.900 780.000 ;
        RECT 311.100 773.400 312.900 780.000 ;
        RECT 314.100 773.400 315.900 779.400 ;
        RECT 317.100 773.400 318.900 780.000 ;
        RECT 216.600 766.050 217.800 767.400 ;
        RECT 216.300 765.000 217.800 766.050 ;
        RECT 221.400 765.300 223.500 767.400 ;
        RECT 216.300 763.050 217.200 765.000 ;
        RECT 209.400 760.050 211.200 761.850 ;
        RECT 215.100 760.950 217.200 763.050 ;
        RECT 218.100 763.500 220.200 763.800 ;
        RECT 218.100 761.700 222.000 763.500 ;
        RECT 121.800 757.950 123.900 760.050 ;
        RECT 139.950 757.950 142.050 760.050 ;
        RECT 142.950 757.950 145.050 760.050 ;
        RECT 145.950 757.950 148.050 760.050 ;
        RECT 148.950 757.950 151.050 760.050 ;
        RECT 163.950 757.950 166.050 760.050 ;
        RECT 166.950 757.950 169.050 760.050 ;
        RECT 169.950 757.950 172.050 760.050 ;
        RECT 184.950 757.950 187.050 760.050 ;
        RECT 187.950 757.950 190.050 760.050 ;
        RECT 190.950 757.950 193.050 760.050 ;
        RECT 209.100 757.950 211.200 760.050 ;
        RECT 215.700 760.800 217.200 760.950 ;
        RECT 215.700 759.900 218.100 760.800 ;
        RECT 80.100 750.600 84.600 751.500 ;
        RECT 80.100 744.600 81.900 750.600 ;
        RECT 87.900 750.000 88.800 752.100 ;
        RECT 92.400 753.000 94.500 753.600 ;
        RECT 92.400 751.500 96.900 753.000 ;
        RECT 119.700 752.700 121.800 753.600 ;
        RECT 95.400 750.600 96.900 751.500 ;
        RECT 83.400 744.000 85.200 749.700 ;
        RECT 87.900 744.600 89.700 750.000 ;
        RECT 92.100 744.000 93.900 749.700 ;
        RECT 95.100 744.600 96.900 750.600 ;
        RECT 116.400 751.800 121.800 752.700 ;
        RECT 116.400 747.600 117.300 751.800 ;
        RECT 123.000 750.600 123.900 757.950 ;
        RECT 140.100 756.150 141.900 757.950 ;
        RECT 143.100 753.600 144.300 757.950 ;
        RECT 146.100 756.150 147.900 757.950 ;
        RECT 164.100 756.150 165.900 757.950 ;
        RECT 140.700 752.700 144.300 753.600 ;
        RECT 167.700 752.700 168.900 757.950 ;
        RECT 169.950 756.150 171.750 757.950 ;
        RECT 185.100 756.150 186.900 757.950 ;
        RECT 188.700 752.700 189.900 757.950 ;
        RECT 190.950 756.150 192.750 757.950 ;
        RECT 213.900 757.200 215.700 759.000 ;
        RECT 213.900 755.100 216.000 757.200 ;
        RECT 216.900 754.200 218.100 759.900 ;
        RECT 219.000 760.050 220.800 760.500 ;
        RECT 239.250 760.050 241.050 761.850 ;
        RECT 242.400 760.050 243.300 767.400 ;
        RECT 245.100 760.050 246.900 761.850 ;
        RECT 260.250 760.050 262.050 761.850 ;
        RECT 263.400 760.050 264.300 767.400 ;
        RECT 266.100 760.050 267.900 761.850 ;
        RECT 284.250 760.050 286.050 761.850 ;
        RECT 291.000 760.050 292.050 767.400 ;
        RECT 298.950 762.450 301.050 766.050 ;
        RECT 298.950 762.000 303.450 762.450 ;
        RECT 296.100 760.050 297.900 761.850 ;
        RECT 299.550 761.550 303.450 762.000 ;
        RECT 219.000 758.700 225.900 760.050 ;
        RECT 223.800 757.950 225.900 758.700 ;
        RECT 238.950 757.950 241.050 760.050 ;
        RECT 241.950 757.950 244.050 760.050 ;
        RECT 244.950 757.950 247.050 760.050 ;
        RECT 259.950 757.950 262.050 760.050 ;
        RECT 262.950 757.950 265.050 760.050 ;
        RECT 265.950 757.950 268.050 760.050 ;
        RECT 283.950 757.950 286.050 760.050 ;
        RECT 286.950 757.950 289.050 760.050 ;
        RECT 289.950 757.950 292.050 760.050 ;
        RECT 140.700 750.600 141.900 752.700 ;
        RECT 164.700 751.800 168.900 752.700 ;
        RECT 185.700 751.800 189.900 752.700 ;
        RECT 113.100 744.600 114.900 747.600 ;
        RECT 116.100 744.600 117.900 747.600 ;
        RECT 113.100 744.000 114.300 744.600 ;
        RECT 119.100 744.000 120.900 750.000 ;
        RECT 122.100 744.600 123.900 750.600 ;
        RECT 140.100 744.600 141.900 750.600 ;
        RECT 143.100 749.700 150.900 751.050 ;
        RECT 143.100 744.600 144.900 749.700 ;
        RECT 146.100 744.000 147.900 748.800 ;
        RECT 149.100 744.600 150.900 749.700 ;
        RECT 164.700 744.600 166.500 751.800 ;
        RECT 169.800 744.000 171.600 750.600 ;
        RECT 185.700 744.600 187.500 751.800 ;
        RECT 211.800 751.500 213.900 752.700 ;
        RECT 215.100 752.100 218.100 754.200 ;
        RECT 219.000 755.400 220.800 757.200 ;
        RECT 223.800 756.150 225.600 757.950 ;
        RECT 219.000 753.300 221.100 755.400 ;
        RECT 219.000 752.400 225.300 753.300 ;
        RECT 209.100 750.600 213.900 751.500 ;
        RECT 216.900 750.600 218.100 752.100 ;
        RECT 224.100 750.600 225.300 752.400 ;
        RECT 190.800 744.000 192.600 750.600 ;
        RECT 209.100 744.600 210.900 750.600 ;
        RECT 212.100 744.000 213.900 749.700 ;
        RECT 216.600 744.600 218.400 750.600 ;
        RECT 221.100 744.000 222.900 749.700 ;
        RECT 224.100 744.600 225.900 750.600 ;
        RECT 242.400 747.600 243.300 757.950 ;
        RECT 263.400 747.600 264.300 757.950 ;
        RECT 287.250 756.150 289.050 757.950 ;
        RECT 291.000 753.300 292.050 757.950 ;
        RECT 292.950 757.950 295.050 760.050 ;
        RECT 295.950 757.950 298.050 760.050 ;
        RECT 292.950 756.150 294.750 757.950 ;
        RECT 302.550 756.450 303.450 761.550 ;
        RECT 314.100 760.050 315.300 773.400 ;
        RECT 335.100 767.400 336.900 779.400 ;
        RECT 338.100 768.300 339.900 779.400 ;
        RECT 341.100 769.200 342.900 780.000 ;
        RECT 344.100 768.300 345.900 779.400 ;
        RECT 359.100 773.400 360.900 780.000 ;
        RECT 362.100 773.400 363.900 779.400 ;
        RECT 365.100 773.400 366.900 780.000 ;
        RECT 338.100 767.400 345.900 768.300 ;
        RECT 335.400 760.050 336.300 767.400 ;
        RECT 337.950 765.450 340.050 766.200 ;
        RECT 343.950 765.450 346.050 766.050 ;
        RECT 337.950 764.550 346.050 765.450 ;
        RECT 337.950 764.100 340.050 764.550 ;
        RECT 343.950 763.950 346.050 764.550 ;
        RECT 340.950 760.050 342.750 761.850 ;
        RECT 362.100 760.050 363.300 773.400 ;
        RECT 380.400 767.400 382.200 780.000 ;
        RECT 385.500 768.900 387.300 779.400 ;
        RECT 388.500 773.400 390.300 780.000 ;
        RECT 404.100 773.400 405.900 779.400 ;
        RECT 407.100 773.400 408.900 780.000 ;
        RECT 388.200 770.100 390.000 771.900 ;
        RECT 385.500 767.400 387.900 768.900 ;
        RECT 380.100 760.050 381.900 761.850 ;
        RECT 386.700 760.050 387.900 767.400 ;
        RECT 404.700 760.050 405.900 773.400 ;
        RECT 422.100 767.400 423.900 779.400 ;
        RECT 425.100 768.000 426.900 780.000 ;
        RECT 428.100 773.400 429.900 779.400 ;
        RECT 431.100 773.400 432.900 780.000 ;
        RECT 407.100 760.050 408.900 761.850 ;
        RECT 422.700 760.050 423.600 767.400 ;
        RECT 426.000 760.050 427.800 761.850 ;
        RECT 310.950 757.950 313.050 760.050 ;
        RECT 313.950 757.950 316.050 760.050 ;
        RECT 316.950 757.950 319.050 760.050 ;
        RECT 334.950 757.950 337.050 760.050 ;
        RECT 337.950 757.950 340.050 760.050 ;
        RECT 340.950 757.950 343.050 760.050 ;
        RECT 343.950 757.950 346.050 760.050 ;
        RECT 358.950 757.950 361.050 760.050 ;
        RECT 361.950 757.950 364.050 760.050 ;
        RECT 364.950 757.950 367.050 760.050 ;
        RECT 379.950 757.950 382.050 760.050 ;
        RECT 382.950 757.950 385.050 760.050 ;
        RECT 385.950 757.950 388.050 760.050 ;
        RECT 388.950 757.950 391.050 760.050 ;
        RECT 403.950 757.950 406.050 760.050 ;
        RECT 406.950 757.950 409.050 760.050 ;
        RECT 422.100 757.950 424.200 760.050 ;
        RECT 425.400 757.950 427.500 760.050 ;
        RECT 307.950 756.450 310.050 757.050 ;
        RECT 302.550 755.550 310.050 756.450 ;
        RECT 311.250 756.150 313.050 757.950 ;
        RECT 307.950 754.950 310.050 755.550 ;
        RECT 287.700 752.100 292.050 753.300 ;
        RECT 314.100 752.700 315.300 757.950 ;
        RECT 317.100 756.150 318.900 757.950 ;
        RECT 287.700 750.600 288.600 752.100 ;
        RECT 314.100 751.800 318.300 752.700 ;
        RECT 239.100 744.000 240.900 747.600 ;
        RECT 242.100 744.600 243.900 747.600 ;
        RECT 245.100 744.000 246.900 747.600 ;
        RECT 260.100 744.000 261.900 747.600 ;
        RECT 263.100 744.600 264.900 747.600 ;
        RECT 266.100 744.000 267.900 747.600 ;
        RECT 284.100 745.500 285.900 750.600 ;
        RECT 287.100 746.400 288.900 750.600 ;
        RECT 290.100 750.000 297.900 750.900 ;
        RECT 290.100 745.500 291.900 750.000 ;
        RECT 284.100 744.600 291.900 745.500 ;
        RECT 293.100 744.000 294.900 749.100 ;
        RECT 296.100 744.600 297.900 750.000 ;
        RECT 311.400 744.000 313.200 750.600 ;
        RECT 316.500 744.600 318.300 751.800 ;
        RECT 335.400 750.600 336.300 757.950 ;
        RECT 337.950 756.150 339.750 757.950 ;
        RECT 344.100 756.150 345.900 757.950 ;
        RECT 359.250 756.150 361.050 757.950 ;
        RECT 362.100 752.700 363.300 757.950 ;
        RECT 365.100 756.150 366.900 757.950 ;
        RECT 383.100 756.150 384.900 757.950 ;
        RECT 386.700 753.600 387.900 757.950 ;
        RECT 389.100 756.150 390.900 757.950 ;
        RECT 386.700 752.700 390.300 753.600 ;
        RECT 362.100 751.800 366.300 752.700 ;
        RECT 335.400 749.400 340.500 750.600 ;
        RECT 335.700 744.000 337.500 747.600 ;
        RECT 338.700 744.600 340.500 749.400 ;
        RECT 343.200 744.000 345.000 750.600 ;
        RECT 359.400 744.000 361.200 750.600 ;
        RECT 364.500 744.600 366.300 751.800 ;
        RECT 380.100 749.700 387.900 751.050 ;
        RECT 380.100 744.600 381.900 749.700 ;
        RECT 383.100 744.000 384.900 748.800 ;
        RECT 386.100 744.600 387.900 749.700 ;
        RECT 389.100 750.600 390.300 752.700 ;
        RECT 389.100 744.600 390.900 750.600 ;
        RECT 404.700 747.600 405.900 757.950 ;
        RECT 406.950 750.450 409.050 751.050 ;
        RECT 412.950 750.450 415.050 751.050 ;
        RECT 406.950 749.550 415.050 750.450 ;
        RECT 406.950 748.950 409.050 749.550 ;
        RECT 412.950 748.950 415.050 749.550 ;
        RECT 422.700 750.600 423.600 757.950 ;
        RECT 429.000 753.300 429.900 773.400 ;
        RECT 446.100 768.600 447.900 779.400 ;
        RECT 449.100 769.500 451.200 780.000 ;
        RECT 446.100 767.400 451.200 768.600 ;
        RECT 453.600 768.300 455.400 779.400 ;
        RECT 458.100 769.500 459.900 780.000 ;
        RECT 461.100 768.300 462.900 779.400 ;
        RECT 479.100 773.400 480.900 780.000 ;
        RECT 482.100 773.400 483.900 779.400 ;
        RECT 449.100 766.500 451.200 767.400 ;
        RECT 452.100 767.400 455.400 768.300 ;
        RECT 452.100 763.050 453.300 767.400 ;
        RECT 458.100 767.100 462.900 768.300 ;
        RECT 458.100 766.200 460.200 767.100 ;
        RECT 454.800 765.300 460.200 766.200 ;
        RECT 454.800 763.500 456.600 765.300 ;
        RECT 451.800 762.300 453.900 763.050 ;
        RECT 446.400 760.050 448.200 761.850 ;
        RECT 451.800 760.950 454.800 762.300 ;
        RECT 430.800 757.950 432.900 760.050 ;
        RECT 446.100 757.950 448.200 760.050 ;
        RECT 451.200 758.100 453.000 759.900 ;
        RECT 430.950 756.150 432.750 757.950 ;
        RECT 450.900 756.000 453.000 758.100 ;
        RECT 453.900 754.200 454.800 760.950 ;
        RECT 456.300 760.200 458.100 762.000 ;
        RECT 456.000 758.100 458.100 760.200 ;
        RECT 460.800 757.800 462.900 760.050 ;
        RECT 479.100 757.950 481.200 760.050 ;
        RECT 460.800 757.200 462.600 757.800 ;
        RECT 456.000 756.000 462.600 757.200 ;
        RECT 479.250 756.150 481.050 757.950 ;
        RECT 456.000 755.100 458.100 756.000 ;
        RECT 424.500 752.400 432.900 753.300 ;
        RECT 424.500 751.500 426.300 752.400 ;
        RECT 422.700 748.800 425.400 750.600 ;
        RECT 404.100 744.600 405.900 747.600 ;
        RECT 407.100 744.000 408.900 747.600 ;
        RECT 423.600 744.600 425.400 748.800 ;
        RECT 426.600 744.000 428.400 750.600 ;
        RECT 431.100 744.600 432.900 752.400 ;
        RECT 448.500 751.500 450.600 753.900 ;
        RECT 451.800 752.100 454.800 754.200 ;
        RECT 455.700 753.300 457.500 755.100 ;
        RECT 446.100 750.600 450.600 751.500 ;
        RECT 446.100 744.600 447.900 750.600 ;
        RECT 453.900 750.000 454.800 752.100 ;
        RECT 458.400 753.000 460.500 753.600 ;
        RECT 482.100 753.300 483.000 773.400 ;
        RECT 485.100 768.000 486.900 780.000 ;
        RECT 488.100 767.400 489.900 779.400 ;
        RECT 503.100 773.400 504.900 780.000 ;
        RECT 506.100 773.400 507.900 779.400 ;
        RECT 509.100 773.400 510.900 780.000 ;
        RECT 524.100 773.400 525.900 780.000 ;
        RECT 527.100 773.400 528.900 779.400 ;
        RECT 530.100 773.400 531.900 780.000 ;
        RECT 545.100 773.400 546.900 780.000 ;
        RECT 548.100 773.400 549.900 779.400 ;
        RECT 551.100 773.400 552.900 780.000 ;
        RECT 566.700 773.400 568.500 780.000 ;
        RECT 484.200 760.050 486.000 761.850 ;
        RECT 488.400 760.050 489.300 767.400 ;
        RECT 506.700 760.050 507.900 773.400 ;
        RECT 508.950 771.450 511.050 772.050 ;
        RECT 523.950 771.450 526.050 772.050 ;
        RECT 508.950 770.550 526.050 771.450 ;
        RECT 508.950 769.950 511.050 770.550 ;
        RECT 523.950 769.950 526.050 770.550 ;
        RECT 527.700 760.050 528.900 773.400 ;
        RECT 548.700 760.050 549.900 773.400 ;
        RECT 567.000 770.100 568.800 771.900 ;
        RECT 569.700 768.900 571.500 779.400 ;
        RECT 569.100 767.400 571.500 768.900 ;
        RECT 574.800 767.400 576.600 780.000 ;
        RECT 593.100 767.400 594.900 780.000 ;
        RECT 598.200 768.600 600.000 779.400 ;
        RECT 596.400 767.400 600.000 768.600 ;
        RECT 614.100 767.400 615.900 779.400 ;
        RECT 617.100 768.000 618.900 780.000 ;
        RECT 620.100 773.400 621.900 779.400 ;
        RECT 623.100 773.400 624.900 780.000 ;
        RECT 569.100 760.050 570.300 767.400 ;
        RECT 575.100 760.050 576.900 761.850 ;
        RECT 593.250 760.050 595.050 761.850 ;
        RECT 596.400 760.050 597.300 767.400 ;
        RECT 599.100 760.050 600.900 761.850 ;
        RECT 614.700 760.050 615.600 767.400 ;
        RECT 618.000 760.050 619.800 761.850 ;
        RECT 484.500 757.950 486.600 760.050 ;
        RECT 487.800 757.950 489.900 760.050 ;
        RECT 502.950 757.950 505.050 760.050 ;
        RECT 505.950 757.950 508.050 760.050 ;
        RECT 508.950 757.950 511.050 760.050 ;
        RECT 523.950 757.950 526.050 760.050 ;
        RECT 526.950 757.950 529.050 760.050 ;
        RECT 529.950 757.950 532.050 760.050 ;
        RECT 544.950 757.950 547.050 760.050 ;
        RECT 547.950 757.950 550.050 760.050 ;
        RECT 550.950 757.950 553.050 760.050 ;
        RECT 565.950 757.950 568.050 760.050 ;
        RECT 568.950 757.950 571.050 760.050 ;
        RECT 571.950 757.950 574.050 760.050 ;
        RECT 574.950 757.950 577.050 760.050 ;
        RECT 592.950 757.950 595.050 760.050 ;
        RECT 595.950 757.950 598.050 760.050 ;
        RECT 598.950 757.950 601.050 760.050 ;
        RECT 614.100 757.950 616.200 760.050 ;
        RECT 617.400 757.950 619.500 760.050 ;
        RECT 458.400 751.500 462.900 753.000 ;
        RECT 461.400 750.600 462.900 751.500 ;
        RECT 449.400 744.000 451.200 749.700 ;
        RECT 453.900 744.600 455.700 750.000 ;
        RECT 458.100 744.000 459.900 749.700 ;
        RECT 461.100 744.600 462.900 750.600 ;
        RECT 479.100 752.400 487.500 753.300 ;
        RECT 479.100 744.600 480.900 752.400 ;
        RECT 485.700 751.500 487.500 752.400 ;
        RECT 488.400 750.600 489.300 757.950 ;
        RECT 503.100 756.150 504.900 757.950 ;
        RECT 506.700 752.700 507.900 757.950 ;
        RECT 508.950 756.150 510.750 757.950 ;
        RECT 524.100 756.150 525.900 757.950 ;
        RECT 527.700 752.700 528.900 757.950 ;
        RECT 529.950 756.150 531.750 757.950 ;
        RECT 545.100 756.150 546.900 757.950 ;
        RECT 548.700 752.700 549.900 757.950 ;
        RECT 550.950 756.150 552.750 757.950 ;
        RECT 566.100 756.150 567.900 757.950 ;
        RECT 569.100 753.600 570.300 757.950 ;
        RECT 572.100 756.150 573.900 757.950 ;
        RECT 483.600 744.000 485.400 750.600 ;
        RECT 486.600 748.800 489.300 750.600 ;
        RECT 503.700 751.800 507.900 752.700 ;
        RECT 524.700 751.800 528.900 752.700 ;
        RECT 545.700 751.800 549.900 752.700 ;
        RECT 566.700 752.700 570.300 753.600 ;
        RECT 586.950 753.450 589.050 754.050 ;
        RECT 592.950 753.450 595.050 754.050 ;
        RECT 486.600 744.600 488.400 748.800 ;
        RECT 503.700 744.600 505.500 751.800 ;
        RECT 508.800 744.000 510.600 750.600 ;
        RECT 524.700 744.600 526.500 751.800 ;
        RECT 529.800 744.000 531.600 750.600 ;
        RECT 545.700 744.600 547.500 751.800 ;
        RECT 566.700 750.600 567.900 752.700 ;
        RECT 586.950 752.550 595.050 753.450 ;
        RECT 586.950 751.950 589.050 752.550 ;
        RECT 592.950 751.950 595.050 752.550 ;
        RECT 550.800 744.000 552.600 750.600 ;
        RECT 566.100 744.600 567.900 750.600 ;
        RECT 569.100 749.700 576.900 751.050 ;
        RECT 569.100 744.600 570.900 749.700 ;
        RECT 572.100 744.000 573.900 748.800 ;
        RECT 575.100 744.600 576.900 749.700 ;
        RECT 596.400 747.600 597.300 757.950 ;
        RECT 614.700 750.600 615.600 757.950 ;
        RECT 621.000 753.300 621.900 773.400 ;
        RECT 641.100 767.400 642.900 779.400 ;
        RECT 644.100 768.300 645.900 779.400 ;
        RECT 647.100 769.200 648.900 780.000 ;
        RECT 650.100 768.300 651.900 779.400 ;
        RECT 668.100 773.400 669.900 779.400 ;
        RECT 671.100 774.000 672.900 780.000 ;
        RECT 644.100 767.400 651.900 768.300 ;
        RECT 669.000 773.100 669.900 773.400 ;
        RECT 674.100 773.400 675.900 779.400 ;
        RECT 677.100 773.400 678.900 780.000 ;
        RECT 695.100 773.400 696.900 780.000 ;
        RECT 698.100 773.400 699.900 779.400 ;
        RECT 713.100 773.400 714.900 780.000 ;
        RECT 716.100 773.400 717.900 779.400 ;
        RECT 719.100 774.000 720.900 780.000 ;
        RECT 674.100 773.100 675.600 773.400 ;
        RECT 669.000 772.200 675.600 773.100 ;
        RECT 641.400 760.050 642.300 767.400 ;
        RECT 646.950 760.050 648.750 761.850 ;
        RECT 669.000 760.050 669.900 772.200 ;
        RECT 690.000 762.450 694.050 763.050 ;
        RECT 674.100 760.050 675.900 761.850 ;
        RECT 689.550 760.950 694.050 762.450 ;
        RECT 622.800 757.950 624.900 760.050 ;
        RECT 640.950 757.950 643.050 760.050 ;
        RECT 643.950 757.950 646.050 760.050 ;
        RECT 646.950 757.950 649.050 760.050 ;
        RECT 649.950 757.950 652.050 760.050 ;
        RECT 667.950 757.950 670.050 760.050 ;
        RECT 670.950 757.950 673.050 760.050 ;
        RECT 673.950 757.950 676.050 760.050 ;
        RECT 676.950 757.950 679.050 760.050 ;
        RECT 622.950 756.150 624.750 757.950 ;
        RECT 616.500 752.400 624.900 753.300 ;
        RECT 616.500 751.500 618.300 752.400 ;
        RECT 614.700 748.800 617.400 750.600 ;
        RECT 593.100 744.000 594.900 747.600 ;
        RECT 596.100 744.600 597.900 747.600 ;
        RECT 599.100 744.000 600.900 747.600 ;
        RECT 615.600 744.600 617.400 748.800 ;
        RECT 618.600 744.000 620.400 750.600 ;
        RECT 623.100 744.600 624.900 752.400 ;
        RECT 641.400 750.600 642.300 757.950 ;
        RECT 643.950 756.150 645.750 757.950 ;
        RECT 650.100 756.150 651.900 757.950 ;
        RECT 669.000 754.200 669.900 757.950 ;
        RECT 671.100 756.150 672.900 757.950 ;
        RECT 677.100 756.150 678.900 757.950 ;
        RECT 679.950 756.450 682.050 757.050 ;
        RECT 689.550 756.450 690.450 760.950 ;
        RECT 695.100 760.050 696.900 761.850 ;
        RECT 698.100 760.050 699.300 773.400 ;
        RECT 716.400 773.100 717.900 773.400 ;
        RECT 722.100 773.400 723.900 779.400 ;
        RECT 740.100 773.400 741.900 780.000 ;
        RECT 743.100 773.400 744.900 779.400 ;
        RECT 722.100 773.100 723.000 773.400 ;
        RECT 716.400 772.200 723.000 773.100 ;
        RECT 700.950 765.450 703.050 766.050 ;
        RECT 718.950 765.450 721.050 766.050 ;
        RECT 700.950 764.550 721.050 765.450 ;
        RECT 700.950 763.950 703.050 764.550 ;
        RECT 718.950 763.950 721.050 764.550 ;
        RECT 716.100 760.050 717.900 761.850 ;
        RECT 722.100 760.050 723.000 772.200 ;
        RECT 733.950 765.450 736.050 766.050 ;
        RECT 739.950 765.450 742.050 766.050 ;
        RECT 733.950 764.550 742.050 765.450 ;
        RECT 733.950 763.950 736.050 764.550 ;
        RECT 739.950 763.950 742.050 764.550 ;
        RECT 694.950 757.950 697.050 760.050 ;
        RECT 697.950 757.950 700.050 760.050 ;
        RECT 712.950 757.950 715.050 760.050 ;
        RECT 715.950 757.950 718.050 760.050 ;
        RECT 718.950 757.950 721.050 760.050 ;
        RECT 721.950 757.950 724.050 760.050 ;
        RECT 740.100 757.950 742.200 760.050 ;
        RECT 679.950 755.550 690.450 756.450 ;
        RECT 679.950 754.950 682.050 755.550 ;
        RECT 669.000 753.000 672.300 754.200 ;
        RECT 641.400 749.400 646.500 750.600 ;
        RECT 641.700 744.000 643.500 747.600 ;
        RECT 644.700 744.600 646.500 749.400 ;
        RECT 649.200 744.000 651.000 750.600 ;
        RECT 670.500 744.600 672.300 753.000 ;
        RECT 677.100 744.000 678.900 753.600 ;
        RECT 698.100 747.600 699.300 757.950 ;
        RECT 713.100 756.150 714.900 757.950 ;
        RECT 719.100 756.150 720.900 757.950 ;
        RECT 722.100 754.200 723.000 757.950 ;
        RECT 740.250 756.150 742.050 757.950 ;
        RECT 695.100 744.000 696.900 747.600 ;
        RECT 698.100 744.600 699.900 747.600 ;
        RECT 713.100 744.000 714.900 753.600 ;
        RECT 719.700 753.000 723.000 754.200 ;
        RECT 743.100 753.300 744.000 773.400 ;
        RECT 746.100 768.000 747.900 780.000 ;
        RECT 749.100 767.400 750.900 779.400 ;
        RECT 764.100 773.400 765.900 780.000 ;
        RECT 767.100 773.400 768.900 779.400 ;
        RECT 770.100 774.000 771.900 780.000 ;
        RECT 767.400 773.100 768.900 773.400 ;
        RECT 773.100 773.400 774.900 779.400 ;
        RECT 773.100 773.100 774.000 773.400 ;
        RECT 767.400 772.200 774.000 773.100 ;
        RECT 745.200 760.050 747.000 761.850 ;
        RECT 749.400 760.050 750.300 767.400 ;
        RECT 757.950 765.450 760.050 766.050 ;
        RECT 769.950 765.450 772.050 766.050 ;
        RECT 757.950 764.550 772.050 765.450 ;
        RECT 757.950 763.950 760.050 764.550 ;
        RECT 769.950 763.950 772.050 764.550 ;
        RECT 767.100 760.050 768.900 761.850 ;
        RECT 773.100 760.050 774.000 772.200 ;
        RECT 788.400 767.400 790.200 780.000 ;
        RECT 793.500 768.900 795.300 779.400 ;
        RECT 796.500 773.400 798.300 780.000 ;
        RECT 815.100 773.400 816.900 780.000 ;
        RECT 818.100 773.400 819.900 779.400 ;
        RECT 821.100 774.000 822.900 780.000 ;
        RECT 818.400 773.100 819.900 773.400 ;
        RECT 824.100 773.400 825.900 779.400 ;
        RECT 839.100 773.400 840.900 780.000 ;
        RECT 842.100 773.400 843.900 779.400 ;
        RECT 845.100 773.400 846.900 780.000 ;
        RECT 824.100 773.100 825.000 773.400 ;
        RECT 818.400 772.200 825.000 773.100 ;
        RECT 796.200 770.100 798.000 771.900 ;
        RECT 793.500 767.400 795.900 768.900 ;
        RECT 788.100 760.050 789.900 761.850 ;
        RECT 794.700 760.050 795.900 767.400 ;
        RECT 818.100 760.050 819.900 761.850 ;
        RECT 824.100 760.050 825.000 772.200 ;
        RECT 842.100 760.050 843.300 773.400 ;
        RECT 860.100 767.400 861.900 779.400 ;
        RECT 863.100 768.000 864.900 780.000 ;
        RECT 866.100 773.400 867.900 779.400 ;
        RECT 869.100 773.400 870.900 780.000 ;
        RECT 844.950 765.450 847.050 766.050 ;
        RECT 856.950 765.450 859.050 766.050 ;
        RECT 844.950 764.550 859.050 765.450 ;
        RECT 844.950 763.950 847.050 764.550 ;
        RECT 856.950 763.950 859.050 764.550 ;
        RECT 860.700 760.050 861.600 767.400 ;
        RECT 864.000 760.050 865.800 761.850 ;
        RECT 745.500 757.950 747.600 760.050 ;
        RECT 748.800 757.950 750.900 760.050 ;
        RECT 763.950 757.950 766.050 760.050 ;
        RECT 766.950 757.950 769.050 760.050 ;
        RECT 769.950 757.950 772.050 760.050 ;
        RECT 772.950 757.950 775.050 760.050 ;
        RECT 787.950 757.950 790.050 760.050 ;
        RECT 790.950 757.950 793.050 760.050 ;
        RECT 793.950 757.950 796.050 760.050 ;
        RECT 796.950 757.950 799.050 760.050 ;
        RECT 814.950 757.950 817.050 760.050 ;
        RECT 817.950 757.950 820.050 760.050 ;
        RECT 820.950 757.950 823.050 760.050 ;
        RECT 823.950 757.950 826.050 760.050 ;
        RECT 838.950 757.950 841.050 760.050 ;
        RECT 841.950 757.950 844.050 760.050 ;
        RECT 844.950 757.950 847.050 760.050 ;
        RECT 860.100 757.950 862.200 760.050 ;
        RECT 863.400 757.950 865.500 760.050 ;
        RECT 719.700 744.600 721.500 753.000 ;
        RECT 740.100 752.400 748.500 753.300 ;
        RECT 740.100 744.600 741.900 752.400 ;
        RECT 746.700 751.500 748.500 752.400 ;
        RECT 749.400 750.600 750.300 757.950 ;
        RECT 764.100 756.150 765.900 757.950 ;
        RECT 770.100 756.150 771.900 757.950 ;
        RECT 773.100 754.200 774.000 757.950 ;
        RECT 791.100 756.150 792.900 757.950 ;
        RECT 744.600 744.000 746.400 750.600 ;
        RECT 747.600 748.800 750.300 750.600 ;
        RECT 747.600 744.600 749.400 748.800 ;
        RECT 764.100 744.000 765.900 753.600 ;
        RECT 770.700 753.000 774.000 754.200 ;
        RECT 794.700 753.600 795.900 757.950 ;
        RECT 797.100 756.150 798.900 757.950 ;
        RECT 799.950 756.450 802.050 757.050 ;
        RECT 805.950 756.450 808.050 757.050 ;
        RECT 799.950 755.550 808.050 756.450 ;
        RECT 815.100 756.150 816.900 757.950 ;
        RECT 821.100 756.150 822.900 757.950 ;
        RECT 799.950 754.950 802.050 755.550 ;
        RECT 805.950 754.950 808.050 755.550 ;
        RECT 824.100 754.200 825.000 757.950 ;
        RECT 839.250 756.150 841.050 757.950 ;
        RECT 770.700 744.600 772.500 753.000 ;
        RECT 794.700 752.700 798.300 753.600 ;
        RECT 788.100 749.700 795.900 751.050 ;
        RECT 788.100 744.600 789.900 749.700 ;
        RECT 791.100 744.000 792.900 748.800 ;
        RECT 794.100 744.600 795.900 749.700 ;
        RECT 797.100 750.600 798.300 752.700 ;
        RECT 797.100 744.600 798.900 750.600 ;
        RECT 815.100 744.000 816.900 753.600 ;
        RECT 821.700 753.000 825.000 754.200 ;
        RECT 821.700 744.600 823.500 753.000 ;
        RECT 842.100 752.700 843.300 757.950 ;
        RECT 845.100 756.150 846.900 757.950 ;
        RECT 842.100 751.800 846.300 752.700 ;
        RECT 839.400 744.000 841.200 750.600 ;
        RECT 844.500 744.600 846.300 751.800 ;
        RECT 860.700 750.600 861.600 757.950 ;
        RECT 867.000 753.300 867.900 773.400 ;
        RECT 887.100 767.400 888.900 779.400 ;
        RECT 890.100 768.300 891.900 779.400 ;
        RECT 893.100 769.200 894.900 780.000 ;
        RECT 896.100 768.300 897.900 779.400 ;
        RECT 914.700 773.400 916.500 780.000 ;
        RECT 915.000 770.100 916.800 771.900 ;
        RECT 917.700 768.900 919.500 779.400 ;
        RECT 890.100 767.400 897.900 768.300 ;
        RECT 917.100 767.400 919.500 768.900 ;
        RECT 922.800 767.400 924.600 780.000 ;
        RECT 941.100 768.300 942.900 779.400 ;
        RECT 944.100 769.200 945.900 780.000 ;
        RECT 947.100 768.300 948.900 779.400 ;
        RECT 941.100 767.400 948.900 768.300 ;
        RECT 950.100 767.400 951.900 779.400 ;
        RECT 968.100 768.300 969.900 779.400 ;
        RECT 971.100 769.200 972.900 780.000 ;
        RECT 974.100 768.300 975.900 779.400 ;
        RECT 968.100 767.400 975.900 768.300 ;
        RECT 977.100 767.400 978.900 779.400 ;
        RECT 992.700 773.400 994.500 780.000 ;
        RECT 993.000 770.100 994.800 771.900 ;
        RECT 995.700 768.900 997.500 779.400 ;
        RECT 995.100 767.400 997.500 768.900 ;
        RECT 1000.800 767.400 1002.600 780.000 ;
        RECT 887.400 760.050 888.300 767.400 ;
        RECT 889.950 765.450 892.050 766.050 ;
        RECT 901.950 765.450 904.050 766.050 ;
        RECT 889.950 764.550 904.050 765.450 ;
        RECT 889.950 763.950 892.050 764.550 ;
        RECT 901.950 763.950 904.050 764.550 ;
        RECT 892.950 760.050 894.750 761.850 ;
        RECT 917.100 760.050 918.300 767.400 ;
        RECT 919.950 765.450 922.050 766.200 ;
        RECT 928.950 765.450 931.050 766.050 ;
        RECT 919.950 764.550 931.050 765.450 ;
        RECT 919.950 764.100 922.050 764.550 ;
        RECT 928.950 763.950 931.050 764.550 ;
        RECT 925.950 762.450 930.000 763.050 ;
        RECT 923.100 760.050 924.900 761.850 ;
        RECT 925.950 760.950 930.450 762.450 ;
        RECT 868.800 757.950 870.900 760.050 ;
        RECT 886.950 757.950 889.050 760.050 ;
        RECT 889.950 757.950 892.050 760.050 ;
        RECT 892.950 757.950 895.050 760.050 ;
        RECT 895.950 757.950 898.050 760.050 ;
        RECT 913.950 757.950 916.050 760.050 ;
        RECT 916.950 757.950 919.050 760.050 ;
        RECT 919.950 757.950 922.050 760.050 ;
        RECT 922.950 757.950 925.050 760.050 ;
        RECT 868.950 756.150 870.750 757.950 ;
        RECT 862.500 752.400 870.900 753.300 ;
        RECT 862.500 751.500 864.300 752.400 ;
        RECT 860.700 748.800 863.400 750.600 ;
        RECT 861.600 744.600 863.400 748.800 ;
        RECT 864.600 744.000 866.400 750.600 ;
        RECT 869.100 744.600 870.900 752.400 ;
        RECT 887.400 750.600 888.300 757.950 ;
        RECT 889.950 756.150 891.750 757.950 ;
        RECT 896.100 756.150 897.900 757.950 ;
        RECT 914.100 756.150 915.900 757.950 ;
        RECT 917.100 753.600 918.300 757.950 ;
        RECT 920.100 756.150 921.900 757.950 ;
        RECT 929.550 757.050 930.450 760.950 ;
        RECT 944.250 760.050 946.050 761.850 ;
        RECT 950.700 760.050 951.600 767.400 ;
        RECT 971.250 760.050 973.050 761.850 ;
        RECT 977.700 760.050 978.600 767.400 ;
        RECT 995.100 760.050 996.300 767.400 ;
        RECT 1001.100 760.050 1002.900 761.850 ;
        RECT 940.950 757.950 943.050 760.050 ;
        RECT 943.950 757.950 946.050 760.050 ;
        RECT 946.950 757.950 949.050 760.050 ;
        RECT 949.950 757.950 952.050 760.050 ;
        RECT 967.950 757.950 970.050 760.050 ;
        RECT 970.950 757.950 973.050 760.050 ;
        RECT 973.950 757.950 976.050 760.050 ;
        RECT 976.950 757.950 979.050 760.050 ;
        RECT 991.950 757.950 994.050 760.050 ;
        RECT 994.950 757.950 997.050 760.050 ;
        RECT 997.950 757.950 1000.050 760.050 ;
        RECT 1000.950 757.950 1003.050 760.050 ;
        RECT 925.950 755.550 930.450 757.050 ;
        RECT 941.100 756.150 942.900 757.950 ;
        RECT 947.250 756.150 949.050 757.950 ;
        RECT 925.950 754.950 930.000 755.550 ;
        RECT 914.700 752.700 918.300 753.600 ;
        RECT 914.700 750.600 915.900 752.700 ;
        RECT 887.400 749.400 892.500 750.600 ;
        RECT 887.700 744.000 889.500 747.600 ;
        RECT 890.700 744.600 892.500 749.400 ;
        RECT 895.200 744.000 897.000 750.600 ;
        RECT 914.100 744.600 915.900 750.600 ;
        RECT 917.100 749.700 924.900 751.050 ;
        RECT 950.700 750.600 951.600 757.950 ;
        RECT 968.100 756.150 969.900 757.950 ;
        RECT 974.250 756.150 976.050 757.950 ;
        RECT 977.700 750.600 978.600 757.950 ;
        RECT 992.100 756.150 993.900 757.950 ;
        RECT 995.100 753.600 996.300 757.950 ;
        RECT 998.100 756.150 999.900 757.950 ;
        RECT 992.700 752.700 996.300 753.600 ;
        RECT 992.700 750.600 993.900 752.700 ;
        RECT 917.100 744.600 918.900 749.700 ;
        RECT 920.100 744.000 921.900 748.800 ;
        RECT 923.100 744.600 924.900 749.700 ;
        RECT 942.000 744.000 943.800 750.600 ;
        RECT 946.500 749.400 951.600 750.600 ;
        RECT 946.500 744.600 948.300 749.400 ;
        RECT 949.500 744.000 951.300 747.600 ;
        RECT 969.000 744.000 970.800 750.600 ;
        RECT 973.500 749.400 978.600 750.600 ;
        RECT 973.500 744.600 975.300 749.400 ;
        RECT 976.500 744.000 978.300 747.600 ;
        RECT 992.100 744.600 993.900 750.600 ;
        RECT 995.100 749.700 1002.900 751.050 ;
        RECT 995.100 744.600 996.900 749.700 ;
        RECT 998.100 744.000 999.900 748.800 ;
        RECT 1001.100 744.600 1002.900 749.700 ;
        RECT 14.400 734.400 16.200 741.000 ;
        RECT 19.500 733.200 21.300 740.400 ;
        RECT 35.100 737.400 36.900 741.000 ;
        RECT 38.100 737.400 39.900 740.400 ;
        RECT 17.100 732.300 21.300 733.200 ;
        RECT 14.250 727.050 16.050 728.850 ;
        RECT 17.100 727.050 18.300 732.300 ;
        RECT 20.100 727.050 21.900 728.850 ;
        RECT 38.100 727.050 39.300 737.400 ;
        RECT 53.400 734.400 55.200 741.000 ;
        RECT 58.500 733.200 60.300 740.400 ;
        RECT 74.400 734.400 76.200 741.000 ;
        RECT 79.500 733.200 81.300 740.400 ;
        RECT 56.100 732.300 60.300 733.200 ;
        RECT 77.100 732.300 81.300 733.200 ;
        RECT 98.700 733.200 100.500 740.400 ;
        RECT 103.800 734.400 105.600 741.000 ;
        RECT 119.100 734.400 120.900 740.400 ;
        RECT 98.700 732.300 102.900 733.200 ;
        RECT 53.250 727.050 55.050 728.850 ;
        RECT 56.100 727.050 57.300 732.300 ;
        RECT 59.100 727.050 60.900 728.850 ;
        RECT 74.250 727.050 76.050 728.850 ;
        RECT 77.100 727.050 78.300 732.300 ;
        RECT 80.100 727.050 81.900 728.850 ;
        RECT 98.100 727.050 99.900 728.850 ;
        RECT 101.700 727.050 102.900 732.300 ;
        RECT 103.950 732.450 106.050 733.050 ;
        RECT 109.950 732.450 112.050 733.050 ;
        RECT 103.950 731.550 112.050 732.450 ;
        RECT 103.950 730.950 106.050 731.550 ;
        RECT 109.950 730.950 112.050 731.550 ;
        RECT 119.700 732.300 120.900 734.400 ;
        RECT 122.100 735.300 123.900 740.400 ;
        RECT 125.100 736.200 126.900 741.000 ;
        RECT 128.100 735.300 129.900 740.400 ;
        RECT 122.100 733.950 129.900 735.300 ;
        RECT 146.400 734.400 148.200 741.000 ;
        RECT 167.100 740.400 168.300 741.000 ;
        RECT 151.500 733.200 153.300 740.400 ;
        RECT 167.100 737.400 168.900 740.400 ;
        RECT 170.100 737.400 171.900 740.400 ;
        RECT 149.100 732.300 153.300 733.200 ;
        RECT 170.400 733.200 171.300 737.400 ;
        RECT 173.100 735.000 174.900 741.000 ;
        RECT 176.100 734.400 177.900 740.400 ;
        RECT 170.400 732.300 175.800 733.200 ;
        RECT 119.700 731.400 123.300 732.300 ;
        RECT 103.950 727.050 105.750 728.850 ;
        RECT 119.100 727.050 120.900 728.850 ;
        RECT 122.100 727.050 123.300 731.400 ;
        RECT 125.100 727.050 126.900 728.850 ;
        RECT 146.250 727.050 148.050 728.850 ;
        RECT 149.100 727.050 150.300 732.300 ;
        RECT 173.700 731.400 175.800 732.300 ;
        RECT 152.100 727.050 153.900 728.850 ;
        RECT 167.400 727.050 169.200 728.850 ;
        RECT 13.950 724.950 16.050 727.050 ;
        RECT 16.950 724.950 19.050 727.050 ;
        RECT 19.950 724.950 22.050 727.050 ;
        RECT 34.950 724.950 37.050 727.050 ;
        RECT 37.950 724.950 40.050 727.050 ;
        RECT 52.950 724.950 55.050 727.050 ;
        RECT 55.950 724.950 58.050 727.050 ;
        RECT 58.950 724.950 61.050 727.050 ;
        RECT 73.950 724.950 76.050 727.050 ;
        RECT 76.950 724.950 79.050 727.050 ;
        RECT 79.950 724.950 82.050 727.050 ;
        RECT 97.950 724.950 100.050 727.050 ;
        RECT 100.950 724.950 103.050 727.050 ;
        RECT 103.950 724.950 106.050 727.050 ;
        RECT 118.950 724.950 121.050 727.050 ;
        RECT 121.950 724.950 124.050 727.050 ;
        RECT 124.950 724.950 127.050 727.050 ;
        RECT 127.950 724.950 130.050 727.050 ;
        RECT 145.950 724.950 148.050 727.050 ;
        RECT 148.950 724.950 151.050 727.050 ;
        RECT 151.950 724.950 154.050 727.050 ;
        RECT 167.100 724.950 169.200 727.050 ;
        RECT 170.400 724.950 172.500 727.050 ;
        RECT 17.100 711.600 18.300 724.950 ;
        RECT 35.100 723.150 36.900 724.950 ;
        RECT 38.100 711.600 39.300 724.950 ;
        RECT 56.100 711.600 57.300 724.950 ;
        RECT 77.100 711.600 78.300 724.950 ;
        RECT 101.700 711.600 102.900 724.950 ;
        RECT 109.950 720.450 112.050 721.050 ;
        RECT 118.950 720.450 121.050 721.050 ;
        RECT 109.950 719.550 121.050 720.450 ;
        RECT 109.950 718.950 112.050 719.550 ;
        RECT 118.950 718.950 121.050 719.550 ;
        RECT 122.100 717.600 123.300 724.950 ;
        RECT 128.100 723.150 129.900 724.950 ;
        RECT 122.100 716.100 124.500 717.600 ;
        RECT 120.000 713.100 121.800 714.900 ;
        RECT 14.100 705.000 15.900 711.600 ;
        RECT 17.100 705.600 18.900 711.600 ;
        RECT 20.100 705.000 21.900 711.600 ;
        RECT 35.100 705.000 36.900 711.600 ;
        RECT 38.100 705.600 39.900 711.600 ;
        RECT 53.100 705.000 54.900 711.600 ;
        RECT 56.100 705.600 57.900 711.600 ;
        RECT 59.100 705.000 60.900 711.600 ;
        RECT 74.100 705.000 75.900 711.600 ;
        RECT 77.100 705.600 78.900 711.600 ;
        RECT 80.100 705.000 81.900 711.600 ;
        RECT 98.100 705.000 99.900 711.600 ;
        RECT 101.100 705.600 102.900 711.600 ;
        RECT 104.100 705.000 105.900 711.600 ;
        RECT 119.700 705.000 121.500 711.600 ;
        RECT 122.700 705.600 124.500 716.100 ;
        RECT 127.800 705.000 129.600 717.600 ;
        RECT 149.100 711.600 150.300 724.950 ;
        RECT 171.000 723.150 172.800 724.950 ;
        RECT 173.700 720.900 174.600 731.400 ;
        RECT 177.000 727.050 177.900 734.400 ;
        RECT 191.100 735.300 192.900 740.400 ;
        RECT 194.100 736.200 195.900 741.000 ;
        RECT 197.100 735.300 198.900 740.400 ;
        RECT 191.100 733.950 198.900 735.300 ;
        RECT 200.100 734.400 201.900 740.400 ;
        RECT 200.100 732.300 201.300 734.400 ;
        RECT 197.700 731.400 201.300 732.300 ;
        RECT 215.100 732.600 216.900 740.400 ;
        RECT 219.600 734.400 221.400 741.000 ;
        RECT 222.600 736.200 224.400 740.400 ;
        RECT 222.600 734.400 225.300 736.200 ;
        RECT 239.100 734.400 240.900 740.400 ;
        RECT 221.700 732.600 223.500 733.500 ;
        RECT 215.100 731.700 223.500 732.600 ;
        RECT 194.100 727.050 195.900 728.850 ;
        RECT 197.700 727.050 198.900 731.400 ;
        RECT 200.100 727.050 201.900 728.850 ;
        RECT 215.250 727.050 217.050 728.850 ;
        RECT 175.800 724.950 177.900 727.050 ;
        RECT 190.950 724.950 193.050 727.050 ;
        RECT 193.950 724.950 196.050 727.050 ;
        RECT 196.950 724.950 199.050 727.050 ;
        RECT 199.950 724.950 202.050 727.050 ;
        RECT 215.100 724.950 217.200 727.050 ;
        RECT 173.100 720.300 174.900 720.900 ;
        RECT 167.100 719.100 174.900 720.300 ;
        RECT 167.100 717.600 168.300 719.100 ;
        RECT 175.800 717.600 177.000 724.950 ;
        RECT 191.100 723.150 192.900 724.950 ;
        RECT 197.700 717.600 198.900 724.950 ;
        RECT 146.100 705.000 147.900 711.600 ;
        RECT 149.100 705.600 150.900 711.600 ;
        RECT 152.100 705.000 153.900 711.600 ;
        RECT 167.100 705.600 168.900 717.600 ;
        RECT 171.600 705.000 173.400 717.600 ;
        RECT 174.600 716.100 177.000 717.600 ;
        RECT 174.600 705.600 176.400 716.100 ;
        RECT 191.400 705.000 193.200 717.600 ;
        RECT 196.500 716.100 198.900 717.600 ;
        RECT 196.500 705.600 198.300 716.100 ;
        RECT 199.200 713.100 201.000 714.900 ;
        RECT 218.100 711.600 219.000 731.700 ;
        RECT 224.400 727.050 225.300 734.400 ;
        RECT 239.700 732.300 240.900 734.400 ;
        RECT 242.100 735.300 243.900 740.400 ;
        RECT 245.100 736.200 246.900 741.000 ;
        RECT 248.100 735.300 249.900 740.400 ;
        RECT 242.100 733.950 249.900 735.300 ;
        RECT 263.100 734.400 264.900 740.400 ;
        RECT 266.100 735.300 267.900 741.000 ;
        RECT 270.600 734.400 272.400 740.400 ;
        RECT 275.100 735.300 276.900 741.000 ;
        RECT 278.100 734.400 279.900 740.400 ;
        RECT 296.100 737.400 297.900 741.000 ;
        RECT 299.100 737.400 300.900 740.400 ;
        RECT 302.100 737.400 303.900 741.000 ;
        RECT 239.700 731.400 243.300 732.300 ;
        RECT 239.100 727.050 240.900 728.850 ;
        RECT 242.100 727.050 243.300 731.400 ;
        RECT 259.950 730.950 262.050 733.050 ;
        RECT 263.700 732.600 264.900 734.400 ;
        RECT 270.900 732.900 272.100 734.400 ;
        RECT 275.100 733.500 279.900 734.400 ;
        RECT 263.700 731.700 270.000 732.600 ;
        RECT 245.100 727.050 246.900 728.850 ;
        RECT 220.500 724.950 222.600 727.050 ;
        RECT 223.800 724.950 225.900 727.050 ;
        RECT 238.950 724.950 241.050 727.050 ;
        RECT 241.950 724.950 244.050 727.050 ;
        RECT 244.950 724.950 247.050 727.050 ;
        RECT 247.950 724.950 250.050 727.050 ;
        RECT 220.200 723.150 222.000 724.950 ;
        RECT 224.400 717.600 225.300 724.950 ;
        RECT 242.100 717.600 243.300 724.950 ;
        RECT 248.100 723.150 249.900 724.950 ;
        RECT 199.500 705.000 201.300 711.600 ;
        RECT 215.100 705.000 216.900 711.600 ;
        RECT 218.100 705.600 219.900 711.600 ;
        RECT 221.100 705.000 222.900 717.000 ;
        RECT 224.100 705.600 225.900 717.600 ;
        RECT 242.100 716.100 244.500 717.600 ;
        RECT 240.000 713.100 241.800 714.900 ;
        RECT 239.700 705.000 241.500 711.600 ;
        RECT 242.700 705.600 244.500 716.100 ;
        RECT 247.800 705.000 249.600 717.600 ;
        RECT 260.550 714.900 261.450 730.950 ;
        RECT 267.900 729.600 270.000 731.700 ;
        RECT 263.400 727.050 265.200 728.850 ;
        RECT 268.200 727.800 270.000 729.600 ;
        RECT 270.900 730.800 273.900 732.900 ;
        RECT 275.100 732.300 277.200 733.500 ;
        RECT 263.100 726.300 265.200 727.050 ;
        RECT 263.100 724.950 270.000 726.300 ;
        RECT 268.200 724.500 270.000 724.950 ;
        RECT 270.900 725.100 272.100 730.800 ;
        RECT 273.000 727.800 275.100 729.900 ;
        RECT 273.300 726.000 275.100 727.800 ;
        RECT 299.400 727.050 300.300 737.400 ;
        RECT 318.600 736.200 320.400 740.400 ;
        RECT 317.700 734.400 320.400 736.200 ;
        RECT 321.600 734.400 323.400 741.000 ;
        RECT 317.700 727.050 318.600 734.400 ;
        RECT 319.500 732.600 321.300 733.500 ;
        RECT 326.100 732.600 327.900 740.400 ;
        RECT 319.500 731.700 327.900 732.600 ;
        RECT 341.700 733.200 343.500 740.400 ;
        RECT 346.800 734.400 348.600 741.000 ;
        RECT 362.700 737.400 364.500 741.000 ;
        RECT 365.700 735.600 367.500 740.400 ;
        RECT 362.400 734.400 367.500 735.600 ;
        RECT 370.200 734.400 372.000 741.000 ;
        RECT 389.100 737.400 390.900 741.000 ;
        RECT 392.100 737.400 393.900 740.400 ;
        RECT 395.100 737.400 396.900 741.000 ;
        RECT 376.950 735.450 379.050 736.050 ;
        RECT 385.950 735.450 388.050 736.050 ;
        RECT 376.950 734.550 388.050 735.450 ;
        RECT 341.700 732.300 345.900 733.200 ;
        RECT 270.900 724.200 273.300 725.100 ;
        RECT 271.800 724.050 273.300 724.200 ;
        RECT 277.800 724.950 279.900 727.050 ;
        RECT 295.950 724.950 298.050 727.050 ;
        RECT 298.950 724.950 301.050 727.050 ;
        RECT 301.950 724.950 304.050 727.050 ;
        RECT 317.100 724.950 319.200 727.050 ;
        RECT 320.400 724.950 322.500 727.050 ;
        RECT 267.000 721.500 270.900 723.300 ;
        RECT 268.800 721.200 270.900 721.500 ;
        RECT 271.800 721.950 273.900 724.050 ;
        RECT 277.800 723.150 279.600 724.950 ;
        RECT 296.250 723.150 298.050 724.950 ;
        RECT 271.800 720.000 272.700 721.950 ;
        RECT 265.500 717.600 267.600 719.700 ;
        RECT 271.200 718.950 272.700 720.000 ;
        RECT 271.200 717.600 272.400 718.950 ;
        RECT 263.100 716.700 267.600 717.600 ;
        RECT 259.950 712.800 262.050 714.900 ;
        RECT 263.100 705.600 264.900 716.700 ;
        RECT 266.100 705.000 267.900 715.500 ;
        RECT 270.600 705.600 272.400 717.600 ;
        RECT 275.100 717.600 277.200 718.500 ;
        RECT 299.400 717.600 300.300 724.950 ;
        RECT 302.100 723.150 303.900 724.950 ;
        RECT 317.700 717.600 318.600 724.950 ;
        RECT 321.000 723.150 322.800 724.950 ;
        RECT 275.100 716.400 279.900 717.600 ;
        RECT 275.100 705.000 276.900 715.500 ;
        RECT 278.100 705.600 279.900 716.400 ;
        RECT 296.100 705.000 297.900 717.600 ;
        RECT 299.400 716.400 303.000 717.600 ;
        RECT 301.200 705.600 303.000 716.400 ;
        RECT 317.100 705.600 318.900 717.600 ;
        RECT 320.100 705.000 321.900 717.000 ;
        RECT 324.000 711.600 324.900 731.700 ;
        RECT 325.950 727.050 327.750 728.850 ;
        RECT 341.100 727.050 342.900 728.850 ;
        RECT 344.700 727.050 345.900 732.300 ;
        RECT 357.000 729.450 361.050 730.050 ;
        RECT 346.950 727.050 348.750 728.850 ;
        RECT 356.550 727.950 361.050 729.450 ;
        RECT 325.800 724.950 327.900 727.050 ;
        RECT 340.950 724.950 343.050 727.050 ;
        RECT 343.950 724.950 346.050 727.050 ;
        RECT 346.950 724.950 349.050 727.050 ;
        RECT 344.700 711.600 345.900 724.950 ;
        RECT 356.550 724.050 357.450 727.950 ;
        RECT 362.400 727.050 363.300 734.400 ;
        RECT 376.950 733.950 379.050 734.550 ;
        RECT 385.950 733.950 388.050 734.550 ;
        RECT 379.950 732.450 382.050 733.050 ;
        RECT 388.950 732.450 391.050 733.050 ;
        RECT 379.950 731.550 391.050 732.450 ;
        RECT 379.950 730.950 382.050 731.550 ;
        RECT 388.950 730.950 391.050 731.550 ;
        RECT 364.950 727.050 366.750 728.850 ;
        RECT 371.100 727.050 372.900 728.850 ;
        RECT 392.400 727.050 393.300 737.400 ;
        RECT 413.100 734.400 414.900 741.000 ;
        RECT 416.100 734.400 417.900 740.400 ;
        RECT 431.700 737.400 433.500 741.000 ;
        RECT 434.700 735.600 436.500 740.400 ;
        RECT 431.400 734.400 436.500 735.600 ;
        RECT 439.200 734.400 441.000 741.000 ;
        RECT 413.100 727.050 414.900 728.850 ;
        RECT 416.100 727.050 417.300 734.400 ;
        RECT 431.400 727.050 432.300 734.400 ;
        RECT 458.700 733.200 460.500 740.400 ;
        RECT 463.800 734.400 465.600 741.000 ;
        RECT 458.700 732.300 462.900 733.200 ;
        RECT 433.950 727.050 435.750 728.850 ;
        RECT 440.100 727.050 441.900 728.850 ;
        RECT 458.100 727.050 459.900 728.850 ;
        RECT 461.700 727.050 462.900 732.300 ;
        RECT 479.100 732.600 480.900 740.400 ;
        RECT 483.600 734.400 485.400 741.000 ;
        RECT 486.600 736.200 488.400 740.400 ;
        RECT 486.600 734.400 489.300 736.200 ;
        RECT 503.700 734.400 505.500 741.000 ;
        RECT 508.200 734.400 510.000 740.400 ;
        RECT 512.700 734.400 514.500 741.000 ;
        RECT 530.100 735.300 531.900 740.400 ;
        RECT 533.100 736.200 534.900 741.000 ;
        RECT 536.100 735.300 537.900 740.400 ;
        RECT 485.700 732.600 487.500 733.500 ;
        RECT 479.100 731.700 487.500 732.600 ;
        RECT 463.950 727.050 465.750 728.850 ;
        RECT 479.250 727.050 481.050 728.850 ;
        RECT 361.950 724.950 364.050 727.050 ;
        RECT 364.950 724.950 367.050 727.050 ;
        RECT 367.950 724.950 370.050 727.050 ;
        RECT 370.950 724.950 373.050 727.050 ;
        RECT 388.950 724.950 391.050 727.050 ;
        RECT 391.950 724.950 394.050 727.050 ;
        RECT 394.950 724.950 397.050 727.050 ;
        RECT 412.950 724.950 415.050 727.050 ;
        RECT 415.950 724.950 418.050 727.050 ;
        RECT 430.950 724.950 433.050 727.050 ;
        RECT 433.950 724.950 436.050 727.050 ;
        RECT 436.950 724.950 439.050 727.050 ;
        RECT 439.950 724.950 442.050 727.050 ;
        RECT 457.950 724.950 460.050 727.050 ;
        RECT 460.950 724.950 463.050 727.050 ;
        RECT 463.950 724.950 466.050 727.050 ;
        RECT 479.100 724.950 481.200 727.050 ;
        RECT 356.550 722.550 361.050 724.050 ;
        RECT 357.000 721.950 361.050 722.550 ;
        RECT 362.400 717.600 363.300 724.950 ;
        RECT 367.950 723.150 369.750 724.950 ;
        RECT 389.250 723.150 391.050 724.950 ;
        RECT 392.400 717.600 393.300 724.950 ;
        RECT 395.100 723.150 396.900 724.950 ;
        RECT 416.100 717.600 417.300 724.950 ;
        RECT 431.400 717.600 432.300 724.950 ;
        RECT 436.950 723.150 438.750 724.950 ;
        RECT 323.100 705.600 324.900 711.600 ;
        RECT 326.100 705.000 327.900 711.600 ;
        RECT 341.100 705.000 342.900 711.600 ;
        RECT 344.100 705.600 345.900 711.600 ;
        RECT 347.100 705.000 348.900 711.600 ;
        RECT 362.100 705.600 363.900 717.600 ;
        RECT 365.100 716.700 372.900 717.600 ;
        RECT 365.100 705.600 366.900 716.700 ;
        RECT 368.100 705.000 369.900 715.800 ;
        RECT 371.100 705.600 372.900 716.700 ;
        RECT 389.100 705.000 390.900 717.600 ;
        RECT 392.400 716.400 396.000 717.600 ;
        RECT 394.200 705.600 396.000 716.400 ;
        RECT 413.100 705.000 414.900 717.600 ;
        RECT 416.100 705.600 417.900 717.600 ;
        RECT 431.100 705.600 432.900 717.600 ;
        RECT 434.100 716.700 441.900 717.600 ;
        RECT 434.100 705.600 435.900 716.700 ;
        RECT 437.100 705.000 438.900 715.800 ;
        RECT 440.100 705.600 441.900 716.700 ;
        RECT 461.700 711.600 462.900 724.950 ;
        RECT 482.100 711.600 483.000 731.700 ;
        RECT 488.400 727.050 489.300 734.400 ;
        RECT 503.250 727.050 505.050 728.850 ;
        RECT 509.100 727.050 510.300 734.400 ;
        RECT 530.100 733.950 537.900 735.300 ;
        RECT 539.100 734.400 540.900 740.400 ;
        RECT 554.400 734.400 556.200 741.000 ;
        RECT 539.100 732.300 540.300 734.400 ;
        RECT 559.500 733.200 561.300 740.400 ;
        RECT 536.700 731.400 540.300 732.300 ;
        RECT 557.100 732.300 561.300 733.200 ;
        RECT 515.100 727.050 516.900 728.850 ;
        RECT 533.100 727.050 534.900 728.850 ;
        RECT 536.700 727.050 537.900 731.400 ;
        RECT 539.100 727.050 540.900 728.850 ;
        RECT 554.250 727.050 556.050 728.850 ;
        RECT 557.100 727.050 558.300 732.300 ;
        RECT 575.100 731.400 576.900 741.000 ;
        RECT 581.700 732.000 583.500 740.400 ;
        RECT 602.100 734.400 603.900 740.400 ;
        RECT 602.700 732.300 603.900 734.400 ;
        RECT 605.100 735.300 606.900 740.400 ;
        RECT 608.100 736.200 609.900 741.000 ;
        RECT 611.100 735.300 612.900 740.400 ;
        RECT 605.100 733.950 612.900 735.300 ;
        RECT 626.100 735.300 627.900 740.400 ;
        RECT 629.100 736.200 630.900 741.000 ;
        RECT 632.100 735.300 633.900 740.400 ;
        RECT 626.100 733.950 633.900 735.300 ;
        RECT 635.100 734.400 636.900 740.400 ;
        RECT 635.100 732.300 636.300 734.400 ;
        RECT 653.700 733.200 655.500 740.400 ;
        RECT 658.800 734.400 660.600 741.000 ;
        RECT 653.700 732.300 657.900 733.200 ;
        RECT 581.700 730.800 585.000 732.000 ;
        RECT 602.700 731.400 606.300 732.300 ;
        RECT 560.100 727.050 561.900 728.850 ;
        RECT 575.100 727.050 576.900 728.850 ;
        RECT 581.100 727.050 582.900 728.850 ;
        RECT 584.100 727.050 585.000 730.800 ;
        RECT 602.100 727.050 603.900 728.850 ;
        RECT 605.100 727.050 606.300 731.400 ;
        RECT 632.700 731.400 636.300 732.300 ;
        RECT 608.100 727.050 609.900 728.850 ;
        RECT 629.100 727.050 630.900 728.850 ;
        RECT 632.700 727.050 633.900 731.400 ;
        RECT 635.100 727.050 636.900 728.850 ;
        RECT 653.100 727.050 654.900 728.850 ;
        RECT 656.700 727.050 657.900 732.300 ;
        RECT 674.100 732.600 675.900 740.400 ;
        RECT 678.600 734.400 680.400 741.000 ;
        RECT 681.600 736.200 683.400 740.400 ;
        RECT 681.600 734.400 684.300 736.200 ;
        RECT 680.700 732.600 682.500 733.500 ;
        RECT 674.100 731.700 682.500 732.600 ;
        RECT 658.950 727.050 660.750 728.850 ;
        RECT 674.250 727.050 676.050 728.850 ;
        RECT 484.500 724.950 486.600 727.050 ;
        RECT 487.800 724.950 489.900 727.050 ;
        RECT 502.950 724.950 505.050 727.050 ;
        RECT 505.950 724.950 508.050 727.050 ;
        RECT 508.950 724.950 511.050 727.050 ;
        RECT 511.950 724.950 514.050 727.050 ;
        RECT 514.950 724.950 517.050 727.050 ;
        RECT 529.950 724.950 532.050 727.050 ;
        RECT 532.950 724.950 535.050 727.050 ;
        RECT 535.950 724.950 538.050 727.050 ;
        RECT 538.950 724.950 541.050 727.050 ;
        RECT 553.950 724.950 556.050 727.050 ;
        RECT 556.950 724.950 559.050 727.050 ;
        RECT 559.950 724.950 562.050 727.050 ;
        RECT 574.950 724.950 577.050 727.050 ;
        RECT 577.950 724.950 580.050 727.050 ;
        RECT 580.950 724.950 583.050 727.050 ;
        RECT 583.950 724.950 586.050 727.050 ;
        RECT 601.950 724.950 604.050 727.050 ;
        RECT 604.950 724.950 607.050 727.050 ;
        RECT 607.950 724.950 610.050 727.050 ;
        RECT 610.950 724.950 613.050 727.050 ;
        RECT 625.950 724.950 628.050 727.050 ;
        RECT 628.950 724.950 631.050 727.050 ;
        RECT 631.950 724.950 634.050 727.050 ;
        RECT 634.950 724.950 637.050 727.050 ;
        RECT 652.950 724.950 655.050 727.050 ;
        RECT 655.950 724.950 658.050 727.050 ;
        RECT 658.950 724.950 661.050 727.050 ;
        RECT 674.100 724.950 676.200 727.050 ;
        RECT 484.200 723.150 486.000 724.950 ;
        RECT 488.400 717.600 489.300 724.950 ;
        RECT 506.250 723.150 508.050 724.950 ;
        RECT 509.100 719.400 510.000 724.950 ;
        RECT 512.100 723.150 513.900 724.950 ;
        RECT 530.100 723.150 531.900 724.950 ;
        RECT 509.100 718.500 513.900 719.400 ;
        RECT 458.100 705.000 459.900 711.600 ;
        RECT 461.100 705.600 462.900 711.600 ;
        RECT 464.100 705.000 465.900 711.600 ;
        RECT 479.100 705.000 480.900 711.600 ;
        RECT 482.100 705.600 483.900 711.600 ;
        RECT 485.100 705.000 486.900 717.000 ;
        RECT 488.100 705.600 489.900 717.600 ;
        RECT 503.100 716.400 510.900 717.300 ;
        RECT 503.100 705.600 504.900 716.400 ;
        RECT 506.100 705.000 507.900 715.500 ;
        RECT 509.100 706.500 510.900 716.400 ;
        RECT 512.100 707.400 513.900 718.500 ;
        RECT 536.700 717.600 537.900 724.950 ;
        RECT 515.100 706.500 516.900 717.600 ;
        RECT 509.100 705.600 516.900 706.500 ;
        RECT 530.400 705.000 532.200 717.600 ;
        RECT 535.500 716.100 537.900 717.600 ;
        RECT 535.500 705.600 537.300 716.100 ;
        RECT 538.200 713.100 540.000 714.900 ;
        RECT 557.100 711.600 558.300 724.950 ;
        RECT 578.100 723.150 579.900 724.950 ;
        RECT 565.950 720.450 568.050 721.050 ;
        RECT 580.950 720.450 583.050 721.050 ;
        RECT 565.950 719.550 583.050 720.450 ;
        RECT 565.950 718.950 568.050 719.550 ;
        RECT 580.950 718.950 583.050 719.550 ;
        RECT 584.100 712.800 585.000 724.950 ;
        RECT 605.100 717.600 606.300 724.950 ;
        RECT 611.100 723.150 612.900 724.950 ;
        RECT 626.100 723.150 627.900 724.950 ;
        RECT 632.700 717.600 633.900 724.950 ;
        RECT 605.100 716.100 607.500 717.600 ;
        RECT 603.000 713.100 604.800 714.900 ;
        RECT 578.400 711.900 585.000 712.800 ;
        RECT 578.400 711.600 579.900 711.900 ;
        RECT 538.500 705.000 540.300 711.600 ;
        RECT 554.100 705.000 555.900 711.600 ;
        RECT 557.100 705.600 558.900 711.600 ;
        RECT 560.100 705.000 561.900 711.600 ;
        RECT 575.100 705.000 576.900 711.600 ;
        RECT 578.100 705.600 579.900 711.600 ;
        RECT 584.100 711.600 585.000 711.900 ;
        RECT 581.100 705.000 582.900 711.000 ;
        RECT 584.100 705.600 585.900 711.600 ;
        RECT 602.700 705.000 604.500 711.600 ;
        RECT 605.700 705.600 607.500 716.100 ;
        RECT 610.800 705.000 612.600 717.600 ;
        RECT 626.400 705.000 628.200 717.600 ;
        RECT 631.500 716.100 633.900 717.600 ;
        RECT 637.950 717.450 640.050 718.050 ;
        RECT 646.950 717.450 649.050 718.050 ;
        RECT 637.950 716.550 649.050 717.450 ;
        RECT 631.500 705.600 633.300 716.100 ;
        RECT 637.950 715.950 640.050 716.550 ;
        RECT 646.950 715.950 649.050 716.550 ;
        RECT 634.200 713.100 636.000 714.900 ;
        RECT 656.700 711.600 657.900 724.950 ;
        RECT 658.950 717.450 661.050 718.050 ;
        RECT 667.950 717.450 670.050 718.050 ;
        RECT 658.950 716.550 670.050 717.450 ;
        RECT 658.950 715.950 661.050 716.550 ;
        RECT 667.950 715.950 670.050 716.550 ;
        RECT 677.100 711.600 678.000 731.700 ;
        RECT 683.400 727.050 684.300 734.400 ;
        RECT 698.700 733.200 700.500 740.400 ;
        RECT 703.800 734.400 705.600 741.000 ;
        RECT 698.700 732.300 702.900 733.200 ;
        RECT 698.100 727.050 699.900 728.850 ;
        RECT 701.700 727.050 702.900 732.300 ;
        RECT 703.950 732.450 706.050 733.050 ;
        RECT 715.950 732.450 718.050 733.050 ;
        RECT 703.950 731.550 718.050 732.450 ;
        RECT 703.950 730.950 706.050 731.550 ;
        RECT 715.950 730.950 718.050 731.550 ;
        RECT 722.100 731.400 723.900 741.000 ;
        RECT 728.700 732.000 730.500 740.400 ;
        RECT 746.700 733.200 748.500 740.400 ;
        RECT 751.800 734.400 753.600 741.000 ;
        RECT 770.700 733.200 772.500 740.400 ;
        RECT 775.800 734.400 777.600 741.000 ;
        RECT 791.100 737.400 792.900 741.000 ;
        RECT 794.100 737.400 795.900 740.400 ;
        RECT 797.100 737.400 798.900 741.000 ;
        RECT 815.100 737.400 816.900 741.000 ;
        RECT 818.100 737.400 819.900 740.400 ;
        RECT 821.100 737.400 822.900 741.000 ;
        RECT 781.950 735.450 784.050 736.050 ;
        RECT 787.950 735.450 790.050 736.050 ;
        RECT 781.950 734.550 790.050 735.450 ;
        RECT 781.950 733.950 784.050 734.550 ;
        RECT 787.950 733.950 790.050 734.550 ;
        RECT 746.700 732.300 750.900 733.200 ;
        RECT 770.700 732.300 774.900 733.200 ;
        RECT 728.700 730.800 732.000 732.000 ;
        RECT 703.950 727.050 705.750 728.850 ;
        RECT 722.100 727.050 723.900 728.850 ;
        RECT 728.100 727.050 729.900 728.850 ;
        RECT 731.100 727.050 732.000 730.800 ;
        RECT 746.100 727.050 747.900 728.850 ;
        RECT 749.700 727.050 750.900 732.300 ;
        RECT 751.950 727.050 753.750 728.850 ;
        RECT 770.100 727.050 771.900 728.850 ;
        RECT 773.700 727.050 774.900 732.300 ;
        RECT 775.950 727.050 777.750 728.850 ;
        RECT 794.700 727.050 795.600 737.400 ;
        RECT 818.700 727.050 819.600 737.400 ;
        RECT 836.100 735.300 837.900 740.400 ;
        RECT 839.100 736.200 840.900 741.000 ;
        RECT 842.100 735.300 843.900 740.400 ;
        RECT 836.100 733.950 843.900 735.300 ;
        RECT 845.100 734.400 846.900 740.400 ;
        RECT 863.100 735.300 864.900 740.400 ;
        RECT 866.100 736.200 867.900 741.000 ;
        RECT 869.100 735.300 870.900 740.400 ;
        RECT 845.100 732.300 846.300 734.400 ;
        RECT 863.100 733.950 870.900 735.300 ;
        RECT 872.100 734.400 873.900 740.400 ;
        RECT 888.000 734.400 889.800 741.000 ;
        RECT 892.500 735.600 894.300 740.400 ;
        RECT 895.500 737.400 897.300 741.000 ;
        RECT 892.500 734.400 897.600 735.600 ;
        RECT 872.100 732.300 873.300 734.400 ;
        RECT 842.700 731.400 846.300 732.300 ;
        RECT 869.700 731.400 873.300 732.300 ;
        RECT 831.000 729.450 835.050 730.050 ;
        RECT 830.550 727.950 835.050 729.450 ;
        RECT 679.500 724.950 681.600 727.050 ;
        RECT 682.800 724.950 684.900 727.050 ;
        RECT 697.950 724.950 700.050 727.050 ;
        RECT 700.950 724.950 703.050 727.050 ;
        RECT 703.950 724.950 706.050 727.050 ;
        RECT 721.950 724.950 724.050 727.050 ;
        RECT 724.950 724.950 727.050 727.050 ;
        RECT 727.950 724.950 730.050 727.050 ;
        RECT 730.950 724.950 733.050 727.050 ;
        RECT 745.950 724.950 748.050 727.050 ;
        RECT 748.950 724.950 751.050 727.050 ;
        RECT 751.950 724.950 754.050 727.050 ;
        RECT 769.950 724.950 772.050 727.050 ;
        RECT 772.950 724.950 775.050 727.050 ;
        RECT 775.950 724.950 778.050 727.050 ;
        RECT 790.950 724.950 793.050 727.050 ;
        RECT 793.950 724.950 796.050 727.050 ;
        RECT 796.950 724.950 799.050 727.050 ;
        RECT 814.950 724.950 817.050 727.050 ;
        RECT 817.950 724.950 820.050 727.050 ;
        RECT 820.950 724.950 823.050 727.050 ;
        RECT 679.200 723.150 681.000 724.950 ;
        RECT 683.400 717.600 684.300 724.950 ;
        RECT 634.500 705.000 636.300 711.600 ;
        RECT 653.100 705.000 654.900 711.600 ;
        RECT 656.100 705.600 657.900 711.600 ;
        RECT 659.100 705.000 660.900 711.600 ;
        RECT 674.100 705.000 675.900 711.600 ;
        RECT 677.100 705.600 678.900 711.600 ;
        RECT 680.100 705.000 681.900 717.000 ;
        RECT 683.100 705.600 684.900 717.600 ;
        RECT 701.700 711.600 702.900 724.950 ;
        RECT 725.100 723.150 726.900 724.950 ;
        RECT 709.950 720.450 712.050 721.050 ;
        RECT 727.950 720.450 730.050 721.050 ;
        RECT 709.950 719.550 730.050 720.450 ;
        RECT 709.950 718.950 712.050 719.550 ;
        RECT 727.950 718.950 730.050 719.550 ;
        RECT 731.100 712.800 732.000 724.950 ;
        RECT 725.400 711.900 732.000 712.800 ;
        RECT 725.400 711.600 726.900 711.900 ;
        RECT 698.100 705.000 699.900 711.600 ;
        RECT 701.100 705.600 702.900 711.600 ;
        RECT 704.100 705.000 705.900 711.600 ;
        RECT 722.100 705.000 723.900 711.600 ;
        RECT 725.100 705.600 726.900 711.600 ;
        RECT 731.100 711.600 732.000 711.900 ;
        RECT 749.700 711.600 750.900 724.950 ;
        RECT 773.700 711.600 774.900 724.950 ;
        RECT 791.100 723.150 792.900 724.950 ;
        RECT 794.700 717.600 795.600 724.950 ;
        RECT 796.950 723.150 798.750 724.950 ;
        RECT 815.100 723.150 816.900 724.950 ;
        RECT 818.700 717.600 819.600 724.950 ;
        RECT 820.950 723.150 822.750 724.950 ;
        RECT 823.950 723.450 826.050 724.050 ;
        RECT 830.550 723.450 831.450 727.950 ;
        RECT 839.100 727.050 840.900 728.850 ;
        RECT 842.700 727.050 843.900 731.400 ;
        RECT 845.100 727.050 846.900 728.850 ;
        RECT 866.100 727.050 867.900 728.850 ;
        RECT 869.700 727.050 870.900 731.400 ;
        RECT 874.950 729.450 879.000 730.050 ;
        RECT 872.100 727.050 873.900 728.850 ;
        RECT 874.950 727.950 879.450 729.450 ;
        RECT 835.950 724.950 838.050 727.050 ;
        RECT 838.950 724.950 841.050 727.050 ;
        RECT 841.950 724.950 844.050 727.050 ;
        RECT 844.950 724.950 847.050 727.050 ;
        RECT 862.950 724.950 865.050 727.050 ;
        RECT 865.950 724.950 868.050 727.050 ;
        RECT 868.950 724.950 871.050 727.050 ;
        RECT 871.950 724.950 874.050 727.050 ;
        RECT 823.950 722.550 831.450 723.450 ;
        RECT 836.100 723.150 837.900 724.950 ;
        RECT 823.950 721.950 826.050 722.550 ;
        RECT 842.700 717.600 843.900 724.950 ;
        RECT 847.950 723.450 850.050 724.050 ;
        RECT 856.950 723.450 859.050 724.050 ;
        RECT 847.950 722.550 859.050 723.450 ;
        RECT 863.100 723.150 864.900 724.950 ;
        RECT 847.950 721.950 850.050 722.550 ;
        RECT 856.950 721.950 859.050 722.550 ;
        RECT 869.700 717.600 870.900 724.950 ;
        RECT 878.550 723.450 879.450 727.950 ;
        RECT 887.100 727.050 888.900 728.850 ;
        RECT 893.250 727.050 895.050 728.850 ;
        RECT 896.700 727.050 897.600 734.400 ;
        RECT 914.100 735.300 915.900 740.400 ;
        RECT 917.100 736.200 918.900 741.000 ;
        RECT 920.100 735.300 921.900 740.400 ;
        RECT 914.100 733.950 921.900 735.300 ;
        RECT 923.100 734.400 924.900 740.400 ;
        RECT 938.100 735.300 939.900 740.400 ;
        RECT 941.100 736.200 942.900 741.000 ;
        RECT 944.100 735.300 945.900 740.400 ;
        RECT 923.100 732.300 924.300 734.400 ;
        RECT 938.100 733.950 945.900 735.300 ;
        RECT 947.100 734.400 948.900 740.400 ;
        RECT 962.100 735.000 963.900 740.400 ;
        RECT 965.100 735.900 966.900 741.000 ;
        RECT 968.100 739.500 975.900 740.400 ;
        RECT 968.100 735.000 969.900 739.500 ;
        RECT 920.700 731.400 924.300 732.300 ;
        RECT 925.950 732.450 928.050 733.050 ;
        RECT 931.950 732.450 934.050 732.900 ;
        RECT 925.950 731.550 934.050 732.450 ;
        RECT 947.100 732.300 948.300 734.400 ;
        RECT 962.100 734.100 969.900 735.000 ;
        RECT 971.100 734.400 972.900 738.600 ;
        RECT 974.100 734.400 975.900 739.500 ;
        RECT 917.100 727.050 918.900 728.850 ;
        RECT 920.700 727.050 921.900 731.400 ;
        RECT 925.950 730.950 928.050 731.550 ;
        RECT 931.950 730.800 934.050 731.550 ;
        RECT 944.700 731.400 948.300 732.300 ;
        RECT 949.950 732.450 952.050 733.050 ;
        RECT 961.950 732.450 964.050 733.050 ;
        RECT 971.400 732.900 972.300 734.400 ;
        RECT 949.950 731.550 964.050 732.450 ;
        RECT 923.100 727.050 924.900 728.850 ;
        RECT 941.100 727.050 942.900 728.850 ;
        RECT 944.700 727.050 945.900 731.400 ;
        RECT 949.950 730.950 952.050 731.550 ;
        RECT 961.950 730.950 964.050 731.550 ;
        RECT 967.950 731.700 972.300 732.900 ;
        RECT 989.700 733.200 991.500 740.400 ;
        RECT 994.800 734.400 996.600 741.000 ;
        RECT 989.700 732.300 993.900 733.200 ;
        RECT 947.100 727.050 948.900 728.850 ;
        RECT 965.250 727.050 967.050 728.850 ;
        RECT 886.950 724.950 889.050 727.050 ;
        RECT 889.950 724.950 892.050 727.050 ;
        RECT 892.950 724.950 895.050 727.050 ;
        RECT 895.950 724.950 898.050 727.050 ;
        RECT 913.950 724.950 916.050 727.050 ;
        RECT 916.950 724.950 919.050 727.050 ;
        RECT 919.950 724.950 922.050 727.050 ;
        RECT 922.950 724.950 925.050 727.050 ;
        RECT 937.950 724.950 940.050 727.050 ;
        RECT 940.950 724.950 943.050 727.050 ;
        RECT 943.950 724.950 946.050 727.050 ;
        RECT 946.950 724.950 949.050 727.050 ;
        RECT 961.950 724.950 964.050 727.050 ;
        RECT 964.950 724.950 967.050 727.050 ;
        RECT 967.950 727.050 969.000 731.700 ;
        RECT 976.950 729.450 981.000 730.050 ;
        RECT 984.000 729.450 988.050 730.050 ;
        RECT 970.950 727.050 972.750 728.850 ;
        RECT 976.950 727.950 981.450 729.450 ;
        RECT 967.950 724.950 970.050 727.050 ;
        RECT 970.950 724.950 973.050 727.050 ;
        RECT 973.950 724.950 976.050 727.050 ;
        RECT 883.950 723.450 886.050 724.050 ;
        RECT 878.550 722.550 886.050 723.450 ;
        RECT 890.250 723.150 892.050 724.950 ;
        RECT 883.950 721.950 886.050 722.550 ;
        RECT 896.700 717.600 897.600 724.950 ;
        RECT 914.100 723.150 915.900 724.950 ;
        RECT 920.700 717.600 921.900 724.950 ;
        RECT 938.100 723.150 939.900 724.950 ;
        RECT 944.700 717.600 945.900 724.950 ;
        RECT 962.100 723.150 963.900 724.950 ;
        RECT 967.950 717.600 969.000 724.950 ;
        RECT 973.950 723.150 975.750 724.950 ;
        RECT 980.550 724.050 981.450 727.950 ;
        RECT 976.950 722.550 981.450 724.050 ;
        RECT 983.550 727.950 988.050 729.450 ;
        RECT 983.550 724.050 984.450 727.950 ;
        RECT 989.100 727.050 990.900 728.850 ;
        RECT 992.700 727.050 993.900 732.300 ;
        RECT 997.950 729.450 1002.000 730.050 ;
        RECT 994.950 727.050 996.750 728.850 ;
        RECT 997.950 727.950 1002.450 729.450 ;
        RECT 988.950 724.950 991.050 727.050 ;
        RECT 991.950 724.950 994.050 727.050 ;
        RECT 994.950 724.950 997.050 727.050 ;
        RECT 983.550 722.550 988.050 724.050 ;
        RECT 976.950 721.950 981.000 722.550 ;
        RECT 984.000 721.950 988.050 722.550 ;
        RECT 792.000 716.400 795.600 717.600 ;
        RECT 728.100 705.000 729.900 711.000 ;
        RECT 731.100 705.600 732.900 711.600 ;
        RECT 746.100 705.000 747.900 711.600 ;
        RECT 749.100 705.600 750.900 711.600 ;
        RECT 752.100 705.000 753.900 711.600 ;
        RECT 770.100 705.000 771.900 711.600 ;
        RECT 773.100 705.600 774.900 711.600 ;
        RECT 776.100 705.000 777.900 711.600 ;
        RECT 792.000 705.600 793.800 716.400 ;
        RECT 797.100 705.000 798.900 717.600 ;
        RECT 816.000 716.400 819.600 717.600 ;
        RECT 816.000 705.600 817.800 716.400 ;
        RECT 821.100 705.000 822.900 717.600 ;
        RECT 836.400 705.000 838.200 717.600 ;
        RECT 841.500 716.100 843.900 717.600 ;
        RECT 841.500 705.600 843.300 716.100 ;
        RECT 844.200 713.100 846.000 714.900 ;
        RECT 844.500 705.000 846.300 711.600 ;
        RECT 863.400 705.000 865.200 717.600 ;
        RECT 868.500 716.100 870.900 717.600 ;
        RECT 887.100 716.700 894.900 717.600 ;
        RECT 868.500 705.600 870.300 716.100 ;
        RECT 871.200 713.100 873.000 714.900 ;
        RECT 871.500 705.000 873.300 711.600 ;
        RECT 887.100 705.600 888.900 716.700 ;
        RECT 890.100 705.000 891.900 715.800 ;
        RECT 893.100 705.600 894.900 716.700 ;
        RECT 896.100 705.600 897.900 717.600 ;
        RECT 914.400 705.000 916.200 717.600 ;
        RECT 919.500 716.100 921.900 717.600 ;
        RECT 919.500 705.600 921.300 716.100 ;
        RECT 922.200 713.100 924.000 714.900 ;
        RECT 922.500 705.000 924.300 711.600 ;
        RECT 938.400 705.000 940.200 717.600 ;
        RECT 943.500 716.100 945.900 717.600 ;
        RECT 943.500 705.600 945.300 716.100 ;
        RECT 946.200 713.100 948.000 714.900 ;
        RECT 946.500 705.000 948.300 711.600 ;
        RECT 962.100 705.000 963.900 717.600 ;
        RECT 966.600 705.600 969.900 717.600 ;
        RECT 972.600 705.000 974.400 717.600 ;
        RECT 992.700 711.600 993.900 724.950 ;
        RECT 1001.550 723.450 1002.450 727.950 ;
        RECT 998.550 722.550 1002.450 723.450 ;
        RECT 998.550 721.050 999.450 722.550 ;
        RECT 996.000 720.750 999.450 721.050 ;
        RECT 994.950 719.550 999.450 720.750 ;
        RECT 994.950 718.950 999.000 719.550 ;
        RECT 994.950 718.650 997.050 718.950 ;
        RECT 989.100 705.000 990.900 711.600 ;
        RECT 992.100 705.600 993.900 711.600 ;
        RECT 995.100 705.000 996.900 711.600 ;
        RECT 2.550 689.400 4.350 701.400 ;
        RECT 5.550 689.400 7.350 702.000 ;
        RECT 10.350 695.400 12.150 701.400 ;
        RECT 14.850 695.400 16.650 702.000 ;
        RECT 10.350 693.300 12.450 695.400 ;
        RECT 17.850 694.500 19.650 701.400 ;
        RECT 20.850 695.400 22.650 702.000 ;
        RECT 16.950 693.450 23.550 694.500 ;
        RECT 16.950 692.700 18.750 693.450 ;
        RECT 21.750 692.700 23.550 693.450 ;
        RECT 25.650 692.400 27.450 701.400 ;
        RECT 9.450 690.600 12.450 692.400 ;
        RECT 13.350 691.800 15.150 692.400 ;
        RECT 13.350 690.900 19.050 691.800 ;
        RECT 25.650 691.500 27.750 692.400 ;
        RECT 13.350 690.600 15.150 690.900 ;
        RECT 11.250 689.700 12.450 690.600 ;
        RECT 2.550 682.050 3.750 689.400 ;
        RECT 11.250 688.800 16.050 689.700 ;
        RECT 4.650 686.100 6.450 686.550 ;
        RECT 10.350 686.100 12.450 686.700 ;
        RECT 4.650 684.900 12.450 686.100 ;
        RECT 4.650 684.750 6.450 684.900 ;
        RECT 10.350 684.600 12.450 684.900 ;
        RECT 2.550 681.750 7.050 682.050 ;
        RECT 2.550 679.950 8.850 681.750 ;
        RECT 2.550 672.600 3.750 679.950 ;
        RECT 15.150 676.200 16.050 688.800 ;
        RECT 18.150 688.800 19.050 690.900 ;
        RECT 19.950 690.300 27.750 691.500 ;
        RECT 19.950 689.700 21.750 690.300 ;
        RECT 31.050 689.400 32.850 702.000 ;
        RECT 34.050 691.200 35.850 701.400 ;
        RECT 34.050 689.400 36.450 691.200 ;
        RECT 50.400 689.400 52.200 702.000 ;
        RECT 55.500 690.900 57.300 701.400 ;
        RECT 58.500 695.400 60.300 702.000 ;
        RECT 77.100 695.400 78.900 702.000 ;
        RECT 80.100 695.400 81.900 701.400 ;
        RECT 83.100 695.400 84.900 702.000 ;
        RECT 58.200 692.100 60.000 693.900 ;
        RECT 55.500 689.400 57.900 690.900 ;
        RECT 18.150 688.500 26.550 688.800 ;
        RECT 35.550 688.500 36.450 689.400 ;
        RECT 18.150 687.900 36.450 688.500 ;
        RECT 24.750 687.300 36.450 687.900 ;
        RECT 24.750 687.000 26.550 687.300 ;
        RECT 22.800 680.400 24.900 682.050 ;
        RECT 22.800 679.200 30.900 680.400 ;
        RECT 31.950 679.950 34.050 682.050 ;
        RECT 29.100 678.600 30.900 679.200 ;
        RECT 26.100 677.400 27.900 678.000 ;
        RECT 32.250 677.400 34.050 679.950 ;
        RECT 26.100 676.200 34.050 677.400 ;
        RECT 15.150 675.000 27.150 676.200 ;
        RECT 15.150 674.400 16.950 675.000 ;
        RECT 26.100 673.200 27.150 675.000 ;
        RECT 2.550 666.600 4.350 672.600 ;
        RECT 5.850 666.000 7.650 672.600 ;
        RECT 10.350 669.600 12.750 671.700 ;
        RECT 22.350 671.550 24.150 672.300 ;
        RECT 19.200 670.500 24.150 671.550 ;
        RECT 25.350 671.400 27.150 673.200 ;
        RECT 35.550 672.600 36.450 687.300 ;
        RECT 50.100 682.050 51.900 683.850 ;
        RECT 56.700 682.050 57.900 689.400 ;
        RECT 80.100 682.050 81.300 695.400 ;
        RECT 101.100 690.300 102.900 701.400 ;
        RECT 104.100 691.500 105.900 702.000 ;
        RECT 108.600 690.300 110.400 701.400 ;
        RECT 112.800 691.500 114.900 702.000 ;
        RECT 116.100 690.600 117.900 701.400 ;
        RECT 101.100 689.100 105.900 690.300 ;
        RECT 108.600 689.400 111.900 690.300 ;
        RECT 103.800 688.200 105.900 689.100 ;
        RECT 103.800 687.300 109.200 688.200 ;
        RECT 107.400 685.500 109.200 687.300 ;
        RECT 110.700 685.050 111.900 689.400 ;
        RECT 112.800 689.400 117.900 690.600 ;
        RECT 131.100 690.600 132.900 701.400 ;
        RECT 134.100 691.500 135.900 702.000 ;
        RECT 131.100 689.400 135.900 690.600 ;
        RECT 112.800 688.500 114.900 689.400 ;
        RECT 133.800 688.500 135.900 689.400 ;
        RECT 138.600 689.400 140.400 701.400 ;
        RECT 143.100 691.500 144.900 702.000 ;
        RECT 146.100 690.300 147.900 701.400 ;
        RECT 161.100 695.400 162.900 702.000 ;
        RECT 164.100 695.400 165.900 701.400 ;
        RECT 179.100 695.400 180.900 702.000 ;
        RECT 182.100 695.400 183.900 701.400 ;
        RECT 185.100 695.400 186.900 702.000 ;
        RECT 203.100 695.400 204.900 702.000 ;
        RECT 206.100 695.400 207.900 701.400 ;
        RECT 209.100 696.000 210.900 702.000 ;
        RECT 143.400 689.400 147.900 690.300 ;
        RECT 138.600 688.050 139.800 689.400 ;
        RECT 138.300 687.000 139.800 688.050 ;
        RECT 143.400 687.300 145.500 689.400 ;
        RECT 138.300 685.050 139.200 687.000 ;
        RECT 110.100 684.300 112.200 685.050 ;
        RECT 105.900 682.200 107.700 684.000 ;
        RECT 109.200 682.950 112.200 684.300 ;
        RECT 49.950 679.950 52.050 682.050 ;
        RECT 52.950 679.950 55.050 682.050 ;
        RECT 55.950 679.950 58.050 682.050 ;
        RECT 58.950 679.950 61.050 682.050 ;
        RECT 76.950 679.950 79.050 682.050 ;
        RECT 79.950 679.950 82.050 682.050 ;
        RECT 82.950 679.950 85.050 682.050 ;
        RECT 53.100 678.150 54.900 679.950 ;
        RECT 56.700 675.600 57.900 679.950 ;
        RECT 59.100 678.150 60.900 679.950 ;
        RECT 77.250 678.150 79.050 679.950 ;
        RECT 56.700 674.700 60.300 675.600 ;
        RECT 19.200 669.600 20.250 670.500 ;
        RECT 28.050 670.200 30.150 671.700 ;
        RECT 26.250 669.600 30.150 670.200 ;
        RECT 10.950 666.600 12.750 669.600 ;
        RECT 15.450 666.000 17.250 669.600 ;
        RECT 18.450 666.600 20.250 669.600 ;
        RECT 21.750 666.000 23.550 669.600 ;
        RECT 26.250 668.700 29.850 669.600 ;
        RECT 26.250 666.600 28.050 668.700 ;
        RECT 31.050 666.000 32.850 672.600 ;
        RECT 34.050 670.800 36.450 672.600 ;
        RECT 50.100 671.700 57.900 673.050 ;
        RECT 34.050 666.600 35.850 670.800 ;
        RECT 50.100 666.600 51.900 671.700 ;
        RECT 53.100 666.000 54.900 670.800 ;
        RECT 56.100 666.600 57.900 671.700 ;
        RECT 59.100 672.600 60.300 674.700 ;
        RECT 80.100 674.700 81.300 679.950 ;
        RECT 83.100 678.150 84.900 679.950 ;
        RECT 101.100 679.800 103.200 682.050 ;
        RECT 105.900 680.100 108.000 682.200 ;
        RECT 101.400 679.200 103.200 679.800 ;
        RECT 101.400 678.000 108.000 679.200 ;
        RECT 105.900 677.100 108.000 678.000 ;
        RECT 103.500 675.000 105.600 675.600 ;
        RECT 106.500 675.300 108.300 677.100 ;
        RECT 109.200 676.200 110.100 682.950 ;
        RECT 115.800 682.050 117.600 683.850 ;
        RECT 131.400 682.050 133.200 683.850 ;
        RECT 137.100 682.950 139.200 685.050 ;
        RECT 140.100 685.500 142.200 685.800 ;
        RECT 140.100 683.700 144.000 685.500 ;
        RECT 111.000 680.100 112.800 681.900 ;
        RECT 111.000 678.000 113.100 680.100 ;
        RECT 115.800 679.950 117.900 682.050 ;
        RECT 131.100 679.950 133.200 682.050 ;
        RECT 137.700 682.800 139.200 682.950 ;
        RECT 137.700 681.900 140.100 682.800 ;
        RECT 135.900 679.200 137.700 681.000 ;
        RECT 135.900 677.100 138.000 679.200 ;
        RECT 138.900 676.200 140.100 681.900 ;
        RECT 141.000 682.050 142.800 682.500 ;
        RECT 161.100 682.050 162.900 683.850 ;
        RECT 164.100 682.050 165.300 695.400 ;
        RECT 182.100 682.050 183.300 695.400 ;
        RECT 206.400 695.100 207.900 695.400 ;
        RECT 212.100 695.400 213.900 701.400 ;
        RECT 212.100 695.100 213.000 695.400 ;
        RECT 206.400 694.200 213.000 695.100 ;
        RECT 206.100 682.050 207.900 683.850 ;
        RECT 212.100 682.050 213.000 694.200 ;
        RECT 227.400 689.400 229.200 702.000 ;
        RECT 232.500 690.900 234.300 701.400 ;
        RECT 235.500 695.400 237.300 702.000 ;
        RECT 251.100 695.400 252.900 702.000 ;
        RECT 254.100 695.400 255.900 701.400 ;
        RECT 257.100 695.400 258.900 702.000 ;
        RECT 272.100 695.400 273.900 702.000 ;
        RECT 275.100 695.400 276.900 701.400 ;
        RECT 235.200 692.100 237.000 693.900 ;
        RECT 232.500 689.400 234.900 690.900 ;
        RECT 227.100 682.050 228.900 683.850 ;
        RECT 233.700 682.050 234.900 689.400 ;
        RECT 254.700 682.050 255.900 695.400 ;
        RECT 141.000 680.700 147.900 682.050 ;
        RECT 145.800 679.950 147.900 680.700 ;
        RECT 160.950 679.950 163.050 682.050 ;
        RECT 163.950 679.950 166.050 682.050 ;
        RECT 178.950 679.950 181.050 682.050 ;
        RECT 181.950 679.950 184.050 682.050 ;
        RECT 184.950 679.950 187.050 682.050 ;
        RECT 202.950 679.950 205.050 682.050 ;
        RECT 205.950 679.950 208.050 682.050 ;
        RECT 208.950 679.950 211.050 682.050 ;
        RECT 211.950 679.950 214.050 682.050 ;
        RECT 226.950 679.950 229.050 682.050 ;
        RECT 229.950 679.950 232.050 682.050 ;
        RECT 232.950 679.950 235.050 682.050 ;
        RECT 235.950 679.950 238.050 682.050 ;
        RECT 250.950 679.950 253.050 682.050 ;
        RECT 253.950 679.950 256.050 682.050 ;
        RECT 256.950 679.950 259.050 682.050 ;
        RECT 272.100 679.950 274.200 682.050 ;
        RECT 80.100 673.800 84.300 674.700 ;
        RECT 59.100 666.600 60.900 672.600 ;
        RECT 77.400 666.000 79.200 672.600 ;
        RECT 82.500 666.600 84.300 673.800 ;
        RECT 101.100 673.500 105.600 675.000 ;
        RECT 109.200 674.100 112.200 676.200 ;
        RECT 101.100 672.600 102.600 673.500 ;
        RECT 101.100 666.600 102.900 672.600 ;
        RECT 109.200 672.000 110.100 674.100 ;
        RECT 113.400 673.500 115.500 675.900 ;
        RECT 133.800 673.500 135.900 674.700 ;
        RECT 137.100 674.100 140.100 676.200 ;
        RECT 141.000 677.400 142.800 679.200 ;
        RECT 145.800 678.150 147.600 679.950 ;
        RECT 141.000 675.300 143.100 677.400 ;
        RECT 141.000 674.400 147.300 675.300 ;
        RECT 113.400 672.600 117.900 673.500 ;
        RECT 104.100 666.000 105.900 671.700 ;
        RECT 108.300 666.600 110.100 672.000 ;
        RECT 112.800 666.000 114.600 671.700 ;
        RECT 116.100 666.600 117.900 672.600 ;
        RECT 131.100 672.600 135.900 673.500 ;
        RECT 138.900 672.600 140.100 674.100 ;
        RECT 146.100 672.600 147.300 674.400 ;
        RECT 131.100 666.600 132.900 672.600 ;
        RECT 134.100 666.000 135.900 671.700 ;
        RECT 138.600 666.600 140.400 672.600 ;
        RECT 143.100 666.000 144.900 671.700 ;
        RECT 146.100 666.600 147.900 672.600 ;
        RECT 164.100 669.600 165.300 679.950 ;
        RECT 179.250 678.150 181.050 679.950 ;
        RECT 182.100 674.700 183.300 679.950 ;
        RECT 185.100 678.150 186.900 679.950 ;
        RECT 203.100 678.150 204.900 679.950 ;
        RECT 209.100 678.150 210.900 679.950 ;
        RECT 212.100 676.200 213.000 679.950 ;
        RECT 230.100 678.150 231.900 679.950 ;
        RECT 182.100 673.800 186.300 674.700 ;
        RECT 161.100 666.000 162.900 669.600 ;
        RECT 164.100 666.600 165.900 669.600 ;
        RECT 179.400 666.000 181.200 672.600 ;
        RECT 184.500 666.600 186.300 673.800 ;
        RECT 203.100 666.000 204.900 675.600 ;
        RECT 209.700 675.000 213.000 676.200 ;
        RECT 233.700 675.600 234.900 679.950 ;
        RECT 236.100 678.150 237.900 679.950 ;
        RECT 251.100 678.150 252.900 679.950 ;
        RECT 209.700 666.600 211.500 675.000 ;
        RECT 233.700 674.700 237.300 675.600 ;
        RECT 254.700 674.700 255.900 679.950 ;
        RECT 256.950 678.150 258.750 679.950 ;
        RECT 272.250 678.150 274.050 679.950 ;
        RECT 275.100 675.300 276.000 695.400 ;
        RECT 278.100 690.000 279.900 702.000 ;
        RECT 281.100 689.400 282.900 701.400 ;
        RECT 296.700 695.400 298.500 702.000 ;
        RECT 297.000 692.100 298.800 693.900 ;
        RECT 299.700 690.900 301.500 701.400 ;
        RECT 299.100 689.400 301.500 690.900 ;
        RECT 304.800 689.400 306.600 702.000 ;
        RECT 320.100 695.400 321.900 701.400 ;
        RECT 323.100 695.400 324.900 702.000 ;
        RECT 341.700 695.400 343.500 702.000 ;
        RECT 277.200 682.050 279.000 683.850 ;
        RECT 281.400 682.050 282.300 689.400 ;
        RECT 299.100 682.050 300.300 689.400 ;
        RECT 305.100 682.050 306.900 683.850 ;
        RECT 320.700 682.050 321.900 695.400 ;
        RECT 342.000 692.100 343.800 693.900 ;
        RECT 344.700 690.900 346.500 701.400 ;
        RECT 344.100 689.400 346.500 690.900 ;
        RECT 349.800 689.400 351.600 702.000 ;
        RECT 365.100 700.500 372.900 701.400 ;
        RECT 365.100 689.400 366.900 700.500 ;
        RECT 323.100 682.050 324.900 683.850 ;
        RECT 344.100 682.050 345.300 689.400 ;
        RECT 368.100 688.500 369.900 699.600 ;
        RECT 371.100 690.600 372.900 700.500 ;
        RECT 374.100 691.500 375.900 702.000 ;
        RECT 377.100 690.600 378.900 701.400 ;
        RECT 392.100 695.400 393.900 701.400 ;
        RECT 395.100 695.400 396.900 702.000 ;
        RECT 371.100 689.700 378.900 690.600 ;
        RECT 368.100 687.600 372.900 688.500 ;
        RECT 352.950 684.450 357.000 685.050 ;
        RECT 350.100 682.050 351.900 683.850 ;
        RECT 352.950 682.950 357.450 684.450 ;
        RECT 277.500 679.950 279.600 682.050 ;
        RECT 280.800 679.950 282.900 682.050 ;
        RECT 295.950 679.950 298.050 682.050 ;
        RECT 298.950 679.950 301.050 682.050 ;
        RECT 301.950 679.950 304.050 682.050 ;
        RECT 304.950 679.950 307.050 682.050 ;
        RECT 319.950 679.950 322.050 682.050 ;
        RECT 322.950 679.950 325.050 682.050 ;
        RECT 340.950 679.950 343.050 682.050 ;
        RECT 343.950 679.950 346.050 682.050 ;
        RECT 346.950 679.950 349.050 682.050 ;
        RECT 349.950 679.950 352.050 682.050 ;
        RECT 356.550 681.450 357.450 682.950 ;
        RECT 368.100 682.050 369.900 683.850 ;
        RECT 372.000 682.050 372.900 687.600 ;
        RECT 373.950 682.050 375.750 683.850 ;
        RECT 392.700 682.050 393.900 695.400 ;
        RECT 410.400 689.400 412.200 702.000 ;
        RECT 415.500 690.900 417.300 701.400 ;
        RECT 418.500 695.400 420.300 702.000 ;
        RECT 418.200 692.100 420.000 693.900 ;
        RECT 415.500 689.400 417.900 690.900 ;
        RECT 437.100 689.400 438.900 701.400 ;
        RECT 440.100 690.000 441.900 702.000 ;
        RECT 443.100 695.400 444.900 701.400 ;
        RECT 446.100 695.400 447.900 702.000 ;
        RECT 395.100 682.050 396.900 683.850 ;
        RECT 410.100 682.050 411.900 683.850 ;
        RECT 416.700 682.050 417.900 689.400 ;
        RECT 437.700 682.050 438.600 689.400 ;
        RECT 441.000 682.050 442.800 683.850 ;
        RECT 356.550 680.550 360.450 681.450 ;
        RECT 227.100 671.700 234.900 673.050 ;
        RECT 227.100 666.600 228.900 671.700 ;
        RECT 230.100 666.000 231.900 670.800 ;
        RECT 233.100 666.600 234.900 671.700 ;
        RECT 236.100 672.600 237.300 674.700 ;
        RECT 251.700 673.800 255.900 674.700 ;
        RECT 272.100 674.400 280.500 675.300 ;
        RECT 236.100 666.600 237.900 672.600 ;
        RECT 251.700 666.600 253.500 673.800 ;
        RECT 256.800 666.000 258.600 672.600 ;
        RECT 272.100 666.600 273.900 674.400 ;
        RECT 278.700 673.500 280.500 674.400 ;
        RECT 281.400 672.600 282.300 679.950 ;
        RECT 296.100 678.150 297.900 679.950 ;
        RECT 299.100 675.600 300.300 679.950 ;
        RECT 302.100 678.150 303.900 679.950 ;
        RECT 296.700 674.700 300.300 675.600 ;
        RECT 296.700 672.600 297.900 674.700 ;
        RECT 276.600 666.000 278.400 672.600 ;
        RECT 279.600 670.800 282.300 672.600 ;
        RECT 279.600 666.600 281.400 670.800 ;
        RECT 296.100 666.600 297.900 672.600 ;
        RECT 299.100 671.700 306.900 673.050 ;
        RECT 299.100 666.600 300.900 671.700 ;
        RECT 302.100 666.000 303.900 670.800 ;
        RECT 305.100 666.600 306.900 671.700 ;
        RECT 320.700 669.600 321.900 679.950 ;
        RECT 341.100 678.150 342.900 679.950 ;
        RECT 344.100 675.600 345.300 679.950 ;
        RECT 347.100 678.150 348.900 679.950 ;
        RECT 359.550 679.050 360.450 680.550 ;
        RECT 364.950 679.950 367.050 682.050 ;
        RECT 367.950 679.950 370.050 682.050 ;
        RECT 370.950 679.950 373.050 682.050 ;
        RECT 373.950 679.950 376.050 682.050 ;
        RECT 376.950 679.950 379.050 682.050 ;
        RECT 391.950 679.950 394.050 682.050 ;
        RECT 394.950 679.950 397.050 682.050 ;
        RECT 409.950 679.950 412.050 682.050 ;
        RECT 412.950 679.950 415.050 682.050 ;
        RECT 415.950 679.950 418.050 682.050 ;
        RECT 418.950 679.950 421.050 682.050 ;
        RECT 437.100 679.950 439.200 682.050 ;
        RECT 440.400 679.950 442.500 682.050 ;
        RECT 359.550 677.550 364.050 679.050 ;
        RECT 365.100 678.150 366.900 679.950 ;
        RECT 360.000 676.950 364.050 677.550 ;
        RECT 341.700 674.700 345.300 675.600 ;
        RECT 341.700 672.600 342.900 674.700 ;
        RECT 320.100 666.600 321.900 669.600 ;
        RECT 323.100 666.000 324.900 669.600 ;
        RECT 341.100 666.600 342.900 672.600 ;
        RECT 344.100 671.700 351.900 673.050 ;
        RECT 371.700 672.600 372.900 679.950 ;
        RECT 376.950 678.150 378.750 679.950 ;
        RECT 373.950 675.450 376.050 676.050 ;
        RECT 385.950 675.450 388.050 676.050 ;
        RECT 373.950 674.550 388.050 675.450 ;
        RECT 373.950 673.950 376.050 674.550 ;
        RECT 385.950 673.950 388.050 674.550 ;
        RECT 344.100 666.600 345.900 671.700 ;
        RECT 347.100 666.000 348.900 670.800 ;
        RECT 350.100 666.600 351.900 671.700 ;
        RECT 367.500 666.000 369.300 672.600 ;
        RECT 372.000 666.600 373.800 672.600 ;
        RECT 376.500 666.000 378.300 672.600 ;
        RECT 392.700 669.600 393.900 679.950 ;
        RECT 413.100 678.150 414.900 679.950 ;
        RECT 416.700 675.600 417.900 679.950 ;
        RECT 419.100 678.150 420.900 679.950 ;
        RECT 416.700 674.700 420.300 675.600 ;
        RECT 410.100 671.700 417.900 673.050 ;
        RECT 392.100 666.600 393.900 669.600 ;
        RECT 395.100 666.000 396.900 669.600 ;
        RECT 410.100 666.600 411.900 671.700 ;
        RECT 413.100 666.000 414.900 670.800 ;
        RECT 416.100 666.600 417.900 671.700 ;
        RECT 419.100 672.600 420.300 674.700 ;
        RECT 437.700 672.600 438.600 679.950 ;
        RECT 444.000 675.300 444.900 695.400 ;
        RECT 461.100 689.400 462.900 702.000 ;
        RECT 466.200 690.600 468.000 701.400 ;
        RECT 485.700 695.400 487.500 702.000 ;
        RECT 486.000 692.100 487.800 693.900 ;
        RECT 488.700 690.900 490.500 701.400 ;
        RECT 464.400 689.400 468.000 690.600 ;
        RECT 488.100 689.400 490.500 690.900 ;
        RECT 493.800 689.400 495.600 702.000 ;
        RECT 509.100 689.400 510.900 702.000 ;
        RECT 514.200 690.600 516.000 701.400 ;
        RECT 533.100 695.400 534.900 701.400 ;
        RECT 536.100 696.000 537.900 702.000 ;
        RECT 512.400 689.400 516.000 690.600 ;
        RECT 534.000 695.100 534.900 695.400 ;
        RECT 539.100 695.400 540.900 701.400 ;
        RECT 542.100 695.400 543.900 702.000 ;
        RECT 539.100 695.100 540.600 695.400 ;
        RECT 534.000 694.200 540.600 695.100 ;
        RECT 461.250 682.050 463.050 683.850 ;
        RECT 464.400 682.050 465.300 689.400 ;
        RECT 467.100 682.050 468.900 683.850 ;
        RECT 488.100 682.050 489.300 689.400 ;
        RECT 494.100 682.050 495.900 683.850 ;
        RECT 509.250 682.050 511.050 683.850 ;
        RECT 512.400 682.050 513.300 689.400 ;
        RECT 514.950 687.450 517.050 688.050 ;
        RECT 520.950 687.450 523.050 687.900 ;
        RECT 514.950 686.550 523.050 687.450 ;
        RECT 514.950 685.950 517.050 686.550 ;
        RECT 520.950 685.800 523.050 686.550 ;
        RECT 515.100 682.050 516.900 683.850 ;
        RECT 534.000 682.050 534.900 694.200 ;
        RECT 560.100 689.400 561.900 701.400 ;
        RECT 563.100 690.300 564.900 701.400 ;
        RECT 566.100 691.200 567.900 702.000 ;
        RECT 569.100 690.300 570.900 701.400 ;
        RECT 563.100 689.400 570.900 690.300 ;
        RECT 585.600 689.400 587.400 702.000 ;
        RECT 590.100 689.400 593.400 701.400 ;
        RECT 596.100 689.400 597.900 702.000 ;
        RECT 611.100 695.400 612.900 702.000 ;
        RECT 614.100 695.400 615.900 701.400 ;
        RECT 617.100 695.400 618.900 702.000 ;
        RECT 635.100 695.400 636.900 702.000 ;
        RECT 638.100 695.400 639.900 701.400 ;
        RECT 541.950 687.450 544.050 688.050 ;
        RECT 556.950 687.450 559.050 688.050 ;
        RECT 541.950 686.550 559.050 687.450 ;
        RECT 541.950 685.950 544.050 686.550 ;
        RECT 556.950 685.950 559.050 686.550 ;
        RECT 539.100 682.050 540.900 683.850 ;
        RECT 560.400 682.050 561.300 689.400 ;
        RECT 565.950 682.050 567.750 683.850 ;
        RECT 584.250 682.050 586.050 683.850 ;
        RECT 591.000 682.050 592.050 689.400 ;
        RECT 596.100 682.050 597.900 683.850 ;
        RECT 614.100 682.050 615.300 695.400 ;
        RECT 635.100 682.050 636.900 683.850 ;
        RECT 638.100 682.050 639.300 695.400 ;
        RECT 654.000 690.600 655.800 701.400 ;
        RECT 654.000 689.400 657.600 690.600 ;
        RECT 659.100 689.400 660.900 702.000 ;
        RECT 677.100 690.600 678.900 701.400 ;
        RECT 680.100 691.500 682.200 702.000 ;
        RECT 677.100 689.400 682.200 690.600 ;
        RECT 684.600 690.300 686.400 701.400 ;
        RECT 689.100 691.500 690.900 702.000 ;
        RECT 692.100 690.300 693.900 701.400 ;
        RECT 653.100 682.050 654.900 683.850 ;
        RECT 656.700 682.050 657.600 689.400 ;
        RECT 680.100 688.500 682.200 689.400 ;
        RECT 683.100 689.400 686.400 690.300 ;
        RECT 658.950 687.450 661.050 688.050 ;
        RECT 664.950 687.450 667.050 688.050 ;
        RECT 658.950 686.550 667.050 687.450 ;
        RECT 658.950 685.950 661.050 686.550 ;
        RECT 664.950 685.950 667.050 686.550 ;
        RECT 683.100 685.050 684.300 689.400 ;
        RECT 689.100 689.100 693.900 690.300 ;
        RECT 710.400 689.400 712.200 702.000 ;
        RECT 715.500 690.900 717.300 701.400 ;
        RECT 718.500 695.400 720.300 702.000 ;
        RECT 718.200 692.100 720.000 693.900 ;
        RECT 715.500 689.400 717.900 690.900 ;
        RECT 737.100 690.300 738.900 701.400 ;
        RECT 740.100 691.200 741.900 702.000 ;
        RECT 743.100 690.300 744.900 701.400 ;
        RECT 737.100 689.400 744.900 690.300 ;
        RECT 746.100 689.400 747.900 701.400 ;
        RECT 761.100 695.400 762.900 701.400 ;
        RECT 764.100 695.400 765.900 702.000 ;
        RECT 689.100 688.200 691.200 689.100 ;
        RECT 685.800 687.300 691.200 688.200 ;
        RECT 685.800 685.500 687.600 687.300 ;
        RECT 682.800 684.300 684.900 685.050 ;
        RECT 658.950 682.050 660.750 683.850 ;
        RECT 677.400 682.050 679.200 683.850 ;
        RECT 682.800 682.950 685.800 684.300 ;
        RECT 445.800 679.950 447.900 682.050 ;
        RECT 460.950 679.950 463.050 682.050 ;
        RECT 463.950 679.950 466.050 682.050 ;
        RECT 466.950 679.950 469.050 682.050 ;
        RECT 484.950 679.950 487.050 682.050 ;
        RECT 487.950 679.950 490.050 682.050 ;
        RECT 490.950 679.950 493.050 682.050 ;
        RECT 493.950 679.950 496.050 682.050 ;
        RECT 508.950 679.950 511.050 682.050 ;
        RECT 511.950 679.950 514.050 682.050 ;
        RECT 514.950 679.950 517.050 682.050 ;
        RECT 532.950 679.950 535.050 682.050 ;
        RECT 535.950 679.950 538.050 682.050 ;
        RECT 538.950 679.950 541.050 682.050 ;
        RECT 541.950 679.950 544.050 682.050 ;
        RECT 559.950 679.950 562.050 682.050 ;
        RECT 562.950 679.950 565.050 682.050 ;
        RECT 565.950 679.950 568.050 682.050 ;
        RECT 568.950 679.950 571.050 682.050 ;
        RECT 583.950 679.950 586.050 682.050 ;
        RECT 586.950 679.950 589.050 682.050 ;
        RECT 589.950 679.950 592.050 682.050 ;
        RECT 445.950 678.150 447.750 679.950 ;
        RECT 439.500 674.400 447.900 675.300 ;
        RECT 439.500 673.500 441.300 674.400 ;
        RECT 419.100 666.600 420.900 672.600 ;
        RECT 437.700 670.800 440.400 672.600 ;
        RECT 438.600 666.600 440.400 670.800 ;
        RECT 441.600 666.000 443.400 672.600 ;
        RECT 446.100 666.600 447.900 674.400 ;
        RECT 464.400 669.600 465.300 679.950 ;
        RECT 485.100 678.150 486.900 679.950 ;
        RECT 488.100 675.600 489.300 679.950 ;
        RECT 491.100 678.150 492.900 679.950 ;
        RECT 485.700 674.700 489.300 675.600 ;
        RECT 485.700 672.600 486.900 674.700 ;
        RECT 461.100 666.000 462.900 669.600 ;
        RECT 464.100 666.600 465.900 669.600 ;
        RECT 467.100 666.000 468.900 669.600 ;
        RECT 485.100 666.600 486.900 672.600 ;
        RECT 488.100 671.700 495.900 673.050 ;
        RECT 488.100 666.600 489.900 671.700 ;
        RECT 491.100 666.000 492.900 670.800 ;
        RECT 494.100 666.600 495.900 671.700 ;
        RECT 512.400 669.600 513.300 679.950 ;
        RECT 534.000 676.200 534.900 679.950 ;
        RECT 536.100 678.150 537.900 679.950 ;
        RECT 542.100 678.150 543.900 679.950 ;
        RECT 534.000 675.000 537.300 676.200 ;
        RECT 509.100 666.000 510.900 669.600 ;
        RECT 512.100 666.600 513.900 669.600 ;
        RECT 515.100 666.000 516.900 669.600 ;
        RECT 535.500 666.600 537.300 675.000 ;
        RECT 542.100 666.000 543.900 675.600 ;
        RECT 560.400 672.600 561.300 679.950 ;
        RECT 562.950 678.150 564.750 679.950 ;
        RECT 569.100 678.150 570.900 679.950 ;
        RECT 587.250 678.150 589.050 679.950 ;
        RECT 591.000 675.300 592.050 679.950 ;
        RECT 592.950 679.950 595.050 682.050 ;
        RECT 595.950 679.950 598.050 682.050 ;
        RECT 610.950 679.950 613.050 682.050 ;
        RECT 613.950 679.950 616.050 682.050 ;
        RECT 616.950 679.950 619.050 682.050 ;
        RECT 634.950 679.950 637.050 682.050 ;
        RECT 637.950 679.950 640.050 682.050 ;
        RECT 652.950 679.950 655.050 682.050 ;
        RECT 655.950 679.950 658.050 682.050 ;
        RECT 658.950 679.950 661.050 682.050 ;
        RECT 677.100 679.950 679.200 682.050 ;
        RECT 682.200 680.100 684.000 681.900 ;
        RECT 592.950 678.150 594.750 679.950 ;
        RECT 611.250 678.150 613.050 679.950 ;
        RECT 587.700 674.100 592.050 675.300 ;
        RECT 614.100 674.700 615.300 679.950 ;
        RECT 617.100 678.150 618.900 679.950 ;
        RECT 587.700 672.600 588.600 674.100 ;
        RECT 614.100 673.800 618.300 674.700 ;
        RECT 560.400 671.400 565.500 672.600 ;
        RECT 560.700 666.000 562.500 669.600 ;
        RECT 563.700 666.600 565.500 671.400 ;
        RECT 568.200 666.000 570.000 672.600 ;
        RECT 584.100 667.500 585.900 672.600 ;
        RECT 587.100 668.400 588.900 672.600 ;
        RECT 590.100 672.000 597.900 672.900 ;
        RECT 590.100 667.500 591.900 672.000 ;
        RECT 584.100 666.600 591.900 667.500 ;
        RECT 593.100 666.000 594.900 671.100 ;
        RECT 596.100 666.600 597.900 672.000 ;
        RECT 611.400 666.000 613.200 672.600 ;
        RECT 616.500 666.600 618.300 673.800 ;
        RECT 638.100 669.600 639.300 679.950 ;
        RECT 656.700 669.600 657.600 679.950 ;
        RECT 661.950 678.450 664.050 679.050 ;
        RECT 667.950 678.450 670.050 679.050 ;
        RECT 661.950 677.550 670.050 678.450 ;
        RECT 681.900 678.000 684.000 680.100 ;
        RECT 661.950 676.950 664.050 677.550 ;
        RECT 667.950 676.950 670.050 677.550 ;
        RECT 684.900 676.200 685.800 682.950 ;
        RECT 687.300 682.200 689.100 684.000 ;
        RECT 687.000 680.100 689.100 682.200 ;
        RECT 710.100 682.050 711.900 683.850 ;
        RECT 716.700 682.050 717.900 689.400 ;
        RECT 721.950 684.450 726.000 685.050 ;
        RECT 721.950 682.950 726.450 684.450 ;
        RECT 691.800 679.800 693.900 682.050 ;
        RECT 709.950 679.950 712.050 682.050 ;
        RECT 712.950 679.950 715.050 682.050 ;
        RECT 715.950 679.950 718.050 682.050 ;
        RECT 718.950 679.950 721.050 682.050 ;
        RECT 691.800 679.200 693.600 679.800 ;
        RECT 687.000 678.000 693.600 679.200 ;
        RECT 713.100 678.150 714.900 679.950 ;
        RECT 687.000 677.100 689.100 678.000 ;
        RECT 679.500 673.500 681.600 675.900 ;
        RECT 682.800 674.100 685.800 676.200 ;
        RECT 686.700 675.300 688.500 677.100 ;
        RECT 716.700 675.600 717.900 679.950 ;
        RECT 719.100 678.150 720.900 679.950 ;
        RECT 725.550 679.050 726.450 682.950 ;
        RECT 740.250 682.050 742.050 683.850 ;
        RECT 746.700 682.050 747.600 689.400 ;
        RECT 761.700 682.050 762.900 695.400 ;
        RECT 782.100 690.300 783.900 701.400 ;
        RECT 785.100 691.200 786.900 702.000 ;
        RECT 788.100 690.300 789.900 701.400 ;
        RECT 782.100 689.400 789.900 690.300 ;
        RECT 791.100 689.400 792.900 701.400 ;
        RECT 806.100 695.400 807.900 702.000 ;
        RECT 809.100 695.400 810.900 701.400 ;
        RECT 812.100 696.000 813.900 702.000 ;
        RECT 809.400 695.100 810.900 695.400 ;
        RECT 815.100 695.400 816.900 701.400 ;
        RECT 830.100 695.400 831.900 702.000 ;
        RECT 833.100 695.400 834.900 701.400 ;
        RECT 815.100 695.100 816.000 695.400 ;
        RECT 809.400 694.200 816.000 695.100 ;
        RECT 769.950 687.450 772.050 688.050 ;
        RECT 781.950 687.450 784.050 688.200 ;
        RECT 769.950 686.550 784.050 687.450 ;
        RECT 769.950 685.950 772.050 686.550 ;
        RECT 781.950 686.100 784.050 686.550 ;
        RECT 764.100 682.050 765.900 683.850 ;
        RECT 785.250 682.050 787.050 683.850 ;
        RECT 791.700 682.050 792.600 689.400 ;
        RECT 793.950 687.450 796.050 688.050 ;
        RECT 811.950 687.450 814.050 688.050 ;
        RECT 793.950 686.550 814.050 687.450 ;
        RECT 793.950 685.950 796.050 686.550 ;
        RECT 811.950 685.950 814.050 686.550 ;
        RECT 809.100 682.050 810.900 683.850 ;
        RECT 815.100 682.050 816.000 694.200 ;
        RECT 828.000 687.450 832.050 688.050 ;
        RECT 827.550 685.950 832.050 687.450 ;
        RECT 827.550 684.450 828.450 685.950 ;
        RECT 824.550 683.550 828.450 684.450 ;
        RECT 736.950 679.950 739.050 682.050 ;
        RECT 739.950 679.950 742.050 682.050 ;
        RECT 742.950 679.950 745.050 682.050 ;
        RECT 745.950 679.950 748.050 682.050 ;
        RECT 760.950 679.950 763.050 682.050 ;
        RECT 763.950 679.950 766.050 682.050 ;
        RECT 781.950 679.950 784.050 682.050 ;
        RECT 784.950 679.950 787.050 682.050 ;
        RECT 787.950 679.950 790.050 682.050 ;
        RECT 790.950 679.950 793.050 682.050 ;
        RECT 805.950 679.950 808.050 682.050 ;
        RECT 808.950 679.950 811.050 682.050 ;
        RECT 811.950 679.950 814.050 682.050 ;
        RECT 814.950 679.950 817.050 682.050 ;
        RECT 721.950 677.550 726.450 679.050 ;
        RECT 737.100 678.150 738.900 679.950 ;
        RECT 743.250 678.150 745.050 679.950 ;
        RECT 721.950 676.950 726.000 677.550 ;
        RECT 677.100 672.600 681.600 673.500 ;
        RECT 635.100 666.000 636.900 669.600 ;
        RECT 638.100 666.600 639.900 669.600 ;
        RECT 653.100 666.000 654.900 669.600 ;
        RECT 656.100 666.600 657.900 669.600 ;
        RECT 659.100 666.000 660.900 669.600 ;
        RECT 677.100 666.600 678.900 672.600 ;
        RECT 684.900 672.000 685.800 674.100 ;
        RECT 689.400 675.000 691.500 675.600 ;
        RECT 689.400 673.500 693.900 675.000 ;
        RECT 716.700 674.700 720.300 675.600 ;
        RECT 692.400 672.600 693.900 673.500 ;
        RECT 680.400 666.000 682.200 671.700 ;
        RECT 684.900 666.600 686.700 672.000 ;
        RECT 689.100 666.000 690.900 671.700 ;
        RECT 692.100 666.600 693.900 672.600 ;
        RECT 710.100 671.700 717.900 673.050 ;
        RECT 710.100 666.600 711.900 671.700 ;
        RECT 713.100 666.000 714.900 670.800 ;
        RECT 716.100 666.600 717.900 671.700 ;
        RECT 719.100 672.600 720.300 674.700 ;
        RECT 746.700 672.600 747.600 679.950 ;
        RECT 719.100 666.600 720.900 672.600 ;
        RECT 738.000 666.000 739.800 672.600 ;
        RECT 742.500 671.400 747.600 672.600 ;
        RECT 742.500 666.600 744.300 671.400 ;
        RECT 761.700 669.600 762.900 679.950 ;
        RECT 766.950 678.450 769.050 679.050 ;
        RECT 772.950 678.450 775.050 679.050 ;
        RECT 766.950 677.550 775.050 678.450 ;
        RECT 782.100 678.150 783.900 679.950 ;
        RECT 788.250 678.150 790.050 679.950 ;
        RECT 766.950 676.950 769.050 677.550 ;
        RECT 772.950 676.950 775.050 677.550 ;
        RECT 791.700 672.600 792.600 679.950 ;
        RECT 806.100 678.150 807.900 679.950 ;
        RECT 812.100 678.150 813.900 679.950 ;
        RECT 815.100 676.200 816.000 679.950 ;
        RECT 824.550 679.050 825.450 683.550 ;
        RECT 830.100 682.050 831.900 683.850 ;
        RECT 833.100 682.050 834.300 695.400 ;
        RECT 848.100 690.300 849.900 701.400 ;
        RECT 851.100 691.200 852.900 702.000 ;
        RECT 854.100 690.300 855.900 701.400 ;
        RECT 848.100 689.400 855.900 690.300 ;
        RECT 857.100 689.400 858.900 701.400 ;
        RECT 872.400 689.400 874.200 702.000 ;
        RECT 877.500 690.900 879.300 701.400 ;
        RECT 880.500 695.400 882.300 702.000 ;
        RECT 880.200 692.100 882.000 693.900 ;
        RECT 877.500 689.400 879.900 690.900 ;
        RECT 896.400 689.400 898.200 702.000 ;
        RECT 901.500 690.900 903.300 701.400 ;
        RECT 904.500 695.400 906.300 702.000 ;
        RECT 920.100 695.400 921.900 701.400 ;
        RECT 923.100 695.400 924.900 702.000 ;
        RECT 931.950 699.450 934.050 700.050 ;
        RECT 937.950 699.450 940.050 699.900 ;
        RECT 931.950 698.550 940.050 699.450 ;
        RECT 931.950 697.950 934.050 698.550 ;
        RECT 937.950 697.800 940.050 698.550 ;
        RECT 904.200 692.100 906.000 693.900 ;
        RECT 901.500 689.400 903.900 690.900 ;
        RECT 851.250 682.050 853.050 683.850 ;
        RECT 857.700 682.050 858.600 689.400 ;
        RECT 867.000 684.450 871.050 685.050 ;
        RECT 866.550 682.950 871.050 684.450 ;
        RECT 829.950 679.950 832.050 682.050 ;
        RECT 832.950 679.950 835.050 682.050 ;
        RECT 847.950 679.950 850.050 682.050 ;
        RECT 850.950 679.950 853.050 682.050 ;
        RECT 853.950 679.950 856.050 682.050 ;
        RECT 856.950 679.950 859.050 682.050 ;
        RECT 824.550 677.550 829.050 679.050 ;
        RECT 825.000 676.950 829.050 677.550 ;
        RECT 745.500 666.000 747.300 669.600 ;
        RECT 761.100 666.600 762.900 669.600 ;
        RECT 764.100 666.000 765.900 669.600 ;
        RECT 783.000 666.000 784.800 672.600 ;
        RECT 787.500 671.400 792.600 672.600 ;
        RECT 787.500 666.600 789.300 671.400 ;
        RECT 790.500 666.000 792.300 669.600 ;
        RECT 806.100 666.000 807.900 675.600 ;
        RECT 812.700 675.000 816.000 676.200 ;
        RECT 817.950 675.450 820.050 676.050 ;
        RECT 823.950 675.450 826.050 676.050 ;
        RECT 812.700 666.600 814.500 675.000 ;
        RECT 817.950 674.550 826.050 675.450 ;
        RECT 817.950 673.950 820.050 674.550 ;
        RECT 823.950 673.950 826.050 674.550 ;
        RECT 833.100 669.600 834.300 679.950 ;
        RECT 848.100 678.150 849.900 679.950 ;
        RECT 854.250 678.150 856.050 679.950 ;
        RECT 857.700 672.600 858.600 679.950 ;
        RECT 859.950 678.450 862.050 679.050 ;
        RECT 866.550 678.450 867.450 682.950 ;
        RECT 872.100 682.050 873.900 683.850 ;
        RECT 878.700 682.050 879.900 689.400 ;
        RECT 896.100 682.050 897.900 683.850 ;
        RECT 902.700 682.050 903.900 689.400 ;
        RECT 904.950 687.450 907.050 688.050 ;
        RECT 910.950 687.450 913.050 688.050 ;
        RECT 904.950 686.550 913.050 687.450 ;
        RECT 904.950 685.950 907.050 686.550 ;
        RECT 910.950 685.950 913.050 686.550 ;
        RECT 920.700 682.050 921.900 695.400 ;
        RECT 941.100 690.300 942.900 701.400 ;
        RECT 944.100 691.200 945.900 702.000 ;
        RECT 947.100 690.300 948.900 701.400 ;
        RECT 941.100 689.400 948.900 690.300 ;
        RECT 950.100 689.400 951.900 701.400 ;
        RECT 965.100 695.400 966.900 702.000 ;
        RECT 968.100 695.400 969.900 701.400 ;
        RECT 955.950 690.450 958.050 690.900 ;
        RECT 964.950 690.450 967.050 691.050 ;
        RECT 955.950 689.550 967.050 690.450 ;
        RECT 931.950 687.450 934.050 688.050 ;
        RECT 946.950 687.450 949.050 688.050 ;
        RECT 931.950 686.550 949.050 687.450 ;
        RECT 931.950 685.950 934.050 686.550 ;
        RECT 946.950 685.950 949.050 686.550 ;
        RECT 923.100 682.050 924.900 683.850 ;
        RECT 944.250 682.050 946.050 683.850 ;
        RECT 950.700 682.050 951.600 689.400 ;
        RECT 955.950 688.800 958.050 689.550 ;
        RECT 964.950 688.950 967.050 689.550 ;
        RECT 965.100 682.050 966.900 683.850 ;
        RECT 968.100 682.050 969.300 695.400 ;
        RECT 983.100 690.300 984.900 701.400 ;
        RECT 986.100 691.200 987.900 702.000 ;
        RECT 989.100 690.300 990.900 701.400 ;
        RECT 983.100 689.400 990.900 690.300 ;
        RECT 992.100 689.400 993.900 701.400 ;
        RECT 986.250 682.050 988.050 683.850 ;
        RECT 992.700 682.050 993.600 689.400 ;
        RECT 871.950 679.950 874.050 682.050 ;
        RECT 874.950 679.950 877.050 682.050 ;
        RECT 877.950 679.950 880.050 682.050 ;
        RECT 880.950 679.950 883.050 682.050 ;
        RECT 895.950 679.950 898.050 682.050 ;
        RECT 898.950 679.950 901.050 682.050 ;
        RECT 901.950 679.950 904.050 682.050 ;
        RECT 904.950 679.950 907.050 682.050 ;
        RECT 919.950 679.950 922.050 682.050 ;
        RECT 922.950 679.950 925.050 682.050 ;
        RECT 934.950 679.950 937.050 682.050 ;
        RECT 940.950 679.950 943.050 682.050 ;
        RECT 943.950 679.950 946.050 682.050 ;
        RECT 946.950 679.950 949.050 682.050 ;
        RECT 949.950 679.950 952.050 682.050 ;
        RECT 859.950 677.550 867.450 678.450 ;
        RECT 875.100 678.150 876.900 679.950 ;
        RECT 859.950 676.950 862.050 677.550 ;
        RECT 878.700 675.600 879.900 679.950 ;
        RECT 881.100 678.150 882.900 679.950 ;
        RECT 899.100 678.150 900.900 679.950 ;
        RECT 902.700 675.600 903.900 679.950 ;
        RECT 905.100 678.150 906.900 679.950 ;
        RECT 878.700 674.700 882.300 675.600 ;
        RECT 902.700 674.700 906.300 675.600 ;
        RECT 830.100 666.000 831.900 669.600 ;
        RECT 833.100 666.600 834.900 669.600 ;
        RECT 849.000 666.000 850.800 672.600 ;
        RECT 853.500 671.400 858.600 672.600 ;
        RECT 872.100 671.700 879.900 673.050 ;
        RECT 853.500 666.600 855.300 671.400 ;
        RECT 856.500 666.000 858.300 669.600 ;
        RECT 872.100 666.600 873.900 671.700 ;
        RECT 875.100 666.000 876.900 670.800 ;
        RECT 878.100 666.600 879.900 671.700 ;
        RECT 881.100 672.600 882.300 674.700 ;
        RECT 881.100 666.600 882.900 672.600 ;
        RECT 896.100 671.700 903.900 673.050 ;
        RECT 896.100 666.600 897.900 671.700 ;
        RECT 899.100 666.000 900.900 670.800 ;
        RECT 902.100 666.600 903.900 671.700 ;
        RECT 905.100 672.600 906.300 674.700 ;
        RECT 905.100 666.600 906.900 672.600 ;
        RECT 920.700 669.600 921.900 679.950 ;
        RECT 925.950 678.450 928.050 679.050 ;
        RECT 931.950 678.450 934.050 679.050 ;
        RECT 925.950 677.550 934.050 678.450 ;
        RECT 925.950 676.950 928.050 677.550 ;
        RECT 931.950 676.950 934.050 677.550 ;
        RECT 935.550 675.450 936.450 679.950 ;
        RECT 941.100 678.150 942.900 679.950 ;
        RECT 947.250 678.150 949.050 679.950 ;
        RECT 946.950 675.450 949.050 676.050 ;
        RECT 935.550 674.550 949.050 675.450 ;
        RECT 946.950 673.950 949.050 674.550 ;
        RECT 950.700 672.600 951.600 679.950 ;
        RECT 952.950 678.450 955.050 679.050 ;
        RECT 958.950 678.450 961.050 682.050 ;
        RECT 964.950 679.950 967.050 682.050 ;
        RECT 967.950 679.950 970.050 682.050 ;
        RECT 982.950 679.950 985.050 682.050 ;
        RECT 985.950 679.950 988.050 682.050 ;
        RECT 988.950 679.950 991.050 682.050 ;
        RECT 991.950 679.950 994.050 682.050 ;
        RECT 952.950 678.000 961.050 678.450 ;
        RECT 952.950 677.550 960.450 678.000 ;
        RECT 952.950 676.950 955.050 677.550 ;
        RECT 920.100 666.600 921.900 669.600 ;
        RECT 923.100 666.000 924.900 669.600 ;
        RECT 942.000 666.000 943.800 672.600 ;
        RECT 946.500 671.400 951.600 672.600 ;
        RECT 946.500 666.600 948.300 671.400 ;
        RECT 968.100 669.600 969.300 679.950 ;
        RECT 973.950 678.450 976.050 679.050 ;
        RECT 979.950 678.450 982.050 679.050 ;
        RECT 973.950 677.550 982.050 678.450 ;
        RECT 983.100 678.150 984.900 679.950 ;
        RECT 989.250 678.150 991.050 679.950 ;
        RECT 973.950 676.950 976.050 677.550 ;
        RECT 979.950 676.950 982.050 677.550 ;
        RECT 970.950 675.450 973.050 676.050 ;
        RECT 988.950 675.450 991.050 676.050 ;
        RECT 970.950 674.550 991.050 675.450 ;
        RECT 970.950 673.950 973.050 674.550 ;
        RECT 988.950 673.950 991.050 674.550 ;
        RECT 973.950 672.450 976.050 673.050 ;
        RECT 979.950 672.450 982.050 673.050 ;
        RECT 992.700 672.600 993.600 679.950 ;
        RECT 997.950 675.450 1000.050 676.050 ;
        RECT 1003.950 675.450 1006.050 676.050 ;
        RECT 997.950 674.550 1006.050 675.450 ;
        RECT 997.950 673.950 1000.050 674.550 ;
        RECT 1003.950 673.950 1006.050 674.550 ;
        RECT 973.950 671.550 982.050 672.450 ;
        RECT 973.950 670.950 976.050 671.550 ;
        RECT 979.950 670.950 982.050 671.550 ;
        RECT 949.500 666.000 951.300 669.600 ;
        RECT 965.100 666.000 966.900 669.600 ;
        RECT 968.100 666.600 969.900 669.600 ;
        RECT 984.000 666.000 985.800 672.600 ;
        RECT 988.500 671.400 993.600 672.600 ;
        RECT 988.500 666.600 990.300 671.400 ;
        RECT 991.500 666.000 993.300 669.600 ;
        RECT 14.100 659.400 15.900 663.000 ;
        RECT 17.100 659.400 18.900 662.400 ;
        RECT 17.100 649.050 18.300 659.400 ;
        RECT 35.400 656.400 37.200 663.000 ;
        RECT 40.500 655.200 42.300 662.400 ;
        RECT 57.000 656.400 58.800 663.000 ;
        RECT 61.500 657.600 63.300 662.400 ;
        RECT 64.500 659.400 66.300 663.000 ;
        RECT 69.150 658.200 70.950 662.400 ;
        RECT 61.500 656.400 66.600 657.600 ;
        RECT 38.100 654.300 42.300 655.200 ;
        RECT 35.250 649.050 37.050 650.850 ;
        RECT 38.100 649.050 39.300 654.300 ;
        RECT 41.100 649.050 42.900 650.850 ;
        RECT 56.100 649.050 57.900 650.850 ;
        RECT 62.250 649.050 64.050 650.850 ;
        RECT 65.700 649.050 66.600 656.400 ;
        RECT 68.550 656.400 70.950 658.200 ;
        RECT 72.150 656.400 73.950 663.000 ;
        RECT 76.950 660.300 78.750 662.400 ;
        RECT 75.150 659.400 78.750 660.300 ;
        RECT 81.450 659.400 83.250 663.000 ;
        RECT 84.750 659.400 86.550 662.400 ;
        RECT 87.750 659.400 89.550 663.000 ;
        RECT 92.250 659.400 94.050 662.400 ;
        RECT 74.850 658.800 78.750 659.400 ;
        RECT 74.850 657.300 76.950 658.800 ;
        RECT 84.750 658.500 85.800 659.400 ;
        RECT 13.950 646.950 16.050 649.050 ;
        RECT 16.950 646.950 19.050 649.050 ;
        RECT 34.950 646.950 37.050 649.050 ;
        RECT 37.950 646.950 40.050 649.050 ;
        RECT 40.950 646.950 43.050 649.050 ;
        RECT 55.950 646.950 58.050 649.050 ;
        RECT 58.950 646.950 61.050 649.050 ;
        RECT 61.950 646.950 64.050 649.050 ;
        RECT 64.950 646.950 67.050 649.050 ;
        RECT 14.100 645.150 15.900 646.950 ;
        RECT 17.100 633.600 18.300 646.950 ;
        RECT 38.100 633.600 39.300 646.950 ;
        RECT 59.250 645.150 61.050 646.950 ;
        RECT 65.700 639.600 66.600 646.950 ;
        RECT 68.550 641.700 69.450 656.400 ;
        RECT 77.850 655.800 79.650 657.600 ;
        RECT 80.850 657.450 85.800 658.500 ;
        RECT 80.850 656.700 82.650 657.450 ;
        RECT 92.250 657.300 94.650 659.400 ;
        RECT 97.350 656.400 99.150 663.000 ;
        RECT 100.650 656.400 102.450 662.400 ;
        RECT 119.100 659.400 120.900 663.000 ;
        RECT 122.100 659.400 123.900 662.400 ;
        RECT 125.100 659.400 126.900 663.000 ;
        RECT 77.850 654.000 78.900 655.800 ;
        RECT 88.050 654.000 89.850 654.600 ;
        RECT 77.850 652.800 89.850 654.000 ;
        RECT 70.950 651.600 78.900 652.800 ;
        RECT 70.950 649.050 72.750 651.600 ;
        RECT 77.100 651.000 78.900 651.600 ;
        RECT 74.100 649.800 75.900 650.400 ;
        RECT 70.950 646.950 73.050 649.050 ;
        RECT 74.100 648.600 82.200 649.800 ;
        RECT 80.100 646.950 82.200 648.600 ;
        RECT 78.450 641.700 80.250 642.000 ;
        RECT 68.550 641.100 80.250 641.700 ;
        RECT 68.550 640.500 86.850 641.100 ;
        RECT 68.550 639.600 69.450 640.500 ;
        RECT 78.450 640.200 86.850 640.500 ;
        RECT 56.100 638.700 63.900 639.600 ;
        RECT 14.100 627.000 15.900 633.600 ;
        RECT 17.100 627.600 18.900 633.600 ;
        RECT 35.100 627.000 36.900 633.600 ;
        RECT 38.100 627.600 39.900 633.600 ;
        RECT 41.100 627.000 42.900 633.600 ;
        RECT 56.100 627.600 57.900 638.700 ;
        RECT 59.100 627.000 60.900 637.800 ;
        RECT 62.100 627.600 63.900 638.700 ;
        RECT 65.100 627.600 66.900 639.600 ;
        RECT 68.550 637.800 70.950 639.600 ;
        RECT 69.150 627.600 70.950 637.800 ;
        RECT 72.150 627.000 73.950 639.600 ;
        RECT 83.250 638.700 85.050 639.300 ;
        RECT 77.250 637.500 85.050 638.700 ;
        RECT 85.950 638.100 86.850 640.200 ;
        RECT 88.950 640.200 89.850 652.800 ;
        RECT 101.250 649.050 102.450 656.400 ;
        RECT 122.700 649.050 123.600 659.400 ;
        RECT 140.100 657.300 141.900 662.400 ;
        RECT 143.100 658.200 144.900 663.000 ;
        RECT 146.100 657.300 147.900 662.400 ;
        RECT 140.100 655.950 147.900 657.300 ;
        RECT 149.100 656.400 150.900 662.400 ;
        RECT 149.100 654.300 150.300 656.400 ;
        RECT 167.700 655.200 169.500 662.400 ;
        RECT 172.800 656.400 174.600 663.000 ;
        RECT 177.150 658.200 178.950 662.400 ;
        RECT 176.550 656.400 178.950 658.200 ;
        RECT 180.150 656.400 181.950 663.000 ;
        RECT 184.950 660.300 186.750 662.400 ;
        RECT 183.150 659.400 186.750 660.300 ;
        RECT 189.450 659.400 191.250 663.000 ;
        RECT 192.750 659.400 194.550 662.400 ;
        RECT 195.750 659.400 197.550 663.000 ;
        RECT 200.250 659.400 202.050 662.400 ;
        RECT 182.850 658.800 186.750 659.400 ;
        RECT 182.850 657.300 184.950 658.800 ;
        RECT 192.750 658.500 193.800 659.400 ;
        RECT 167.700 654.300 171.900 655.200 ;
        RECT 146.700 653.400 150.300 654.300 ;
        RECT 127.950 651.450 132.000 652.050 ;
        RECT 127.950 649.950 132.450 651.450 ;
        RECT 96.150 647.250 102.450 649.050 ;
        RECT 97.950 646.950 102.450 647.250 ;
        RECT 118.950 646.950 121.050 649.050 ;
        RECT 121.950 646.950 124.050 649.050 ;
        RECT 124.950 646.950 127.050 649.050 ;
        RECT 131.550 648.450 132.450 649.950 ;
        RECT 143.100 649.050 144.900 650.850 ;
        RECT 146.700 649.050 147.900 653.400 ;
        RECT 149.100 649.050 150.900 650.850 ;
        RECT 167.100 649.050 168.900 650.850 ;
        RECT 170.700 649.050 171.900 654.300 ;
        RECT 172.950 649.050 174.750 650.850 ;
        RECT 131.550 647.550 135.450 648.450 ;
        RECT 92.550 644.100 94.650 644.400 ;
        RECT 98.550 644.100 100.350 644.250 ;
        RECT 92.550 642.900 100.350 644.100 ;
        RECT 92.550 642.300 94.650 642.900 ;
        RECT 98.550 642.450 100.350 642.900 ;
        RECT 88.950 639.300 93.750 640.200 ;
        RECT 101.250 639.600 102.450 646.950 ;
        RECT 119.100 645.150 120.900 646.950 ;
        RECT 122.700 639.600 123.600 646.950 ;
        RECT 124.950 645.150 126.750 646.950 ;
        RECT 134.550 646.050 135.450 647.550 ;
        RECT 139.950 646.950 142.050 649.050 ;
        RECT 142.950 646.950 145.050 649.050 ;
        RECT 145.950 646.950 148.050 649.050 ;
        RECT 148.950 646.950 151.050 649.050 ;
        RECT 166.950 646.950 169.050 649.050 ;
        RECT 169.950 646.950 172.050 649.050 ;
        RECT 172.950 646.950 175.050 649.050 ;
        RECT 134.550 644.550 139.050 646.050 ;
        RECT 140.100 645.150 141.900 646.950 ;
        RECT 135.000 643.950 139.050 644.550 ;
        RECT 124.950 642.450 127.050 643.050 ;
        RECT 133.950 642.450 136.050 643.050 ;
        RECT 124.950 641.550 136.050 642.450 ;
        RECT 124.950 640.950 127.050 641.550 ;
        RECT 133.950 640.950 136.050 641.550 ;
        RECT 146.700 639.600 147.900 646.950 ;
        RECT 92.550 638.400 93.750 639.300 ;
        RECT 89.850 638.100 91.650 638.400 ;
        RECT 77.250 636.600 79.350 637.500 ;
        RECT 85.950 637.200 91.650 638.100 ;
        RECT 89.850 636.600 91.650 637.200 ;
        RECT 92.550 636.600 95.550 638.400 ;
        RECT 77.550 627.600 79.350 636.600 ;
        RECT 81.450 635.550 83.250 636.300 ;
        RECT 86.250 635.550 88.050 636.300 ;
        RECT 81.450 634.500 88.050 635.550 ;
        RECT 82.350 627.000 84.150 633.600 ;
        RECT 85.350 627.600 87.150 634.500 ;
        RECT 92.550 633.600 94.650 635.700 ;
        RECT 88.350 627.000 90.150 633.600 ;
        RECT 92.850 627.600 94.650 633.600 ;
        RECT 97.650 627.000 99.450 639.600 ;
        RECT 100.650 627.600 102.450 639.600 ;
        RECT 120.000 638.400 123.600 639.600 ;
        RECT 120.000 627.600 121.800 638.400 ;
        RECT 125.100 627.000 126.900 639.600 ;
        RECT 140.400 627.000 142.200 639.600 ;
        RECT 145.500 638.100 147.900 639.600 ;
        RECT 145.500 627.600 147.300 638.100 ;
        RECT 148.200 635.100 150.000 636.900 ;
        RECT 170.700 633.600 171.900 646.950 ;
        RECT 176.550 641.700 177.450 656.400 ;
        RECT 185.850 655.800 187.650 657.600 ;
        RECT 188.850 657.450 193.800 658.500 ;
        RECT 188.850 656.700 190.650 657.450 ;
        RECT 200.250 657.300 202.650 659.400 ;
        RECT 205.350 656.400 207.150 663.000 ;
        RECT 208.650 656.400 210.450 662.400 ;
        RECT 185.850 654.000 186.900 655.800 ;
        RECT 196.050 654.000 197.850 654.600 ;
        RECT 185.850 652.800 197.850 654.000 ;
        RECT 178.950 651.600 186.900 652.800 ;
        RECT 178.950 649.050 180.750 651.600 ;
        RECT 185.100 651.000 186.900 651.600 ;
        RECT 182.100 649.800 183.900 650.400 ;
        RECT 178.950 646.950 181.050 649.050 ;
        RECT 182.100 648.600 190.200 649.800 ;
        RECT 188.100 646.950 190.200 648.600 ;
        RECT 186.450 641.700 188.250 642.000 ;
        RECT 176.550 641.100 188.250 641.700 ;
        RECT 176.550 640.500 194.850 641.100 ;
        RECT 176.550 639.600 177.450 640.500 ;
        RECT 186.450 640.200 194.850 640.500 ;
        RECT 176.550 637.800 178.950 639.600 ;
        RECT 148.500 627.000 150.300 633.600 ;
        RECT 167.100 627.000 168.900 633.600 ;
        RECT 170.100 627.600 171.900 633.600 ;
        RECT 173.100 627.000 174.900 633.600 ;
        RECT 177.150 627.600 178.950 637.800 ;
        RECT 180.150 627.000 181.950 639.600 ;
        RECT 191.250 638.700 193.050 639.300 ;
        RECT 185.250 637.500 193.050 638.700 ;
        RECT 193.950 638.100 194.850 640.200 ;
        RECT 196.950 640.200 197.850 652.800 ;
        RECT 209.250 649.050 210.450 656.400 ;
        RECT 224.100 656.400 225.900 662.400 ;
        RECT 227.100 657.300 228.900 663.000 ;
        RECT 231.600 656.400 233.400 662.400 ;
        RECT 236.100 657.300 237.900 663.000 ;
        RECT 239.100 656.400 240.900 662.400 ;
        RECT 257.100 656.400 258.900 662.400 ;
        RECT 224.100 655.500 228.900 656.400 ;
        RECT 226.800 654.300 228.900 655.500 ;
        RECT 231.900 654.900 233.100 656.400 ;
        RECT 230.100 652.800 233.100 654.900 ;
        RECT 239.100 654.600 240.300 656.400 ;
        RECT 228.900 649.800 231.000 651.900 ;
        RECT 204.150 647.250 210.450 649.050 ;
        RECT 205.950 646.950 210.450 647.250 ;
        RECT 224.100 646.950 226.200 649.050 ;
        RECT 228.900 648.000 230.700 649.800 ;
        RECT 231.900 647.100 233.100 652.800 ;
        RECT 234.000 653.700 240.300 654.600 ;
        RECT 257.700 654.300 258.900 656.400 ;
        RECT 260.100 657.300 261.900 662.400 ;
        RECT 263.100 658.200 264.900 663.000 ;
        RECT 266.100 657.300 267.900 662.400 ;
        RECT 284.100 659.400 285.900 663.000 ;
        RECT 287.100 659.400 288.900 662.400 ;
        RECT 290.100 659.400 291.900 663.000 ;
        RECT 260.100 655.950 267.900 657.300 ;
        RECT 234.000 651.600 236.100 653.700 ;
        RECT 257.700 653.400 261.300 654.300 ;
        RECT 234.000 649.800 235.800 651.600 ;
        RECT 238.800 649.050 240.600 650.850 ;
        RECT 257.100 649.050 258.900 650.850 ;
        RECT 260.100 649.050 261.300 653.400 ;
        RECT 263.100 649.050 264.900 650.850 ;
        RECT 287.400 649.050 288.300 659.400 ;
        RECT 293.550 656.400 295.350 662.400 ;
        RECT 296.850 656.400 298.650 663.000 ;
        RECT 301.950 659.400 303.750 662.400 ;
        RECT 306.450 659.400 308.250 663.000 ;
        RECT 309.450 659.400 311.250 662.400 ;
        RECT 312.750 659.400 314.550 663.000 ;
        RECT 317.250 660.300 319.050 662.400 ;
        RECT 317.250 659.400 320.850 660.300 ;
        RECT 301.350 657.300 303.750 659.400 ;
        RECT 310.200 658.500 311.250 659.400 ;
        RECT 317.250 658.800 321.150 659.400 ;
        RECT 310.200 657.450 315.150 658.500 ;
        RECT 313.350 656.700 315.150 657.450 ;
        RECT 293.550 649.050 294.750 656.400 ;
        RECT 316.350 655.800 318.150 657.600 ;
        RECT 319.050 657.300 321.150 658.800 ;
        RECT 322.050 656.400 323.850 663.000 ;
        RECT 325.050 658.200 326.850 662.400 ;
        RECT 325.050 656.400 327.450 658.200 ;
        RECT 344.400 656.400 346.200 663.000 ;
        RECT 306.150 654.000 307.950 654.600 ;
        RECT 317.100 654.000 318.150 655.800 ;
        RECT 306.150 652.800 318.150 654.000 ;
        RECT 238.800 648.300 240.900 649.050 ;
        RECT 200.550 644.100 202.650 644.400 ;
        RECT 206.550 644.100 208.350 644.250 ;
        RECT 200.550 642.900 208.350 644.100 ;
        RECT 200.550 642.300 202.650 642.900 ;
        RECT 206.550 642.450 208.350 642.900 ;
        RECT 196.950 639.300 201.750 640.200 ;
        RECT 209.250 639.600 210.450 646.950 ;
        RECT 224.400 645.150 226.200 646.950 ;
        RECT 230.700 646.200 233.100 647.100 ;
        RECT 234.000 646.950 240.900 648.300 ;
        RECT 256.950 646.950 259.050 649.050 ;
        RECT 259.950 646.950 262.050 649.050 ;
        RECT 262.950 646.950 265.050 649.050 ;
        RECT 265.950 646.950 268.050 649.050 ;
        RECT 283.950 646.950 286.050 649.050 ;
        RECT 286.950 646.950 289.050 649.050 ;
        RECT 289.950 646.950 292.050 649.050 ;
        RECT 293.550 647.250 299.850 649.050 ;
        RECT 293.550 646.950 298.050 647.250 ;
        RECT 234.000 646.500 235.800 646.950 ;
        RECT 230.700 646.050 232.200 646.200 ;
        RECT 230.100 643.950 232.200 646.050 ;
        RECT 231.300 642.000 232.200 643.950 ;
        RECT 233.100 643.500 237.000 645.300 ;
        RECT 233.100 643.200 235.200 643.500 ;
        RECT 231.300 640.950 232.800 642.000 ;
        RECT 226.800 639.600 228.900 640.500 ;
        RECT 200.550 638.400 201.750 639.300 ;
        RECT 197.850 638.100 199.650 638.400 ;
        RECT 185.250 636.600 187.350 637.500 ;
        RECT 193.950 637.200 199.650 638.100 ;
        RECT 197.850 636.600 199.650 637.200 ;
        RECT 200.550 636.600 203.550 638.400 ;
        RECT 185.550 627.600 187.350 636.600 ;
        RECT 189.450 635.550 191.250 636.300 ;
        RECT 194.250 635.550 196.050 636.300 ;
        RECT 189.450 634.500 196.050 635.550 ;
        RECT 190.350 627.000 192.150 633.600 ;
        RECT 193.350 627.600 195.150 634.500 ;
        RECT 200.550 633.600 202.650 635.700 ;
        RECT 196.350 627.000 198.150 633.600 ;
        RECT 200.850 627.600 202.650 633.600 ;
        RECT 205.650 627.000 207.450 639.600 ;
        RECT 208.650 627.600 210.450 639.600 ;
        RECT 224.100 638.400 228.900 639.600 ;
        RECT 231.600 639.600 232.800 640.950 ;
        RECT 236.400 639.600 238.500 641.700 ;
        RECT 260.100 639.600 261.300 646.950 ;
        RECT 266.100 645.150 267.900 646.950 ;
        RECT 284.250 645.150 286.050 646.950 ;
        RECT 287.400 639.600 288.300 646.950 ;
        RECT 290.100 645.150 291.900 646.950 ;
        RECT 293.550 639.600 294.750 646.950 ;
        RECT 295.650 644.100 297.450 644.250 ;
        RECT 301.350 644.100 303.450 644.400 ;
        RECT 295.650 642.900 303.450 644.100 ;
        RECT 295.650 642.450 297.450 642.900 ;
        RECT 301.350 642.300 303.450 642.900 ;
        RECT 306.150 640.200 307.050 652.800 ;
        RECT 317.100 651.600 325.050 652.800 ;
        RECT 317.100 651.000 318.900 651.600 ;
        RECT 320.100 649.800 321.900 650.400 ;
        RECT 313.800 648.600 321.900 649.800 ;
        RECT 323.250 649.050 325.050 651.600 ;
        RECT 313.800 646.950 315.900 648.600 ;
        RECT 322.950 646.950 325.050 649.050 ;
        RECT 315.750 641.700 317.550 642.000 ;
        RECT 326.550 641.700 327.450 656.400 ;
        RECT 349.500 655.200 351.300 662.400 ;
        RECT 354.150 658.200 355.950 662.400 ;
        RECT 328.950 654.450 331.050 655.050 ;
        RECT 343.950 654.450 346.050 655.050 ;
        RECT 328.950 653.550 346.050 654.450 ;
        RECT 328.950 652.950 331.050 653.550 ;
        RECT 343.950 652.950 346.050 653.550 ;
        RECT 347.100 654.300 351.300 655.200 ;
        RECT 353.550 656.400 355.950 658.200 ;
        RECT 357.150 656.400 358.950 663.000 ;
        RECT 361.950 660.300 363.750 662.400 ;
        RECT 360.150 659.400 363.750 660.300 ;
        RECT 366.450 659.400 368.250 663.000 ;
        RECT 369.750 659.400 371.550 662.400 ;
        RECT 372.750 659.400 374.550 663.000 ;
        RECT 377.250 659.400 379.050 662.400 ;
        RECT 359.850 658.800 363.750 659.400 ;
        RECT 359.850 657.300 361.950 658.800 ;
        RECT 369.750 658.500 370.800 659.400 ;
        RECT 344.250 649.050 346.050 650.850 ;
        RECT 347.100 649.050 348.300 654.300 ;
        RECT 350.100 649.050 351.900 650.850 ;
        RECT 343.950 646.950 346.050 649.050 ;
        RECT 346.950 646.950 349.050 649.050 ;
        RECT 349.950 646.950 352.050 649.050 ;
        RECT 315.750 641.100 327.450 641.700 ;
        RECT 224.100 627.600 225.900 638.400 ;
        RECT 227.100 627.000 228.900 637.500 ;
        RECT 231.600 627.600 233.400 639.600 ;
        RECT 236.400 638.700 240.900 639.600 ;
        RECT 236.100 627.000 237.900 637.500 ;
        RECT 239.100 627.600 240.900 638.700 ;
        RECT 260.100 638.100 262.500 639.600 ;
        RECT 258.000 635.100 259.800 636.900 ;
        RECT 257.700 627.000 259.500 633.600 ;
        RECT 260.700 627.600 262.500 638.100 ;
        RECT 265.800 627.000 267.600 639.600 ;
        RECT 284.100 627.000 285.900 639.600 ;
        RECT 287.400 638.400 291.000 639.600 ;
        RECT 289.200 627.600 291.000 638.400 ;
        RECT 293.550 627.600 295.350 639.600 ;
        RECT 296.550 627.000 298.350 639.600 ;
        RECT 302.250 639.300 307.050 640.200 ;
        RECT 309.150 640.500 327.450 641.100 ;
        RECT 309.150 640.200 317.550 640.500 ;
        RECT 302.250 638.400 303.450 639.300 ;
        RECT 300.450 636.600 303.450 638.400 ;
        RECT 304.350 638.100 306.150 638.400 ;
        RECT 309.150 638.100 310.050 640.200 ;
        RECT 326.550 639.600 327.450 640.500 ;
        RECT 304.350 637.200 310.050 638.100 ;
        RECT 310.950 638.700 312.750 639.300 ;
        RECT 310.950 637.500 318.750 638.700 ;
        RECT 304.350 636.600 306.150 637.200 ;
        RECT 316.650 636.600 318.750 637.500 ;
        RECT 301.350 633.600 303.450 635.700 ;
        RECT 307.950 635.550 309.750 636.300 ;
        RECT 312.750 635.550 314.550 636.300 ;
        RECT 307.950 634.500 314.550 635.550 ;
        RECT 301.350 627.600 303.150 633.600 ;
        RECT 305.850 627.000 307.650 633.600 ;
        RECT 308.850 627.600 310.650 634.500 ;
        RECT 311.850 627.000 313.650 633.600 ;
        RECT 316.650 627.600 318.450 636.600 ;
        RECT 322.050 627.000 323.850 639.600 ;
        RECT 325.050 637.800 327.450 639.600 ;
        RECT 325.050 627.600 326.850 637.800 ;
        RECT 347.100 633.600 348.300 646.950 ;
        RECT 353.550 641.700 354.450 656.400 ;
        RECT 362.850 655.800 364.650 657.600 ;
        RECT 365.850 657.450 370.800 658.500 ;
        RECT 365.850 656.700 367.650 657.450 ;
        RECT 377.250 657.300 379.650 659.400 ;
        RECT 382.350 656.400 384.150 663.000 ;
        RECT 385.650 656.400 387.450 662.400 ;
        RECT 390.150 658.200 391.950 662.400 ;
        RECT 362.850 654.000 363.900 655.800 ;
        RECT 373.050 654.000 374.850 654.600 ;
        RECT 362.850 652.800 374.850 654.000 ;
        RECT 355.950 651.600 363.900 652.800 ;
        RECT 355.950 649.050 357.750 651.600 ;
        RECT 362.100 651.000 363.900 651.600 ;
        RECT 359.100 649.800 360.900 650.400 ;
        RECT 355.950 646.950 358.050 649.050 ;
        RECT 359.100 648.600 367.200 649.800 ;
        RECT 365.100 646.950 367.200 648.600 ;
        RECT 363.450 641.700 365.250 642.000 ;
        RECT 353.550 641.100 365.250 641.700 ;
        RECT 353.550 640.500 371.850 641.100 ;
        RECT 353.550 639.600 354.450 640.500 ;
        RECT 363.450 640.200 371.850 640.500 ;
        RECT 353.550 637.800 355.950 639.600 ;
        RECT 344.100 627.000 345.900 633.600 ;
        RECT 347.100 627.600 348.900 633.600 ;
        RECT 350.100 627.000 351.900 633.600 ;
        RECT 354.150 627.600 355.950 637.800 ;
        RECT 357.150 627.000 358.950 639.600 ;
        RECT 368.250 638.700 370.050 639.300 ;
        RECT 362.250 637.500 370.050 638.700 ;
        RECT 370.950 638.100 371.850 640.200 ;
        RECT 373.950 640.200 374.850 652.800 ;
        RECT 386.250 649.050 387.450 656.400 ;
        RECT 381.150 647.250 387.450 649.050 ;
        RECT 382.950 646.950 387.450 647.250 ;
        RECT 377.550 644.100 379.650 644.400 ;
        RECT 383.550 644.100 385.350 644.250 ;
        RECT 377.550 642.900 385.350 644.100 ;
        RECT 377.550 642.300 379.650 642.900 ;
        RECT 383.550 642.450 385.350 642.900 ;
        RECT 373.950 639.300 378.750 640.200 ;
        RECT 386.250 639.600 387.450 646.950 ;
        RECT 377.550 638.400 378.750 639.300 ;
        RECT 374.850 638.100 376.650 638.400 ;
        RECT 362.250 636.600 364.350 637.500 ;
        RECT 370.950 637.200 376.650 638.100 ;
        RECT 374.850 636.600 376.650 637.200 ;
        RECT 377.550 636.600 380.550 638.400 ;
        RECT 362.550 627.600 364.350 636.600 ;
        RECT 366.450 635.550 368.250 636.300 ;
        RECT 371.250 635.550 373.050 636.300 ;
        RECT 366.450 634.500 373.050 635.550 ;
        RECT 367.350 627.000 369.150 633.600 ;
        RECT 370.350 627.600 372.150 634.500 ;
        RECT 377.550 633.600 379.650 635.700 ;
        RECT 373.350 627.000 375.150 633.600 ;
        RECT 377.850 627.600 379.650 633.600 ;
        RECT 382.650 627.000 384.450 639.600 ;
        RECT 385.650 627.600 387.450 639.600 ;
        RECT 389.550 656.400 391.950 658.200 ;
        RECT 393.150 656.400 394.950 663.000 ;
        RECT 397.950 660.300 399.750 662.400 ;
        RECT 396.150 659.400 399.750 660.300 ;
        RECT 402.450 659.400 404.250 663.000 ;
        RECT 405.750 659.400 407.550 662.400 ;
        RECT 408.750 659.400 410.550 663.000 ;
        RECT 413.250 659.400 415.050 662.400 ;
        RECT 395.850 658.800 399.750 659.400 ;
        RECT 395.850 657.300 397.950 658.800 ;
        RECT 405.750 658.500 406.800 659.400 ;
        RECT 389.550 641.700 390.450 656.400 ;
        RECT 398.850 655.800 400.650 657.600 ;
        RECT 401.850 657.450 406.800 658.500 ;
        RECT 401.850 656.700 403.650 657.450 ;
        RECT 413.250 657.300 415.650 659.400 ;
        RECT 418.350 656.400 420.150 663.000 ;
        RECT 421.650 656.400 423.450 662.400 ;
        RECT 437.100 656.400 438.900 662.400 ;
        RECT 398.850 654.000 399.900 655.800 ;
        RECT 409.050 654.000 410.850 654.600 ;
        RECT 398.850 652.800 410.850 654.000 ;
        RECT 391.950 651.600 399.900 652.800 ;
        RECT 391.950 649.050 393.750 651.600 ;
        RECT 398.100 651.000 399.900 651.600 ;
        RECT 395.100 649.800 396.900 650.400 ;
        RECT 391.950 646.950 394.050 649.050 ;
        RECT 395.100 648.600 403.200 649.800 ;
        RECT 401.100 646.950 403.200 648.600 ;
        RECT 399.450 641.700 401.250 642.000 ;
        RECT 389.550 641.100 401.250 641.700 ;
        RECT 389.550 640.500 407.850 641.100 ;
        RECT 389.550 639.600 390.450 640.500 ;
        RECT 399.450 640.200 407.850 640.500 ;
        RECT 389.550 637.800 391.950 639.600 ;
        RECT 390.150 627.600 391.950 637.800 ;
        RECT 393.150 627.000 394.950 639.600 ;
        RECT 404.250 638.700 406.050 639.300 ;
        RECT 398.250 637.500 406.050 638.700 ;
        RECT 406.950 638.100 407.850 640.200 ;
        RECT 409.950 640.200 410.850 652.800 ;
        RECT 422.250 649.050 423.450 656.400 ;
        RECT 437.700 654.300 438.900 656.400 ;
        RECT 440.100 657.300 441.900 662.400 ;
        RECT 443.100 658.200 444.900 663.000 ;
        RECT 446.100 657.300 447.900 662.400 ;
        RECT 440.100 655.950 447.900 657.300 ;
        RECT 461.400 656.400 463.200 663.000 ;
        RECT 466.500 655.200 468.300 662.400 ;
        RECT 464.100 654.300 468.300 655.200 ;
        RECT 437.700 653.400 441.300 654.300 ;
        RECT 437.100 649.050 438.900 650.850 ;
        RECT 440.100 649.050 441.300 653.400 ;
        RECT 443.100 649.050 444.900 650.850 ;
        RECT 461.250 649.050 463.050 650.850 ;
        RECT 464.100 649.050 465.300 654.300 ;
        RECT 485.100 653.400 486.900 663.000 ;
        RECT 491.700 654.000 493.500 662.400 ;
        RECT 512.100 657.300 513.900 662.400 ;
        RECT 515.100 658.200 516.900 663.000 ;
        RECT 518.100 657.300 519.900 662.400 ;
        RECT 512.100 655.950 519.900 657.300 ;
        RECT 521.100 656.400 522.900 662.400 ;
        RECT 521.100 654.300 522.300 656.400 ;
        RECT 491.700 652.800 495.000 654.000 ;
        RECT 467.100 649.050 468.900 650.850 ;
        RECT 485.100 649.050 486.900 650.850 ;
        RECT 491.100 649.050 492.900 650.850 ;
        RECT 494.100 649.050 495.000 652.800 ;
        RECT 518.700 653.400 522.300 654.300 ;
        RECT 536.100 654.600 537.900 662.400 ;
        RECT 540.600 656.400 542.400 663.000 ;
        RECT 543.600 658.200 545.400 662.400 ;
        RECT 543.600 656.400 546.300 658.200 ;
        RECT 561.000 656.400 562.800 663.000 ;
        RECT 565.500 657.600 567.300 662.400 ;
        RECT 568.500 659.400 570.300 663.000 ;
        RECT 565.500 656.400 570.600 657.600 ;
        RECT 587.100 656.400 588.900 663.000 ;
        RECT 590.100 656.400 591.900 662.400 ;
        RECT 608.100 656.400 609.900 662.400 ;
        RECT 611.100 657.300 612.900 663.000 ;
        RECT 615.600 656.400 617.400 662.400 ;
        RECT 620.100 657.300 621.900 663.000 ;
        RECT 623.100 656.400 624.900 662.400 ;
        RECT 638.100 656.400 639.900 662.400 ;
        RECT 542.700 654.600 544.500 655.500 ;
        RECT 536.100 653.700 544.500 654.600 ;
        RECT 515.100 649.050 516.900 650.850 ;
        RECT 518.700 649.050 519.900 653.400 ;
        RECT 521.100 649.050 522.900 650.850 ;
        RECT 536.250 649.050 538.050 650.850 ;
        RECT 417.150 647.250 423.450 649.050 ;
        RECT 418.950 646.950 423.450 647.250 ;
        RECT 436.950 646.950 439.050 649.050 ;
        RECT 439.950 646.950 442.050 649.050 ;
        RECT 442.950 646.950 445.050 649.050 ;
        RECT 445.950 646.950 448.050 649.050 ;
        RECT 460.950 646.950 463.050 649.050 ;
        RECT 463.950 646.950 466.050 649.050 ;
        RECT 466.950 646.950 469.050 649.050 ;
        RECT 484.950 646.950 487.050 649.050 ;
        RECT 487.950 646.950 490.050 649.050 ;
        RECT 490.950 646.950 493.050 649.050 ;
        RECT 493.950 646.950 496.050 649.050 ;
        RECT 511.950 646.950 514.050 649.050 ;
        RECT 514.950 646.950 517.050 649.050 ;
        RECT 517.950 646.950 520.050 649.050 ;
        RECT 520.950 646.950 523.050 649.050 ;
        RECT 536.100 646.950 538.200 649.050 ;
        RECT 413.550 644.100 415.650 644.400 ;
        RECT 419.550 644.100 421.350 644.250 ;
        RECT 413.550 642.900 421.350 644.100 ;
        RECT 413.550 642.300 415.650 642.900 ;
        RECT 419.550 642.450 421.350 642.900 ;
        RECT 409.950 639.300 414.750 640.200 ;
        RECT 422.250 639.600 423.450 646.950 ;
        RECT 413.550 638.400 414.750 639.300 ;
        RECT 410.850 638.100 412.650 638.400 ;
        RECT 398.250 636.600 400.350 637.500 ;
        RECT 406.950 637.200 412.650 638.100 ;
        RECT 410.850 636.600 412.650 637.200 ;
        RECT 413.550 636.600 416.550 638.400 ;
        RECT 398.550 627.600 400.350 636.600 ;
        RECT 402.450 635.550 404.250 636.300 ;
        RECT 407.250 635.550 409.050 636.300 ;
        RECT 402.450 634.500 409.050 635.550 ;
        RECT 403.350 627.000 405.150 633.600 ;
        RECT 406.350 627.600 408.150 634.500 ;
        RECT 413.550 633.600 415.650 635.700 ;
        RECT 409.350 627.000 411.150 633.600 ;
        RECT 413.850 627.600 415.650 633.600 ;
        RECT 418.650 627.000 420.450 639.600 ;
        RECT 421.650 627.600 423.450 639.600 ;
        RECT 440.100 639.600 441.300 646.950 ;
        RECT 446.100 645.150 447.900 646.950 ;
        RECT 440.100 638.100 442.500 639.600 ;
        RECT 438.000 635.100 439.800 636.900 ;
        RECT 437.700 627.000 439.500 633.600 ;
        RECT 440.700 627.600 442.500 638.100 ;
        RECT 445.800 627.000 447.600 639.600 ;
        RECT 464.100 633.600 465.300 646.950 ;
        RECT 488.100 645.150 489.900 646.950 ;
        RECT 494.100 634.800 495.000 646.950 ;
        RECT 512.100 645.150 513.900 646.950 ;
        RECT 518.700 639.600 519.900 646.950 ;
        RECT 488.400 633.900 495.000 634.800 ;
        RECT 488.400 633.600 489.900 633.900 ;
        RECT 461.100 627.000 462.900 633.600 ;
        RECT 464.100 627.600 465.900 633.600 ;
        RECT 467.100 627.000 468.900 633.600 ;
        RECT 485.100 627.000 486.900 633.600 ;
        RECT 488.100 627.600 489.900 633.600 ;
        RECT 494.100 633.600 495.000 633.900 ;
        RECT 491.100 627.000 492.900 633.000 ;
        RECT 494.100 627.600 495.900 633.600 ;
        RECT 512.400 627.000 514.200 639.600 ;
        RECT 517.500 638.100 519.900 639.600 ;
        RECT 517.500 627.600 519.300 638.100 ;
        RECT 520.200 635.100 522.000 636.900 ;
        RECT 539.100 633.600 540.000 653.700 ;
        RECT 545.400 649.050 546.300 656.400 ;
        RECT 560.100 649.050 561.900 650.850 ;
        RECT 566.250 649.050 568.050 650.850 ;
        RECT 569.700 649.050 570.600 656.400 ;
        RECT 587.100 649.050 588.900 650.850 ;
        RECT 590.100 649.050 591.300 656.400 ;
        RECT 608.700 654.600 609.900 656.400 ;
        RECT 615.900 654.900 617.100 656.400 ;
        RECT 620.100 655.500 624.900 656.400 ;
        RECT 608.700 653.700 615.000 654.600 ;
        RECT 612.900 651.600 615.000 653.700 ;
        RECT 608.400 649.050 610.200 650.850 ;
        RECT 613.200 649.800 615.000 651.600 ;
        RECT 615.900 652.800 618.900 654.900 ;
        RECT 620.100 654.300 622.200 655.500 ;
        RECT 638.700 654.300 639.900 656.400 ;
        RECT 641.100 657.300 642.900 662.400 ;
        RECT 644.100 658.200 645.900 663.000 ;
        RECT 647.100 657.300 648.900 662.400 ;
        RECT 641.100 655.950 648.900 657.300 ;
        RECT 662.100 654.600 663.900 662.400 ;
        RECT 666.600 656.400 668.400 663.000 ;
        RECT 669.600 658.200 671.400 662.400 ;
        RECT 686.100 659.400 687.900 663.000 ;
        RECT 689.100 659.400 690.900 662.400 ;
        RECT 692.100 659.400 693.900 663.000 ;
        RECT 669.600 656.400 672.300 658.200 ;
        RECT 668.700 654.600 670.500 655.500 ;
        RECT 638.700 653.400 642.300 654.300 ;
        RECT 662.100 653.700 670.500 654.600 ;
        RECT 541.500 646.950 543.600 649.050 ;
        RECT 544.800 646.950 546.900 649.050 ;
        RECT 559.950 646.950 562.050 649.050 ;
        RECT 562.950 646.950 565.050 649.050 ;
        RECT 565.950 646.950 568.050 649.050 ;
        RECT 568.950 646.950 571.050 649.050 ;
        RECT 586.950 646.950 589.050 649.050 ;
        RECT 589.950 646.950 592.050 649.050 ;
        RECT 608.100 648.300 610.200 649.050 ;
        RECT 608.100 646.950 615.000 648.300 ;
        RECT 541.200 645.150 543.000 646.950 ;
        RECT 545.400 639.600 546.300 646.950 ;
        RECT 563.250 645.150 565.050 646.950 ;
        RECT 569.700 639.600 570.600 646.950 ;
        RECT 590.100 639.600 591.300 646.950 ;
        RECT 613.200 646.500 615.000 646.950 ;
        RECT 615.900 647.100 617.100 652.800 ;
        RECT 618.000 649.800 620.100 651.900 ;
        RECT 618.300 648.000 620.100 649.800 ;
        RECT 638.100 649.050 639.900 650.850 ;
        RECT 641.100 649.050 642.300 653.400 ;
        RECT 644.100 649.050 645.900 650.850 ;
        RECT 662.250 649.050 664.050 650.850 ;
        RECT 615.900 646.200 618.300 647.100 ;
        RECT 616.800 646.050 618.300 646.200 ;
        RECT 622.800 646.950 624.900 649.050 ;
        RECT 637.950 646.950 640.050 649.050 ;
        RECT 640.950 646.950 643.050 649.050 ;
        RECT 643.950 646.950 646.050 649.050 ;
        RECT 646.950 646.950 649.050 649.050 ;
        RECT 662.100 646.950 664.200 649.050 ;
        RECT 612.000 643.500 615.900 645.300 ;
        RECT 613.800 643.200 615.900 643.500 ;
        RECT 616.800 643.950 618.900 646.050 ;
        RECT 622.800 645.150 624.600 646.950 ;
        RECT 616.800 642.000 617.700 643.950 ;
        RECT 610.500 639.600 612.600 641.700 ;
        RECT 616.200 640.950 617.700 642.000 ;
        RECT 616.200 639.600 617.400 640.950 ;
        RECT 520.500 627.000 522.300 633.600 ;
        RECT 536.100 627.000 537.900 633.600 ;
        RECT 539.100 627.600 540.900 633.600 ;
        RECT 542.100 627.000 543.900 639.000 ;
        RECT 545.100 627.600 546.900 639.600 ;
        RECT 560.100 638.700 567.900 639.600 ;
        RECT 560.100 627.600 561.900 638.700 ;
        RECT 563.100 627.000 564.900 637.800 ;
        RECT 566.100 627.600 567.900 638.700 ;
        RECT 569.100 627.600 570.900 639.600 ;
        RECT 587.100 627.000 588.900 639.600 ;
        RECT 590.100 627.600 591.900 639.600 ;
        RECT 608.100 638.700 612.600 639.600 ;
        RECT 608.100 627.600 609.900 638.700 ;
        RECT 611.100 627.000 612.900 637.500 ;
        RECT 615.600 627.600 617.400 639.600 ;
        RECT 620.100 639.600 622.200 640.500 ;
        RECT 641.100 639.600 642.300 646.950 ;
        RECT 647.100 645.150 648.900 646.950 ;
        RECT 643.950 642.450 646.050 643.050 ;
        RECT 658.950 642.450 661.050 643.050 ;
        RECT 643.950 641.550 661.050 642.450 ;
        RECT 643.950 640.950 646.050 641.550 ;
        RECT 658.950 640.950 661.050 641.550 ;
        RECT 620.100 638.400 624.900 639.600 ;
        RECT 620.100 627.000 621.900 637.500 ;
        RECT 623.100 627.600 624.900 638.400 ;
        RECT 641.100 638.100 643.500 639.600 ;
        RECT 639.000 635.100 640.800 636.900 ;
        RECT 638.700 627.000 640.500 633.600 ;
        RECT 641.700 627.600 643.500 638.100 ;
        RECT 646.800 627.000 648.600 639.600 ;
        RECT 665.100 633.600 666.000 653.700 ;
        RECT 671.400 649.050 672.300 656.400 ;
        RECT 689.700 649.050 690.600 659.400 ;
        RECT 710.700 655.200 712.500 662.400 ;
        RECT 715.800 656.400 717.600 663.000 ;
        RECT 731.700 655.200 733.500 662.400 ;
        RECT 736.800 656.400 738.600 663.000 ;
        RECT 710.700 654.300 714.900 655.200 ;
        RECT 731.700 654.300 735.900 655.200 ;
        RECT 710.100 649.050 711.900 650.850 ;
        RECT 713.700 649.050 714.900 654.300 ;
        RECT 715.950 649.050 717.750 650.850 ;
        RECT 731.100 649.050 732.900 650.850 ;
        RECT 734.700 649.050 735.900 654.300 ;
        RECT 755.100 653.400 756.900 663.000 ;
        RECT 761.700 654.000 763.500 662.400 ;
        RECT 779.700 659.400 781.500 663.000 ;
        RECT 782.700 657.600 784.500 662.400 ;
        RECT 779.400 656.400 784.500 657.600 ;
        RECT 787.200 656.400 789.000 663.000 ;
        RECT 769.950 654.450 772.050 655.050 ;
        RECT 775.950 654.450 778.050 655.050 ;
        RECT 761.700 652.800 765.000 654.000 ;
        RECT 769.950 653.550 778.050 654.450 ;
        RECT 769.950 652.950 772.050 653.550 ;
        RECT 775.950 652.950 778.050 653.550 ;
        RECT 736.950 649.050 738.750 650.850 ;
        RECT 755.100 649.050 756.900 650.850 ;
        RECT 761.100 649.050 762.900 650.850 ;
        RECT 764.100 649.050 765.000 652.800 ;
        RECT 779.400 649.050 780.300 656.400 ;
        RECT 803.100 653.400 804.900 663.000 ;
        RECT 809.700 654.000 811.500 662.400 ;
        RECT 809.700 652.800 813.000 654.000 ;
        RECT 827.100 653.400 828.900 663.000 ;
        RECT 833.700 654.000 835.500 662.400 ;
        RECT 833.700 652.800 837.000 654.000 ;
        RECT 854.100 653.400 855.900 663.000 ;
        RECT 860.700 654.000 862.500 662.400 ;
        RECT 879.000 656.400 880.800 663.000 ;
        RECT 883.500 657.600 885.300 662.400 ;
        RECT 886.500 659.400 888.300 663.000 ;
        RECT 889.950 660.450 892.050 661.050 ;
        RECT 895.950 660.450 898.050 661.050 ;
        RECT 889.950 659.550 898.050 660.450 ;
        RECT 889.950 658.950 892.050 659.550 ;
        RECT 895.950 658.950 898.050 659.550 ;
        RECT 883.500 656.400 888.600 657.600 ;
        RECT 860.700 652.800 864.000 654.000 ;
        RECT 781.950 649.050 783.750 650.850 ;
        RECT 788.100 649.050 789.900 650.850 ;
        RECT 803.100 649.050 804.900 650.850 ;
        RECT 809.100 649.050 810.900 650.850 ;
        RECT 812.100 649.050 813.000 652.800 ;
        RECT 827.100 649.050 828.900 650.850 ;
        RECT 833.100 649.050 834.900 650.850 ;
        RECT 836.100 649.050 837.000 652.800 ;
        RECT 854.100 649.050 855.900 650.850 ;
        RECT 860.100 649.050 861.900 650.850 ;
        RECT 863.100 649.050 864.000 652.800 ;
        RECT 874.950 651.450 877.050 652.050 ;
        RECT 869.550 650.550 877.050 651.450 ;
        RECT 667.500 646.950 669.600 649.050 ;
        RECT 670.800 646.950 672.900 649.050 ;
        RECT 685.950 646.950 688.050 649.050 ;
        RECT 688.950 646.950 691.050 649.050 ;
        RECT 691.950 646.950 694.050 649.050 ;
        RECT 709.950 646.950 712.050 649.050 ;
        RECT 712.950 646.950 715.050 649.050 ;
        RECT 715.950 646.950 718.050 649.050 ;
        RECT 730.950 646.950 733.050 649.050 ;
        RECT 733.950 646.950 736.050 649.050 ;
        RECT 736.950 646.950 739.050 649.050 ;
        RECT 754.950 646.950 757.050 649.050 ;
        RECT 757.950 646.950 760.050 649.050 ;
        RECT 760.950 646.950 763.050 649.050 ;
        RECT 763.950 646.950 766.050 649.050 ;
        RECT 778.950 646.950 781.050 649.050 ;
        RECT 781.950 646.950 784.050 649.050 ;
        RECT 784.950 646.950 787.050 649.050 ;
        RECT 787.950 646.950 790.050 649.050 ;
        RECT 802.950 646.950 805.050 649.050 ;
        RECT 805.950 646.950 808.050 649.050 ;
        RECT 808.950 646.950 811.050 649.050 ;
        RECT 811.950 646.950 814.050 649.050 ;
        RECT 826.950 646.950 829.050 649.050 ;
        RECT 829.950 646.950 832.050 649.050 ;
        RECT 832.950 646.950 835.050 649.050 ;
        RECT 835.950 646.950 838.050 649.050 ;
        RECT 853.950 646.950 856.050 649.050 ;
        RECT 856.950 646.950 859.050 649.050 ;
        RECT 859.950 646.950 862.050 649.050 ;
        RECT 862.950 646.950 865.050 649.050 ;
        RECT 667.200 645.150 669.000 646.950 ;
        RECT 671.400 639.600 672.300 646.950 ;
        RECT 686.100 645.150 687.900 646.950 ;
        RECT 689.700 639.600 690.600 646.950 ;
        RECT 691.950 645.150 693.750 646.950 ;
        RECT 662.100 627.000 663.900 633.600 ;
        RECT 665.100 627.600 666.900 633.600 ;
        RECT 668.100 627.000 669.900 639.000 ;
        RECT 671.100 627.600 672.900 639.600 ;
        RECT 687.000 638.400 690.600 639.600 ;
        RECT 687.000 627.600 688.800 638.400 ;
        RECT 692.100 627.000 693.900 639.600 ;
        RECT 713.700 633.600 714.900 646.950 ;
        RECT 734.700 633.600 735.900 646.950 ;
        RECT 758.100 645.150 759.900 646.950 ;
        RECT 736.950 642.450 739.050 643.050 ;
        RECT 748.950 642.450 751.050 643.050 ;
        RECT 736.950 641.550 751.050 642.450 ;
        RECT 736.950 640.950 739.050 641.550 ;
        RECT 748.950 640.950 751.050 641.550 ;
        RECT 764.100 634.800 765.000 646.950 ;
        RECT 779.400 639.600 780.300 646.950 ;
        RECT 784.950 645.150 786.750 646.950 ;
        RECT 796.950 645.450 801.000 646.050 ;
        RECT 796.950 643.950 801.450 645.450 ;
        RECT 806.100 645.150 807.900 646.950 ;
        RECT 781.950 642.450 784.050 643.050 ;
        RECT 800.550 642.450 801.450 643.950 ;
        RECT 808.950 642.450 811.050 643.050 ;
        RECT 781.950 641.550 811.050 642.450 ;
        RECT 781.950 640.950 784.050 641.550 ;
        RECT 808.950 640.950 811.050 641.550 ;
        RECT 758.400 633.900 765.000 634.800 ;
        RECT 758.400 633.600 759.900 633.900 ;
        RECT 710.100 627.000 711.900 633.600 ;
        RECT 713.100 627.600 714.900 633.600 ;
        RECT 716.100 627.000 717.900 633.600 ;
        RECT 731.100 627.000 732.900 633.600 ;
        RECT 734.100 627.600 735.900 633.600 ;
        RECT 737.100 627.000 738.900 633.600 ;
        RECT 755.100 627.000 756.900 633.600 ;
        RECT 758.100 627.600 759.900 633.600 ;
        RECT 764.100 633.600 765.000 633.900 ;
        RECT 761.100 627.000 762.900 633.000 ;
        RECT 764.100 627.600 765.900 633.600 ;
        RECT 779.100 627.600 780.900 639.600 ;
        RECT 782.100 638.700 789.900 639.600 ;
        RECT 782.100 627.600 783.900 638.700 ;
        RECT 785.100 627.000 786.900 637.800 ;
        RECT 788.100 627.600 789.900 638.700 ;
        RECT 793.950 639.450 796.050 640.050 ;
        RECT 808.950 639.450 811.050 639.900 ;
        RECT 793.950 638.550 811.050 639.450 ;
        RECT 793.950 637.950 796.050 638.550 ;
        RECT 808.950 637.800 811.050 638.550 ;
        RECT 812.100 634.800 813.000 646.950 ;
        RECT 830.100 645.150 831.900 646.950 ;
        RECT 836.100 634.800 837.000 646.950 ;
        RECT 857.100 645.150 858.900 646.950 ;
        RECT 863.100 634.800 864.000 646.950 ;
        RECT 869.550 646.050 870.450 650.550 ;
        RECT 874.950 649.950 877.050 650.550 ;
        RECT 878.100 649.050 879.900 650.850 ;
        RECT 884.250 649.050 886.050 650.850 ;
        RECT 887.700 649.050 888.600 656.400 ;
        RECT 907.500 654.000 909.300 662.400 ;
        RECT 906.000 652.800 909.300 654.000 ;
        RECT 914.100 653.400 915.900 663.000 ;
        RECT 930.000 656.400 931.800 663.000 ;
        RECT 934.500 657.600 936.300 662.400 ;
        RECT 937.500 659.400 939.300 663.000 ;
        RECT 934.500 656.400 939.600 657.600 ;
        RECT 956.100 656.400 957.900 662.400 ;
        RECT 934.950 654.450 937.050 655.050 ;
        RECT 926.550 653.550 937.050 654.450 ;
        RECT 889.950 651.450 894.000 652.050 ;
        RECT 889.950 649.950 894.450 651.450 ;
        RECT 865.950 644.550 870.450 646.050 ;
        RECT 871.950 646.050 874.050 649.050 ;
        RECT 877.950 646.950 880.050 649.050 ;
        RECT 880.950 646.950 883.050 649.050 ;
        RECT 883.950 646.950 886.050 649.050 ;
        RECT 886.950 646.950 889.050 649.050 ;
        RECT 871.950 645.000 877.050 646.050 ;
        RECT 881.250 645.150 883.050 646.950 ;
        RECT 872.550 644.550 877.050 645.000 ;
        RECT 865.950 643.950 870.000 644.550 ;
        RECT 873.000 643.950 877.050 644.550 ;
        RECT 887.700 639.600 888.600 646.950 ;
        RECT 893.550 646.050 894.450 649.950 ;
        RECT 906.000 649.050 906.900 652.800 ;
        RECT 926.550 651.450 927.450 653.550 ;
        RECT 934.950 652.950 937.050 653.550 ;
        RECT 908.100 649.050 909.900 650.850 ;
        RECT 914.100 649.050 915.900 650.850 ;
        RECT 923.550 650.550 927.450 651.450 ;
        RECT 904.950 646.950 907.050 649.050 ;
        RECT 907.950 646.950 910.050 649.050 ;
        RECT 910.950 646.950 913.050 649.050 ;
        RECT 913.950 646.950 916.050 649.050 ;
        RECT 889.950 644.550 894.450 646.050 ;
        RECT 889.950 643.950 894.000 644.550 ;
        RECT 806.400 633.900 813.000 634.800 ;
        RECT 806.400 633.600 807.900 633.900 ;
        RECT 803.100 627.000 804.900 633.600 ;
        RECT 806.100 627.600 807.900 633.600 ;
        RECT 812.100 633.600 813.000 633.900 ;
        RECT 830.400 633.900 837.000 634.800 ;
        RECT 830.400 633.600 831.900 633.900 ;
        RECT 809.100 627.000 810.900 633.000 ;
        RECT 812.100 627.600 813.900 633.600 ;
        RECT 827.100 627.000 828.900 633.600 ;
        RECT 830.100 627.600 831.900 633.600 ;
        RECT 836.100 633.600 837.000 633.900 ;
        RECT 857.400 633.900 864.000 634.800 ;
        RECT 857.400 633.600 858.900 633.900 ;
        RECT 833.100 627.000 834.900 633.000 ;
        RECT 836.100 627.600 837.900 633.600 ;
        RECT 854.100 627.000 855.900 633.600 ;
        RECT 857.100 627.600 858.900 633.600 ;
        RECT 863.100 633.600 864.000 633.900 ;
        RECT 878.100 638.700 885.900 639.600 ;
        RECT 860.100 627.000 861.900 633.000 ;
        RECT 863.100 627.600 864.900 633.600 ;
        RECT 878.100 627.600 879.900 638.700 ;
        RECT 881.100 627.000 882.900 637.800 ;
        RECT 884.100 627.600 885.900 638.700 ;
        RECT 887.100 627.600 888.900 639.600 ;
        RECT 906.000 634.800 906.900 646.950 ;
        RECT 911.100 645.150 912.900 646.950 ;
        RECT 923.550 646.050 924.450 650.550 ;
        RECT 929.100 649.050 930.900 650.850 ;
        RECT 935.250 649.050 937.050 650.850 ;
        RECT 938.700 649.050 939.600 656.400 ;
        RECT 956.700 654.300 957.900 656.400 ;
        RECT 959.100 657.300 960.900 662.400 ;
        RECT 962.100 658.200 963.900 663.000 ;
        RECT 965.100 657.300 966.900 662.400 ;
        RECT 967.950 660.450 970.050 661.050 ;
        RECT 967.950 659.550 975.450 660.450 ;
        RECT 967.950 658.950 970.050 659.550 ;
        RECT 959.100 655.950 966.900 657.300 ;
        RECT 956.700 653.400 960.300 654.300 ;
        RECT 943.950 651.450 946.050 652.050 ;
        RECT 952.950 651.450 955.050 652.050 ;
        RECT 943.950 650.550 955.050 651.450 ;
        RECT 943.950 649.950 946.050 650.550 ;
        RECT 952.950 649.950 955.050 650.550 ;
        RECT 956.100 649.050 957.900 650.850 ;
        RECT 959.100 649.050 960.300 653.400 ;
        RECT 962.100 649.050 963.900 650.850 ;
        RECT 928.950 646.950 931.050 649.050 ;
        RECT 931.950 646.950 934.050 649.050 ;
        RECT 934.950 646.950 937.050 649.050 ;
        RECT 937.950 646.950 940.050 649.050 ;
        RECT 955.950 646.950 958.050 649.050 ;
        RECT 958.950 646.950 961.050 649.050 ;
        RECT 961.950 646.950 964.050 649.050 ;
        RECT 964.950 646.950 967.050 649.050 ;
        RECT 923.550 644.550 928.050 646.050 ;
        RECT 932.250 645.150 934.050 646.950 ;
        RECT 924.000 643.950 928.050 644.550 ;
        RECT 907.950 642.450 910.050 643.050 ;
        RECT 916.950 642.450 919.050 643.050 ;
        RECT 934.950 642.450 937.050 643.050 ;
        RECT 907.950 641.550 937.050 642.450 ;
        RECT 907.950 640.950 910.050 641.550 ;
        RECT 916.950 640.950 919.050 641.550 ;
        RECT 934.950 640.950 937.050 641.550 ;
        RECT 938.700 639.600 939.600 646.950 ;
        RECT 955.950 642.450 958.050 643.050 ;
        RECT 941.550 641.550 958.050 642.450 ;
        RECT 929.100 638.700 936.900 639.600 ;
        RECT 906.000 633.900 912.600 634.800 ;
        RECT 906.000 633.600 906.900 633.900 ;
        RECT 905.100 627.600 906.900 633.600 ;
        RECT 911.100 633.600 912.600 633.900 ;
        RECT 908.100 627.000 909.900 633.000 ;
        RECT 911.100 627.600 912.900 633.600 ;
        RECT 914.100 627.000 915.900 633.600 ;
        RECT 929.100 627.600 930.900 638.700 ;
        RECT 932.100 627.000 933.900 637.800 ;
        RECT 935.100 627.600 936.900 638.700 ;
        RECT 938.100 627.600 939.900 639.600 ;
        RECT 941.550 636.450 942.450 641.550 ;
        RECT 955.950 640.950 958.050 641.550 ;
        RECT 943.950 639.450 946.050 640.050 ;
        RECT 952.950 639.450 955.050 640.050 ;
        RECT 943.950 638.550 955.050 639.450 ;
        RECT 943.950 637.950 946.050 638.550 ;
        RECT 952.950 637.950 955.050 638.550 ;
        RECT 959.100 639.600 960.300 646.950 ;
        RECT 965.100 645.150 966.900 646.950 ;
        RECT 974.550 645.450 975.450 659.550 ;
        RECT 980.100 656.400 981.900 662.400 ;
        RECT 980.700 654.300 981.900 656.400 ;
        RECT 983.100 657.300 984.900 662.400 ;
        RECT 986.100 658.200 987.900 663.000 ;
        RECT 989.100 657.300 990.900 662.400 ;
        RECT 1004.700 659.400 1006.500 663.000 ;
        RECT 1007.700 657.600 1009.500 662.400 ;
        RECT 983.100 655.950 990.900 657.300 ;
        RECT 1004.400 656.400 1009.500 657.600 ;
        RECT 1012.200 656.400 1014.000 663.000 ;
        RECT 980.700 653.400 984.300 654.300 ;
        RECT 980.100 649.050 981.900 650.850 ;
        RECT 983.100 649.050 984.300 653.400 ;
        RECT 999.000 651.450 1003.050 652.050 ;
        RECT 986.100 649.050 987.900 650.850 ;
        RECT 998.550 649.950 1003.050 651.450 ;
        RECT 979.950 646.950 982.050 649.050 ;
        RECT 982.950 646.950 985.050 649.050 ;
        RECT 985.950 646.950 988.050 649.050 ;
        RECT 988.950 646.950 991.050 649.050 ;
        RECT 974.550 644.550 978.450 645.450 ;
        RECT 977.550 643.050 978.450 644.550 ;
        RECT 977.550 642.750 981.000 643.050 ;
        RECT 977.550 641.550 982.050 642.750 ;
        RECT 978.000 640.950 982.050 641.550 ;
        RECT 979.950 640.650 982.050 640.950 ;
        RECT 983.100 639.600 984.300 646.950 ;
        RECT 989.100 645.150 990.900 646.950 ;
        RECT 998.550 643.050 999.450 649.950 ;
        RECT 1004.400 649.050 1005.300 656.400 ;
        RECT 1006.950 649.050 1008.750 650.850 ;
        RECT 1013.100 649.050 1014.900 650.850 ;
        RECT 1003.950 646.950 1006.050 649.050 ;
        RECT 1006.950 646.950 1009.050 649.050 ;
        RECT 1009.950 646.950 1012.050 649.050 ;
        RECT 1012.950 646.950 1015.050 649.050 ;
        RECT 997.950 640.950 1000.050 643.050 ;
        RECT 1004.400 639.600 1005.300 646.950 ;
        RECT 1009.950 645.150 1011.750 646.950 ;
        RECT 959.100 638.100 961.500 639.600 ;
        RECT 949.950 636.450 952.050 636.900 ;
        RECT 941.550 635.550 952.050 636.450 ;
        RECT 949.950 634.800 952.050 635.550 ;
        RECT 957.000 635.100 958.800 636.900 ;
        RECT 956.700 627.000 958.500 633.600 ;
        RECT 959.700 627.600 961.500 638.100 ;
        RECT 964.800 627.000 966.600 639.600 ;
        RECT 983.100 638.100 985.500 639.600 ;
        RECT 981.000 635.100 982.800 636.900 ;
        RECT 980.700 627.000 982.500 633.600 ;
        RECT 983.700 627.600 985.500 638.100 ;
        RECT 988.800 627.000 990.600 639.600 ;
        RECT 1004.100 627.600 1005.900 639.600 ;
        RECT 1007.100 638.700 1014.900 639.600 ;
        RECT 1007.100 627.600 1008.900 638.700 ;
        RECT 1010.100 627.000 1011.900 637.800 ;
        RECT 1013.100 627.600 1014.900 638.700 ;
        RECT 2.550 611.400 4.350 623.400 ;
        RECT 5.550 611.400 7.350 624.000 ;
        RECT 10.350 617.400 12.150 623.400 ;
        RECT 14.850 617.400 16.650 624.000 ;
        RECT 10.350 615.300 12.450 617.400 ;
        RECT 17.850 616.500 19.650 623.400 ;
        RECT 20.850 617.400 22.650 624.000 ;
        RECT 16.950 615.450 23.550 616.500 ;
        RECT 16.950 614.700 18.750 615.450 ;
        RECT 21.750 614.700 23.550 615.450 ;
        RECT 25.650 614.400 27.450 623.400 ;
        RECT 9.450 612.600 12.450 614.400 ;
        RECT 13.350 613.800 15.150 614.400 ;
        RECT 13.350 612.900 19.050 613.800 ;
        RECT 25.650 613.500 27.750 614.400 ;
        RECT 13.350 612.600 15.150 612.900 ;
        RECT 11.250 611.700 12.450 612.600 ;
        RECT 2.550 604.050 3.750 611.400 ;
        RECT 11.250 610.800 16.050 611.700 ;
        RECT 4.650 608.100 6.450 608.550 ;
        RECT 10.350 608.100 12.450 608.700 ;
        RECT 4.650 606.900 12.450 608.100 ;
        RECT 4.650 606.750 6.450 606.900 ;
        RECT 10.350 606.600 12.450 606.900 ;
        RECT 2.550 603.750 7.050 604.050 ;
        RECT 2.550 601.950 8.850 603.750 ;
        RECT 2.550 594.600 3.750 601.950 ;
        RECT 15.150 598.200 16.050 610.800 ;
        RECT 18.150 610.800 19.050 612.900 ;
        RECT 19.950 612.300 27.750 613.500 ;
        RECT 19.950 611.700 21.750 612.300 ;
        RECT 31.050 611.400 32.850 624.000 ;
        RECT 34.050 613.200 35.850 623.400 ;
        RECT 34.050 611.400 36.450 613.200 ;
        RECT 50.400 611.400 52.200 624.000 ;
        RECT 55.500 612.900 57.300 623.400 ;
        RECT 58.500 617.400 60.300 624.000 ;
        RECT 58.200 614.100 60.000 615.900 ;
        RECT 55.500 611.400 57.900 612.900 ;
        RECT 74.400 611.400 76.200 624.000 ;
        RECT 79.500 612.900 81.300 623.400 ;
        RECT 82.500 617.400 84.300 624.000 ;
        RECT 82.200 614.100 84.000 615.900 ;
        RECT 87.150 613.200 88.950 623.400 ;
        RECT 79.500 611.400 81.900 612.900 ;
        RECT 18.150 610.500 26.550 610.800 ;
        RECT 35.550 610.500 36.450 611.400 ;
        RECT 18.150 609.900 36.450 610.500 ;
        RECT 24.750 609.300 36.450 609.900 ;
        RECT 24.750 609.000 26.550 609.300 ;
        RECT 22.800 602.400 24.900 604.050 ;
        RECT 22.800 601.200 30.900 602.400 ;
        RECT 31.950 601.950 34.050 604.050 ;
        RECT 29.100 600.600 30.900 601.200 ;
        RECT 26.100 599.400 27.900 600.000 ;
        RECT 32.250 599.400 34.050 601.950 ;
        RECT 26.100 598.200 34.050 599.400 ;
        RECT 15.150 597.000 27.150 598.200 ;
        RECT 15.150 596.400 16.950 597.000 ;
        RECT 26.100 595.200 27.150 597.000 ;
        RECT 2.550 588.600 4.350 594.600 ;
        RECT 5.850 588.000 7.650 594.600 ;
        RECT 10.350 591.600 12.750 593.700 ;
        RECT 22.350 593.550 24.150 594.300 ;
        RECT 19.200 592.500 24.150 593.550 ;
        RECT 25.350 593.400 27.150 595.200 ;
        RECT 35.550 594.600 36.450 609.300 ;
        RECT 50.100 604.050 51.900 605.850 ;
        RECT 56.700 604.050 57.900 611.400 ;
        RECT 74.100 604.050 75.900 605.850 ;
        RECT 80.700 604.050 81.900 611.400 ;
        RECT 86.550 611.400 88.950 613.200 ;
        RECT 90.150 611.400 91.950 624.000 ;
        RECT 95.550 614.400 97.350 623.400 ;
        RECT 100.350 617.400 102.150 624.000 ;
        RECT 103.350 616.500 105.150 623.400 ;
        RECT 106.350 617.400 108.150 624.000 ;
        RECT 110.850 617.400 112.650 623.400 ;
        RECT 99.450 615.450 106.050 616.500 ;
        RECT 99.450 614.700 101.250 615.450 ;
        RECT 104.250 614.700 106.050 615.450 ;
        RECT 110.550 615.300 112.650 617.400 ;
        RECT 95.250 613.500 97.350 614.400 ;
        RECT 107.850 613.800 109.650 614.400 ;
        RECT 95.250 612.300 103.050 613.500 ;
        RECT 101.250 611.700 103.050 612.300 ;
        RECT 103.950 612.900 109.650 613.800 ;
        RECT 86.550 610.500 87.450 611.400 ;
        RECT 103.950 610.800 104.850 612.900 ;
        RECT 107.850 612.600 109.650 612.900 ;
        RECT 110.550 612.600 113.550 614.400 ;
        RECT 110.550 611.700 111.750 612.600 ;
        RECT 96.450 610.500 104.850 610.800 ;
        RECT 86.550 609.900 104.850 610.500 ;
        RECT 106.950 610.800 111.750 611.700 ;
        RECT 115.650 611.400 117.450 624.000 ;
        RECT 118.650 611.400 120.450 623.400 ;
        RECT 137.100 617.400 138.900 624.000 ;
        RECT 140.100 617.400 141.900 623.400 ;
        RECT 143.100 617.400 144.900 624.000 ;
        RECT 86.550 609.300 98.250 609.900 ;
        RECT 49.950 601.950 52.050 604.050 ;
        RECT 52.950 601.950 55.050 604.050 ;
        RECT 55.950 601.950 58.050 604.050 ;
        RECT 58.950 601.950 61.050 604.050 ;
        RECT 73.950 601.950 76.050 604.050 ;
        RECT 76.950 601.950 79.050 604.050 ;
        RECT 79.950 601.950 82.050 604.050 ;
        RECT 82.950 601.950 85.050 604.050 ;
        RECT 53.100 600.150 54.900 601.950 ;
        RECT 56.700 597.600 57.900 601.950 ;
        RECT 59.100 600.150 60.900 601.950 ;
        RECT 77.100 600.150 78.900 601.950 ;
        RECT 80.700 597.600 81.900 601.950 ;
        RECT 83.100 600.150 84.900 601.950 ;
        RECT 56.700 596.700 60.300 597.600 ;
        RECT 80.700 596.700 84.300 597.600 ;
        RECT 19.200 591.600 20.250 592.500 ;
        RECT 28.050 592.200 30.150 593.700 ;
        RECT 26.250 591.600 30.150 592.200 ;
        RECT 10.950 588.600 12.750 591.600 ;
        RECT 15.450 588.000 17.250 591.600 ;
        RECT 18.450 588.600 20.250 591.600 ;
        RECT 21.750 588.000 23.550 591.600 ;
        RECT 26.250 590.700 29.850 591.600 ;
        RECT 26.250 588.600 28.050 590.700 ;
        RECT 31.050 588.000 32.850 594.600 ;
        RECT 34.050 592.800 36.450 594.600 ;
        RECT 50.100 593.700 57.900 595.050 ;
        RECT 34.050 588.600 35.850 592.800 ;
        RECT 50.100 588.600 51.900 593.700 ;
        RECT 53.100 588.000 54.900 592.800 ;
        RECT 56.100 588.600 57.900 593.700 ;
        RECT 59.100 594.600 60.300 596.700 ;
        RECT 59.100 588.600 60.900 594.600 ;
        RECT 74.100 593.700 81.900 595.050 ;
        RECT 74.100 588.600 75.900 593.700 ;
        RECT 77.100 588.000 78.900 592.800 ;
        RECT 80.100 588.600 81.900 593.700 ;
        RECT 83.100 594.600 84.300 596.700 ;
        RECT 86.550 594.600 87.450 609.300 ;
        RECT 96.450 609.000 98.250 609.300 ;
        RECT 88.950 601.950 91.050 604.050 ;
        RECT 98.100 602.400 100.200 604.050 ;
        RECT 88.950 599.400 90.750 601.950 ;
        RECT 92.100 601.200 100.200 602.400 ;
        RECT 92.100 600.600 93.900 601.200 ;
        RECT 95.100 599.400 96.900 600.000 ;
        RECT 88.950 598.200 96.900 599.400 ;
        RECT 106.950 598.200 107.850 610.800 ;
        RECT 110.550 608.100 112.650 608.700 ;
        RECT 116.550 608.100 118.350 608.550 ;
        RECT 110.550 606.900 118.350 608.100 ;
        RECT 110.550 606.600 112.650 606.900 ;
        RECT 116.550 606.750 118.350 606.900 ;
        RECT 119.250 604.050 120.450 611.400 ;
        RECT 140.100 604.050 141.300 617.400 ;
        RECT 161.100 611.400 162.900 624.000 ;
        RECT 164.100 610.500 165.900 623.400 ;
        RECT 167.100 611.400 168.900 624.000 ;
        RECT 170.100 610.500 171.900 623.400 ;
        RECT 173.100 611.400 174.900 624.000 ;
        RECT 176.100 610.500 177.900 623.400 ;
        RECT 179.100 611.400 180.900 624.000 ;
        RECT 182.100 610.500 183.900 623.400 ;
        RECT 185.100 611.400 186.900 624.000 ;
        RECT 189.150 613.200 190.950 623.400 ;
        RECT 188.550 611.400 190.950 613.200 ;
        RECT 192.150 611.400 193.950 624.000 ;
        RECT 197.550 614.400 199.350 623.400 ;
        RECT 202.350 617.400 204.150 624.000 ;
        RECT 205.350 616.500 207.150 623.400 ;
        RECT 208.350 617.400 210.150 624.000 ;
        RECT 212.850 617.400 214.650 623.400 ;
        RECT 201.450 615.450 208.050 616.500 ;
        RECT 201.450 614.700 203.250 615.450 ;
        RECT 206.250 614.700 208.050 615.450 ;
        RECT 212.550 615.300 214.650 617.400 ;
        RECT 197.250 613.500 199.350 614.400 ;
        RECT 209.850 613.800 211.650 614.400 ;
        RECT 197.250 612.300 205.050 613.500 ;
        RECT 203.250 611.700 205.050 612.300 ;
        RECT 205.950 612.900 211.650 613.800 ;
        RECT 163.050 609.300 165.900 610.500 ;
        RECT 168.000 609.300 171.900 610.500 ;
        RECT 174.000 609.300 177.900 610.500 ;
        RECT 180.000 609.300 183.900 610.500 ;
        RECT 188.550 610.500 189.450 611.400 ;
        RECT 205.950 610.800 206.850 612.900 ;
        RECT 209.850 612.600 211.650 612.900 ;
        RECT 212.550 612.600 215.550 614.400 ;
        RECT 212.550 611.700 213.750 612.600 ;
        RECT 198.450 610.500 206.850 610.800 ;
        RECT 188.550 609.900 206.850 610.500 ;
        RECT 208.950 610.800 213.750 611.700 ;
        RECT 217.650 611.400 219.450 624.000 ;
        RECT 220.650 611.400 222.450 623.400 ;
        RECT 236.100 617.400 237.900 624.000 ;
        RECT 239.100 617.400 240.900 623.400 ;
        RECT 188.550 609.300 200.250 609.900 ;
        RECT 163.050 604.050 164.100 609.300 ;
        RECT 115.950 603.750 120.450 604.050 ;
        RECT 114.150 601.950 120.450 603.750 ;
        RECT 136.950 601.950 139.050 604.050 ;
        RECT 139.950 601.950 142.050 604.050 ;
        RECT 142.950 601.950 145.050 604.050 ;
        RECT 163.050 601.950 166.200 604.050 ;
        RECT 95.850 597.000 107.850 598.200 ;
        RECT 95.850 595.200 96.900 597.000 ;
        RECT 106.050 596.400 107.850 597.000 ;
        RECT 83.100 588.600 84.900 594.600 ;
        RECT 86.550 592.800 88.950 594.600 ;
        RECT 87.150 588.600 88.950 592.800 ;
        RECT 90.150 588.000 91.950 594.600 ;
        RECT 92.850 592.200 94.950 593.700 ;
        RECT 95.850 593.400 97.650 595.200 ;
        RECT 119.250 594.600 120.450 601.950 ;
        RECT 137.250 600.150 139.050 601.950 ;
        RECT 140.100 596.700 141.300 601.950 ;
        RECT 143.100 600.150 144.900 601.950 ;
        RECT 163.050 596.700 164.100 601.950 ;
        RECT 165.000 598.800 166.800 599.400 ;
        RECT 168.000 598.800 169.200 609.300 ;
        RECT 165.000 597.600 169.200 598.800 ;
        RECT 171.000 598.800 172.800 599.400 ;
        RECT 174.000 598.800 175.200 609.300 ;
        RECT 171.000 597.600 175.200 598.800 ;
        RECT 177.000 598.800 178.800 599.400 ;
        RECT 180.000 598.800 181.200 609.300 ;
        RECT 182.100 601.950 184.200 604.050 ;
        RECT 182.400 600.150 184.200 601.950 ;
        RECT 177.000 597.600 181.200 598.800 ;
        RECT 168.000 596.700 169.200 597.600 ;
        RECT 174.000 596.700 175.200 597.600 ;
        RECT 180.000 596.700 181.200 597.600 ;
        RECT 140.100 595.800 144.300 596.700 ;
        RECT 98.850 593.550 100.650 594.300 ;
        RECT 98.850 592.500 103.800 593.550 ;
        RECT 92.850 591.600 96.750 592.200 ;
        RECT 102.750 591.600 103.800 592.500 ;
        RECT 110.250 591.600 112.650 593.700 ;
        RECT 93.150 590.700 96.750 591.600 ;
        RECT 94.950 588.600 96.750 590.700 ;
        RECT 99.450 588.000 101.250 591.600 ;
        RECT 102.750 588.600 104.550 591.600 ;
        RECT 105.750 588.000 107.550 591.600 ;
        RECT 110.250 588.600 112.050 591.600 ;
        RECT 115.350 588.000 117.150 594.600 ;
        RECT 118.650 588.600 120.450 594.600 ;
        RECT 137.400 588.000 139.200 594.600 ;
        RECT 142.500 588.600 144.300 595.800 ;
        RECT 163.050 595.500 165.900 596.700 ;
        RECT 168.000 595.500 171.900 596.700 ;
        RECT 174.000 595.500 177.900 596.700 ;
        RECT 180.000 595.500 183.900 596.700 ;
        RECT 161.100 588.000 162.900 594.600 ;
        RECT 164.100 588.600 165.900 595.500 ;
        RECT 167.100 588.000 168.900 594.600 ;
        RECT 170.100 588.600 171.900 595.500 ;
        RECT 173.100 588.000 174.900 594.600 ;
        RECT 176.100 588.600 177.900 595.500 ;
        RECT 179.100 588.000 180.900 594.600 ;
        RECT 182.100 588.600 183.900 595.500 ;
        RECT 188.550 594.600 189.450 609.300 ;
        RECT 198.450 609.000 200.250 609.300 ;
        RECT 190.950 601.950 193.050 604.050 ;
        RECT 200.100 602.400 202.200 604.050 ;
        RECT 190.950 599.400 192.750 601.950 ;
        RECT 194.100 601.200 202.200 602.400 ;
        RECT 194.100 600.600 195.900 601.200 ;
        RECT 197.100 599.400 198.900 600.000 ;
        RECT 190.950 598.200 198.900 599.400 ;
        RECT 208.950 598.200 209.850 610.800 ;
        RECT 212.550 608.100 214.650 608.700 ;
        RECT 218.550 608.100 220.350 608.550 ;
        RECT 212.550 606.900 220.350 608.100 ;
        RECT 212.550 606.600 214.650 606.900 ;
        RECT 218.550 606.750 220.350 606.900 ;
        RECT 221.250 604.050 222.450 611.400 ;
        RECT 236.100 604.050 237.900 605.850 ;
        RECT 239.100 604.050 240.300 617.400 ;
        RECT 254.100 612.600 255.900 623.400 ;
        RECT 257.100 613.500 258.900 624.000 ;
        RECT 260.100 622.500 267.900 623.400 ;
        RECT 260.100 612.600 261.900 622.500 ;
        RECT 254.100 611.700 261.900 612.600 ;
        RECT 263.100 610.500 264.900 621.600 ;
        RECT 266.100 611.400 267.900 622.500 ;
        RECT 281.100 611.400 282.900 623.400 ;
        RECT 284.100 612.000 285.900 624.000 ;
        RECT 287.100 617.400 288.900 623.400 ;
        RECT 290.100 617.400 291.900 624.000 ;
        RECT 260.100 609.600 264.900 610.500 ;
        RECT 257.250 604.050 259.050 605.850 ;
        RECT 260.100 604.050 261.000 609.600 ;
        RECT 263.100 604.050 264.900 605.850 ;
        RECT 281.700 604.050 282.600 611.400 ;
        RECT 285.000 604.050 286.800 605.850 ;
        RECT 217.950 603.750 222.450 604.050 ;
        RECT 216.150 601.950 222.450 603.750 ;
        RECT 235.950 601.950 238.050 604.050 ;
        RECT 238.950 601.950 241.050 604.050 ;
        RECT 253.950 601.950 256.050 604.050 ;
        RECT 256.950 601.950 259.050 604.050 ;
        RECT 259.950 601.950 262.050 604.050 ;
        RECT 262.950 601.950 265.050 604.050 ;
        RECT 265.950 601.950 268.050 604.050 ;
        RECT 281.100 601.950 283.200 604.050 ;
        RECT 284.400 601.950 286.500 604.050 ;
        RECT 197.850 597.000 209.850 598.200 ;
        RECT 197.850 595.200 198.900 597.000 ;
        RECT 208.050 596.400 209.850 597.000 ;
        RECT 185.100 588.000 186.900 594.600 ;
        RECT 188.550 592.800 190.950 594.600 ;
        RECT 189.150 588.600 190.950 592.800 ;
        RECT 192.150 588.000 193.950 594.600 ;
        RECT 194.850 592.200 196.950 593.700 ;
        RECT 197.850 593.400 199.650 595.200 ;
        RECT 221.250 594.600 222.450 601.950 ;
        RECT 200.850 593.550 202.650 594.300 ;
        RECT 200.850 592.500 205.800 593.550 ;
        RECT 194.850 591.600 198.750 592.200 ;
        RECT 204.750 591.600 205.800 592.500 ;
        RECT 212.250 591.600 214.650 593.700 ;
        RECT 195.150 590.700 198.750 591.600 ;
        RECT 196.950 588.600 198.750 590.700 ;
        RECT 201.450 588.000 203.250 591.600 ;
        RECT 204.750 588.600 206.550 591.600 ;
        RECT 207.750 588.000 209.550 591.600 ;
        RECT 212.250 588.600 214.050 591.600 ;
        RECT 217.350 588.000 219.150 594.600 ;
        RECT 220.650 588.600 222.450 594.600 ;
        RECT 239.100 591.600 240.300 601.950 ;
        RECT 254.250 600.150 256.050 601.950 ;
        RECT 260.100 594.600 261.300 601.950 ;
        RECT 266.100 600.150 267.900 601.950 ;
        RECT 281.700 594.600 282.600 601.950 ;
        RECT 288.000 597.300 288.900 617.400 ;
        RECT 293.550 611.400 295.350 623.400 ;
        RECT 296.550 611.400 298.350 624.000 ;
        RECT 301.350 617.400 303.150 623.400 ;
        RECT 305.850 617.400 307.650 624.000 ;
        RECT 301.350 615.300 303.450 617.400 ;
        RECT 308.850 616.500 310.650 623.400 ;
        RECT 311.850 617.400 313.650 624.000 ;
        RECT 307.950 615.450 314.550 616.500 ;
        RECT 307.950 614.700 309.750 615.450 ;
        RECT 312.750 614.700 314.550 615.450 ;
        RECT 316.650 614.400 318.450 623.400 ;
        RECT 300.450 612.600 303.450 614.400 ;
        RECT 304.350 613.800 306.150 614.400 ;
        RECT 304.350 612.900 310.050 613.800 ;
        RECT 316.650 613.500 318.750 614.400 ;
        RECT 304.350 612.600 306.150 612.900 ;
        RECT 302.250 611.700 303.450 612.600 ;
        RECT 293.550 604.050 294.750 611.400 ;
        RECT 302.250 610.800 307.050 611.700 ;
        RECT 295.650 608.100 297.450 608.550 ;
        RECT 301.350 608.100 303.450 608.700 ;
        RECT 295.650 606.900 303.450 608.100 ;
        RECT 295.650 606.750 297.450 606.900 ;
        RECT 301.350 606.600 303.450 606.900 ;
        RECT 289.800 601.950 291.900 604.050 ;
        RECT 293.550 603.750 298.050 604.050 ;
        RECT 293.550 601.950 299.850 603.750 ;
        RECT 289.950 600.150 291.750 601.950 ;
        RECT 283.500 596.400 291.900 597.300 ;
        RECT 283.500 595.500 285.300 596.400 ;
        RECT 236.100 588.000 237.900 591.600 ;
        RECT 239.100 588.600 240.900 591.600 ;
        RECT 254.700 588.000 256.500 594.600 ;
        RECT 259.200 588.600 261.000 594.600 ;
        RECT 263.700 588.000 265.500 594.600 ;
        RECT 281.700 592.800 284.400 594.600 ;
        RECT 282.600 588.600 284.400 592.800 ;
        RECT 285.600 588.000 287.400 594.600 ;
        RECT 290.100 588.600 291.900 596.400 ;
        RECT 293.550 594.600 294.750 601.950 ;
        RECT 306.150 598.200 307.050 610.800 ;
        RECT 309.150 610.800 310.050 612.900 ;
        RECT 310.950 612.300 318.750 613.500 ;
        RECT 310.950 611.700 312.750 612.300 ;
        RECT 322.050 611.400 323.850 624.000 ;
        RECT 325.050 613.200 326.850 623.400 ;
        RECT 341.100 617.400 342.900 624.000 ;
        RECT 344.100 617.400 345.900 623.400 ;
        RECT 325.050 611.400 327.450 613.200 ;
        RECT 309.150 610.500 317.550 610.800 ;
        RECT 326.550 610.500 327.450 611.400 ;
        RECT 309.150 609.900 327.450 610.500 ;
        RECT 315.750 609.300 327.450 609.900 ;
        RECT 315.750 609.000 317.550 609.300 ;
        RECT 313.800 602.400 315.900 604.050 ;
        RECT 313.800 601.200 321.900 602.400 ;
        RECT 322.950 601.950 325.050 604.050 ;
        RECT 320.100 600.600 321.900 601.200 ;
        RECT 317.100 599.400 318.900 600.000 ;
        RECT 323.250 599.400 325.050 601.950 ;
        RECT 317.100 598.200 325.050 599.400 ;
        RECT 306.150 597.000 318.150 598.200 ;
        RECT 306.150 596.400 307.950 597.000 ;
        RECT 317.100 595.200 318.150 597.000 ;
        RECT 293.550 588.600 295.350 594.600 ;
        RECT 296.850 588.000 298.650 594.600 ;
        RECT 301.350 591.600 303.750 593.700 ;
        RECT 313.350 593.550 315.150 594.300 ;
        RECT 310.200 592.500 315.150 593.550 ;
        RECT 316.350 593.400 318.150 595.200 ;
        RECT 326.550 594.600 327.450 609.300 ;
        RECT 341.100 604.050 342.900 605.850 ;
        RECT 344.100 604.050 345.300 617.400 ;
        RECT 347.550 611.400 349.350 623.400 ;
        RECT 350.550 611.400 352.350 624.000 ;
        RECT 355.350 617.400 357.150 623.400 ;
        RECT 359.850 617.400 361.650 624.000 ;
        RECT 355.350 615.300 357.450 617.400 ;
        RECT 362.850 616.500 364.650 623.400 ;
        RECT 365.850 617.400 367.650 624.000 ;
        RECT 361.950 615.450 368.550 616.500 ;
        RECT 361.950 614.700 363.750 615.450 ;
        RECT 366.750 614.700 368.550 615.450 ;
        RECT 370.650 614.400 372.450 623.400 ;
        RECT 354.450 612.600 357.450 614.400 ;
        RECT 358.350 613.800 360.150 614.400 ;
        RECT 358.350 612.900 364.050 613.800 ;
        RECT 370.650 613.500 372.750 614.400 ;
        RECT 358.350 612.600 360.150 612.900 ;
        RECT 356.250 611.700 357.450 612.600 ;
        RECT 347.550 604.050 348.750 611.400 ;
        RECT 356.250 610.800 361.050 611.700 ;
        RECT 349.650 608.100 351.450 608.550 ;
        RECT 355.350 608.100 357.450 608.700 ;
        RECT 349.650 606.900 357.450 608.100 ;
        RECT 349.650 606.750 351.450 606.900 ;
        RECT 355.350 606.600 357.450 606.900 ;
        RECT 340.950 601.950 343.050 604.050 ;
        RECT 343.950 601.950 346.050 604.050 ;
        RECT 347.550 603.750 352.050 604.050 ;
        RECT 347.550 601.950 353.850 603.750 ;
        RECT 310.200 591.600 311.250 592.500 ;
        RECT 319.050 592.200 321.150 593.700 ;
        RECT 317.250 591.600 321.150 592.200 ;
        RECT 301.950 588.600 303.750 591.600 ;
        RECT 306.450 588.000 308.250 591.600 ;
        RECT 309.450 588.600 311.250 591.600 ;
        RECT 312.750 588.000 314.550 591.600 ;
        RECT 317.250 590.700 320.850 591.600 ;
        RECT 317.250 588.600 319.050 590.700 ;
        RECT 322.050 588.000 323.850 594.600 ;
        RECT 325.050 592.800 327.450 594.600 ;
        RECT 325.050 588.600 326.850 592.800 ;
        RECT 344.100 591.600 345.300 601.950 ;
        RECT 347.550 594.600 348.750 601.950 ;
        RECT 360.150 598.200 361.050 610.800 ;
        RECT 363.150 610.800 364.050 612.900 ;
        RECT 364.950 612.300 372.750 613.500 ;
        RECT 364.950 611.700 366.750 612.300 ;
        RECT 376.050 611.400 377.850 624.000 ;
        RECT 379.050 613.200 380.850 623.400 ;
        RECT 379.050 611.400 381.450 613.200 ;
        RECT 398.400 611.400 400.200 624.000 ;
        RECT 403.500 612.900 405.300 623.400 ;
        RECT 406.500 617.400 408.300 624.000 ;
        RECT 406.200 614.100 408.000 615.900 ;
        RECT 403.500 611.400 405.900 612.900 ;
        RECT 422.400 611.400 424.200 624.000 ;
        RECT 427.500 612.900 429.300 623.400 ;
        RECT 430.500 617.400 432.300 624.000 ;
        RECT 449.100 617.400 450.900 624.000 ;
        RECT 452.100 617.400 453.900 623.400 ;
        RECT 455.100 617.400 456.900 624.000 ;
        RECT 473.100 617.400 474.900 624.000 ;
        RECT 476.100 617.400 477.900 623.400 ;
        RECT 479.100 617.400 480.900 624.000 ;
        RECT 430.200 614.100 432.000 615.900 ;
        RECT 427.500 611.400 429.900 612.900 ;
        RECT 363.150 610.500 371.550 610.800 ;
        RECT 380.550 610.500 381.450 611.400 ;
        RECT 363.150 609.900 381.450 610.500 ;
        RECT 369.750 609.300 381.450 609.900 ;
        RECT 369.750 609.000 371.550 609.300 ;
        RECT 367.800 602.400 369.900 604.050 ;
        RECT 367.800 601.200 375.900 602.400 ;
        RECT 376.950 601.950 379.050 604.050 ;
        RECT 374.100 600.600 375.900 601.200 ;
        RECT 371.100 599.400 372.900 600.000 ;
        RECT 377.250 599.400 379.050 601.950 ;
        RECT 371.100 598.200 379.050 599.400 ;
        RECT 360.150 597.000 372.150 598.200 ;
        RECT 360.150 596.400 361.950 597.000 ;
        RECT 371.100 595.200 372.150 597.000 ;
        RECT 341.100 588.000 342.900 591.600 ;
        RECT 344.100 588.600 345.900 591.600 ;
        RECT 347.550 588.600 349.350 594.600 ;
        RECT 350.850 588.000 352.650 594.600 ;
        RECT 355.350 591.600 357.750 593.700 ;
        RECT 367.350 593.550 369.150 594.300 ;
        RECT 364.200 592.500 369.150 593.550 ;
        RECT 370.350 593.400 372.150 595.200 ;
        RECT 380.550 594.600 381.450 609.300 ;
        RECT 398.100 604.050 399.900 605.850 ;
        RECT 404.700 604.050 405.900 611.400 ;
        RECT 422.100 604.050 423.900 605.850 ;
        RECT 428.700 604.050 429.900 611.400 ;
        RECT 452.100 604.050 453.300 617.400 ;
        RECT 476.700 604.050 477.900 617.400 ;
        RECT 497.100 611.400 498.900 623.400 ;
        RECT 500.100 613.200 501.900 624.000 ;
        RECT 503.100 617.400 504.900 623.400 ;
        RECT 497.100 604.050 498.300 611.400 ;
        RECT 503.700 610.500 504.900 617.400 ;
        RECT 499.200 609.600 504.900 610.500 ;
        RECT 521.100 617.400 522.900 623.400 ;
        RECT 521.100 610.500 522.300 617.400 ;
        RECT 524.100 613.200 525.900 624.000 ;
        RECT 527.100 611.400 528.900 623.400 ;
        RECT 542.400 611.400 544.200 624.000 ;
        RECT 547.500 612.900 549.300 623.400 ;
        RECT 550.500 617.400 552.300 624.000 ;
        RECT 569.100 617.400 570.900 624.000 ;
        RECT 572.100 617.400 573.900 623.400 ;
        RECT 575.100 617.400 576.900 624.000 ;
        RECT 590.100 617.400 591.900 624.000 ;
        RECT 593.100 617.400 594.900 623.400 ;
        RECT 596.100 617.400 597.900 624.000 ;
        RECT 550.200 614.100 552.000 615.900 ;
        RECT 547.500 611.400 549.900 612.900 ;
        RECT 521.100 609.600 526.800 610.500 ;
        RECT 499.200 608.700 501.000 609.600 ;
        RECT 397.950 601.950 400.050 604.050 ;
        RECT 400.950 601.950 403.050 604.050 ;
        RECT 403.950 601.950 406.050 604.050 ;
        RECT 406.950 601.950 409.050 604.050 ;
        RECT 421.950 601.950 424.050 604.050 ;
        RECT 424.950 601.950 427.050 604.050 ;
        RECT 427.950 601.950 430.050 604.050 ;
        RECT 430.950 601.950 433.050 604.050 ;
        RECT 448.950 601.950 451.050 604.050 ;
        RECT 451.950 601.950 454.050 604.050 ;
        RECT 454.950 601.950 457.050 604.050 ;
        RECT 472.950 601.950 475.050 604.050 ;
        RECT 475.950 601.950 478.050 604.050 ;
        RECT 478.950 601.950 481.050 604.050 ;
        RECT 497.100 601.950 499.200 604.050 ;
        RECT 401.100 600.150 402.900 601.950 ;
        RECT 404.700 597.600 405.900 601.950 ;
        RECT 407.100 600.150 408.900 601.950 ;
        RECT 425.100 600.150 426.900 601.950 ;
        RECT 428.700 597.600 429.900 601.950 ;
        RECT 431.100 600.150 432.900 601.950 ;
        RECT 449.250 600.150 451.050 601.950 ;
        RECT 404.700 596.700 408.300 597.600 ;
        RECT 428.700 596.700 432.300 597.600 ;
        RECT 364.200 591.600 365.250 592.500 ;
        RECT 373.050 592.200 375.150 593.700 ;
        RECT 371.250 591.600 375.150 592.200 ;
        RECT 355.950 588.600 357.750 591.600 ;
        RECT 360.450 588.000 362.250 591.600 ;
        RECT 363.450 588.600 365.250 591.600 ;
        RECT 366.750 588.000 368.550 591.600 ;
        RECT 371.250 590.700 374.850 591.600 ;
        RECT 371.250 588.600 373.050 590.700 ;
        RECT 376.050 588.000 377.850 594.600 ;
        RECT 379.050 592.800 381.450 594.600 ;
        RECT 398.100 593.700 405.900 595.050 ;
        RECT 379.050 588.600 380.850 592.800 ;
        RECT 398.100 588.600 399.900 593.700 ;
        RECT 401.100 588.000 402.900 592.800 ;
        RECT 404.100 588.600 405.900 593.700 ;
        RECT 407.100 594.600 408.300 596.700 ;
        RECT 407.100 588.600 408.900 594.600 ;
        RECT 422.100 593.700 429.900 595.050 ;
        RECT 422.100 588.600 423.900 593.700 ;
        RECT 425.100 588.000 426.900 592.800 ;
        RECT 428.100 588.600 429.900 593.700 ;
        RECT 431.100 594.600 432.300 596.700 ;
        RECT 452.100 596.700 453.300 601.950 ;
        RECT 455.100 600.150 456.900 601.950 ;
        RECT 473.100 600.150 474.900 601.950 ;
        RECT 476.700 596.700 477.900 601.950 ;
        RECT 478.950 600.150 480.750 601.950 ;
        RECT 452.100 595.800 456.300 596.700 ;
        RECT 431.100 588.600 432.900 594.600 ;
        RECT 449.400 588.000 451.200 594.600 ;
        RECT 454.500 588.600 456.300 595.800 ;
        RECT 473.700 595.800 477.900 596.700 ;
        RECT 473.700 588.600 475.500 595.800 ;
        RECT 497.100 594.600 498.300 601.950 ;
        RECT 500.100 597.300 501.000 608.700 ;
        RECT 525.000 608.700 526.800 609.600 ;
        RECT 502.800 604.050 504.600 605.850 ;
        RECT 502.500 601.950 504.600 604.050 ;
        RECT 521.400 604.050 523.200 605.850 ;
        RECT 521.400 601.950 523.500 604.050 ;
        RECT 499.200 596.400 501.000 597.300 ;
        RECT 525.000 597.300 525.900 608.700 ;
        RECT 527.700 604.050 528.900 611.400 ;
        RECT 542.100 604.050 543.900 605.850 ;
        RECT 548.700 604.050 549.900 611.400 ;
        RECT 550.950 612.450 553.050 613.050 ;
        RECT 568.950 612.450 571.050 613.050 ;
        RECT 550.950 611.550 571.050 612.450 ;
        RECT 550.950 610.950 553.050 611.550 ;
        RECT 568.950 610.950 571.050 611.550 ;
        RECT 550.950 609.450 553.050 609.900 ;
        RECT 556.950 609.450 559.050 609.900 ;
        RECT 550.950 608.550 559.050 609.450 ;
        RECT 550.950 607.800 553.050 608.550 ;
        RECT 556.950 607.800 559.050 608.550 ;
        RECT 572.700 604.050 573.900 617.400 ;
        RECT 574.950 615.450 577.050 616.050 ;
        RECT 586.950 615.450 589.050 616.050 ;
        RECT 574.950 614.550 589.050 615.450 ;
        RECT 574.950 613.950 577.050 614.550 ;
        RECT 586.950 613.950 589.050 614.550 ;
        RECT 585.000 606.450 589.050 607.050 ;
        RECT 584.550 604.950 589.050 606.450 ;
        RECT 526.800 601.950 528.900 604.050 ;
        RECT 541.950 601.950 544.050 604.050 ;
        RECT 544.950 601.950 547.050 604.050 ;
        RECT 547.950 601.950 550.050 604.050 ;
        RECT 550.950 601.950 553.050 604.050 ;
        RECT 568.950 601.950 571.050 604.050 ;
        RECT 571.950 601.950 574.050 604.050 ;
        RECT 574.950 601.950 577.050 604.050 ;
        RECT 525.000 596.400 526.800 597.300 ;
        RECT 499.200 595.500 504.900 596.400 ;
        RECT 478.800 588.000 480.600 594.600 ;
        RECT 497.100 588.600 498.900 594.600 ;
        RECT 500.100 588.000 501.900 594.600 ;
        RECT 503.700 591.600 504.900 595.500 ;
        RECT 503.100 588.600 504.900 591.600 ;
        RECT 521.100 595.500 526.800 596.400 ;
        RECT 521.100 591.600 522.300 595.500 ;
        RECT 527.700 594.600 528.900 601.950 ;
        RECT 545.100 600.150 546.900 601.950 ;
        RECT 548.700 597.600 549.900 601.950 ;
        RECT 551.100 600.150 552.900 601.950 ;
        RECT 569.100 600.150 570.900 601.950 ;
        RECT 548.700 596.700 552.300 597.600 ;
        RECT 572.700 596.700 573.900 601.950 ;
        RECT 574.950 600.150 576.750 601.950 ;
        RECT 584.550 597.900 585.450 604.950 ;
        RECT 593.100 604.050 594.300 617.400 ;
        RECT 611.400 611.400 613.200 624.000 ;
        RECT 616.500 612.900 618.300 623.400 ;
        RECT 619.500 617.400 621.300 624.000 ;
        RECT 635.100 617.400 636.900 624.000 ;
        RECT 638.100 617.400 639.900 623.400 ;
        RECT 641.100 617.400 642.900 624.000 ;
        RECT 656.100 617.400 657.900 624.000 ;
        RECT 659.100 617.400 660.900 623.400 ;
        RECT 662.100 618.000 663.900 624.000 ;
        RECT 619.200 614.100 621.000 615.900 ;
        RECT 616.500 611.400 618.900 612.900 ;
        RECT 611.100 604.050 612.900 605.850 ;
        RECT 617.700 604.050 618.900 611.400 ;
        RECT 633.000 609.450 637.050 610.050 ;
        RECT 632.550 607.950 637.050 609.450 ;
        RECT 632.550 606.450 633.450 607.950 ;
        RECT 629.550 605.550 633.450 606.450 ;
        RECT 589.950 601.950 592.050 604.050 ;
        RECT 592.950 601.950 595.050 604.050 ;
        RECT 595.950 601.950 598.050 604.050 ;
        RECT 610.950 601.950 613.050 604.050 ;
        RECT 613.950 601.950 616.050 604.050 ;
        RECT 616.950 601.950 619.050 604.050 ;
        RECT 619.950 601.950 622.050 604.050 ;
        RECT 590.250 600.150 592.050 601.950 ;
        RECT 521.100 588.600 522.900 591.600 ;
        RECT 524.100 588.000 525.900 594.600 ;
        RECT 527.100 588.600 528.900 594.600 ;
        RECT 529.950 594.450 532.050 595.050 ;
        RECT 535.950 594.450 538.050 595.050 ;
        RECT 529.950 593.550 538.050 594.450 ;
        RECT 529.950 592.950 532.050 593.550 ;
        RECT 535.950 592.950 538.050 593.550 ;
        RECT 542.100 593.700 549.900 595.050 ;
        RECT 542.100 588.600 543.900 593.700 ;
        RECT 545.100 588.000 546.900 592.800 ;
        RECT 548.100 588.600 549.900 593.700 ;
        RECT 551.100 594.600 552.300 596.700 ;
        RECT 569.700 595.800 573.900 596.700 ;
        RECT 583.950 595.800 586.050 597.900 ;
        RECT 593.100 596.700 594.300 601.950 ;
        RECT 596.100 600.150 597.900 601.950 ;
        RECT 614.100 600.150 615.900 601.950 ;
        RECT 617.700 597.600 618.900 601.950 ;
        RECT 620.100 600.150 621.900 601.950 ;
        RECT 629.550 601.050 630.450 605.550 ;
        RECT 638.100 604.050 639.300 617.400 ;
        RECT 659.400 617.100 660.900 617.400 ;
        RECT 665.100 617.400 666.900 623.400 ;
        RECT 665.100 617.100 666.000 617.400 ;
        RECT 659.400 616.200 666.000 617.100 ;
        RECT 659.100 604.050 660.900 605.850 ;
        RECT 665.100 604.050 666.000 616.200 ;
        RECT 680.100 612.300 681.900 623.400 ;
        RECT 683.100 613.200 684.900 624.000 ;
        RECT 686.100 612.300 687.900 623.400 ;
        RECT 680.100 611.400 687.900 612.300 ;
        RECT 689.100 611.400 690.900 623.400 ;
        RECT 707.100 617.400 708.900 624.000 ;
        RECT 710.100 617.400 711.900 623.400 ;
        RECT 713.100 617.400 714.900 624.000 ;
        RECT 728.700 617.400 730.500 624.000 ;
        RECT 675.000 606.450 679.050 607.050 ;
        RECT 674.550 604.950 679.050 606.450 ;
        RECT 634.950 601.950 637.050 604.050 ;
        RECT 637.950 601.950 640.050 604.050 ;
        RECT 640.950 601.950 643.050 604.050 ;
        RECT 655.950 601.950 658.050 604.050 ;
        RECT 658.950 601.950 661.050 604.050 ;
        RECT 661.950 601.950 664.050 604.050 ;
        RECT 664.950 601.950 667.050 604.050 ;
        RECT 629.550 599.550 634.050 601.050 ;
        RECT 635.250 600.150 637.050 601.950 ;
        RECT 630.000 598.950 634.050 599.550 ;
        RECT 617.700 596.700 621.300 597.600 ;
        RECT 593.100 595.800 597.300 596.700 ;
        RECT 551.100 588.600 552.900 594.600 ;
        RECT 569.700 588.600 571.500 595.800 ;
        RECT 574.800 588.000 576.600 594.600 ;
        RECT 590.400 588.000 592.200 594.600 ;
        RECT 595.500 588.600 597.300 595.800 ;
        RECT 611.100 593.700 618.900 595.050 ;
        RECT 611.100 588.600 612.900 593.700 ;
        RECT 614.100 588.000 615.900 592.800 ;
        RECT 617.100 588.600 618.900 593.700 ;
        RECT 620.100 594.600 621.300 596.700 ;
        RECT 625.950 597.450 628.050 598.050 ;
        RECT 634.950 597.450 637.050 598.050 ;
        RECT 625.950 596.550 637.050 597.450 ;
        RECT 625.950 595.950 628.050 596.550 ;
        RECT 634.950 595.950 637.050 596.550 ;
        RECT 638.100 596.700 639.300 601.950 ;
        RECT 641.100 600.150 642.900 601.950 ;
        RECT 656.100 600.150 657.900 601.950 ;
        RECT 662.100 600.150 663.900 601.950 ;
        RECT 665.100 598.200 666.000 601.950 ;
        RECT 638.100 595.800 642.300 596.700 ;
        RECT 620.100 588.600 621.900 594.600 ;
        RECT 635.400 588.000 637.200 594.600 ;
        RECT 640.500 588.600 642.300 595.800 ;
        RECT 656.100 588.000 657.900 597.600 ;
        RECT 662.700 597.000 666.000 598.200 ;
        RECT 674.550 597.450 675.450 604.950 ;
        RECT 683.250 604.050 685.050 605.850 ;
        RECT 689.700 604.050 690.600 611.400 ;
        RECT 710.700 604.050 711.900 617.400 ;
        RECT 729.000 614.100 730.800 615.900 ;
        RECT 731.700 612.900 733.500 623.400 ;
        RECT 731.100 611.400 733.500 612.900 ;
        RECT 736.800 611.400 738.600 624.000 ;
        RECT 752.400 611.400 754.200 624.000 ;
        RECT 757.500 612.900 759.300 623.400 ;
        RECT 760.500 617.400 762.300 624.000 ;
        RECT 776.100 617.400 777.900 624.000 ;
        RECT 779.100 617.400 780.900 623.400 ;
        RECT 782.100 617.400 783.900 624.000 ;
        RECT 800.100 617.400 801.900 624.000 ;
        RECT 803.100 617.400 804.900 623.400 ;
        RECT 821.100 617.400 822.900 624.000 ;
        RECT 824.100 617.400 825.900 623.400 ;
        RECT 827.100 618.000 828.900 624.000 ;
        RECT 760.200 614.100 762.000 615.900 ;
        RECT 757.500 611.400 759.900 612.900 ;
        RECT 731.100 604.050 732.300 611.400 ;
        RECT 745.950 609.450 748.050 610.050 ;
        RECT 754.950 609.450 757.050 610.050 ;
        RECT 745.950 608.550 757.050 609.450 ;
        RECT 745.950 607.950 748.050 608.550 ;
        RECT 754.950 607.950 757.050 608.550 ;
        RECT 737.100 604.050 738.900 605.850 ;
        RECT 752.100 604.050 753.900 605.850 ;
        RECT 758.700 604.050 759.900 611.400 ;
        RECT 779.100 604.050 780.300 617.400 ;
        RECT 800.100 604.050 801.900 605.850 ;
        RECT 803.100 604.050 804.300 617.400 ;
        RECT 824.400 617.100 825.900 617.400 ;
        RECT 830.100 617.400 831.900 623.400 ;
        RECT 830.100 617.100 831.000 617.400 ;
        RECT 824.400 616.200 831.000 617.100 ;
        RECT 824.100 604.050 825.900 605.850 ;
        RECT 830.100 604.050 831.000 616.200 ;
        RECT 845.100 612.300 846.900 623.400 ;
        RECT 848.100 613.200 849.900 624.000 ;
        RECT 851.100 612.300 852.900 623.400 ;
        RECT 845.100 611.400 852.900 612.300 ;
        RECT 854.100 611.400 855.900 623.400 ;
        RECT 869.100 617.400 870.900 624.000 ;
        RECT 872.100 617.400 873.900 623.400 ;
        RECT 875.100 617.400 876.900 624.000 ;
        RECT 890.100 617.400 891.900 624.000 ;
        RECT 893.100 617.400 894.900 623.400 ;
        RECT 896.100 618.000 897.900 624.000 ;
        RECT 848.250 604.050 850.050 605.850 ;
        RECT 854.700 604.050 855.600 611.400 ;
        RECT 872.100 604.050 873.300 617.400 ;
        RECT 893.400 617.100 894.900 617.400 ;
        RECT 899.100 617.400 900.900 623.400 ;
        RECT 899.100 617.100 900.000 617.400 ;
        RECT 893.400 616.200 900.000 617.100 ;
        RECT 874.950 609.450 877.050 610.200 ;
        RECT 874.950 608.550 885.450 609.450 ;
        RECT 874.950 608.100 877.050 608.550 ;
        RECT 679.950 601.950 682.050 604.050 ;
        RECT 682.950 601.950 685.050 604.050 ;
        RECT 685.950 601.950 688.050 604.050 ;
        RECT 688.950 601.950 691.050 604.050 ;
        RECT 706.950 601.950 709.050 604.050 ;
        RECT 709.950 601.950 712.050 604.050 ;
        RECT 712.950 601.950 715.050 604.050 ;
        RECT 727.950 601.950 730.050 604.050 ;
        RECT 730.950 601.950 733.050 604.050 ;
        RECT 733.950 601.950 736.050 604.050 ;
        RECT 736.950 601.950 739.050 604.050 ;
        RECT 751.950 601.950 754.050 604.050 ;
        RECT 754.950 601.950 757.050 604.050 ;
        RECT 757.950 601.950 760.050 604.050 ;
        RECT 760.950 601.950 763.050 604.050 ;
        RECT 775.950 601.950 778.050 604.050 ;
        RECT 778.950 601.950 781.050 604.050 ;
        RECT 781.950 601.950 784.050 604.050 ;
        RECT 799.950 601.950 802.050 604.050 ;
        RECT 802.950 601.950 805.050 604.050 ;
        RECT 820.950 601.950 823.050 604.050 ;
        RECT 823.950 601.950 826.050 604.050 ;
        RECT 826.950 601.950 829.050 604.050 ;
        RECT 829.950 601.950 832.050 604.050 ;
        RECT 844.950 601.950 847.050 604.050 ;
        RECT 847.950 601.950 850.050 604.050 ;
        RECT 850.950 601.950 853.050 604.050 ;
        RECT 853.950 601.950 856.050 604.050 ;
        RECT 868.950 601.950 871.050 604.050 ;
        RECT 871.950 601.950 874.050 604.050 ;
        RECT 874.950 601.950 877.050 604.050 ;
        RECT 680.100 600.150 681.900 601.950 ;
        RECT 686.250 600.150 688.050 601.950 ;
        RECT 679.950 597.450 682.050 598.050 ;
        RECT 662.700 588.600 664.500 597.000 ;
        RECT 674.550 596.550 682.050 597.450 ;
        RECT 679.950 595.950 682.050 596.550 ;
        RECT 689.700 594.600 690.600 601.950 ;
        RECT 707.100 600.150 708.900 601.950 ;
        RECT 710.700 596.700 711.900 601.950 ;
        RECT 712.950 600.150 714.750 601.950 ;
        RECT 728.100 600.150 729.900 601.950 ;
        RECT 681.000 588.000 682.800 594.600 ;
        RECT 685.500 593.400 690.600 594.600 ;
        RECT 707.700 595.800 711.900 596.700 ;
        RECT 712.950 597.450 715.050 598.050 ;
        RECT 721.950 597.450 724.050 598.050 ;
        RECT 731.100 597.600 732.300 601.950 ;
        RECT 734.100 600.150 735.900 601.950 ;
        RECT 755.100 600.150 756.900 601.950 ;
        RECT 712.950 596.550 724.050 597.450 ;
        RECT 712.950 595.950 715.050 596.550 ;
        RECT 721.950 595.950 724.050 596.550 ;
        RECT 728.700 596.700 732.300 597.600 ;
        RECT 758.700 597.600 759.900 601.950 ;
        RECT 761.100 600.150 762.900 601.950 ;
        RECT 776.250 600.150 778.050 601.950 ;
        RECT 758.700 596.700 762.300 597.600 ;
        RECT 685.500 588.600 687.300 593.400 ;
        RECT 688.500 588.000 690.300 591.600 ;
        RECT 707.700 588.600 709.500 595.800 ;
        RECT 728.700 594.600 729.900 596.700 ;
        RECT 712.800 588.000 714.600 594.600 ;
        RECT 728.100 588.600 729.900 594.600 ;
        RECT 731.100 593.700 738.900 595.050 ;
        RECT 731.100 588.600 732.900 593.700 ;
        RECT 734.100 588.000 735.900 592.800 ;
        RECT 737.100 588.600 738.900 593.700 ;
        RECT 752.100 593.700 759.900 595.050 ;
        RECT 752.100 588.600 753.900 593.700 ;
        RECT 755.100 588.000 756.900 592.800 ;
        RECT 758.100 588.600 759.900 593.700 ;
        RECT 761.100 594.600 762.300 596.700 ;
        RECT 779.100 596.700 780.300 601.950 ;
        RECT 782.100 600.150 783.900 601.950 ;
        RECT 779.100 595.800 783.300 596.700 ;
        RECT 761.100 588.600 762.900 594.600 ;
        RECT 776.400 588.000 778.200 594.600 ;
        RECT 781.500 588.600 783.300 595.800 ;
        RECT 803.100 591.600 804.300 601.950 ;
        RECT 821.100 600.150 822.900 601.950 ;
        RECT 827.100 600.150 828.900 601.950 ;
        RECT 830.100 598.200 831.000 601.950 ;
        RECT 845.100 600.150 846.900 601.950 ;
        RECT 851.250 600.150 853.050 601.950 ;
        RECT 800.100 588.000 801.900 591.600 ;
        RECT 803.100 588.600 804.900 591.600 ;
        RECT 821.100 588.000 822.900 597.600 ;
        RECT 827.700 597.000 831.000 598.200 ;
        RECT 827.700 588.600 829.500 597.000 ;
        RECT 854.700 594.600 855.600 601.950 ;
        RECT 869.250 600.150 871.050 601.950 ;
        RECT 872.100 596.700 873.300 601.950 ;
        RECT 875.100 600.150 876.900 601.950 ;
        RECT 884.550 601.050 885.450 608.550 ;
        RECT 893.100 604.050 894.900 605.850 ;
        RECT 899.100 604.050 900.000 616.200 ;
        RECT 917.100 611.400 918.900 623.400 ;
        RECT 920.100 612.000 921.900 624.000 ;
        RECT 923.100 617.400 924.900 623.400 ;
        RECT 926.100 617.400 927.900 624.000 ;
        RECT 941.100 617.400 942.900 624.000 ;
        RECT 944.100 617.400 945.900 623.400 ;
        RECT 947.100 618.000 948.900 624.000 ;
        RECT 917.700 604.050 918.600 611.400 ;
        RECT 921.000 604.050 922.800 605.850 ;
        RECT 889.950 601.950 892.050 604.050 ;
        RECT 892.950 601.950 895.050 604.050 ;
        RECT 895.950 601.950 898.050 604.050 ;
        RECT 898.950 601.950 901.050 604.050 ;
        RECT 917.100 601.950 919.200 604.050 ;
        RECT 920.400 601.950 922.500 604.050 ;
        RECT 884.550 599.550 889.050 601.050 ;
        RECT 890.100 600.150 891.900 601.950 ;
        RECT 896.100 600.150 897.900 601.950 ;
        RECT 885.000 598.950 889.050 599.550 ;
        RECT 899.100 598.200 900.000 601.950 ;
        RECT 872.100 595.800 876.300 596.700 ;
        RECT 846.000 588.000 847.800 594.600 ;
        RECT 850.500 593.400 855.600 594.600 ;
        RECT 850.500 588.600 852.300 593.400 ;
        RECT 853.500 588.000 855.300 591.600 ;
        RECT 869.400 588.000 871.200 594.600 ;
        RECT 874.500 588.600 876.300 595.800 ;
        RECT 890.100 588.000 891.900 597.600 ;
        RECT 896.700 597.000 900.000 598.200 ;
        RECT 896.700 588.600 898.500 597.000 ;
        RECT 917.700 594.600 918.600 601.950 ;
        RECT 924.000 597.300 924.900 617.400 ;
        RECT 944.400 617.100 945.900 617.400 ;
        RECT 950.100 617.400 951.900 623.400 ;
        RECT 950.100 617.100 951.000 617.400 ;
        RECT 944.400 616.200 951.000 617.100 ;
        RECT 934.950 609.450 937.050 610.050 ;
        RECT 946.950 609.450 949.050 610.200 ;
        RECT 934.950 608.550 949.050 609.450 ;
        RECT 934.950 607.950 937.050 608.550 ;
        RECT 946.950 608.100 949.050 608.550 ;
        RECT 944.100 604.050 945.900 605.850 ;
        RECT 950.100 604.050 951.000 616.200 ;
        RECT 968.400 611.400 970.200 624.000 ;
        RECT 973.500 612.900 975.300 623.400 ;
        RECT 976.500 617.400 978.300 624.000 ;
        RECT 992.100 617.400 993.900 624.000 ;
        RECT 995.100 617.400 996.900 623.400 ;
        RECT 998.100 618.000 999.900 624.000 ;
        RECT 995.400 617.100 996.900 617.400 ;
        RECT 1001.100 617.400 1002.900 623.400 ;
        RECT 1001.100 617.100 1002.000 617.400 ;
        RECT 995.400 616.200 1002.000 617.100 ;
        RECT 976.200 614.100 978.000 615.900 ;
        RECT 973.500 611.400 975.900 612.900 ;
        RECT 968.100 604.050 969.900 605.850 ;
        RECT 974.700 604.050 975.900 611.400 ;
        RECT 979.950 606.450 984.000 607.050 ;
        RECT 979.950 604.950 984.450 606.450 ;
        RECT 925.800 601.950 927.900 604.050 ;
        RECT 940.950 601.950 943.050 604.050 ;
        RECT 943.950 601.950 946.050 604.050 ;
        RECT 946.950 601.950 949.050 604.050 ;
        RECT 949.950 601.950 952.050 604.050 ;
        RECT 967.950 601.950 970.050 604.050 ;
        RECT 970.950 601.950 973.050 604.050 ;
        RECT 973.950 601.950 976.050 604.050 ;
        RECT 976.950 601.950 979.050 604.050 ;
        RECT 925.950 600.150 927.750 601.950 ;
        RECT 941.100 600.150 942.900 601.950 ;
        RECT 947.100 600.150 948.900 601.950 ;
        RECT 950.100 598.200 951.000 601.950 ;
        RECT 955.950 600.450 958.050 601.050 ;
        RECT 964.950 600.450 967.050 601.050 ;
        RECT 955.950 599.550 967.050 600.450 ;
        RECT 971.100 600.150 972.900 601.950 ;
        RECT 955.950 598.950 958.050 599.550 ;
        RECT 964.950 598.950 967.050 599.550 ;
        RECT 919.500 596.400 927.900 597.300 ;
        RECT 919.500 595.500 921.300 596.400 ;
        RECT 917.700 592.800 920.400 594.600 ;
        RECT 918.600 588.600 920.400 592.800 ;
        RECT 921.600 588.000 923.400 594.600 ;
        RECT 926.100 588.600 927.900 596.400 ;
        RECT 941.100 588.000 942.900 597.600 ;
        RECT 947.700 597.000 951.000 598.200 ;
        RECT 974.700 597.600 975.900 601.950 ;
        RECT 977.100 600.150 978.900 601.950 ;
        RECT 983.550 600.450 984.450 604.950 ;
        RECT 995.100 604.050 996.900 605.850 ;
        RECT 1001.100 604.050 1002.000 616.200 ;
        RECT 991.950 601.950 994.050 604.050 ;
        RECT 994.950 601.950 997.050 604.050 ;
        RECT 997.950 601.950 1000.050 604.050 ;
        RECT 1000.950 601.950 1003.050 604.050 ;
        RECT 988.950 600.450 991.050 601.050 ;
        RECT 983.550 599.550 991.050 600.450 ;
        RECT 992.100 600.150 993.900 601.950 ;
        RECT 998.100 600.150 999.900 601.950 ;
        RECT 988.950 598.950 991.050 599.550 ;
        RECT 1001.100 598.200 1002.000 601.950 ;
        RECT 947.700 588.600 949.500 597.000 ;
        RECT 974.700 596.700 978.300 597.600 ;
        RECT 968.100 593.700 975.900 595.050 ;
        RECT 968.100 588.600 969.900 593.700 ;
        RECT 971.100 588.000 972.900 592.800 ;
        RECT 974.100 588.600 975.900 593.700 ;
        RECT 977.100 594.600 978.300 596.700 ;
        RECT 977.100 588.600 978.900 594.600 ;
        RECT 992.100 588.000 993.900 597.600 ;
        RECT 998.700 597.000 1002.000 598.200 ;
        RECT 998.700 588.600 1000.500 597.000 ;
        RECT 17.400 578.400 19.200 585.000 ;
        RECT 22.500 577.200 24.300 584.400 ;
        RECT 41.100 578.400 42.900 585.000 ;
        RECT 44.100 577.500 45.900 584.400 ;
        RECT 47.100 578.400 48.900 585.000 ;
        RECT 50.100 577.500 51.900 584.400 ;
        RECT 53.100 578.400 54.900 585.000 ;
        RECT 56.100 577.500 57.900 584.400 ;
        RECT 59.100 578.400 60.900 585.000 ;
        RECT 62.100 577.500 63.900 584.400 ;
        RECT 65.100 578.400 66.900 585.000 ;
        RECT 69.150 580.200 70.950 584.400 ;
        RECT 68.550 578.400 70.950 580.200 ;
        RECT 72.150 578.400 73.950 585.000 ;
        RECT 76.950 582.300 78.750 584.400 ;
        RECT 75.150 581.400 78.750 582.300 ;
        RECT 81.450 581.400 83.250 585.000 ;
        RECT 84.750 581.400 86.550 584.400 ;
        RECT 87.750 581.400 89.550 585.000 ;
        RECT 92.250 581.400 94.050 584.400 ;
        RECT 74.850 580.800 78.750 581.400 ;
        RECT 74.850 579.300 76.950 580.800 ;
        RECT 84.750 580.500 85.800 581.400 ;
        RECT 20.100 576.300 24.300 577.200 ;
        RECT 43.050 576.300 45.900 577.500 ;
        RECT 48.000 576.300 51.900 577.500 ;
        RECT 54.000 576.300 57.900 577.500 ;
        RECT 60.000 576.300 63.900 577.500 ;
        RECT 17.250 571.050 19.050 572.850 ;
        RECT 20.100 571.050 21.300 576.300 ;
        RECT 23.100 571.050 24.900 572.850 ;
        RECT 43.050 571.050 44.100 576.300 ;
        RECT 48.000 575.400 49.200 576.300 ;
        RECT 54.000 575.400 55.200 576.300 ;
        RECT 60.000 575.400 61.200 576.300 ;
        RECT 45.000 574.200 49.200 575.400 ;
        RECT 45.000 573.600 46.800 574.200 ;
        RECT 16.950 568.950 19.050 571.050 ;
        RECT 19.950 568.950 22.050 571.050 ;
        RECT 22.950 568.950 25.050 571.050 ;
        RECT 43.050 568.950 46.200 571.050 ;
        RECT 20.100 555.600 21.300 568.950 ;
        RECT 43.050 563.700 44.100 568.950 ;
        RECT 48.000 563.700 49.200 574.200 ;
        RECT 51.000 574.200 55.200 575.400 ;
        RECT 51.000 573.600 52.800 574.200 ;
        RECT 54.000 563.700 55.200 574.200 ;
        RECT 57.000 574.200 61.200 575.400 ;
        RECT 57.000 573.600 58.800 574.200 ;
        RECT 60.000 563.700 61.200 574.200 ;
        RECT 62.400 571.050 64.200 572.850 ;
        RECT 62.100 568.950 64.200 571.050 ;
        RECT 68.550 563.700 69.450 578.400 ;
        RECT 77.850 577.800 79.650 579.600 ;
        RECT 80.850 579.450 85.800 580.500 ;
        RECT 80.850 578.700 82.650 579.450 ;
        RECT 92.250 579.300 94.650 581.400 ;
        RECT 97.350 578.400 99.150 585.000 ;
        RECT 100.650 578.400 102.450 584.400 ;
        RECT 77.850 576.000 78.900 577.800 ;
        RECT 88.050 576.000 89.850 576.600 ;
        RECT 77.850 574.800 89.850 576.000 ;
        RECT 70.950 573.600 78.900 574.800 ;
        RECT 70.950 571.050 72.750 573.600 ;
        RECT 77.100 573.000 78.900 573.600 ;
        RECT 74.100 571.800 75.900 572.400 ;
        RECT 70.950 568.950 73.050 571.050 ;
        RECT 74.100 570.600 82.200 571.800 ;
        RECT 80.100 568.950 82.200 570.600 ;
        RECT 78.450 563.700 80.250 564.000 ;
        RECT 43.050 562.500 45.900 563.700 ;
        RECT 48.000 562.500 51.900 563.700 ;
        RECT 54.000 562.500 57.900 563.700 ;
        RECT 60.000 562.500 63.900 563.700 ;
        RECT 17.100 549.000 18.900 555.600 ;
        RECT 20.100 549.600 21.900 555.600 ;
        RECT 23.100 549.000 24.900 555.600 ;
        RECT 41.100 549.000 42.900 561.600 ;
        RECT 44.100 549.600 45.900 562.500 ;
        RECT 47.100 549.000 48.900 561.600 ;
        RECT 50.100 549.600 51.900 562.500 ;
        RECT 53.100 549.000 54.900 561.600 ;
        RECT 56.100 549.600 57.900 562.500 ;
        RECT 59.100 549.000 60.900 561.600 ;
        RECT 62.100 549.600 63.900 562.500 ;
        RECT 68.550 563.100 80.250 563.700 ;
        RECT 68.550 562.500 86.850 563.100 ;
        RECT 68.550 561.600 69.450 562.500 ;
        RECT 78.450 562.200 86.850 562.500 ;
        RECT 65.100 549.000 66.900 561.600 ;
        RECT 68.550 559.800 70.950 561.600 ;
        RECT 69.150 549.600 70.950 559.800 ;
        RECT 72.150 549.000 73.950 561.600 ;
        RECT 83.250 560.700 85.050 561.300 ;
        RECT 77.250 559.500 85.050 560.700 ;
        RECT 85.950 560.100 86.850 562.200 ;
        RECT 88.950 562.200 89.850 574.800 ;
        RECT 101.250 571.050 102.450 578.400 ;
        RECT 96.150 569.250 102.450 571.050 ;
        RECT 97.950 568.950 102.450 569.250 ;
        RECT 92.550 566.100 94.650 566.400 ;
        RECT 98.550 566.100 100.350 566.250 ;
        RECT 92.550 564.900 100.350 566.100 ;
        RECT 92.550 564.300 94.650 564.900 ;
        RECT 98.550 564.450 100.350 564.900 ;
        RECT 88.950 561.300 93.750 562.200 ;
        RECT 101.250 561.600 102.450 568.950 ;
        RECT 92.550 560.400 93.750 561.300 ;
        RECT 89.850 560.100 91.650 560.400 ;
        RECT 77.250 558.600 79.350 559.500 ;
        RECT 85.950 559.200 91.650 560.100 ;
        RECT 89.850 558.600 91.650 559.200 ;
        RECT 92.550 558.600 95.550 560.400 ;
        RECT 77.550 549.600 79.350 558.600 ;
        RECT 81.450 557.550 83.250 558.300 ;
        RECT 86.250 557.550 88.050 558.300 ;
        RECT 81.450 556.500 88.050 557.550 ;
        RECT 82.350 549.000 84.150 555.600 ;
        RECT 85.350 549.600 87.150 556.500 ;
        RECT 92.550 555.600 94.650 557.700 ;
        RECT 88.350 549.000 90.150 555.600 ;
        RECT 92.850 549.600 94.650 555.600 ;
        RECT 97.650 549.000 99.450 561.600 ;
        RECT 100.650 549.600 102.450 561.600 ;
        RECT 104.550 578.400 106.350 584.400 ;
        RECT 107.850 578.400 109.650 585.000 ;
        RECT 112.950 581.400 114.750 584.400 ;
        RECT 117.450 581.400 119.250 585.000 ;
        RECT 120.450 581.400 122.250 584.400 ;
        RECT 123.750 581.400 125.550 585.000 ;
        RECT 128.250 582.300 130.050 584.400 ;
        RECT 128.250 581.400 131.850 582.300 ;
        RECT 112.350 579.300 114.750 581.400 ;
        RECT 121.200 580.500 122.250 581.400 ;
        RECT 128.250 580.800 132.150 581.400 ;
        RECT 121.200 579.450 126.150 580.500 ;
        RECT 124.350 578.700 126.150 579.450 ;
        RECT 104.550 571.050 105.750 578.400 ;
        RECT 127.350 577.800 129.150 579.600 ;
        RECT 130.050 579.300 132.150 580.800 ;
        RECT 133.050 578.400 134.850 585.000 ;
        RECT 136.050 580.200 137.850 584.400 ;
        RECT 152.100 581.400 153.900 585.000 ;
        RECT 155.100 581.400 156.900 584.400 ;
        RECT 158.100 581.400 159.900 585.000 ;
        RECT 136.050 578.400 138.450 580.200 ;
        RECT 117.150 576.000 118.950 576.600 ;
        RECT 128.100 576.000 129.150 577.800 ;
        RECT 117.150 574.800 129.150 576.000 ;
        RECT 104.550 569.250 110.850 571.050 ;
        RECT 104.550 568.950 109.050 569.250 ;
        RECT 104.550 561.600 105.750 568.950 ;
        RECT 106.650 566.100 108.450 566.250 ;
        RECT 112.350 566.100 114.450 566.400 ;
        RECT 106.650 564.900 114.450 566.100 ;
        RECT 106.650 564.450 108.450 564.900 ;
        RECT 112.350 564.300 114.450 564.900 ;
        RECT 117.150 562.200 118.050 574.800 ;
        RECT 128.100 573.600 136.050 574.800 ;
        RECT 128.100 573.000 129.900 573.600 ;
        RECT 131.100 571.800 132.900 572.400 ;
        RECT 124.800 570.600 132.900 571.800 ;
        RECT 134.250 571.050 136.050 573.600 ;
        RECT 124.800 568.950 126.900 570.600 ;
        RECT 133.950 568.950 136.050 571.050 ;
        RECT 126.750 563.700 128.550 564.000 ;
        RECT 137.550 563.700 138.450 578.400 ;
        RECT 155.400 571.050 156.300 581.400 ;
        RECT 176.400 578.400 178.200 585.000 ;
        RECT 181.500 577.200 183.300 584.400 ;
        RECT 197.100 578.400 198.900 584.400 ;
        RECT 179.100 576.300 183.300 577.200 ;
        RECT 197.700 576.300 198.900 578.400 ;
        RECT 200.100 579.300 201.900 584.400 ;
        RECT 203.100 580.200 204.900 585.000 ;
        RECT 206.100 579.300 207.900 584.400 ;
        RECT 221.100 581.400 222.900 585.000 ;
        RECT 224.100 581.400 225.900 584.400 ;
        RECT 200.100 577.950 207.900 579.300 ;
        RECT 176.250 571.050 178.050 572.850 ;
        RECT 179.100 571.050 180.300 576.300 ;
        RECT 197.700 575.400 201.300 576.300 ;
        RECT 182.100 571.050 183.900 572.850 ;
        RECT 197.100 571.050 198.900 572.850 ;
        RECT 200.100 571.050 201.300 575.400 ;
        RECT 203.100 571.050 204.900 572.850 ;
        RECT 224.100 571.050 225.300 581.400 ;
        RECT 239.100 579.300 240.900 584.400 ;
        RECT 242.100 580.200 243.900 585.000 ;
        RECT 245.100 579.300 246.900 584.400 ;
        RECT 239.100 577.950 246.900 579.300 ;
        RECT 248.100 578.400 249.900 584.400 ;
        RECT 266.400 578.400 268.200 585.000 ;
        RECT 248.100 576.300 249.300 578.400 ;
        RECT 271.500 577.200 273.300 584.400 ;
        RECT 290.400 578.400 292.200 585.000 ;
        RECT 295.500 577.200 297.300 584.400 ;
        RECT 300.150 580.200 301.950 584.400 ;
        RECT 245.700 575.400 249.300 576.300 ;
        RECT 269.100 576.300 273.300 577.200 ;
        RECT 293.100 576.300 297.300 577.200 ;
        RECT 299.550 578.400 301.950 580.200 ;
        RECT 303.150 578.400 304.950 585.000 ;
        RECT 307.950 582.300 309.750 584.400 ;
        RECT 306.150 581.400 309.750 582.300 ;
        RECT 312.450 581.400 314.250 585.000 ;
        RECT 315.750 581.400 317.550 584.400 ;
        RECT 318.750 581.400 320.550 585.000 ;
        RECT 323.250 581.400 325.050 584.400 ;
        RECT 305.850 580.800 309.750 581.400 ;
        RECT 305.850 579.300 307.950 580.800 ;
        RECT 315.750 580.500 316.800 581.400 ;
        RECT 242.100 571.050 243.900 572.850 ;
        RECT 245.700 571.050 246.900 575.400 ;
        RECT 248.100 571.050 249.900 572.850 ;
        RECT 266.250 571.050 268.050 572.850 ;
        RECT 269.100 571.050 270.300 576.300 ;
        RECT 272.100 571.050 273.900 572.850 ;
        RECT 290.250 571.050 292.050 572.850 ;
        RECT 293.100 571.050 294.300 576.300 ;
        RECT 296.100 571.050 297.900 572.850 ;
        RECT 151.950 568.950 154.050 571.050 ;
        RECT 154.950 568.950 157.050 571.050 ;
        RECT 157.950 568.950 160.050 571.050 ;
        RECT 175.950 568.950 178.050 571.050 ;
        RECT 178.950 568.950 181.050 571.050 ;
        RECT 181.950 568.950 184.050 571.050 ;
        RECT 196.950 568.950 199.050 571.050 ;
        RECT 199.950 568.950 202.050 571.050 ;
        RECT 202.950 568.950 205.050 571.050 ;
        RECT 205.950 568.950 208.050 571.050 ;
        RECT 220.950 568.950 223.050 571.050 ;
        RECT 223.950 568.950 226.050 571.050 ;
        RECT 238.950 568.950 241.050 571.050 ;
        RECT 241.950 568.950 244.050 571.050 ;
        RECT 244.950 568.950 247.050 571.050 ;
        RECT 247.950 568.950 250.050 571.050 ;
        RECT 265.950 568.950 268.050 571.050 ;
        RECT 268.950 568.950 271.050 571.050 ;
        RECT 271.950 568.950 274.050 571.050 ;
        RECT 289.950 568.950 292.050 571.050 ;
        RECT 292.950 568.950 295.050 571.050 ;
        RECT 295.950 568.950 298.050 571.050 ;
        RECT 152.250 567.150 154.050 568.950 ;
        RECT 126.750 563.100 138.450 563.700 ;
        RECT 104.550 549.600 106.350 561.600 ;
        RECT 107.550 549.000 109.350 561.600 ;
        RECT 113.250 561.300 118.050 562.200 ;
        RECT 120.150 562.500 138.450 563.100 ;
        RECT 120.150 562.200 128.550 562.500 ;
        RECT 113.250 560.400 114.450 561.300 ;
        RECT 111.450 558.600 114.450 560.400 ;
        RECT 115.350 560.100 117.150 560.400 ;
        RECT 120.150 560.100 121.050 562.200 ;
        RECT 137.550 561.600 138.450 562.500 ;
        RECT 155.400 561.600 156.300 568.950 ;
        RECT 158.100 567.150 159.900 568.950 ;
        RECT 115.350 559.200 121.050 560.100 ;
        RECT 121.950 560.700 123.750 561.300 ;
        RECT 121.950 559.500 129.750 560.700 ;
        RECT 115.350 558.600 117.150 559.200 ;
        RECT 127.650 558.600 129.750 559.500 ;
        RECT 112.350 555.600 114.450 557.700 ;
        RECT 118.950 557.550 120.750 558.300 ;
        RECT 123.750 557.550 125.550 558.300 ;
        RECT 118.950 556.500 125.550 557.550 ;
        RECT 112.350 549.600 114.150 555.600 ;
        RECT 116.850 549.000 118.650 555.600 ;
        RECT 119.850 549.600 121.650 556.500 ;
        RECT 122.850 549.000 124.650 555.600 ;
        RECT 127.650 549.600 129.450 558.600 ;
        RECT 133.050 549.000 134.850 561.600 ;
        RECT 136.050 559.800 138.450 561.600 ;
        RECT 136.050 549.600 137.850 559.800 ;
        RECT 152.100 549.000 153.900 561.600 ;
        RECT 155.400 560.400 159.000 561.600 ;
        RECT 157.200 549.600 159.000 560.400 ;
        RECT 179.100 555.600 180.300 568.950 ;
        RECT 181.950 564.450 184.050 565.050 ;
        RECT 187.950 564.450 190.050 565.050 ;
        RECT 181.950 563.550 190.050 564.450 ;
        RECT 181.950 562.950 184.050 563.550 ;
        RECT 187.950 562.950 190.050 563.550 ;
        RECT 200.100 561.600 201.300 568.950 ;
        RECT 206.100 567.150 207.900 568.950 ;
        RECT 221.100 567.150 222.900 568.950 ;
        RECT 200.100 560.100 202.500 561.600 ;
        RECT 198.000 557.100 199.800 558.900 ;
        RECT 176.100 549.000 177.900 555.600 ;
        RECT 179.100 549.600 180.900 555.600 ;
        RECT 182.100 549.000 183.900 555.600 ;
        RECT 197.700 549.000 199.500 555.600 ;
        RECT 200.700 549.600 202.500 560.100 ;
        RECT 205.800 549.000 207.600 561.600 ;
        RECT 224.100 555.600 225.300 568.950 ;
        RECT 239.100 567.150 240.900 568.950 ;
        RECT 245.700 561.600 246.900 568.950 ;
        RECT 221.100 549.000 222.900 555.600 ;
        RECT 224.100 549.600 225.900 555.600 ;
        RECT 239.400 549.000 241.200 561.600 ;
        RECT 244.500 560.100 246.900 561.600 ;
        RECT 244.500 549.600 246.300 560.100 ;
        RECT 247.200 557.100 249.000 558.900 ;
        RECT 269.100 555.600 270.300 568.950 ;
        RECT 293.100 555.600 294.300 568.950 ;
        RECT 299.550 563.700 300.450 578.400 ;
        RECT 308.850 577.800 310.650 579.600 ;
        RECT 311.850 579.450 316.800 580.500 ;
        RECT 311.850 578.700 313.650 579.450 ;
        RECT 323.250 579.300 325.650 581.400 ;
        RECT 328.350 578.400 330.150 585.000 ;
        RECT 331.650 578.400 333.450 584.400 ;
        RECT 347.100 581.400 348.900 585.000 ;
        RECT 350.100 581.400 351.900 584.400 ;
        RECT 308.850 576.000 309.900 577.800 ;
        RECT 319.050 576.000 320.850 576.600 ;
        RECT 308.850 574.800 320.850 576.000 ;
        RECT 301.950 573.600 309.900 574.800 ;
        RECT 301.950 571.050 303.750 573.600 ;
        RECT 308.100 573.000 309.900 573.600 ;
        RECT 305.100 571.800 306.900 572.400 ;
        RECT 301.950 568.950 304.050 571.050 ;
        RECT 305.100 570.600 313.200 571.800 ;
        RECT 311.100 568.950 313.200 570.600 ;
        RECT 309.450 563.700 311.250 564.000 ;
        RECT 299.550 563.100 311.250 563.700 ;
        RECT 299.550 562.500 317.850 563.100 ;
        RECT 299.550 561.600 300.450 562.500 ;
        RECT 309.450 562.200 317.850 562.500 ;
        RECT 299.550 559.800 301.950 561.600 ;
        RECT 247.500 549.000 249.300 555.600 ;
        RECT 266.100 549.000 267.900 555.600 ;
        RECT 269.100 549.600 270.900 555.600 ;
        RECT 272.100 549.000 273.900 555.600 ;
        RECT 290.100 549.000 291.900 555.600 ;
        RECT 293.100 549.600 294.900 555.600 ;
        RECT 296.100 549.000 297.900 555.600 ;
        RECT 300.150 549.600 301.950 559.800 ;
        RECT 303.150 549.000 304.950 561.600 ;
        RECT 314.250 560.700 316.050 561.300 ;
        RECT 308.250 559.500 316.050 560.700 ;
        RECT 316.950 560.100 317.850 562.200 ;
        RECT 319.950 562.200 320.850 574.800 ;
        RECT 332.250 571.050 333.450 578.400 ;
        RECT 337.950 579.450 340.050 580.050 ;
        RECT 346.950 579.450 349.050 580.050 ;
        RECT 337.950 578.550 349.050 579.450 ;
        RECT 337.950 577.950 340.050 578.550 ;
        RECT 346.950 577.950 349.050 578.550 ;
        RECT 350.100 571.050 351.300 581.400 ;
        RECT 365.100 579.300 366.900 584.400 ;
        RECT 368.100 580.200 369.900 585.000 ;
        RECT 371.100 579.300 372.900 584.400 ;
        RECT 365.100 577.950 372.900 579.300 ;
        RECT 374.100 578.400 375.900 584.400 ;
        RECT 378.150 580.200 379.950 584.400 ;
        RECT 377.550 578.400 379.950 580.200 ;
        RECT 381.150 578.400 382.950 585.000 ;
        RECT 385.950 582.300 387.750 584.400 ;
        RECT 384.150 581.400 387.750 582.300 ;
        RECT 390.450 581.400 392.250 585.000 ;
        RECT 393.750 581.400 395.550 584.400 ;
        RECT 396.750 581.400 398.550 585.000 ;
        RECT 401.250 581.400 403.050 584.400 ;
        RECT 383.850 580.800 387.750 581.400 ;
        RECT 383.850 579.300 385.950 580.800 ;
        RECT 393.750 580.500 394.800 581.400 ;
        RECT 374.100 576.300 375.300 578.400 ;
        RECT 371.700 575.400 375.300 576.300 ;
        RECT 368.100 571.050 369.900 572.850 ;
        RECT 371.700 571.050 372.900 575.400 ;
        RECT 374.100 571.050 375.900 572.850 ;
        RECT 327.150 569.250 333.450 571.050 ;
        RECT 328.950 568.950 333.450 569.250 ;
        RECT 346.950 568.950 349.050 571.050 ;
        RECT 349.950 568.950 352.050 571.050 ;
        RECT 364.950 568.950 367.050 571.050 ;
        RECT 367.950 568.950 370.050 571.050 ;
        RECT 370.950 568.950 373.050 571.050 ;
        RECT 373.950 568.950 376.050 571.050 ;
        RECT 323.550 566.100 325.650 566.400 ;
        RECT 329.550 566.100 331.350 566.250 ;
        RECT 323.550 564.900 331.350 566.100 ;
        RECT 323.550 564.300 325.650 564.900 ;
        RECT 329.550 564.450 331.350 564.900 ;
        RECT 319.950 561.300 324.750 562.200 ;
        RECT 332.250 561.600 333.450 568.950 ;
        RECT 347.100 567.150 348.900 568.950 ;
        RECT 323.550 560.400 324.750 561.300 ;
        RECT 320.850 560.100 322.650 560.400 ;
        RECT 308.250 558.600 310.350 559.500 ;
        RECT 316.950 559.200 322.650 560.100 ;
        RECT 320.850 558.600 322.650 559.200 ;
        RECT 323.550 558.600 326.550 560.400 ;
        RECT 308.550 549.600 310.350 558.600 ;
        RECT 312.450 557.550 314.250 558.300 ;
        RECT 317.250 557.550 319.050 558.300 ;
        RECT 312.450 556.500 319.050 557.550 ;
        RECT 313.350 549.000 315.150 555.600 ;
        RECT 316.350 549.600 318.150 556.500 ;
        RECT 323.550 555.600 325.650 557.700 ;
        RECT 319.350 549.000 321.150 555.600 ;
        RECT 323.850 549.600 325.650 555.600 ;
        RECT 328.650 549.000 330.450 561.600 ;
        RECT 331.650 549.600 333.450 561.600 ;
        RECT 350.100 555.600 351.300 568.950 ;
        RECT 365.100 567.150 366.900 568.950 ;
        RECT 371.700 561.600 372.900 568.950 ;
        RECT 347.100 549.000 348.900 555.600 ;
        RECT 350.100 549.600 351.900 555.600 ;
        RECT 365.400 549.000 367.200 561.600 ;
        RECT 370.500 560.100 372.900 561.600 ;
        RECT 377.550 563.700 378.450 578.400 ;
        RECT 386.850 577.800 388.650 579.600 ;
        RECT 389.850 579.450 394.800 580.500 ;
        RECT 389.850 578.700 391.650 579.450 ;
        RECT 401.250 579.300 403.650 581.400 ;
        RECT 406.350 578.400 408.150 585.000 ;
        RECT 409.650 578.400 411.450 584.400 ;
        RECT 428.400 578.400 430.200 585.000 ;
        RECT 386.850 576.000 387.900 577.800 ;
        RECT 397.050 576.000 398.850 576.600 ;
        RECT 386.850 574.800 398.850 576.000 ;
        RECT 379.950 573.600 387.900 574.800 ;
        RECT 379.950 571.050 381.750 573.600 ;
        RECT 386.100 573.000 387.900 573.600 ;
        RECT 383.100 571.800 384.900 572.400 ;
        RECT 379.950 568.950 382.050 571.050 ;
        RECT 383.100 570.600 391.200 571.800 ;
        RECT 389.100 568.950 391.200 570.600 ;
        RECT 387.450 563.700 389.250 564.000 ;
        RECT 377.550 563.100 389.250 563.700 ;
        RECT 377.550 562.500 395.850 563.100 ;
        RECT 377.550 561.600 378.450 562.500 ;
        RECT 387.450 562.200 395.850 562.500 ;
        RECT 370.500 549.600 372.300 560.100 ;
        RECT 377.550 559.800 379.950 561.600 ;
        RECT 373.200 557.100 375.000 558.900 ;
        RECT 373.500 549.000 375.300 555.600 ;
        RECT 378.150 549.600 379.950 559.800 ;
        RECT 381.150 549.000 382.950 561.600 ;
        RECT 392.250 560.700 394.050 561.300 ;
        RECT 386.250 559.500 394.050 560.700 ;
        RECT 394.950 560.100 395.850 562.200 ;
        RECT 397.950 562.200 398.850 574.800 ;
        RECT 410.250 571.050 411.450 578.400 ;
        RECT 433.500 577.200 435.300 584.400 ;
        RECT 431.100 576.300 435.300 577.200 ;
        RECT 437.550 578.400 439.350 584.400 ;
        RECT 440.850 578.400 442.650 585.000 ;
        RECT 445.950 581.400 447.750 584.400 ;
        RECT 450.450 581.400 452.250 585.000 ;
        RECT 453.450 581.400 455.250 584.400 ;
        RECT 456.750 581.400 458.550 585.000 ;
        RECT 461.250 582.300 463.050 584.400 ;
        RECT 461.250 581.400 464.850 582.300 ;
        RECT 445.350 579.300 447.750 581.400 ;
        RECT 454.200 580.500 455.250 581.400 ;
        RECT 461.250 580.800 465.150 581.400 ;
        RECT 454.200 579.450 459.150 580.500 ;
        RECT 457.350 578.700 459.150 579.450 ;
        RECT 428.250 571.050 430.050 572.850 ;
        RECT 431.100 571.050 432.300 576.300 ;
        RECT 434.100 571.050 435.900 572.850 ;
        RECT 437.550 571.050 438.750 578.400 ;
        RECT 460.350 577.800 462.150 579.600 ;
        RECT 463.050 579.300 465.150 580.800 ;
        RECT 466.050 578.400 467.850 585.000 ;
        RECT 469.050 580.200 470.850 584.400 ;
        RECT 474.150 580.200 475.950 584.400 ;
        RECT 469.050 578.400 471.450 580.200 ;
        RECT 450.150 576.000 451.950 576.600 ;
        RECT 461.100 576.000 462.150 577.800 ;
        RECT 450.150 574.800 462.150 576.000 ;
        RECT 405.150 569.250 411.450 571.050 ;
        RECT 406.950 568.950 411.450 569.250 ;
        RECT 427.950 568.950 430.050 571.050 ;
        RECT 430.950 568.950 433.050 571.050 ;
        RECT 433.950 568.950 436.050 571.050 ;
        RECT 437.550 569.250 443.850 571.050 ;
        RECT 437.550 568.950 442.050 569.250 ;
        RECT 401.550 566.100 403.650 566.400 ;
        RECT 407.550 566.100 409.350 566.250 ;
        RECT 401.550 564.900 409.350 566.100 ;
        RECT 401.550 564.300 403.650 564.900 ;
        RECT 407.550 564.450 409.350 564.900 ;
        RECT 397.950 561.300 402.750 562.200 ;
        RECT 410.250 561.600 411.450 568.950 ;
        RECT 401.550 560.400 402.750 561.300 ;
        RECT 398.850 560.100 400.650 560.400 ;
        RECT 386.250 558.600 388.350 559.500 ;
        RECT 394.950 559.200 400.650 560.100 ;
        RECT 398.850 558.600 400.650 559.200 ;
        RECT 401.550 558.600 404.550 560.400 ;
        RECT 386.550 549.600 388.350 558.600 ;
        RECT 390.450 557.550 392.250 558.300 ;
        RECT 395.250 557.550 397.050 558.300 ;
        RECT 390.450 556.500 397.050 557.550 ;
        RECT 391.350 549.000 393.150 555.600 ;
        RECT 394.350 549.600 396.150 556.500 ;
        RECT 401.550 555.600 403.650 557.700 ;
        RECT 397.350 549.000 399.150 555.600 ;
        RECT 401.850 549.600 403.650 555.600 ;
        RECT 406.650 549.000 408.450 561.600 ;
        RECT 409.650 549.600 411.450 561.600 ;
        RECT 431.100 555.600 432.300 568.950 ;
        RECT 437.550 561.600 438.750 568.950 ;
        RECT 439.650 566.100 441.450 566.250 ;
        RECT 445.350 566.100 447.450 566.400 ;
        RECT 439.650 564.900 447.450 566.100 ;
        RECT 439.650 564.450 441.450 564.900 ;
        RECT 445.350 564.300 447.450 564.900 ;
        RECT 450.150 562.200 451.050 574.800 ;
        RECT 461.100 573.600 469.050 574.800 ;
        RECT 461.100 573.000 462.900 573.600 ;
        RECT 464.100 571.800 465.900 572.400 ;
        RECT 457.800 570.600 465.900 571.800 ;
        RECT 467.250 571.050 469.050 573.600 ;
        RECT 457.800 568.950 459.900 570.600 ;
        RECT 466.950 568.950 469.050 571.050 ;
        RECT 459.750 563.700 461.550 564.000 ;
        RECT 470.550 563.700 471.450 578.400 ;
        RECT 459.750 563.100 471.450 563.700 ;
        RECT 428.100 549.000 429.900 555.600 ;
        RECT 431.100 549.600 432.900 555.600 ;
        RECT 434.100 549.000 435.900 555.600 ;
        RECT 437.550 549.600 439.350 561.600 ;
        RECT 440.550 549.000 442.350 561.600 ;
        RECT 446.250 561.300 451.050 562.200 ;
        RECT 453.150 562.500 471.450 563.100 ;
        RECT 453.150 562.200 461.550 562.500 ;
        RECT 446.250 560.400 447.450 561.300 ;
        RECT 444.450 558.600 447.450 560.400 ;
        RECT 448.350 560.100 450.150 560.400 ;
        RECT 453.150 560.100 454.050 562.200 ;
        RECT 470.550 561.600 471.450 562.500 ;
        RECT 448.350 559.200 454.050 560.100 ;
        RECT 454.950 560.700 456.750 561.300 ;
        RECT 454.950 559.500 462.750 560.700 ;
        RECT 448.350 558.600 450.150 559.200 ;
        RECT 460.650 558.600 462.750 559.500 ;
        RECT 445.350 555.600 447.450 557.700 ;
        RECT 451.950 557.550 453.750 558.300 ;
        RECT 456.750 557.550 458.550 558.300 ;
        RECT 451.950 556.500 458.550 557.550 ;
        RECT 445.350 549.600 447.150 555.600 ;
        RECT 449.850 549.000 451.650 555.600 ;
        RECT 452.850 549.600 454.650 556.500 ;
        RECT 455.850 549.000 457.650 555.600 ;
        RECT 460.650 549.600 462.450 558.600 ;
        RECT 466.050 549.000 467.850 561.600 ;
        RECT 469.050 559.800 471.450 561.600 ;
        RECT 473.550 578.400 475.950 580.200 ;
        RECT 477.150 578.400 478.950 585.000 ;
        RECT 481.950 582.300 483.750 584.400 ;
        RECT 480.150 581.400 483.750 582.300 ;
        RECT 486.450 581.400 488.250 585.000 ;
        RECT 489.750 581.400 491.550 584.400 ;
        RECT 492.750 581.400 494.550 585.000 ;
        RECT 497.250 581.400 499.050 584.400 ;
        RECT 479.850 580.800 483.750 581.400 ;
        RECT 479.850 579.300 481.950 580.800 ;
        RECT 489.750 580.500 490.800 581.400 ;
        RECT 473.550 563.700 474.450 578.400 ;
        RECT 482.850 577.800 484.650 579.600 ;
        RECT 485.850 579.450 490.800 580.500 ;
        RECT 485.850 578.700 487.650 579.450 ;
        RECT 497.250 579.300 499.650 581.400 ;
        RECT 502.350 578.400 504.150 585.000 ;
        RECT 505.650 578.400 507.450 584.400 ;
        RECT 521.100 581.400 522.900 585.000 ;
        RECT 524.100 581.400 525.900 584.400 ;
        RECT 482.850 576.000 483.900 577.800 ;
        RECT 493.050 576.000 494.850 576.600 ;
        RECT 482.850 574.800 494.850 576.000 ;
        RECT 475.950 573.600 483.900 574.800 ;
        RECT 475.950 571.050 477.750 573.600 ;
        RECT 482.100 573.000 483.900 573.600 ;
        RECT 479.100 571.800 480.900 572.400 ;
        RECT 475.950 568.950 478.050 571.050 ;
        RECT 479.100 570.600 487.200 571.800 ;
        RECT 485.100 568.950 487.200 570.600 ;
        RECT 483.450 563.700 485.250 564.000 ;
        RECT 473.550 563.100 485.250 563.700 ;
        RECT 473.550 562.500 491.850 563.100 ;
        RECT 473.550 561.600 474.450 562.500 ;
        RECT 483.450 562.200 491.850 562.500 ;
        RECT 473.550 559.800 475.950 561.600 ;
        RECT 469.050 549.600 470.850 559.800 ;
        RECT 474.150 549.600 475.950 559.800 ;
        RECT 477.150 549.000 478.950 561.600 ;
        RECT 488.250 560.700 490.050 561.300 ;
        RECT 482.250 559.500 490.050 560.700 ;
        RECT 490.950 560.100 491.850 562.200 ;
        RECT 493.950 562.200 494.850 574.800 ;
        RECT 506.250 571.050 507.450 578.400 ;
        RECT 524.100 571.050 525.300 581.400 ;
        RECT 539.100 575.400 540.900 585.000 ;
        RECT 545.700 576.000 547.500 584.400 ;
        RECT 563.400 578.400 565.200 585.000 ;
        RECT 568.500 577.200 570.300 584.400 ;
        RECT 566.100 576.300 570.300 577.200 ;
        RECT 587.700 577.200 589.500 584.400 ;
        RECT 592.800 578.400 594.600 585.000 ;
        RECT 597.150 580.200 598.950 584.400 ;
        RECT 596.550 578.400 598.950 580.200 ;
        RECT 600.150 578.400 601.950 585.000 ;
        RECT 604.950 582.300 606.750 584.400 ;
        RECT 603.150 581.400 606.750 582.300 ;
        RECT 609.450 581.400 611.250 585.000 ;
        RECT 612.750 581.400 614.550 584.400 ;
        RECT 615.750 581.400 617.550 585.000 ;
        RECT 620.250 581.400 622.050 584.400 ;
        RECT 602.850 580.800 606.750 581.400 ;
        RECT 602.850 579.300 604.950 580.800 ;
        RECT 612.750 580.500 613.800 581.400 ;
        RECT 587.700 576.300 591.900 577.200 ;
        RECT 545.700 574.800 549.000 576.000 ;
        RECT 539.100 571.050 540.900 572.850 ;
        RECT 545.100 571.050 546.900 572.850 ;
        RECT 548.100 571.050 549.000 574.800 ;
        RECT 563.250 571.050 565.050 572.850 ;
        RECT 566.100 571.050 567.300 576.300 ;
        RECT 582.000 573.450 586.050 574.050 ;
        RECT 569.100 571.050 570.900 572.850 ;
        RECT 581.550 571.950 586.050 573.450 ;
        RECT 501.150 569.250 507.450 571.050 ;
        RECT 502.950 568.950 507.450 569.250 ;
        RECT 520.950 568.950 523.050 571.050 ;
        RECT 523.950 568.950 526.050 571.050 ;
        RECT 538.950 568.950 541.050 571.050 ;
        RECT 541.950 568.950 544.050 571.050 ;
        RECT 544.950 568.950 547.050 571.050 ;
        RECT 547.950 568.950 550.050 571.050 ;
        RECT 562.950 568.950 565.050 571.050 ;
        RECT 565.950 568.950 568.050 571.050 ;
        RECT 568.950 568.950 571.050 571.050 ;
        RECT 497.550 566.100 499.650 566.400 ;
        RECT 503.550 566.100 505.350 566.250 ;
        RECT 497.550 564.900 505.350 566.100 ;
        RECT 497.550 564.300 499.650 564.900 ;
        RECT 503.550 564.450 505.350 564.900 ;
        RECT 493.950 561.300 498.750 562.200 ;
        RECT 506.250 561.600 507.450 568.950 ;
        RECT 521.100 567.150 522.900 568.950 ;
        RECT 497.550 560.400 498.750 561.300 ;
        RECT 494.850 560.100 496.650 560.400 ;
        RECT 482.250 558.600 484.350 559.500 ;
        RECT 490.950 559.200 496.650 560.100 ;
        RECT 494.850 558.600 496.650 559.200 ;
        RECT 497.550 558.600 500.550 560.400 ;
        RECT 482.550 549.600 484.350 558.600 ;
        RECT 486.450 557.550 488.250 558.300 ;
        RECT 491.250 557.550 493.050 558.300 ;
        RECT 486.450 556.500 493.050 557.550 ;
        RECT 487.350 549.000 489.150 555.600 ;
        RECT 490.350 549.600 492.150 556.500 ;
        RECT 497.550 555.600 499.650 557.700 ;
        RECT 493.350 549.000 495.150 555.600 ;
        RECT 497.850 549.600 499.650 555.600 ;
        RECT 502.650 549.000 504.450 561.600 ;
        RECT 505.650 549.600 507.450 561.600 ;
        RECT 524.100 555.600 525.300 568.950 ;
        RECT 542.100 567.150 543.900 568.950 ;
        RECT 526.950 564.450 529.050 565.050 ;
        RECT 544.950 564.450 547.050 565.050 ;
        RECT 526.950 563.550 547.050 564.450 ;
        RECT 526.950 562.950 529.050 563.550 ;
        RECT 544.950 562.950 547.050 563.550 ;
        RECT 548.100 556.800 549.000 568.950 ;
        RECT 550.950 564.450 553.050 565.050 ;
        RECT 562.950 564.450 565.050 565.050 ;
        RECT 550.950 563.550 565.050 564.450 ;
        RECT 550.950 562.950 553.050 563.550 ;
        RECT 562.950 562.950 565.050 563.550 ;
        RECT 542.400 555.900 549.000 556.800 ;
        RECT 542.400 555.600 543.900 555.900 ;
        RECT 521.100 549.000 522.900 555.600 ;
        RECT 524.100 549.600 525.900 555.600 ;
        RECT 539.100 549.000 540.900 555.600 ;
        RECT 542.100 549.600 543.900 555.600 ;
        RECT 548.100 555.600 549.000 555.900 ;
        RECT 566.100 555.600 567.300 568.950 ;
        RECT 571.950 567.450 574.050 568.050 ;
        RECT 581.550 567.450 582.450 571.950 ;
        RECT 587.100 571.050 588.900 572.850 ;
        RECT 590.700 571.050 591.900 576.300 ;
        RECT 592.950 571.050 594.750 572.850 ;
        RECT 586.950 568.950 589.050 571.050 ;
        RECT 589.950 568.950 592.050 571.050 ;
        RECT 592.950 568.950 595.050 571.050 ;
        RECT 571.950 566.550 582.450 567.450 ;
        RECT 571.950 565.950 574.050 566.550 ;
        RECT 590.700 555.600 591.900 568.950 ;
        RECT 596.550 563.700 597.450 578.400 ;
        RECT 605.850 577.800 607.650 579.600 ;
        RECT 608.850 579.450 613.800 580.500 ;
        RECT 608.850 578.700 610.650 579.450 ;
        RECT 620.250 579.300 622.650 581.400 ;
        RECT 625.350 578.400 627.150 585.000 ;
        RECT 628.650 578.400 630.450 584.400 ;
        RECT 605.850 576.000 606.900 577.800 ;
        RECT 616.050 576.000 617.850 576.600 ;
        RECT 605.850 574.800 617.850 576.000 ;
        RECT 598.950 573.600 606.900 574.800 ;
        RECT 598.950 571.050 600.750 573.600 ;
        RECT 605.100 573.000 606.900 573.600 ;
        RECT 602.100 571.800 603.900 572.400 ;
        RECT 598.950 568.950 601.050 571.050 ;
        RECT 602.100 570.600 610.200 571.800 ;
        RECT 608.100 568.950 610.200 570.600 ;
        RECT 606.450 563.700 608.250 564.000 ;
        RECT 596.550 563.100 608.250 563.700 ;
        RECT 596.550 562.500 614.850 563.100 ;
        RECT 596.550 561.600 597.450 562.500 ;
        RECT 606.450 562.200 614.850 562.500 ;
        RECT 596.550 559.800 598.950 561.600 ;
        RECT 545.100 549.000 546.900 555.000 ;
        RECT 548.100 549.600 549.900 555.600 ;
        RECT 563.100 549.000 564.900 555.600 ;
        RECT 566.100 549.600 567.900 555.600 ;
        RECT 569.100 549.000 570.900 555.600 ;
        RECT 587.100 549.000 588.900 555.600 ;
        RECT 590.100 549.600 591.900 555.600 ;
        RECT 593.100 549.000 594.900 555.600 ;
        RECT 597.150 549.600 598.950 559.800 ;
        RECT 600.150 549.000 601.950 561.600 ;
        RECT 611.250 560.700 613.050 561.300 ;
        RECT 605.250 559.500 613.050 560.700 ;
        RECT 613.950 560.100 614.850 562.200 ;
        RECT 616.950 562.200 617.850 574.800 ;
        RECT 629.250 571.050 630.450 578.400 ;
        RECT 644.700 577.200 646.500 584.400 ;
        RECT 649.800 578.400 651.600 585.000 ;
        RECT 669.000 578.400 670.800 585.000 ;
        RECT 673.500 579.600 675.300 584.400 ;
        RECT 676.500 581.400 678.300 585.000 ;
        RECT 673.500 578.400 678.600 579.600 ;
        RECT 644.700 576.300 648.900 577.200 ;
        RECT 644.100 571.050 645.900 572.850 ;
        RECT 647.700 571.050 648.900 576.300 ;
        RECT 649.950 571.050 651.750 572.850 ;
        RECT 668.100 571.050 669.900 572.850 ;
        RECT 674.250 571.050 676.050 572.850 ;
        RECT 677.700 571.050 678.600 578.400 ;
        RECT 692.100 575.400 693.900 585.000 ;
        RECT 698.700 576.000 700.500 584.400 ;
        RECT 716.700 577.200 718.500 584.400 ;
        RECT 721.800 578.400 723.600 585.000 ;
        RECT 737.700 581.400 739.500 585.000 ;
        RECT 740.700 579.600 742.500 584.400 ;
        RECT 737.400 578.400 742.500 579.600 ;
        RECT 745.200 578.400 747.000 585.000 ;
        RECT 716.700 576.300 720.900 577.200 ;
        RECT 698.700 574.800 702.000 576.000 ;
        RECT 679.950 573.450 684.000 574.050 ;
        RECT 679.950 571.950 684.450 573.450 ;
        RECT 624.150 569.250 630.450 571.050 ;
        RECT 625.950 568.950 630.450 569.250 ;
        RECT 643.950 568.950 646.050 571.050 ;
        RECT 646.950 568.950 649.050 571.050 ;
        RECT 649.950 568.950 652.050 571.050 ;
        RECT 667.950 568.950 670.050 571.050 ;
        RECT 670.950 568.950 673.050 571.050 ;
        RECT 673.950 568.950 676.050 571.050 ;
        RECT 676.950 568.950 679.050 571.050 ;
        RECT 620.550 566.100 622.650 566.400 ;
        RECT 626.550 566.100 628.350 566.250 ;
        RECT 620.550 564.900 628.350 566.100 ;
        RECT 620.550 564.300 622.650 564.900 ;
        RECT 626.550 564.450 628.350 564.900 ;
        RECT 616.950 561.300 621.750 562.200 ;
        RECT 629.250 561.600 630.450 568.950 ;
        RECT 620.550 560.400 621.750 561.300 ;
        RECT 617.850 560.100 619.650 560.400 ;
        RECT 605.250 558.600 607.350 559.500 ;
        RECT 613.950 559.200 619.650 560.100 ;
        RECT 617.850 558.600 619.650 559.200 ;
        RECT 620.550 558.600 623.550 560.400 ;
        RECT 605.550 549.600 607.350 558.600 ;
        RECT 609.450 557.550 611.250 558.300 ;
        RECT 614.250 557.550 616.050 558.300 ;
        RECT 609.450 556.500 616.050 557.550 ;
        RECT 610.350 549.000 612.150 555.600 ;
        RECT 613.350 549.600 615.150 556.500 ;
        RECT 620.550 555.600 622.650 557.700 ;
        RECT 616.350 549.000 618.150 555.600 ;
        RECT 620.850 549.600 622.650 555.600 ;
        RECT 625.650 549.000 627.450 561.600 ;
        RECT 628.650 549.600 630.450 561.600 ;
        RECT 647.700 555.600 648.900 568.950 ;
        RECT 671.250 567.150 673.050 568.950 ;
        RECT 677.700 561.600 678.600 568.950 ;
        RECT 683.550 567.450 684.450 571.950 ;
        RECT 692.100 571.050 693.900 572.850 ;
        RECT 698.100 571.050 699.900 572.850 ;
        RECT 701.100 571.050 702.000 574.800 ;
        RECT 711.000 573.450 715.050 574.050 ;
        RECT 710.550 571.950 715.050 573.450 ;
        RECT 691.950 568.950 694.050 571.050 ;
        RECT 694.950 568.950 697.050 571.050 ;
        RECT 697.950 568.950 700.050 571.050 ;
        RECT 700.950 568.950 703.050 571.050 ;
        RECT 688.950 567.450 691.050 568.050 ;
        RECT 683.550 566.550 691.050 567.450 ;
        RECT 695.100 567.150 696.900 568.950 ;
        RECT 688.950 565.950 691.050 566.550 ;
        RECT 679.950 564.450 682.050 565.050 ;
        RECT 697.950 564.450 700.050 565.050 ;
        RECT 679.950 563.550 700.050 564.450 ;
        RECT 679.950 562.950 682.050 563.550 ;
        RECT 697.950 562.950 700.050 563.550 ;
        RECT 668.100 560.700 675.900 561.600 ;
        RECT 644.100 549.000 645.900 555.600 ;
        RECT 647.100 549.600 648.900 555.600 ;
        RECT 650.100 549.000 651.900 555.600 ;
        RECT 668.100 549.600 669.900 560.700 ;
        RECT 671.100 549.000 672.900 559.800 ;
        RECT 674.100 549.600 675.900 560.700 ;
        RECT 677.100 549.600 678.900 561.600 ;
        RECT 701.100 556.800 702.000 568.950 ;
        RECT 710.550 568.050 711.450 571.950 ;
        RECT 716.100 571.050 717.900 572.850 ;
        RECT 719.700 571.050 720.900 576.300 ;
        RECT 721.950 571.050 723.750 572.850 ;
        RECT 737.400 571.050 738.300 578.400 ;
        RECT 748.950 573.450 751.050 576.900 ;
        RECT 761.100 575.400 762.900 585.000 ;
        RECT 767.700 576.000 769.500 584.400 ;
        RECT 785.100 576.600 786.900 584.400 ;
        RECT 789.600 578.400 791.400 585.000 ;
        RECT 792.600 580.200 794.400 584.400 ;
        RECT 792.600 578.400 795.300 580.200 ;
        RECT 791.700 576.600 793.500 577.500 ;
        RECT 767.700 574.800 771.000 576.000 ;
        RECT 785.100 575.700 793.500 576.600 ;
        RECT 748.950 573.000 756.450 573.450 ;
        RECT 739.950 571.050 741.750 572.850 ;
        RECT 746.100 571.050 747.900 572.850 ;
        RECT 749.550 572.550 756.450 573.000 ;
        RECT 715.950 568.950 718.050 571.050 ;
        RECT 718.950 568.950 721.050 571.050 ;
        RECT 721.950 568.950 724.050 571.050 ;
        RECT 736.950 568.950 739.050 571.050 ;
        RECT 739.950 568.950 742.050 571.050 ;
        RECT 742.950 568.950 745.050 571.050 ;
        RECT 745.950 568.950 748.050 571.050 ;
        RECT 710.550 566.550 715.050 568.050 ;
        RECT 711.000 565.950 715.050 566.550 ;
        RECT 703.950 564.450 706.050 565.050 ;
        RECT 715.950 564.450 718.050 565.050 ;
        RECT 703.950 563.550 718.050 564.450 ;
        RECT 703.950 562.950 706.050 563.550 ;
        RECT 715.950 562.950 718.050 563.550 ;
        RECT 695.400 555.900 702.000 556.800 ;
        RECT 695.400 555.600 696.900 555.900 ;
        RECT 692.100 549.000 693.900 555.600 ;
        RECT 695.100 549.600 696.900 555.600 ;
        RECT 701.100 555.600 702.000 555.900 ;
        RECT 719.700 555.600 720.900 568.950 ;
        RECT 737.400 561.600 738.300 568.950 ;
        RECT 742.950 567.150 744.750 568.950 ;
        RECT 755.550 568.050 756.450 572.550 ;
        RECT 761.100 571.050 762.900 572.850 ;
        RECT 767.100 571.050 768.900 572.850 ;
        RECT 770.100 571.050 771.000 574.800 ;
        RECT 785.250 571.050 787.050 572.850 ;
        RECT 760.950 568.950 763.050 571.050 ;
        RECT 763.950 568.950 766.050 571.050 ;
        RECT 766.950 568.950 769.050 571.050 ;
        RECT 769.950 568.950 772.050 571.050 ;
        RECT 785.100 568.950 787.200 571.050 ;
        RECT 755.550 566.550 760.050 568.050 ;
        RECT 764.100 567.150 765.900 568.950 ;
        RECT 756.000 565.950 760.050 566.550 ;
        RECT 698.100 549.000 699.900 555.000 ;
        RECT 701.100 549.600 702.900 555.600 ;
        RECT 716.100 549.000 717.900 555.600 ;
        RECT 719.100 549.600 720.900 555.600 ;
        RECT 722.100 549.000 723.900 555.600 ;
        RECT 737.100 549.600 738.900 561.600 ;
        RECT 740.100 560.700 747.900 561.600 ;
        RECT 740.100 549.600 741.900 560.700 ;
        RECT 743.100 549.000 744.900 559.800 ;
        RECT 746.100 549.600 747.900 560.700 ;
        RECT 770.100 556.800 771.000 568.950 ;
        RECT 764.400 555.900 771.000 556.800 ;
        RECT 764.400 555.600 765.900 555.900 ;
        RECT 761.100 549.000 762.900 555.600 ;
        RECT 764.100 549.600 765.900 555.600 ;
        RECT 770.100 555.600 771.000 555.900 ;
        RECT 788.100 555.600 789.000 575.700 ;
        RECT 794.400 571.050 795.300 578.400 ;
        RECT 812.100 579.300 813.900 584.400 ;
        RECT 815.100 580.200 816.900 585.000 ;
        RECT 818.100 579.300 819.900 584.400 ;
        RECT 812.100 577.950 819.900 579.300 ;
        RECT 821.100 578.400 822.900 584.400 ;
        RECT 836.100 579.300 837.900 584.400 ;
        RECT 839.100 580.200 840.900 585.000 ;
        RECT 842.100 579.300 843.900 584.400 ;
        RECT 821.100 576.300 822.300 578.400 ;
        RECT 836.100 577.950 843.900 579.300 ;
        RECT 845.100 578.400 846.900 584.400 ;
        RECT 860.100 579.300 861.900 584.400 ;
        RECT 863.100 580.200 864.900 585.000 ;
        RECT 866.100 579.300 867.900 584.400 ;
        RECT 845.100 576.300 846.300 578.400 ;
        RECT 860.100 577.950 867.900 579.300 ;
        RECT 869.100 578.400 870.900 584.400 ;
        RECT 869.100 576.300 870.300 578.400 ;
        RECT 887.700 577.200 889.500 584.400 ;
        RECT 892.800 578.400 894.600 585.000 ;
        RECT 908.100 581.400 909.900 584.400 ;
        RECT 911.100 581.400 912.900 585.000 ;
        RECT 887.700 576.300 891.900 577.200 ;
        RECT 818.700 575.400 822.300 576.300 ;
        RECT 842.700 575.400 846.300 576.300 ;
        RECT 866.700 575.400 870.300 576.300 ;
        RECT 815.100 571.050 816.900 572.850 ;
        RECT 818.700 571.050 819.900 575.400 ;
        RECT 821.100 571.050 822.900 572.850 ;
        RECT 839.100 571.050 840.900 572.850 ;
        RECT 842.700 571.050 843.900 575.400 ;
        RECT 845.100 571.050 846.900 572.850 ;
        RECT 863.100 571.050 864.900 572.850 ;
        RECT 866.700 571.050 867.900 575.400 ;
        RECT 871.950 573.450 876.000 574.050 ;
        RECT 869.100 571.050 870.900 572.850 ;
        RECT 871.950 571.950 876.450 573.450 ;
        RECT 790.500 568.950 792.600 571.050 ;
        RECT 793.800 568.950 795.900 571.050 ;
        RECT 811.950 568.950 814.050 571.050 ;
        RECT 814.950 568.950 817.050 571.050 ;
        RECT 817.950 568.950 820.050 571.050 ;
        RECT 820.950 568.950 823.050 571.050 ;
        RECT 835.950 568.950 838.050 571.050 ;
        RECT 838.950 568.950 841.050 571.050 ;
        RECT 841.950 568.950 844.050 571.050 ;
        RECT 844.950 568.950 847.050 571.050 ;
        RECT 859.950 568.950 862.050 571.050 ;
        RECT 862.950 568.950 865.050 571.050 ;
        RECT 865.950 568.950 868.050 571.050 ;
        RECT 868.950 568.950 871.050 571.050 ;
        RECT 790.200 567.150 792.000 568.950 ;
        RECT 794.400 561.600 795.300 568.950 ;
        RECT 812.100 567.150 813.900 568.950 ;
        RECT 818.700 561.600 819.900 568.950 ;
        RECT 836.100 567.150 837.900 568.950 ;
        RECT 842.700 561.600 843.900 568.950 ;
        RECT 860.100 567.150 861.900 568.950 ;
        RECT 866.700 561.600 867.900 568.950 ;
        RECT 875.550 567.450 876.450 571.950 ;
        RECT 887.100 571.050 888.900 572.850 ;
        RECT 890.700 571.050 891.900 576.300 ;
        RECT 892.950 571.050 894.750 572.850 ;
        RECT 908.700 571.050 909.900 581.400 ;
        RECT 926.100 575.400 927.900 585.000 ;
        RECT 932.700 576.000 934.500 584.400 ;
        RECT 953.700 581.400 955.500 585.000 ;
        RECT 956.700 579.600 958.500 584.400 ;
        RECT 953.400 578.400 958.500 579.600 ;
        RECT 961.200 578.400 963.000 585.000 ;
        RECT 932.700 574.800 936.000 576.000 ;
        RECT 926.100 571.050 927.900 572.850 ;
        RECT 932.100 571.050 933.900 572.850 ;
        RECT 935.100 571.050 936.000 574.800 ;
        RECT 948.000 573.450 952.050 574.050 ;
        RECT 947.550 571.950 952.050 573.450 ;
        RECT 886.950 568.950 889.050 571.050 ;
        RECT 889.950 568.950 892.050 571.050 ;
        RECT 892.950 568.950 895.050 571.050 ;
        RECT 907.950 568.950 910.050 571.050 ;
        RECT 910.950 568.950 913.050 571.050 ;
        RECT 925.950 568.950 928.050 571.050 ;
        RECT 928.950 568.950 931.050 571.050 ;
        RECT 931.950 568.950 934.050 571.050 ;
        RECT 934.950 568.950 937.050 571.050 ;
        RECT 947.550 570.450 948.450 571.950 ;
        RECT 953.400 571.050 954.300 578.400 ;
        RECT 979.500 576.000 981.300 584.400 ;
        RECT 978.000 574.800 981.300 576.000 ;
        RECT 986.100 575.400 987.900 585.000 ;
        RECT 1001.100 575.400 1002.900 585.000 ;
        RECT 1007.700 576.000 1009.500 584.400 ;
        RECT 1007.700 574.800 1011.000 576.000 ;
        RECT 955.950 571.050 957.750 572.850 ;
        RECT 962.100 571.050 963.900 572.850 ;
        RECT 978.000 571.050 978.900 574.800 ;
        RECT 988.950 573.450 993.000 574.050 ;
        RECT 996.000 573.450 1000.050 574.050 ;
        RECT 980.100 571.050 981.900 572.850 ;
        RECT 986.100 571.050 987.900 572.850 ;
        RECT 988.950 571.950 993.450 573.450 ;
        RECT 941.550 569.550 948.450 570.450 ;
        RECT 883.950 567.450 886.050 568.050 ;
        RECT 875.550 566.550 886.050 567.450 ;
        RECT 883.950 565.950 886.050 566.550 ;
        RECT 767.100 549.000 768.900 555.000 ;
        RECT 770.100 549.600 771.900 555.600 ;
        RECT 785.100 549.000 786.900 555.600 ;
        RECT 788.100 549.600 789.900 555.600 ;
        RECT 791.100 549.000 792.900 561.000 ;
        RECT 794.100 549.600 795.900 561.600 ;
        RECT 812.400 549.000 814.200 561.600 ;
        RECT 817.500 560.100 819.900 561.600 ;
        RECT 817.500 549.600 819.300 560.100 ;
        RECT 820.200 557.100 822.000 558.900 ;
        RECT 820.500 549.000 822.300 555.600 ;
        RECT 836.400 549.000 838.200 561.600 ;
        RECT 841.500 560.100 843.900 561.600 ;
        RECT 841.500 549.600 843.300 560.100 ;
        RECT 844.200 557.100 846.000 558.900 ;
        RECT 844.500 549.000 846.300 555.600 ;
        RECT 860.400 549.000 862.200 561.600 ;
        RECT 865.500 560.100 867.900 561.600 ;
        RECT 865.500 549.600 867.300 560.100 ;
        RECT 868.200 557.100 870.000 558.900 ;
        RECT 890.700 555.600 891.900 568.950 ;
        RECT 908.700 555.600 909.900 568.950 ;
        RECT 911.100 567.150 912.900 568.950 ;
        RECT 929.100 567.150 930.900 568.950 ;
        RECT 919.950 564.450 922.050 565.050 ;
        RECT 931.950 564.450 934.050 565.050 ;
        RECT 919.950 563.550 934.050 564.450 ;
        RECT 919.950 562.950 922.050 563.550 ;
        RECT 931.950 562.950 934.050 563.550 ;
        RECT 935.100 556.800 936.000 568.950 ;
        RECT 941.550 568.050 942.450 569.550 ;
        RECT 952.950 568.950 955.050 571.050 ;
        RECT 955.950 568.950 958.050 571.050 ;
        RECT 958.950 568.950 961.050 571.050 ;
        RECT 961.950 568.950 964.050 571.050 ;
        RECT 976.950 568.950 979.050 571.050 ;
        RECT 979.950 568.950 982.050 571.050 ;
        RECT 982.950 568.950 985.050 571.050 ;
        RECT 985.950 568.950 988.050 571.050 ;
        RECT 937.950 566.550 942.450 568.050 ;
        RECT 943.950 567.450 946.050 568.050 ;
        RECT 949.950 567.450 952.050 568.050 ;
        RECT 943.950 566.550 952.050 567.450 ;
        RECT 937.950 565.950 942.000 566.550 ;
        RECT 943.950 565.950 946.050 566.550 ;
        RECT 949.950 565.950 952.050 566.550 ;
        RECT 953.400 561.600 954.300 568.950 ;
        RECT 958.950 567.150 960.750 568.950 ;
        RECT 929.400 555.900 936.000 556.800 ;
        RECT 929.400 555.600 930.900 555.900 ;
        RECT 868.500 549.000 870.300 555.600 ;
        RECT 887.100 549.000 888.900 555.600 ;
        RECT 890.100 549.600 891.900 555.600 ;
        RECT 893.100 549.000 894.900 555.600 ;
        RECT 908.100 549.600 909.900 555.600 ;
        RECT 911.100 549.000 912.900 555.600 ;
        RECT 926.100 549.000 927.900 555.600 ;
        RECT 929.100 549.600 930.900 555.600 ;
        RECT 935.100 555.600 936.000 555.900 ;
        RECT 932.100 549.000 933.900 555.000 ;
        RECT 935.100 549.600 936.900 555.600 ;
        RECT 953.100 549.600 954.900 561.600 ;
        RECT 956.100 560.700 963.900 561.600 ;
        RECT 956.100 549.600 957.900 560.700 ;
        RECT 959.100 549.000 960.900 559.800 ;
        RECT 962.100 549.600 963.900 560.700 ;
        RECT 978.000 556.800 978.900 568.950 ;
        RECT 983.100 567.150 984.900 568.950 ;
        RECT 992.550 565.050 993.450 571.950 ;
        RECT 995.550 571.950 1000.050 573.450 ;
        RECT 991.950 562.950 994.050 565.050 ;
        RECT 995.550 564.450 996.450 571.950 ;
        RECT 1001.100 571.050 1002.900 572.850 ;
        RECT 1007.100 571.050 1008.900 572.850 ;
        RECT 1010.100 571.050 1011.000 574.800 ;
        RECT 1000.950 568.950 1003.050 571.050 ;
        RECT 1003.950 568.950 1006.050 571.050 ;
        RECT 1006.950 568.950 1009.050 571.050 ;
        RECT 1009.950 568.950 1012.050 571.050 ;
        RECT 1004.100 567.150 1005.900 568.950 ;
        RECT 1000.950 564.450 1003.050 565.050 ;
        RECT 995.550 563.550 1003.050 564.450 ;
        RECT 1000.950 562.950 1003.050 563.550 ;
        RECT 1010.100 556.800 1011.000 568.950 ;
        RECT 978.000 555.900 984.600 556.800 ;
        RECT 978.000 555.600 978.900 555.900 ;
        RECT 977.100 549.600 978.900 555.600 ;
        RECT 983.100 555.600 984.600 555.900 ;
        RECT 1004.400 555.900 1011.000 556.800 ;
        RECT 1004.400 555.600 1005.900 555.900 ;
        RECT 980.100 549.000 981.900 555.000 ;
        RECT 983.100 549.600 984.900 555.600 ;
        RECT 986.100 549.000 987.900 555.600 ;
        RECT 1001.100 549.000 1002.900 555.600 ;
        RECT 1004.100 549.600 1005.900 555.600 ;
        RECT 1010.100 555.600 1011.000 555.900 ;
        RECT 1007.100 549.000 1008.900 555.000 ;
        RECT 1010.100 549.600 1011.900 555.600 ;
        RECT 14.100 533.400 15.900 545.400 ;
        RECT 17.100 535.200 18.900 546.000 ;
        RECT 20.100 539.400 21.900 545.400 ;
        RECT 35.100 539.400 36.900 546.000 ;
        RECT 38.100 539.400 39.900 545.400 ;
        RECT 53.100 539.400 54.900 546.000 ;
        RECT 56.100 539.400 57.900 545.400 ;
        RECT 59.100 539.400 60.900 546.000 ;
        RECT 74.700 539.400 76.500 546.000 ;
        RECT 14.100 526.050 15.300 533.400 ;
        RECT 20.700 532.500 21.900 539.400 ;
        RECT 16.200 531.600 21.900 532.500 ;
        RECT 16.200 530.700 18.000 531.600 ;
        RECT 14.100 523.950 16.200 526.050 ;
        RECT 14.100 516.600 15.300 523.950 ;
        RECT 17.100 519.300 18.000 530.700 ;
        RECT 19.800 526.050 21.600 527.850 ;
        RECT 35.100 526.050 36.900 527.850 ;
        RECT 38.100 526.050 39.300 539.400 ;
        RECT 56.700 526.050 57.900 539.400 ;
        RECT 75.000 536.100 76.800 537.900 ;
        RECT 77.700 534.900 79.500 545.400 ;
        RECT 77.100 533.400 79.500 534.900 ;
        RECT 82.800 533.400 84.600 546.000 ;
        RECT 98.400 533.400 100.200 546.000 ;
        RECT 103.500 534.900 105.300 545.400 ;
        RECT 106.500 539.400 108.300 546.000 ;
        RECT 125.700 539.400 127.500 546.000 ;
        RECT 106.200 536.100 108.000 537.900 ;
        RECT 126.000 536.100 127.800 537.900 ;
        RECT 128.700 534.900 130.500 545.400 ;
        RECT 103.500 533.400 105.900 534.900 ;
        RECT 77.100 526.050 78.300 533.400 ;
        RECT 82.950 531.450 85.050 532.050 ;
        RECT 88.950 531.450 91.050 532.050 ;
        RECT 82.950 530.550 91.050 531.450 ;
        RECT 82.950 529.950 85.050 530.550 ;
        RECT 88.950 529.950 91.050 530.550 ;
        RECT 83.100 526.050 84.900 527.850 ;
        RECT 98.100 526.050 99.900 527.850 ;
        RECT 104.700 526.050 105.900 533.400 ;
        RECT 128.100 533.400 130.500 534.900 ;
        RECT 133.800 533.400 135.600 546.000 ;
        RECT 149.100 539.400 150.900 546.000 ;
        RECT 152.100 539.400 153.900 545.400 ;
        RECT 167.100 539.400 168.900 545.400 ;
        RECT 170.100 540.000 171.900 546.000 ;
        RECT 128.100 526.050 129.300 533.400 ;
        RECT 134.100 526.050 135.900 527.850 ;
        RECT 149.100 526.050 150.900 527.850 ;
        RECT 152.100 526.050 153.300 539.400 ;
        RECT 168.000 539.100 168.900 539.400 ;
        RECT 173.100 539.400 174.900 545.400 ;
        RECT 176.100 539.400 177.900 546.000 ;
        RECT 173.100 539.100 174.600 539.400 ;
        RECT 168.000 538.200 174.600 539.100 ;
        RECT 159.000 528.450 163.050 529.050 ;
        RECT 158.550 526.950 163.050 528.450 ;
        RECT 19.500 523.950 21.600 526.050 ;
        RECT 34.950 523.950 37.050 526.050 ;
        RECT 37.950 523.950 40.050 526.050 ;
        RECT 52.950 523.950 55.050 526.050 ;
        RECT 55.950 523.950 58.050 526.050 ;
        RECT 58.950 523.950 61.050 526.050 ;
        RECT 16.200 518.400 18.000 519.300 ;
        RECT 16.200 517.500 21.900 518.400 ;
        RECT 14.100 510.600 15.900 516.600 ;
        RECT 17.100 510.000 18.900 516.600 ;
        RECT 20.700 513.600 21.900 517.500 ;
        RECT 38.100 513.600 39.300 523.950 ;
        RECT 53.100 522.150 54.900 523.950 ;
        RECT 56.700 518.700 57.900 523.950 ;
        RECT 58.950 522.150 60.750 523.950 ;
        RECT 64.950 523.050 67.050 526.050 ;
        RECT 73.950 523.950 76.050 526.050 ;
        RECT 76.950 523.950 79.050 526.050 ;
        RECT 79.950 523.950 82.050 526.050 ;
        RECT 82.950 523.950 85.050 526.050 ;
        RECT 97.950 523.950 100.050 526.050 ;
        RECT 100.950 523.950 103.050 526.050 ;
        RECT 103.950 523.950 106.050 526.050 ;
        RECT 106.950 523.950 109.050 526.050 ;
        RECT 124.950 523.950 127.050 526.050 ;
        RECT 127.950 523.950 130.050 526.050 ;
        RECT 130.950 523.950 133.050 526.050 ;
        RECT 133.950 523.950 136.050 526.050 ;
        RECT 148.950 523.950 151.050 526.050 ;
        RECT 151.950 523.950 154.050 526.050 ;
        RECT 61.950 522.000 67.050 523.050 ;
        RECT 74.100 522.150 75.900 523.950 ;
        RECT 61.950 521.550 66.450 522.000 ;
        RECT 61.950 520.950 66.000 521.550 ;
        RECT 77.100 519.600 78.300 523.950 ;
        RECT 80.100 522.150 81.900 523.950 ;
        RECT 101.100 522.150 102.900 523.950 ;
        RECT 53.700 517.800 57.900 518.700 ;
        RECT 74.700 518.700 78.300 519.600 ;
        RECT 104.700 519.600 105.900 523.950 ;
        RECT 107.100 522.150 108.900 523.950 ;
        RECT 125.100 522.150 126.900 523.950 ;
        RECT 128.100 519.600 129.300 523.950 ;
        RECT 131.100 522.150 132.900 523.950 ;
        RECT 104.700 518.700 108.300 519.600 ;
        RECT 20.100 510.600 21.900 513.600 ;
        RECT 35.100 510.000 36.900 513.600 ;
        RECT 38.100 510.600 39.900 513.600 ;
        RECT 53.700 510.600 55.500 517.800 ;
        RECT 74.700 516.600 75.900 518.700 ;
        RECT 58.800 510.000 60.600 516.600 ;
        RECT 74.100 510.600 75.900 516.600 ;
        RECT 77.100 515.700 84.900 517.050 ;
        RECT 77.100 510.600 78.900 515.700 ;
        RECT 80.100 510.000 81.900 514.800 ;
        RECT 83.100 510.600 84.900 515.700 ;
        RECT 98.100 515.700 105.900 517.050 ;
        RECT 98.100 510.600 99.900 515.700 ;
        RECT 101.100 510.000 102.900 514.800 ;
        RECT 104.100 510.600 105.900 515.700 ;
        RECT 107.100 516.600 108.300 518.700 ;
        RECT 125.700 518.700 129.300 519.600 ;
        RECT 125.700 516.600 126.900 518.700 ;
        RECT 107.100 510.600 108.900 516.600 ;
        RECT 125.100 510.600 126.900 516.600 ;
        RECT 128.100 515.700 135.900 517.050 ;
        RECT 128.100 510.600 129.900 515.700 ;
        RECT 131.100 510.000 132.900 514.800 ;
        RECT 134.100 510.600 135.900 515.700 ;
        RECT 152.100 513.600 153.300 523.950 ;
        RECT 158.550 523.050 159.450 526.950 ;
        RECT 168.000 526.050 168.900 538.200 ;
        RECT 180.150 535.200 181.950 545.400 ;
        RECT 179.550 533.400 181.950 535.200 ;
        RECT 183.150 533.400 184.950 546.000 ;
        RECT 188.550 536.400 190.350 545.400 ;
        RECT 193.350 539.400 195.150 546.000 ;
        RECT 196.350 538.500 198.150 545.400 ;
        RECT 199.350 539.400 201.150 546.000 ;
        RECT 203.850 539.400 205.650 545.400 ;
        RECT 192.450 537.450 199.050 538.500 ;
        RECT 192.450 536.700 194.250 537.450 ;
        RECT 197.250 536.700 199.050 537.450 ;
        RECT 203.550 537.300 205.650 539.400 ;
        RECT 188.250 535.500 190.350 536.400 ;
        RECT 200.850 535.800 202.650 536.400 ;
        RECT 188.250 534.300 196.050 535.500 ;
        RECT 194.250 533.700 196.050 534.300 ;
        RECT 196.950 534.900 202.650 535.800 ;
        RECT 179.550 532.500 180.450 533.400 ;
        RECT 196.950 532.800 197.850 534.900 ;
        RECT 200.850 534.600 202.650 534.900 ;
        RECT 203.550 534.600 206.550 536.400 ;
        RECT 203.550 533.700 204.750 534.600 ;
        RECT 189.450 532.500 197.850 532.800 ;
        RECT 179.550 531.900 197.850 532.500 ;
        RECT 199.950 532.800 204.750 533.700 ;
        RECT 208.650 533.400 210.450 546.000 ;
        RECT 211.650 533.400 213.450 545.400 ;
        RECT 230.400 533.400 232.200 546.000 ;
        RECT 235.500 534.900 237.300 545.400 ;
        RECT 238.500 539.400 240.300 546.000 ;
        RECT 254.100 539.400 255.900 546.000 ;
        RECT 257.100 539.400 258.900 545.400 ;
        RECT 260.100 539.400 261.900 546.000 ;
        RECT 238.200 536.100 240.000 537.900 ;
        RECT 235.500 533.400 237.900 534.900 ;
        RECT 179.550 531.300 191.250 531.900 ;
        RECT 173.100 526.050 174.900 527.850 ;
        RECT 166.950 523.950 169.050 526.050 ;
        RECT 169.950 523.950 172.050 526.050 ;
        RECT 172.950 523.950 175.050 526.050 ;
        RECT 175.950 523.950 178.050 526.050 ;
        RECT 154.950 521.550 159.450 523.050 ;
        RECT 154.950 520.950 159.000 521.550 ;
        RECT 168.000 520.200 168.900 523.950 ;
        RECT 170.100 522.150 171.900 523.950 ;
        RECT 176.100 522.150 177.900 523.950 ;
        RECT 157.950 519.450 160.050 520.050 ;
        RECT 163.950 519.450 166.050 520.050 ;
        RECT 157.950 518.550 166.050 519.450 ;
        RECT 168.000 519.000 171.300 520.200 ;
        RECT 157.950 517.950 160.050 518.550 ;
        RECT 163.950 517.950 166.050 518.550 ;
        RECT 149.100 510.000 150.900 513.600 ;
        RECT 152.100 510.600 153.900 513.600 ;
        RECT 169.500 510.600 171.300 519.000 ;
        RECT 176.100 510.000 177.900 519.600 ;
        RECT 179.550 516.600 180.450 531.300 ;
        RECT 189.450 531.000 191.250 531.300 ;
        RECT 181.950 523.950 184.050 526.050 ;
        RECT 191.100 524.400 193.200 526.050 ;
        RECT 181.950 521.400 183.750 523.950 ;
        RECT 185.100 523.200 193.200 524.400 ;
        RECT 185.100 522.600 186.900 523.200 ;
        RECT 188.100 521.400 189.900 522.000 ;
        RECT 181.950 520.200 189.900 521.400 ;
        RECT 199.950 520.200 200.850 532.800 ;
        RECT 203.550 530.100 205.650 530.700 ;
        RECT 209.550 530.100 211.350 530.550 ;
        RECT 203.550 528.900 211.350 530.100 ;
        RECT 203.550 528.600 205.650 528.900 ;
        RECT 209.550 528.750 211.350 528.900 ;
        RECT 212.250 526.050 213.450 533.400 ;
        RECT 230.100 526.050 231.900 527.850 ;
        RECT 236.700 526.050 237.900 533.400 ;
        RECT 238.950 531.450 241.050 532.050 ;
        RECT 244.950 531.450 247.050 532.050 ;
        RECT 238.950 530.550 247.050 531.450 ;
        RECT 238.950 529.950 241.050 530.550 ;
        RECT 244.950 529.950 247.050 530.550 ;
        RECT 257.700 526.050 258.900 539.400 ;
        RECT 275.400 533.400 277.200 546.000 ;
        RECT 280.500 534.900 282.300 545.400 ;
        RECT 283.500 539.400 285.300 546.000 ;
        RECT 299.100 539.400 300.900 545.400 ;
        RECT 302.100 539.400 303.900 546.000 ;
        RECT 283.200 536.100 285.000 537.900 ;
        RECT 280.500 533.400 282.900 534.900 ;
        RECT 275.100 526.050 276.900 527.850 ;
        RECT 281.700 526.050 282.900 533.400 ;
        RECT 299.700 526.050 300.900 539.400 ;
        RECT 317.100 533.400 318.900 546.000 ;
        RECT 320.100 532.500 321.900 545.400 ;
        RECT 323.100 533.400 324.900 546.000 ;
        RECT 326.100 532.500 327.900 545.400 ;
        RECT 329.100 533.400 330.900 546.000 ;
        RECT 332.100 532.500 333.900 545.400 ;
        RECT 335.100 533.400 336.900 546.000 ;
        RECT 338.100 532.500 339.900 545.400 ;
        RECT 341.100 533.400 342.900 546.000 ;
        RECT 359.100 539.400 360.900 546.000 ;
        RECT 362.100 539.400 363.900 545.400 ;
        RECT 365.100 539.400 366.900 546.000 ;
        RECT 383.100 539.400 384.900 546.000 ;
        RECT 386.100 539.400 387.900 545.400 ;
        RECT 389.100 539.400 390.900 546.000 ;
        RECT 404.100 539.400 405.900 545.400 ;
        RECT 407.100 539.400 408.900 546.000 ;
        RECT 320.100 531.300 324.000 532.500 ;
        RECT 326.100 531.300 330.000 532.500 ;
        RECT 332.100 531.300 336.000 532.500 ;
        RECT 338.100 531.300 340.950 532.500 ;
        RECT 302.100 526.050 303.900 527.850 ;
        RECT 208.950 525.750 213.450 526.050 ;
        RECT 207.150 523.950 213.450 525.750 ;
        RECT 229.950 523.950 232.050 526.050 ;
        RECT 232.950 523.950 235.050 526.050 ;
        RECT 235.950 523.950 238.050 526.050 ;
        RECT 238.950 523.950 241.050 526.050 ;
        RECT 253.950 523.950 256.050 526.050 ;
        RECT 256.950 523.950 259.050 526.050 ;
        RECT 259.950 523.950 262.050 526.050 ;
        RECT 274.950 523.950 277.050 526.050 ;
        RECT 277.950 523.950 280.050 526.050 ;
        RECT 280.950 523.950 283.050 526.050 ;
        RECT 283.950 523.950 286.050 526.050 ;
        RECT 298.950 523.950 301.050 526.050 ;
        RECT 301.950 523.950 304.050 526.050 ;
        RECT 319.800 523.950 321.900 526.050 ;
        RECT 188.850 519.000 200.850 520.200 ;
        RECT 188.850 517.200 189.900 519.000 ;
        RECT 199.050 518.400 200.850 519.000 ;
        RECT 179.550 514.800 181.950 516.600 ;
        RECT 180.150 510.600 181.950 514.800 ;
        RECT 183.150 510.000 184.950 516.600 ;
        RECT 185.850 514.200 187.950 515.700 ;
        RECT 188.850 515.400 190.650 517.200 ;
        RECT 212.250 516.600 213.450 523.950 ;
        RECT 233.100 522.150 234.900 523.950 ;
        RECT 236.700 519.600 237.900 523.950 ;
        RECT 239.100 522.150 240.900 523.950 ;
        RECT 254.100 522.150 255.900 523.950 ;
        RECT 236.700 518.700 240.300 519.600 ;
        RECT 257.700 518.700 258.900 523.950 ;
        RECT 259.950 522.150 261.750 523.950 ;
        RECT 278.100 522.150 279.900 523.950 ;
        RECT 281.700 519.600 282.900 523.950 ;
        RECT 284.100 522.150 285.900 523.950 ;
        RECT 281.700 518.700 285.300 519.600 ;
        RECT 191.850 515.550 193.650 516.300 ;
        RECT 191.850 514.500 196.800 515.550 ;
        RECT 185.850 513.600 189.750 514.200 ;
        RECT 195.750 513.600 196.800 514.500 ;
        RECT 203.250 513.600 205.650 515.700 ;
        RECT 186.150 512.700 189.750 513.600 ;
        RECT 187.950 510.600 189.750 512.700 ;
        RECT 192.450 510.000 194.250 513.600 ;
        RECT 195.750 510.600 197.550 513.600 ;
        RECT 198.750 510.000 200.550 513.600 ;
        RECT 203.250 510.600 205.050 513.600 ;
        RECT 208.350 510.000 210.150 516.600 ;
        RECT 211.650 510.600 213.450 516.600 ;
        RECT 230.100 515.700 237.900 517.050 ;
        RECT 230.100 510.600 231.900 515.700 ;
        RECT 233.100 510.000 234.900 514.800 ;
        RECT 236.100 510.600 237.900 515.700 ;
        RECT 239.100 516.600 240.300 518.700 ;
        RECT 254.700 517.800 258.900 518.700 ;
        RECT 239.100 510.600 240.900 516.600 ;
        RECT 254.700 510.600 256.500 517.800 ;
        RECT 259.800 510.000 261.600 516.600 ;
        RECT 275.100 515.700 282.900 517.050 ;
        RECT 275.100 510.600 276.900 515.700 ;
        RECT 278.100 510.000 279.900 514.800 ;
        RECT 281.100 510.600 282.900 515.700 ;
        RECT 284.100 516.600 285.300 518.700 ;
        RECT 284.100 510.600 285.900 516.600 ;
        RECT 299.700 513.600 300.900 523.950 ;
        RECT 319.800 522.150 321.600 523.950 ;
        RECT 322.800 520.800 324.000 531.300 ;
        RECT 325.200 520.800 327.000 521.400 ;
        RECT 322.800 519.600 327.000 520.800 ;
        RECT 328.800 520.800 330.000 531.300 ;
        RECT 331.200 520.800 333.000 521.400 ;
        RECT 328.800 519.600 333.000 520.800 ;
        RECT 334.800 520.800 336.000 531.300 ;
        RECT 339.900 526.050 340.950 531.300 ;
        RECT 362.100 526.050 363.300 539.400 ;
        RECT 386.100 526.050 387.300 539.400 ;
        RECT 404.700 526.050 405.900 539.400 ;
        RECT 422.400 533.400 424.200 546.000 ;
        RECT 427.500 534.900 429.300 545.400 ;
        RECT 430.500 539.400 432.300 546.000 ;
        RECT 430.200 536.100 432.000 537.900 ;
        RECT 427.500 533.400 429.900 534.900 ;
        RECT 417.000 528.450 421.050 529.050 ;
        RECT 407.100 526.050 408.900 527.850 ;
        RECT 416.550 526.950 421.050 528.450 ;
        RECT 337.800 523.950 340.950 526.050 ;
        RECT 358.950 523.950 361.050 526.050 ;
        RECT 361.950 523.950 364.050 526.050 ;
        RECT 364.950 523.950 367.050 526.050 ;
        RECT 382.950 523.950 385.050 526.050 ;
        RECT 385.950 523.950 388.050 526.050 ;
        RECT 388.950 523.950 391.050 526.050 ;
        RECT 403.950 523.950 406.050 526.050 ;
        RECT 406.950 523.950 409.050 526.050 ;
        RECT 337.200 520.800 339.000 521.400 ;
        RECT 334.800 519.600 339.000 520.800 ;
        RECT 322.800 518.700 324.000 519.600 ;
        RECT 328.800 518.700 330.000 519.600 ;
        RECT 334.800 518.700 336.000 519.600 ;
        RECT 339.900 518.700 340.950 523.950 ;
        RECT 359.250 522.150 361.050 523.950 ;
        RECT 320.100 517.500 324.000 518.700 ;
        RECT 326.100 517.500 330.000 518.700 ;
        RECT 332.100 517.500 336.000 518.700 ;
        RECT 338.100 517.500 340.950 518.700 ;
        RECT 362.100 518.700 363.300 523.950 ;
        RECT 365.100 522.150 366.900 523.950 ;
        RECT 383.250 522.150 385.050 523.950 ;
        RECT 386.100 518.700 387.300 523.950 ;
        RECT 389.100 522.150 390.900 523.950 ;
        RECT 362.100 517.800 366.300 518.700 ;
        RECT 386.100 517.800 390.300 518.700 ;
        RECT 299.100 510.600 300.900 513.600 ;
        RECT 302.100 510.000 303.900 513.600 ;
        RECT 317.100 510.000 318.900 516.600 ;
        RECT 320.100 510.600 321.900 517.500 ;
        RECT 323.100 510.000 324.900 516.600 ;
        RECT 326.100 510.600 327.900 517.500 ;
        RECT 329.100 510.000 330.900 516.600 ;
        RECT 332.100 510.600 333.900 517.500 ;
        RECT 335.100 510.000 336.900 516.600 ;
        RECT 338.100 510.600 339.900 517.500 ;
        RECT 341.100 510.000 342.900 516.600 ;
        RECT 359.400 510.000 361.200 516.600 ;
        RECT 364.500 510.600 366.300 517.800 ;
        RECT 383.400 510.000 385.200 516.600 ;
        RECT 388.500 510.600 390.300 517.800 ;
        RECT 404.700 513.600 405.900 523.950 ;
        RECT 416.550 523.050 417.450 526.950 ;
        RECT 422.100 526.050 423.900 527.850 ;
        RECT 428.700 526.050 429.900 533.400 ;
        RECT 434.550 533.400 436.350 545.400 ;
        RECT 437.550 533.400 439.350 546.000 ;
        RECT 442.350 539.400 444.150 545.400 ;
        RECT 446.850 539.400 448.650 546.000 ;
        RECT 442.350 537.300 444.450 539.400 ;
        RECT 449.850 538.500 451.650 545.400 ;
        RECT 452.850 539.400 454.650 546.000 ;
        RECT 448.950 537.450 455.550 538.500 ;
        RECT 448.950 536.700 450.750 537.450 ;
        RECT 453.750 536.700 455.550 537.450 ;
        RECT 457.650 536.400 459.450 545.400 ;
        RECT 441.450 534.600 444.450 536.400 ;
        RECT 445.350 535.800 447.150 536.400 ;
        RECT 445.350 534.900 451.050 535.800 ;
        RECT 457.650 535.500 459.750 536.400 ;
        RECT 445.350 534.600 447.150 534.900 ;
        RECT 443.250 533.700 444.450 534.600 ;
        RECT 434.550 526.050 435.750 533.400 ;
        RECT 443.250 532.800 448.050 533.700 ;
        RECT 436.650 530.100 438.450 530.550 ;
        RECT 442.350 530.100 444.450 530.700 ;
        RECT 436.650 528.900 444.450 530.100 ;
        RECT 436.650 528.750 438.450 528.900 ;
        RECT 442.350 528.600 444.450 528.900 ;
        RECT 421.950 523.950 424.050 526.050 ;
        RECT 424.950 523.950 427.050 526.050 ;
        RECT 427.950 523.950 430.050 526.050 ;
        RECT 430.950 523.950 433.050 526.050 ;
        RECT 434.550 525.750 439.050 526.050 ;
        RECT 434.550 523.950 440.850 525.750 ;
        RECT 416.550 521.550 421.050 523.050 ;
        RECT 425.100 522.150 426.900 523.950 ;
        RECT 417.000 520.950 421.050 521.550 ;
        RECT 428.700 519.600 429.900 523.950 ;
        RECT 431.100 522.150 432.900 523.950 ;
        RECT 428.700 518.700 432.300 519.600 ;
        RECT 422.100 515.700 429.900 517.050 ;
        RECT 404.100 510.600 405.900 513.600 ;
        RECT 407.100 510.000 408.900 513.600 ;
        RECT 422.100 510.600 423.900 515.700 ;
        RECT 425.100 510.000 426.900 514.800 ;
        RECT 428.100 510.600 429.900 515.700 ;
        RECT 431.100 516.600 432.300 518.700 ;
        RECT 434.550 516.600 435.750 523.950 ;
        RECT 447.150 520.200 448.050 532.800 ;
        RECT 450.150 532.800 451.050 534.900 ;
        RECT 451.950 534.300 459.750 535.500 ;
        RECT 451.950 533.700 453.750 534.300 ;
        RECT 463.050 533.400 464.850 546.000 ;
        RECT 466.050 535.200 467.850 545.400 ;
        RECT 466.050 533.400 468.450 535.200 ;
        RECT 482.400 533.400 484.200 546.000 ;
        RECT 487.500 534.900 489.300 545.400 ;
        RECT 490.500 539.400 492.300 546.000 ;
        RECT 506.100 539.400 507.900 546.000 ;
        RECT 509.100 539.400 510.900 545.400 ;
        RECT 512.100 539.400 513.900 546.000 ;
        RECT 527.100 539.400 528.900 545.400 ;
        RECT 530.100 539.400 531.900 546.000 ;
        RECT 490.200 536.100 492.000 537.900 ;
        RECT 493.950 537.450 496.050 538.050 ;
        RECT 499.950 537.450 502.050 538.050 ;
        RECT 493.950 536.550 502.050 537.450 ;
        RECT 493.950 535.950 496.050 536.550 ;
        RECT 499.950 535.950 502.050 536.550 ;
        RECT 487.500 533.400 489.900 534.900 ;
        RECT 450.150 532.500 458.550 532.800 ;
        RECT 467.550 532.500 468.450 533.400 ;
        RECT 450.150 531.900 468.450 532.500 ;
        RECT 456.750 531.300 468.450 531.900 ;
        RECT 456.750 531.000 458.550 531.300 ;
        RECT 454.800 524.400 456.900 526.050 ;
        RECT 454.800 523.200 462.900 524.400 ;
        RECT 463.950 523.950 466.050 526.050 ;
        RECT 461.100 522.600 462.900 523.200 ;
        RECT 458.100 521.400 459.900 522.000 ;
        RECT 464.250 521.400 466.050 523.950 ;
        RECT 458.100 520.200 466.050 521.400 ;
        RECT 447.150 519.000 459.150 520.200 ;
        RECT 447.150 518.400 448.950 519.000 ;
        RECT 458.100 517.200 459.150 519.000 ;
        RECT 431.100 510.600 432.900 516.600 ;
        RECT 434.550 510.600 436.350 516.600 ;
        RECT 437.850 510.000 439.650 516.600 ;
        RECT 442.350 513.600 444.750 515.700 ;
        RECT 454.350 515.550 456.150 516.300 ;
        RECT 451.200 514.500 456.150 515.550 ;
        RECT 457.350 515.400 459.150 517.200 ;
        RECT 467.550 516.600 468.450 531.300 ;
        RECT 482.100 526.050 483.900 527.850 ;
        RECT 488.700 526.050 489.900 533.400 ;
        RECT 509.100 526.050 510.300 539.400 ;
        RECT 527.700 526.050 528.900 539.400 ;
        RECT 533.550 533.400 535.350 545.400 ;
        RECT 536.550 533.400 538.350 546.000 ;
        RECT 541.350 539.400 543.150 545.400 ;
        RECT 545.850 539.400 547.650 546.000 ;
        RECT 541.350 537.300 543.450 539.400 ;
        RECT 548.850 538.500 550.650 545.400 ;
        RECT 551.850 539.400 553.650 546.000 ;
        RECT 547.950 537.450 554.550 538.500 ;
        RECT 547.950 536.700 549.750 537.450 ;
        RECT 552.750 536.700 554.550 537.450 ;
        RECT 556.650 536.400 558.450 545.400 ;
        RECT 540.450 534.600 543.450 536.400 ;
        RECT 544.350 535.800 546.150 536.400 ;
        RECT 544.350 534.900 550.050 535.800 ;
        RECT 556.650 535.500 558.750 536.400 ;
        RECT 544.350 534.600 546.150 534.900 ;
        RECT 542.250 533.700 543.450 534.600 ;
        RECT 530.100 526.050 531.900 527.850 ;
        RECT 533.550 526.050 534.750 533.400 ;
        RECT 542.250 532.800 547.050 533.700 ;
        RECT 535.650 530.100 537.450 530.550 ;
        RECT 541.350 530.100 543.450 530.700 ;
        RECT 535.650 528.900 543.450 530.100 ;
        RECT 535.650 528.750 537.450 528.900 ;
        RECT 541.350 528.600 543.450 528.900 ;
        RECT 481.950 523.950 484.050 526.050 ;
        RECT 484.950 523.950 487.050 526.050 ;
        RECT 487.950 523.950 490.050 526.050 ;
        RECT 490.950 523.950 493.050 526.050 ;
        RECT 505.950 523.950 508.050 526.050 ;
        RECT 508.950 523.950 511.050 526.050 ;
        RECT 511.950 523.950 514.050 526.050 ;
        RECT 526.950 523.950 529.050 526.050 ;
        RECT 529.950 523.950 532.050 526.050 ;
        RECT 533.550 525.750 538.050 526.050 ;
        RECT 533.550 523.950 539.850 525.750 ;
        RECT 485.100 522.150 486.900 523.950 ;
        RECT 488.700 519.600 489.900 523.950 ;
        RECT 491.100 522.150 492.900 523.950 ;
        RECT 506.250 522.150 508.050 523.950 ;
        RECT 488.700 518.700 492.300 519.600 ;
        RECT 451.200 513.600 452.250 514.500 ;
        RECT 460.050 514.200 462.150 515.700 ;
        RECT 458.250 513.600 462.150 514.200 ;
        RECT 442.950 510.600 444.750 513.600 ;
        RECT 447.450 510.000 449.250 513.600 ;
        RECT 450.450 510.600 452.250 513.600 ;
        RECT 453.750 510.000 455.550 513.600 ;
        RECT 458.250 512.700 461.850 513.600 ;
        RECT 458.250 510.600 460.050 512.700 ;
        RECT 463.050 510.000 464.850 516.600 ;
        RECT 466.050 514.800 468.450 516.600 ;
        RECT 482.100 515.700 489.900 517.050 ;
        RECT 466.050 510.600 467.850 514.800 ;
        RECT 482.100 510.600 483.900 515.700 ;
        RECT 485.100 510.000 486.900 514.800 ;
        RECT 488.100 510.600 489.900 515.700 ;
        RECT 491.100 516.600 492.300 518.700 ;
        RECT 496.950 519.450 499.050 520.050 ;
        RECT 505.950 519.450 508.050 520.050 ;
        RECT 496.950 518.550 508.050 519.450 ;
        RECT 496.950 517.950 499.050 518.550 ;
        RECT 505.950 517.950 508.050 518.550 ;
        RECT 509.100 518.700 510.300 523.950 ;
        RECT 512.100 522.150 513.900 523.950 ;
        RECT 509.100 517.800 513.300 518.700 ;
        RECT 491.100 510.600 492.900 516.600 ;
        RECT 506.400 510.000 508.200 516.600 ;
        RECT 511.500 510.600 513.300 517.800 ;
        RECT 527.700 513.600 528.900 523.950 ;
        RECT 533.550 516.600 534.750 523.950 ;
        RECT 546.150 520.200 547.050 532.800 ;
        RECT 549.150 532.800 550.050 534.900 ;
        RECT 550.950 534.300 558.750 535.500 ;
        RECT 550.950 533.700 552.750 534.300 ;
        RECT 562.050 533.400 563.850 546.000 ;
        RECT 565.050 535.200 566.850 545.400 ;
        RECT 565.050 533.400 567.450 535.200 ;
        RECT 581.100 533.400 582.900 546.000 ;
        RECT 584.100 533.400 585.900 545.400 ;
        RECT 599.100 539.400 600.900 546.000 ;
        RECT 602.100 539.400 603.900 545.400 ;
        RECT 605.100 539.400 606.900 546.000 ;
        RECT 620.100 539.400 621.900 546.000 ;
        RECT 623.100 539.400 624.900 545.400 ;
        RECT 626.100 539.400 627.900 546.000 ;
        RECT 549.150 532.500 557.550 532.800 ;
        RECT 566.550 532.500 567.450 533.400 ;
        RECT 549.150 531.900 567.450 532.500 ;
        RECT 555.750 531.300 567.450 531.900 ;
        RECT 555.750 531.000 557.550 531.300 ;
        RECT 553.800 524.400 555.900 526.050 ;
        RECT 553.800 523.200 561.900 524.400 ;
        RECT 562.950 523.950 565.050 526.050 ;
        RECT 560.100 522.600 561.900 523.200 ;
        RECT 557.100 521.400 558.900 522.000 ;
        RECT 563.250 521.400 565.050 523.950 ;
        RECT 557.100 520.200 565.050 521.400 ;
        RECT 546.150 519.000 558.150 520.200 ;
        RECT 546.150 518.400 547.950 519.000 ;
        RECT 557.100 517.200 558.150 519.000 ;
        RECT 527.100 510.600 528.900 513.600 ;
        RECT 530.100 510.000 531.900 513.600 ;
        RECT 533.550 510.600 535.350 516.600 ;
        RECT 536.850 510.000 538.650 516.600 ;
        RECT 541.350 513.600 543.750 515.700 ;
        RECT 553.350 515.550 555.150 516.300 ;
        RECT 550.200 514.500 555.150 515.550 ;
        RECT 556.350 515.400 558.150 517.200 ;
        RECT 566.550 516.600 567.450 531.300 ;
        RECT 584.100 526.050 585.300 533.400 ;
        RECT 602.100 526.050 603.300 539.400 ;
        RECT 623.700 526.050 624.900 539.400 ;
        RECT 644.100 534.300 645.900 545.400 ;
        RECT 647.100 535.200 648.900 546.000 ;
        RECT 650.100 534.300 651.900 545.400 ;
        RECT 644.100 533.400 651.900 534.300 ;
        RECT 653.100 533.400 654.900 545.400 ;
        RECT 671.400 533.400 673.200 546.000 ;
        RECT 676.500 534.900 678.300 545.400 ;
        RECT 679.500 539.400 681.300 546.000 ;
        RECT 698.100 539.400 699.900 546.000 ;
        RECT 701.100 539.400 702.900 545.400 ;
        RECT 704.100 540.000 705.900 546.000 ;
        RECT 701.400 539.100 702.900 539.400 ;
        RECT 707.100 539.400 708.900 545.400 ;
        RECT 707.100 539.100 708.000 539.400 ;
        RECT 701.400 538.200 708.000 539.100 ;
        RECT 679.200 536.100 681.000 537.900 ;
        RECT 676.500 533.400 678.900 534.900 ;
        RECT 647.250 526.050 649.050 527.850 ;
        RECT 653.700 526.050 654.600 533.400 ;
        RECT 671.100 526.050 672.900 527.850 ;
        RECT 677.700 526.050 678.900 533.400 ;
        RECT 691.950 531.450 694.050 532.050 ;
        RECT 703.950 531.450 706.050 532.050 ;
        RECT 691.950 530.550 706.050 531.450 ;
        RECT 691.950 529.950 694.050 530.550 ;
        RECT 703.950 529.950 706.050 530.550 ;
        RECT 701.100 526.050 702.900 527.850 ;
        RECT 707.100 526.050 708.000 538.200 ;
        RECT 722.100 534.300 723.900 545.400 ;
        RECT 725.100 535.200 726.900 546.000 ;
        RECT 728.100 534.300 729.900 545.400 ;
        RECT 722.100 533.400 729.900 534.300 ;
        RECT 731.100 533.400 732.900 545.400 ;
        RECT 746.100 539.400 747.900 546.000 ;
        RECT 749.100 539.400 750.900 545.400 ;
        RECT 712.950 531.450 715.050 532.050 ;
        RECT 721.950 531.450 724.050 532.050 ;
        RECT 712.950 530.550 724.050 531.450 ;
        RECT 712.950 529.950 715.050 530.550 ;
        RECT 721.950 529.950 724.050 530.550 ;
        RECT 725.250 526.050 727.050 527.850 ;
        RECT 731.700 526.050 732.600 533.400 ;
        RECT 746.100 526.050 747.900 527.850 ;
        RECT 749.100 526.050 750.300 539.400 ;
        RECT 767.400 533.400 769.200 546.000 ;
        RECT 772.500 534.900 774.300 545.400 ;
        RECT 775.500 539.400 777.300 546.000 ;
        RECT 775.200 536.100 777.000 537.900 ;
        RECT 772.500 533.400 774.900 534.900 ;
        RECT 791.400 533.400 793.200 546.000 ;
        RECT 796.500 534.900 798.300 545.400 ;
        RECT 799.500 539.400 801.300 546.000 ;
        RECT 815.100 539.400 816.900 546.000 ;
        RECT 818.100 539.400 819.900 545.400 ;
        RECT 821.100 540.000 822.900 546.000 ;
        RECT 818.400 539.100 819.900 539.400 ;
        RECT 824.100 539.400 825.900 545.400 ;
        RECT 839.100 539.400 840.900 546.000 ;
        RECT 842.100 539.400 843.900 545.400 ;
        RECT 845.100 540.000 846.900 546.000 ;
        RECT 824.100 539.100 825.000 539.400 ;
        RECT 818.400 538.200 825.000 539.100 ;
        RECT 842.400 539.100 843.900 539.400 ;
        RECT 848.100 539.400 849.900 545.400 ;
        RECT 863.100 539.400 864.900 546.000 ;
        RECT 866.100 539.400 867.900 545.400 ;
        RECT 869.100 540.000 870.900 546.000 ;
        RECT 848.100 539.100 849.000 539.400 ;
        RECT 842.400 538.200 849.000 539.100 ;
        RECT 866.400 539.100 867.900 539.400 ;
        RECT 872.100 539.400 873.900 545.400 ;
        RECT 887.100 539.400 888.900 545.400 ;
        RECT 890.100 540.000 891.900 546.000 ;
        RECT 872.100 539.100 873.000 539.400 ;
        RECT 866.400 538.200 873.000 539.100 ;
        RECT 799.200 536.100 801.000 537.900 ;
        RECT 796.500 533.400 798.900 534.900 ;
        RECT 767.100 526.050 768.900 527.850 ;
        RECT 773.700 526.050 774.900 533.400 ;
        RECT 781.950 531.450 784.050 532.050 ;
        RECT 793.950 531.450 796.050 532.050 ;
        RECT 781.950 530.550 796.050 531.450 ;
        RECT 781.950 529.950 784.050 530.550 ;
        RECT 793.950 529.950 796.050 530.550 ;
        RECT 791.100 526.050 792.900 527.850 ;
        RECT 797.700 526.050 798.900 533.400 ;
        RECT 818.100 526.050 819.900 527.850 ;
        RECT 824.100 526.050 825.000 538.200 ;
        RECT 826.950 528.450 831.000 529.050 ;
        RECT 826.950 526.950 831.450 528.450 ;
        RECT 580.950 523.950 583.050 526.050 ;
        RECT 583.950 523.950 586.050 526.050 ;
        RECT 598.950 523.950 601.050 526.050 ;
        RECT 601.950 523.950 604.050 526.050 ;
        RECT 604.950 523.950 607.050 526.050 ;
        RECT 619.950 523.950 622.050 526.050 ;
        RECT 622.950 523.950 625.050 526.050 ;
        RECT 625.950 523.950 628.050 526.050 ;
        RECT 643.950 523.950 646.050 526.050 ;
        RECT 646.950 523.950 649.050 526.050 ;
        RECT 649.950 523.950 652.050 526.050 ;
        RECT 652.950 523.950 655.050 526.050 ;
        RECT 670.950 523.950 673.050 526.050 ;
        RECT 673.950 523.950 676.050 526.050 ;
        RECT 676.950 523.950 679.050 526.050 ;
        RECT 679.950 523.950 682.050 526.050 ;
        RECT 697.950 523.950 700.050 526.050 ;
        RECT 700.950 523.950 703.050 526.050 ;
        RECT 703.950 523.950 706.050 526.050 ;
        RECT 706.950 523.950 709.050 526.050 ;
        RECT 721.950 523.950 724.050 526.050 ;
        RECT 724.950 523.950 727.050 526.050 ;
        RECT 727.950 523.950 730.050 526.050 ;
        RECT 730.950 523.950 733.050 526.050 ;
        RECT 745.950 523.950 748.050 526.050 ;
        RECT 748.950 523.950 751.050 526.050 ;
        RECT 766.950 523.950 769.050 526.050 ;
        RECT 769.950 523.950 772.050 526.050 ;
        RECT 772.950 523.950 775.050 526.050 ;
        RECT 775.950 523.950 778.050 526.050 ;
        RECT 790.950 523.950 793.050 526.050 ;
        RECT 793.950 523.950 796.050 526.050 ;
        RECT 796.950 523.950 799.050 526.050 ;
        RECT 799.950 523.950 802.050 526.050 ;
        RECT 814.950 523.950 817.050 526.050 ;
        RECT 817.950 523.950 820.050 526.050 ;
        RECT 820.950 523.950 823.050 526.050 ;
        RECT 823.950 523.950 826.050 526.050 ;
        RECT 581.100 522.150 582.900 523.950 ;
        RECT 584.100 516.600 585.300 523.950 ;
        RECT 599.250 522.150 601.050 523.950 ;
        RECT 602.100 518.700 603.300 523.950 ;
        RECT 605.100 522.150 606.900 523.950 ;
        RECT 620.100 522.150 621.900 523.950 ;
        RECT 623.700 518.700 624.900 523.950 ;
        RECT 625.950 522.150 627.750 523.950 ;
        RECT 644.100 522.150 645.900 523.950 ;
        RECT 650.250 522.150 652.050 523.950 ;
        RECT 602.100 517.800 606.300 518.700 ;
        RECT 550.200 513.600 551.250 514.500 ;
        RECT 559.050 514.200 561.150 515.700 ;
        RECT 557.250 513.600 561.150 514.200 ;
        RECT 541.950 510.600 543.750 513.600 ;
        RECT 546.450 510.000 548.250 513.600 ;
        RECT 549.450 510.600 551.250 513.600 ;
        RECT 552.750 510.000 554.550 513.600 ;
        RECT 557.250 512.700 560.850 513.600 ;
        RECT 557.250 510.600 559.050 512.700 ;
        RECT 562.050 510.000 563.850 516.600 ;
        RECT 565.050 514.800 567.450 516.600 ;
        RECT 565.050 510.600 566.850 514.800 ;
        RECT 581.100 510.000 582.900 516.600 ;
        RECT 584.100 510.600 585.900 516.600 ;
        RECT 599.400 510.000 601.200 516.600 ;
        RECT 604.500 510.600 606.300 517.800 ;
        RECT 620.700 517.800 624.900 518.700 ;
        RECT 625.950 519.450 628.050 520.050 ;
        RECT 646.950 519.450 649.050 520.050 ;
        RECT 625.950 518.550 649.050 519.450 ;
        RECT 625.950 517.950 628.050 518.550 ;
        RECT 646.950 517.950 649.050 518.550 ;
        RECT 620.700 510.600 622.500 517.800 ;
        RECT 653.700 516.600 654.600 523.950 ;
        RECT 674.100 522.150 675.900 523.950 ;
        RECT 677.700 519.600 678.900 523.950 ;
        RECT 680.100 522.150 681.900 523.950 ;
        RECT 698.100 522.150 699.900 523.950 ;
        RECT 704.100 522.150 705.900 523.950 ;
        RECT 707.100 520.200 708.000 523.950 ;
        RECT 722.100 522.150 723.900 523.950 ;
        RECT 728.250 522.150 730.050 523.950 ;
        RECT 677.700 518.700 681.300 519.600 ;
        RECT 625.800 510.000 627.600 516.600 ;
        RECT 645.000 510.000 646.800 516.600 ;
        RECT 649.500 515.400 654.600 516.600 ;
        RECT 671.100 515.700 678.900 517.050 ;
        RECT 649.500 510.600 651.300 515.400 ;
        RECT 652.500 510.000 654.300 513.600 ;
        RECT 671.100 510.600 672.900 515.700 ;
        RECT 674.100 510.000 675.900 514.800 ;
        RECT 677.100 510.600 678.900 515.700 ;
        RECT 680.100 516.600 681.300 518.700 ;
        RECT 680.100 510.600 681.900 516.600 ;
        RECT 698.100 510.000 699.900 519.600 ;
        RECT 704.700 519.000 708.000 520.200 ;
        RECT 704.700 510.600 706.500 519.000 ;
        RECT 731.700 516.600 732.600 523.950 ;
        RECT 723.000 510.000 724.800 516.600 ;
        RECT 727.500 515.400 732.600 516.600 ;
        RECT 727.500 510.600 729.300 515.400 ;
        RECT 749.100 513.600 750.300 523.950 ;
        RECT 757.950 522.450 760.050 523.050 ;
        RECT 763.950 522.450 766.050 523.050 ;
        RECT 757.950 521.550 766.050 522.450 ;
        RECT 770.100 522.150 771.900 523.950 ;
        RECT 757.950 520.950 760.050 521.550 ;
        RECT 763.950 520.950 766.050 521.550 ;
        RECT 773.700 519.600 774.900 523.950 ;
        RECT 776.100 522.150 777.900 523.950 ;
        RECT 794.100 522.150 795.900 523.950 ;
        RECT 797.700 519.600 798.900 523.950 ;
        RECT 800.100 522.150 801.900 523.950 ;
        RECT 815.100 522.150 816.900 523.950 ;
        RECT 821.100 522.150 822.900 523.950 ;
        RECT 824.100 520.200 825.000 523.950 ;
        RECT 830.550 523.050 831.450 526.950 ;
        RECT 842.100 526.050 843.900 527.850 ;
        RECT 848.100 526.050 849.000 538.200 ;
        RECT 866.100 526.050 867.900 527.850 ;
        RECT 872.100 526.050 873.000 538.200 ;
        RECT 888.000 539.100 888.900 539.400 ;
        RECT 893.100 539.400 894.900 545.400 ;
        RECT 896.100 539.400 897.900 546.000 ;
        RECT 911.100 539.400 912.900 545.400 ;
        RECT 914.100 540.000 915.900 546.000 ;
        RECT 893.100 539.100 894.600 539.400 ;
        RECT 888.000 538.200 894.600 539.100 ;
        RECT 912.000 539.100 912.900 539.400 ;
        RECT 917.100 539.400 918.900 545.400 ;
        RECT 920.100 539.400 921.900 546.000 ;
        RECT 938.100 539.400 939.900 546.000 ;
        RECT 941.100 539.400 942.900 545.400 ;
        RECT 917.100 539.100 918.600 539.400 ;
        RECT 912.000 538.200 918.600 539.100 ;
        RECT 882.000 528.450 886.050 529.050 ;
        RECT 881.550 526.950 886.050 528.450 ;
        RECT 838.950 523.950 841.050 526.050 ;
        RECT 841.950 523.950 844.050 526.050 ;
        RECT 844.950 523.950 847.050 526.050 ;
        RECT 847.950 523.950 850.050 526.050 ;
        RECT 862.950 523.950 865.050 526.050 ;
        RECT 865.950 523.950 868.050 526.050 ;
        RECT 868.950 523.950 871.050 526.050 ;
        RECT 871.950 523.950 874.050 526.050 ;
        RECT 826.950 521.550 831.450 523.050 ;
        RECT 839.100 522.150 840.900 523.950 ;
        RECT 845.100 522.150 846.900 523.950 ;
        RECT 826.950 520.950 831.000 521.550 ;
        RECT 848.100 520.200 849.000 523.950 ;
        RECT 863.100 522.150 864.900 523.950 ;
        RECT 869.100 522.150 870.900 523.950 ;
        RECT 872.100 520.200 873.000 523.950 ;
        RECT 773.700 518.700 777.300 519.600 ;
        RECT 797.700 518.700 801.300 519.600 ;
        RECT 767.100 515.700 774.900 517.050 ;
        RECT 730.500 510.000 732.300 513.600 ;
        RECT 746.100 510.000 747.900 513.600 ;
        RECT 749.100 510.600 750.900 513.600 ;
        RECT 767.100 510.600 768.900 515.700 ;
        RECT 770.100 510.000 771.900 514.800 ;
        RECT 773.100 510.600 774.900 515.700 ;
        RECT 776.100 516.600 777.300 518.700 ;
        RECT 776.100 510.600 777.900 516.600 ;
        RECT 791.100 515.700 798.900 517.050 ;
        RECT 791.100 510.600 792.900 515.700 ;
        RECT 794.100 510.000 795.900 514.800 ;
        RECT 797.100 510.600 798.900 515.700 ;
        RECT 800.100 516.600 801.300 518.700 ;
        RECT 800.100 510.600 801.900 516.600 ;
        RECT 815.100 510.000 816.900 519.600 ;
        RECT 821.700 519.000 825.000 520.200 ;
        RECT 821.700 510.600 823.500 519.000 ;
        RECT 839.100 510.000 840.900 519.600 ;
        RECT 845.700 519.000 849.000 520.200 ;
        RECT 845.700 510.600 847.500 519.000 ;
        RECT 863.100 510.000 864.900 519.600 ;
        RECT 869.700 519.000 873.000 520.200 ;
        RECT 874.950 519.450 877.050 519.900 ;
        RECT 881.550 519.450 882.450 526.950 ;
        RECT 888.000 526.050 888.900 538.200 ;
        RECT 904.950 529.950 907.050 532.050 ;
        RECT 893.100 526.050 894.900 527.850 ;
        RECT 886.950 523.950 889.050 526.050 ;
        RECT 889.950 523.950 892.050 526.050 ;
        RECT 892.950 523.950 895.050 526.050 ;
        RECT 895.950 523.950 898.050 526.050 ;
        RECT 869.700 510.600 871.500 519.000 ;
        RECT 874.950 518.550 882.450 519.450 ;
        RECT 888.000 520.200 888.900 523.950 ;
        RECT 890.100 522.150 891.900 523.950 ;
        RECT 896.100 522.150 897.900 523.950 ;
        RECT 898.950 522.450 901.050 523.050 ;
        RECT 905.550 522.450 906.450 529.950 ;
        RECT 912.000 526.050 912.900 538.200 ;
        RECT 933.000 528.450 937.050 529.050 ;
        RECT 917.100 526.050 918.900 527.850 ;
        RECT 932.550 526.950 937.050 528.450 ;
        RECT 910.950 523.950 913.050 526.050 ;
        RECT 913.950 523.950 916.050 526.050 ;
        RECT 916.950 523.950 919.050 526.050 ;
        RECT 919.950 523.950 922.050 526.050 ;
        RECT 898.950 521.550 906.450 522.450 ;
        RECT 898.950 520.950 901.050 521.550 ;
        RECT 912.000 520.200 912.900 523.950 ;
        RECT 914.100 522.150 915.900 523.950 ;
        RECT 920.100 522.150 921.900 523.950 ;
        RECT 922.950 522.450 925.050 523.050 ;
        RECT 932.550 522.450 933.450 526.950 ;
        RECT 938.100 526.050 939.900 527.850 ;
        RECT 941.100 526.050 942.300 539.400 ;
        RECT 956.100 533.400 957.900 545.400 ;
        RECT 959.100 534.300 960.900 545.400 ;
        RECT 962.100 535.200 963.900 546.000 ;
        RECT 965.100 534.300 966.900 545.400 ;
        RECT 983.100 539.400 984.900 545.400 ;
        RECT 986.100 539.400 987.900 546.000 ;
        RECT 959.100 533.400 966.900 534.300 ;
        RECT 956.400 526.050 957.300 533.400 ;
        RECT 961.950 526.050 963.750 527.850 ;
        RECT 983.700 526.050 984.900 539.400 ;
        RECT 1001.400 533.400 1003.200 546.000 ;
        RECT 1006.500 534.900 1008.300 545.400 ;
        RECT 1009.500 539.400 1011.300 546.000 ;
        RECT 1009.200 536.100 1011.000 537.900 ;
        RECT 1006.500 533.400 1008.900 534.900 ;
        RECT 986.100 526.050 987.900 527.850 ;
        RECT 1001.100 526.050 1002.900 527.850 ;
        RECT 1007.700 526.050 1008.900 533.400 ;
        RECT 937.950 523.950 940.050 526.050 ;
        RECT 940.950 523.950 943.050 526.050 ;
        RECT 955.950 523.950 958.050 526.050 ;
        RECT 958.950 523.950 961.050 526.050 ;
        RECT 961.950 523.950 964.050 526.050 ;
        RECT 964.950 523.950 967.050 526.050 ;
        RECT 982.950 523.950 985.050 526.050 ;
        RECT 985.950 523.950 988.050 526.050 ;
        RECT 1000.950 523.950 1003.050 526.050 ;
        RECT 1003.950 523.950 1006.050 526.050 ;
        RECT 1006.950 523.950 1009.050 526.050 ;
        RECT 1009.950 523.950 1012.050 526.050 ;
        RECT 922.950 521.550 933.450 522.450 ;
        RECT 922.950 520.950 925.050 521.550 ;
        RECT 888.000 519.000 891.300 520.200 ;
        RECT 874.950 517.800 877.050 518.550 ;
        RECT 877.950 516.450 880.050 517.050 ;
        RECT 883.950 516.450 886.050 517.050 ;
        RECT 877.950 515.550 886.050 516.450 ;
        RECT 877.950 514.950 880.050 515.550 ;
        RECT 883.950 514.950 886.050 515.550 ;
        RECT 889.500 510.600 891.300 519.000 ;
        RECT 896.100 510.000 897.900 519.600 ;
        RECT 912.000 519.000 915.300 520.200 ;
        RECT 913.500 510.600 915.300 519.000 ;
        RECT 920.100 510.000 921.900 519.600 ;
        RECT 941.100 513.600 942.300 523.950 ;
        RECT 946.950 522.450 949.050 523.050 ;
        RECT 952.950 522.450 955.050 523.050 ;
        RECT 946.950 521.550 955.050 522.450 ;
        RECT 946.950 520.950 949.050 521.550 ;
        RECT 952.950 520.950 955.050 521.550 ;
        RECT 956.400 516.600 957.300 523.950 ;
        RECT 958.950 522.150 960.750 523.950 ;
        RECT 965.100 522.150 966.900 523.950 ;
        RECT 956.400 515.400 961.500 516.600 ;
        RECT 938.100 510.000 939.900 513.600 ;
        RECT 941.100 510.600 942.900 513.600 ;
        RECT 956.700 510.000 958.500 513.600 ;
        RECT 959.700 510.600 961.500 515.400 ;
        RECT 964.200 510.000 966.000 516.600 ;
        RECT 983.700 513.600 984.900 523.950 ;
        RECT 1004.100 522.150 1005.900 523.950 ;
        RECT 1007.700 519.600 1008.900 523.950 ;
        RECT 1010.100 522.150 1011.900 523.950 ;
        RECT 1007.700 518.700 1011.300 519.600 ;
        RECT 1001.100 515.700 1008.900 517.050 ;
        RECT 983.100 510.600 984.900 513.600 ;
        RECT 986.100 510.000 987.900 513.600 ;
        RECT 1001.100 510.600 1002.900 515.700 ;
        RECT 1004.100 510.000 1005.900 514.800 ;
        RECT 1007.100 510.600 1008.900 515.700 ;
        RECT 1010.100 516.600 1011.300 518.700 ;
        RECT 1010.100 510.600 1011.900 516.600 ;
        RECT 14.100 500.400 15.900 506.400 ;
        RECT 17.100 500.400 18.900 507.000 ;
        RECT 20.100 503.400 21.900 506.400 ;
        RECT 14.100 493.050 15.300 500.400 ;
        RECT 20.700 499.500 21.900 503.400 ;
        RECT 35.100 500.400 36.900 507.000 ;
        RECT 16.200 498.600 21.900 499.500 ;
        RECT 38.100 499.500 39.900 506.400 ;
        RECT 41.100 500.400 42.900 507.000 ;
        RECT 44.100 499.500 45.900 506.400 ;
        RECT 47.100 500.400 48.900 507.000 ;
        RECT 50.100 499.500 51.900 506.400 ;
        RECT 53.100 500.400 54.900 507.000 ;
        RECT 56.100 499.500 57.900 506.400 ;
        RECT 59.100 500.400 60.900 507.000 ;
        RECT 63.150 502.200 64.950 506.400 ;
        RECT 62.550 500.400 64.950 502.200 ;
        RECT 66.150 500.400 67.950 507.000 ;
        RECT 70.950 504.300 72.750 506.400 ;
        RECT 69.150 503.400 72.750 504.300 ;
        RECT 75.450 503.400 77.250 507.000 ;
        RECT 78.750 503.400 80.550 506.400 ;
        RECT 81.750 503.400 83.550 507.000 ;
        RECT 86.250 503.400 88.050 506.400 ;
        RECT 68.850 502.800 72.750 503.400 ;
        RECT 68.850 501.300 70.950 502.800 ;
        RECT 78.750 502.500 79.800 503.400 ;
        RECT 16.200 497.700 18.000 498.600 ;
        RECT 38.100 498.300 42.000 499.500 ;
        RECT 44.100 498.300 48.000 499.500 ;
        RECT 50.100 498.300 54.000 499.500 ;
        RECT 56.100 498.300 58.950 499.500 ;
        RECT 14.100 490.950 16.200 493.050 ;
        RECT 14.100 483.600 15.300 490.950 ;
        RECT 17.100 486.300 18.000 497.700 ;
        RECT 40.800 497.400 42.000 498.300 ;
        RECT 46.800 497.400 48.000 498.300 ;
        RECT 52.800 497.400 54.000 498.300 ;
        RECT 40.800 496.200 45.000 497.400 ;
        RECT 37.800 493.050 39.600 494.850 ;
        RECT 19.500 490.950 21.600 493.050 ;
        RECT 37.800 490.950 39.900 493.050 ;
        RECT 19.800 489.150 21.600 490.950 ;
        RECT 16.200 485.400 18.000 486.300 ;
        RECT 40.800 485.700 42.000 496.200 ;
        RECT 43.200 495.600 45.000 496.200 ;
        RECT 46.800 496.200 51.000 497.400 ;
        RECT 46.800 485.700 48.000 496.200 ;
        RECT 49.200 495.600 51.000 496.200 ;
        RECT 52.800 496.200 57.000 497.400 ;
        RECT 52.800 485.700 54.000 496.200 ;
        RECT 55.200 495.600 57.000 496.200 ;
        RECT 57.900 493.050 58.950 498.300 ;
        RECT 55.800 490.950 58.950 493.050 ;
        RECT 57.900 485.700 58.950 490.950 ;
        RECT 16.200 484.500 21.900 485.400 ;
        RECT 14.100 471.600 15.900 483.600 ;
        RECT 17.100 471.000 18.900 481.800 ;
        RECT 20.700 477.600 21.900 484.500 ;
        RECT 38.100 484.500 42.000 485.700 ;
        RECT 44.100 484.500 48.000 485.700 ;
        RECT 50.100 484.500 54.000 485.700 ;
        RECT 56.100 484.500 58.950 485.700 ;
        RECT 62.550 485.700 63.450 500.400 ;
        RECT 71.850 499.800 73.650 501.600 ;
        RECT 74.850 501.450 79.800 502.500 ;
        RECT 74.850 500.700 76.650 501.450 ;
        RECT 86.250 501.300 88.650 503.400 ;
        RECT 91.350 500.400 93.150 507.000 ;
        RECT 94.650 500.400 96.450 506.400 ;
        RECT 99.150 502.200 100.950 506.400 ;
        RECT 71.850 498.000 72.900 499.800 ;
        RECT 82.050 498.000 83.850 498.600 ;
        RECT 71.850 496.800 83.850 498.000 ;
        RECT 64.950 495.600 72.900 496.800 ;
        RECT 64.950 493.050 66.750 495.600 ;
        RECT 71.100 495.000 72.900 495.600 ;
        RECT 68.100 493.800 69.900 494.400 ;
        RECT 64.950 490.950 67.050 493.050 ;
        RECT 68.100 492.600 76.200 493.800 ;
        RECT 74.100 490.950 76.200 492.600 ;
        RECT 72.450 485.700 74.250 486.000 ;
        RECT 62.550 485.100 74.250 485.700 ;
        RECT 62.550 484.500 80.850 485.100 ;
        RECT 20.100 471.600 21.900 477.600 ;
        RECT 35.100 471.000 36.900 483.600 ;
        RECT 38.100 471.600 39.900 484.500 ;
        RECT 41.100 471.000 42.900 483.600 ;
        RECT 44.100 471.600 45.900 484.500 ;
        RECT 47.100 471.000 48.900 483.600 ;
        RECT 50.100 471.600 51.900 484.500 ;
        RECT 53.100 471.000 54.900 483.600 ;
        RECT 56.100 471.600 57.900 484.500 ;
        RECT 62.550 483.600 63.450 484.500 ;
        RECT 72.450 484.200 80.850 484.500 ;
        RECT 59.100 471.000 60.900 483.600 ;
        RECT 62.550 481.800 64.950 483.600 ;
        RECT 63.150 471.600 64.950 481.800 ;
        RECT 66.150 471.000 67.950 483.600 ;
        RECT 77.250 482.700 79.050 483.300 ;
        RECT 71.250 481.500 79.050 482.700 ;
        RECT 79.950 482.100 80.850 484.200 ;
        RECT 82.950 484.200 83.850 496.800 ;
        RECT 95.250 493.050 96.450 500.400 ;
        RECT 90.150 491.250 96.450 493.050 ;
        RECT 91.950 490.950 96.450 491.250 ;
        RECT 86.550 488.100 88.650 488.400 ;
        RECT 92.550 488.100 94.350 488.250 ;
        RECT 86.550 486.900 94.350 488.100 ;
        RECT 86.550 486.300 88.650 486.900 ;
        RECT 92.550 486.450 94.350 486.900 ;
        RECT 82.950 483.300 87.750 484.200 ;
        RECT 95.250 483.600 96.450 490.950 ;
        RECT 86.550 482.400 87.750 483.300 ;
        RECT 83.850 482.100 85.650 482.400 ;
        RECT 71.250 480.600 73.350 481.500 ;
        RECT 79.950 481.200 85.650 482.100 ;
        RECT 83.850 480.600 85.650 481.200 ;
        RECT 86.550 480.600 89.550 482.400 ;
        RECT 71.550 471.600 73.350 480.600 ;
        RECT 75.450 479.550 77.250 480.300 ;
        RECT 80.250 479.550 82.050 480.300 ;
        RECT 75.450 478.500 82.050 479.550 ;
        RECT 76.350 471.000 78.150 477.600 ;
        RECT 79.350 471.600 81.150 478.500 ;
        RECT 86.550 477.600 88.650 479.700 ;
        RECT 82.350 471.000 84.150 477.600 ;
        RECT 86.850 471.600 88.650 477.600 ;
        RECT 91.650 471.000 93.450 483.600 ;
        RECT 94.650 471.600 96.450 483.600 ;
        RECT 98.550 500.400 100.950 502.200 ;
        RECT 102.150 500.400 103.950 507.000 ;
        RECT 106.950 504.300 108.750 506.400 ;
        RECT 105.150 503.400 108.750 504.300 ;
        RECT 111.450 503.400 113.250 507.000 ;
        RECT 114.750 503.400 116.550 506.400 ;
        RECT 117.750 503.400 119.550 507.000 ;
        RECT 122.250 503.400 124.050 506.400 ;
        RECT 104.850 502.800 108.750 503.400 ;
        RECT 104.850 501.300 106.950 502.800 ;
        RECT 114.750 502.500 115.800 503.400 ;
        RECT 98.550 485.700 99.450 500.400 ;
        RECT 107.850 499.800 109.650 501.600 ;
        RECT 110.850 501.450 115.800 502.500 ;
        RECT 110.850 500.700 112.650 501.450 ;
        RECT 122.250 501.300 124.650 503.400 ;
        RECT 127.350 500.400 129.150 507.000 ;
        RECT 130.650 500.400 132.450 506.400 ;
        RECT 149.100 503.400 150.900 507.000 ;
        RECT 152.100 503.400 153.900 506.400 ;
        RECT 155.100 503.400 156.900 507.000 ;
        RECT 107.850 498.000 108.900 499.800 ;
        RECT 118.050 498.000 119.850 498.600 ;
        RECT 107.850 496.800 119.850 498.000 ;
        RECT 100.950 495.600 108.900 496.800 ;
        RECT 100.950 493.050 102.750 495.600 ;
        RECT 107.100 495.000 108.900 495.600 ;
        RECT 104.100 493.800 105.900 494.400 ;
        RECT 100.950 490.950 103.050 493.050 ;
        RECT 104.100 492.600 112.200 493.800 ;
        RECT 110.100 490.950 112.200 492.600 ;
        RECT 108.450 485.700 110.250 486.000 ;
        RECT 98.550 485.100 110.250 485.700 ;
        RECT 98.550 484.500 116.850 485.100 ;
        RECT 98.550 483.600 99.450 484.500 ;
        RECT 108.450 484.200 116.850 484.500 ;
        RECT 98.550 481.800 100.950 483.600 ;
        RECT 99.150 471.600 100.950 481.800 ;
        RECT 102.150 471.000 103.950 483.600 ;
        RECT 113.250 482.700 115.050 483.300 ;
        RECT 107.250 481.500 115.050 482.700 ;
        RECT 115.950 482.100 116.850 484.200 ;
        RECT 118.950 484.200 119.850 496.800 ;
        RECT 131.250 493.050 132.450 500.400 ;
        RECT 152.700 493.050 153.600 503.400 ;
        RECT 170.100 500.400 171.900 506.400 ;
        RECT 173.100 500.400 174.900 507.000 ;
        RECT 188.100 500.400 189.900 507.000 ;
        RECT 191.100 500.400 192.900 506.400 ;
        RECT 206.100 500.400 207.900 506.400 ;
        RECT 157.950 495.450 162.000 496.050 ;
        RECT 157.950 495.000 162.450 495.450 ;
        RECT 157.950 493.950 163.050 495.000 ;
        RECT 126.150 491.250 132.450 493.050 ;
        RECT 127.950 490.950 132.450 491.250 ;
        RECT 148.950 490.950 151.050 493.050 ;
        RECT 151.950 490.950 154.050 493.050 ;
        RECT 154.950 490.950 157.050 493.050 ;
        RECT 122.550 488.100 124.650 488.400 ;
        RECT 128.550 488.100 130.350 488.250 ;
        RECT 122.550 486.900 130.350 488.100 ;
        RECT 122.550 486.300 124.650 486.900 ;
        RECT 128.550 486.450 130.350 486.900 ;
        RECT 118.950 483.300 123.750 484.200 ;
        RECT 131.250 483.600 132.450 490.950 ;
        RECT 149.100 489.150 150.900 490.950 ;
        RECT 152.700 483.600 153.600 490.950 ;
        RECT 154.950 489.150 156.750 490.950 ;
        RECT 160.950 490.800 163.050 493.950 ;
        RECT 170.700 493.050 171.900 500.400 ;
        RECT 173.100 493.050 174.900 494.850 ;
        RECT 188.100 493.050 189.900 494.850 ;
        RECT 191.100 493.050 192.300 500.400 ;
        RECT 206.700 498.300 207.900 500.400 ;
        RECT 209.100 501.300 210.900 506.400 ;
        RECT 212.100 502.200 213.900 507.000 ;
        RECT 215.100 501.300 216.900 506.400 ;
        RECT 209.100 499.950 216.900 501.300 ;
        RECT 230.100 501.300 231.900 506.400 ;
        RECT 233.100 502.200 234.900 507.000 ;
        RECT 236.100 501.300 237.900 506.400 ;
        RECT 230.100 499.950 237.900 501.300 ;
        RECT 239.100 500.400 240.900 506.400 ;
        RECT 243.150 502.200 244.950 506.400 ;
        RECT 242.550 500.400 244.950 502.200 ;
        RECT 246.150 500.400 247.950 507.000 ;
        RECT 250.950 504.300 252.750 506.400 ;
        RECT 249.150 503.400 252.750 504.300 ;
        RECT 255.450 503.400 257.250 507.000 ;
        RECT 258.750 503.400 260.550 506.400 ;
        RECT 261.750 503.400 263.550 507.000 ;
        RECT 266.250 503.400 268.050 506.400 ;
        RECT 248.850 502.800 252.750 503.400 ;
        RECT 248.850 501.300 250.950 502.800 ;
        RECT 258.750 502.500 259.800 503.400 ;
        RECT 239.100 498.300 240.300 500.400 ;
        RECT 206.700 497.400 210.300 498.300 ;
        RECT 206.100 493.050 207.900 494.850 ;
        RECT 209.100 493.050 210.300 497.400 ;
        RECT 236.700 497.400 240.300 498.300 ;
        RECT 212.100 493.050 213.900 494.850 ;
        RECT 233.100 493.050 234.900 494.850 ;
        RECT 236.700 493.050 237.900 497.400 ;
        RECT 239.100 493.050 240.900 494.850 ;
        RECT 169.950 490.950 172.050 493.050 ;
        RECT 172.950 490.950 175.050 493.050 ;
        RECT 187.950 490.950 190.050 493.050 ;
        RECT 190.950 490.950 193.050 493.050 ;
        RECT 205.950 490.950 208.050 493.050 ;
        RECT 208.950 490.950 211.050 493.050 ;
        RECT 211.950 490.950 214.050 493.050 ;
        RECT 214.950 490.950 217.050 493.050 ;
        RECT 229.950 490.950 232.050 493.050 ;
        RECT 232.950 490.950 235.050 493.050 ;
        RECT 235.950 490.950 238.050 493.050 ;
        RECT 238.950 490.950 241.050 493.050 ;
        RECT 170.700 483.600 171.900 490.950 ;
        RECT 191.100 483.600 192.300 490.950 ;
        RECT 209.100 483.600 210.300 490.950 ;
        RECT 215.100 489.150 216.900 490.950 ;
        RECT 230.100 489.150 231.900 490.950 ;
        RECT 236.700 483.600 237.900 490.950 ;
        RECT 122.550 482.400 123.750 483.300 ;
        RECT 119.850 482.100 121.650 482.400 ;
        RECT 107.250 480.600 109.350 481.500 ;
        RECT 115.950 481.200 121.650 482.100 ;
        RECT 119.850 480.600 121.650 481.200 ;
        RECT 122.550 480.600 125.550 482.400 ;
        RECT 107.550 471.600 109.350 480.600 ;
        RECT 111.450 479.550 113.250 480.300 ;
        RECT 116.250 479.550 118.050 480.300 ;
        RECT 111.450 478.500 118.050 479.550 ;
        RECT 112.350 471.000 114.150 477.600 ;
        RECT 115.350 471.600 117.150 478.500 ;
        RECT 122.550 477.600 124.650 479.700 ;
        RECT 118.350 471.000 120.150 477.600 ;
        RECT 122.850 471.600 124.650 477.600 ;
        RECT 127.650 471.000 129.450 483.600 ;
        RECT 130.650 471.600 132.450 483.600 ;
        RECT 150.000 482.400 153.600 483.600 ;
        RECT 150.000 471.600 151.800 482.400 ;
        RECT 155.100 471.000 156.900 483.600 ;
        RECT 170.100 471.600 171.900 483.600 ;
        RECT 173.100 471.000 174.900 483.600 ;
        RECT 188.100 471.000 189.900 483.600 ;
        RECT 191.100 471.600 192.900 483.600 ;
        RECT 209.100 482.100 211.500 483.600 ;
        RECT 207.000 479.100 208.800 480.900 ;
        RECT 206.700 471.000 208.500 477.600 ;
        RECT 209.700 471.600 211.500 482.100 ;
        RECT 214.800 471.000 216.600 483.600 ;
        RECT 230.400 471.000 232.200 483.600 ;
        RECT 235.500 482.100 237.900 483.600 ;
        RECT 242.550 485.700 243.450 500.400 ;
        RECT 251.850 499.800 253.650 501.600 ;
        RECT 254.850 501.450 259.800 502.500 ;
        RECT 254.850 500.700 256.650 501.450 ;
        RECT 266.250 501.300 268.650 503.400 ;
        RECT 271.350 500.400 273.150 507.000 ;
        RECT 274.650 500.400 276.450 506.400 ;
        RECT 279.150 502.200 280.950 506.400 ;
        RECT 251.850 498.000 252.900 499.800 ;
        RECT 262.050 498.000 263.850 498.600 ;
        RECT 251.850 496.800 263.850 498.000 ;
        RECT 244.950 495.600 252.900 496.800 ;
        RECT 244.950 493.050 246.750 495.600 ;
        RECT 251.100 495.000 252.900 495.600 ;
        RECT 248.100 493.800 249.900 494.400 ;
        RECT 244.950 490.950 247.050 493.050 ;
        RECT 248.100 492.600 256.200 493.800 ;
        RECT 254.100 490.950 256.200 492.600 ;
        RECT 252.450 485.700 254.250 486.000 ;
        RECT 242.550 485.100 254.250 485.700 ;
        RECT 242.550 484.500 260.850 485.100 ;
        RECT 242.550 483.600 243.450 484.500 ;
        RECT 252.450 484.200 260.850 484.500 ;
        RECT 235.500 471.600 237.300 482.100 ;
        RECT 242.550 481.800 244.950 483.600 ;
        RECT 238.200 479.100 240.000 480.900 ;
        RECT 238.500 471.000 240.300 477.600 ;
        RECT 243.150 471.600 244.950 481.800 ;
        RECT 246.150 471.000 247.950 483.600 ;
        RECT 257.250 482.700 259.050 483.300 ;
        RECT 251.250 481.500 259.050 482.700 ;
        RECT 259.950 482.100 260.850 484.200 ;
        RECT 262.950 484.200 263.850 496.800 ;
        RECT 275.250 493.050 276.450 500.400 ;
        RECT 270.150 491.250 276.450 493.050 ;
        RECT 271.950 490.950 276.450 491.250 ;
        RECT 266.550 488.100 268.650 488.400 ;
        RECT 272.550 488.100 274.350 488.250 ;
        RECT 266.550 486.900 274.350 488.100 ;
        RECT 266.550 486.300 268.650 486.900 ;
        RECT 272.550 486.450 274.350 486.900 ;
        RECT 262.950 483.300 267.750 484.200 ;
        RECT 275.250 483.600 276.450 490.950 ;
        RECT 266.550 482.400 267.750 483.300 ;
        RECT 263.850 482.100 265.650 482.400 ;
        RECT 251.250 480.600 253.350 481.500 ;
        RECT 259.950 481.200 265.650 482.100 ;
        RECT 263.850 480.600 265.650 481.200 ;
        RECT 266.550 480.600 269.550 482.400 ;
        RECT 251.550 471.600 253.350 480.600 ;
        RECT 255.450 479.550 257.250 480.300 ;
        RECT 260.250 479.550 262.050 480.300 ;
        RECT 255.450 478.500 262.050 479.550 ;
        RECT 256.350 471.000 258.150 477.600 ;
        RECT 259.350 471.600 261.150 478.500 ;
        RECT 266.550 477.600 268.650 479.700 ;
        RECT 262.350 471.000 264.150 477.600 ;
        RECT 266.850 471.600 268.650 477.600 ;
        RECT 271.650 471.000 273.450 483.600 ;
        RECT 274.650 471.600 276.450 483.600 ;
        RECT 278.550 500.400 280.950 502.200 ;
        RECT 282.150 500.400 283.950 507.000 ;
        RECT 286.950 504.300 288.750 506.400 ;
        RECT 285.150 503.400 288.750 504.300 ;
        RECT 291.450 503.400 293.250 507.000 ;
        RECT 294.750 503.400 296.550 506.400 ;
        RECT 297.750 503.400 299.550 507.000 ;
        RECT 302.250 503.400 304.050 506.400 ;
        RECT 284.850 502.800 288.750 503.400 ;
        RECT 284.850 501.300 286.950 502.800 ;
        RECT 294.750 502.500 295.800 503.400 ;
        RECT 278.550 485.700 279.450 500.400 ;
        RECT 287.850 499.800 289.650 501.600 ;
        RECT 290.850 501.450 295.800 502.500 ;
        RECT 290.850 500.700 292.650 501.450 ;
        RECT 302.250 501.300 304.650 503.400 ;
        RECT 307.350 500.400 309.150 507.000 ;
        RECT 310.650 500.400 312.450 506.400 ;
        RECT 287.850 498.000 288.900 499.800 ;
        RECT 298.050 498.000 299.850 498.600 ;
        RECT 287.850 496.800 299.850 498.000 ;
        RECT 280.950 495.600 288.900 496.800 ;
        RECT 280.950 493.050 282.750 495.600 ;
        RECT 287.100 495.000 288.900 495.600 ;
        RECT 284.100 493.800 285.900 494.400 ;
        RECT 280.950 490.950 283.050 493.050 ;
        RECT 284.100 492.600 292.200 493.800 ;
        RECT 290.100 490.950 292.200 492.600 ;
        RECT 288.450 485.700 290.250 486.000 ;
        RECT 278.550 485.100 290.250 485.700 ;
        RECT 278.550 484.500 296.850 485.100 ;
        RECT 278.550 483.600 279.450 484.500 ;
        RECT 288.450 484.200 296.850 484.500 ;
        RECT 278.550 481.800 280.950 483.600 ;
        RECT 279.150 471.600 280.950 481.800 ;
        RECT 282.150 471.000 283.950 483.600 ;
        RECT 293.250 482.700 295.050 483.300 ;
        RECT 287.250 481.500 295.050 482.700 ;
        RECT 295.950 482.100 296.850 484.200 ;
        RECT 298.950 484.200 299.850 496.800 ;
        RECT 311.250 493.050 312.450 500.400 ;
        RECT 326.100 501.300 327.900 506.400 ;
        RECT 329.100 502.200 330.900 507.000 ;
        RECT 332.100 501.300 333.900 506.400 ;
        RECT 326.100 499.950 333.900 501.300 ;
        RECT 335.100 500.400 336.900 506.400 ;
        RECT 339.150 502.200 340.950 506.400 ;
        RECT 338.550 500.400 340.950 502.200 ;
        RECT 342.150 500.400 343.950 507.000 ;
        RECT 346.950 504.300 348.750 506.400 ;
        RECT 345.150 503.400 348.750 504.300 ;
        RECT 351.450 503.400 353.250 507.000 ;
        RECT 354.750 503.400 356.550 506.400 ;
        RECT 357.750 503.400 359.550 507.000 ;
        RECT 362.250 503.400 364.050 506.400 ;
        RECT 344.850 502.800 348.750 503.400 ;
        RECT 344.850 501.300 346.950 502.800 ;
        RECT 354.750 502.500 355.800 503.400 ;
        RECT 335.100 498.300 336.300 500.400 ;
        RECT 332.700 497.400 336.300 498.300 ;
        RECT 329.100 493.050 330.900 494.850 ;
        RECT 332.700 493.050 333.900 497.400 ;
        RECT 335.100 493.050 336.900 494.850 ;
        RECT 306.150 491.250 312.450 493.050 ;
        RECT 307.950 490.950 312.450 491.250 ;
        RECT 325.950 490.950 328.050 493.050 ;
        RECT 328.950 490.950 331.050 493.050 ;
        RECT 331.950 490.950 334.050 493.050 ;
        RECT 334.950 490.950 337.050 493.050 ;
        RECT 302.550 488.100 304.650 488.400 ;
        RECT 308.550 488.100 310.350 488.250 ;
        RECT 302.550 486.900 310.350 488.100 ;
        RECT 302.550 486.300 304.650 486.900 ;
        RECT 308.550 486.450 310.350 486.900 ;
        RECT 298.950 483.300 303.750 484.200 ;
        RECT 311.250 483.600 312.450 490.950 ;
        RECT 326.100 489.150 327.900 490.950 ;
        RECT 332.700 483.600 333.900 490.950 ;
        RECT 302.550 482.400 303.750 483.300 ;
        RECT 299.850 482.100 301.650 482.400 ;
        RECT 287.250 480.600 289.350 481.500 ;
        RECT 295.950 481.200 301.650 482.100 ;
        RECT 299.850 480.600 301.650 481.200 ;
        RECT 302.550 480.600 305.550 482.400 ;
        RECT 287.550 471.600 289.350 480.600 ;
        RECT 291.450 479.550 293.250 480.300 ;
        RECT 296.250 479.550 298.050 480.300 ;
        RECT 291.450 478.500 298.050 479.550 ;
        RECT 292.350 471.000 294.150 477.600 ;
        RECT 295.350 471.600 297.150 478.500 ;
        RECT 302.550 477.600 304.650 479.700 ;
        RECT 298.350 471.000 300.150 477.600 ;
        RECT 302.850 471.600 304.650 477.600 ;
        RECT 307.650 471.000 309.450 483.600 ;
        RECT 310.650 471.600 312.450 483.600 ;
        RECT 326.400 471.000 328.200 483.600 ;
        RECT 331.500 482.100 333.900 483.600 ;
        RECT 338.550 485.700 339.450 500.400 ;
        RECT 347.850 499.800 349.650 501.600 ;
        RECT 350.850 501.450 355.800 502.500 ;
        RECT 350.850 500.700 352.650 501.450 ;
        RECT 362.250 501.300 364.650 503.400 ;
        RECT 367.350 500.400 369.150 507.000 ;
        RECT 370.650 500.400 372.450 506.400 ;
        RECT 386.100 500.400 387.900 506.400 ;
        RECT 347.850 498.000 348.900 499.800 ;
        RECT 358.050 498.000 359.850 498.600 ;
        RECT 347.850 496.800 359.850 498.000 ;
        RECT 340.950 495.600 348.900 496.800 ;
        RECT 340.950 493.050 342.750 495.600 ;
        RECT 347.100 495.000 348.900 495.600 ;
        RECT 344.100 493.800 345.900 494.400 ;
        RECT 340.950 490.950 343.050 493.050 ;
        RECT 344.100 492.600 352.200 493.800 ;
        RECT 350.100 490.950 352.200 492.600 ;
        RECT 348.450 485.700 350.250 486.000 ;
        RECT 338.550 485.100 350.250 485.700 ;
        RECT 338.550 484.500 356.850 485.100 ;
        RECT 338.550 483.600 339.450 484.500 ;
        RECT 348.450 484.200 356.850 484.500 ;
        RECT 331.500 471.600 333.300 482.100 ;
        RECT 338.550 481.800 340.950 483.600 ;
        RECT 334.200 479.100 336.000 480.900 ;
        RECT 334.500 471.000 336.300 477.600 ;
        RECT 339.150 471.600 340.950 481.800 ;
        RECT 342.150 471.000 343.950 483.600 ;
        RECT 353.250 482.700 355.050 483.300 ;
        RECT 347.250 481.500 355.050 482.700 ;
        RECT 355.950 482.100 356.850 484.200 ;
        RECT 358.950 484.200 359.850 496.800 ;
        RECT 371.250 493.050 372.450 500.400 ;
        RECT 386.700 498.300 387.900 500.400 ;
        RECT 389.100 501.300 390.900 506.400 ;
        RECT 392.100 502.200 393.900 507.000 ;
        RECT 395.100 501.300 396.900 506.400 ;
        RECT 389.100 499.950 396.900 501.300 ;
        RECT 410.100 500.400 411.900 506.400 ;
        RECT 413.100 500.400 414.900 507.000 ;
        RECT 416.100 503.400 417.900 506.400 ;
        RECT 386.700 497.400 390.300 498.300 ;
        RECT 386.100 493.050 387.900 494.850 ;
        RECT 389.100 493.050 390.300 497.400 ;
        RECT 392.100 493.050 393.900 494.850 ;
        RECT 410.100 493.050 411.300 500.400 ;
        RECT 416.700 499.500 417.900 503.400 ;
        RECT 431.100 501.300 432.900 506.400 ;
        RECT 434.100 502.200 435.900 507.000 ;
        RECT 437.100 501.300 438.900 506.400 ;
        RECT 431.100 499.950 438.900 501.300 ;
        RECT 440.100 500.400 441.900 506.400 ;
        RECT 455.400 500.400 457.200 507.000 ;
        RECT 412.200 498.600 417.900 499.500 ;
        RECT 412.200 497.700 414.000 498.600 ;
        RECT 440.100 498.300 441.300 500.400 ;
        RECT 460.500 499.200 462.300 506.400 ;
        RECT 366.150 491.250 372.450 493.050 ;
        RECT 367.950 490.950 372.450 491.250 ;
        RECT 385.950 490.950 388.050 493.050 ;
        RECT 388.950 490.950 391.050 493.050 ;
        RECT 391.950 490.950 394.050 493.050 ;
        RECT 394.950 490.950 397.050 493.050 ;
        RECT 410.100 490.950 412.200 493.050 ;
        RECT 362.550 488.100 364.650 488.400 ;
        RECT 368.550 488.100 370.350 488.250 ;
        RECT 362.550 486.900 370.350 488.100 ;
        RECT 362.550 486.300 364.650 486.900 ;
        RECT 368.550 486.450 370.350 486.900 ;
        RECT 358.950 483.300 363.750 484.200 ;
        RECT 371.250 483.600 372.450 490.950 ;
        RECT 362.550 482.400 363.750 483.300 ;
        RECT 359.850 482.100 361.650 482.400 ;
        RECT 347.250 480.600 349.350 481.500 ;
        RECT 355.950 481.200 361.650 482.100 ;
        RECT 359.850 480.600 361.650 481.200 ;
        RECT 362.550 480.600 365.550 482.400 ;
        RECT 347.550 471.600 349.350 480.600 ;
        RECT 351.450 479.550 353.250 480.300 ;
        RECT 356.250 479.550 358.050 480.300 ;
        RECT 351.450 478.500 358.050 479.550 ;
        RECT 352.350 471.000 354.150 477.600 ;
        RECT 355.350 471.600 357.150 478.500 ;
        RECT 362.550 477.600 364.650 479.700 ;
        RECT 358.350 471.000 360.150 477.600 ;
        RECT 362.850 471.600 364.650 477.600 ;
        RECT 367.650 471.000 369.450 483.600 ;
        RECT 370.650 471.600 372.450 483.600 ;
        RECT 389.100 483.600 390.300 490.950 ;
        RECT 395.100 489.150 396.900 490.950 ;
        RECT 410.100 483.600 411.300 490.950 ;
        RECT 413.100 486.300 414.000 497.700 ;
        RECT 437.700 497.400 441.300 498.300 ;
        RECT 458.100 498.300 462.300 499.200 ;
        RECT 476.100 500.400 477.900 506.400 ;
        RECT 479.100 500.400 480.900 507.000 ;
        RECT 482.100 503.400 483.900 506.400 ;
        RECT 434.100 493.050 435.900 494.850 ;
        RECT 437.700 493.050 438.900 497.400 ;
        RECT 440.100 493.050 441.900 494.850 ;
        RECT 455.250 493.050 457.050 494.850 ;
        RECT 458.100 493.050 459.300 498.300 ;
        RECT 461.100 493.050 462.900 494.850 ;
        RECT 476.100 493.050 477.300 500.400 ;
        RECT 482.700 499.500 483.900 503.400 ;
        RECT 478.200 498.600 483.900 499.500 ;
        RECT 500.100 503.400 501.900 506.400 ;
        RECT 500.100 499.500 501.300 503.400 ;
        RECT 503.100 500.400 504.900 507.000 ;
        RECT 506.100 500.400 507.900 506.400 ;
        RECT 521.100 500.400 522.900 507.000 ;
        RECT 524.100 500.400 525.900 506.400 ;
        RECT 527.100 500.400 528.900 507.000 ;
        RECT 530.100 500.400 531.900 506.400 ;
        RECT 533.100 500.400 534.900 507.000 ;
        RECT 551.100 503.400 552.900 506.400 ;
        RECT 554.100 503.400 555.900 507.000 ;
        RECT 500.100 498.600 505.800 499.500 ;
        RECT 478.200 497.700 480.000 498.600 ;
        RECT 415.500 490.950 417.600 493.050 ;
        RECT 430.950 490.950 433.050 493.050 ;
        RECT 433.950 490.950 436.050 493.050 ;
        RECT 436.950 490.950 439.050 493.050 ;
        RECT 439.950 490.950 442.050 493.050 ;
        RECT 454.950 490.950 457.050 493.050 ;
        RECT 457.950 490.950 460.050 493.050 ;
        RECT 460.950 490.950 463.050 493.050 ;
        RECT 476.100 490.950 478.200 493.050 ;
        RECT 415.800 489.150 417.600 490.950 ;
        RECT 431.100 489.150 432.900 490.950 ;
        RECT 412.200 485.400 414.000 486.300 ;
        RECT 412.200 484.500 417.900 485.400 ;
        RECT 389.100 482.100 391.500 483.600 ;
        RECT 387.000 479.100 388.800 480.900 ;
        RECT 386.700 471.000 388.500 477.600 ;
        RECT 389.700 471.600 391.500 482.100 ;
        RECT 394.800 471.000 396.600 483.600 ;
        RECT 410.100 471.600 411.900 483.600 ;
        RECT 413.100 471.000 414.900 481.800 ;
        RECT 416.700 477.600 417.900 484.500 ;
        RECT 437.700 483.600 438.900 490.950 ;
        RECT 416.100 471.600 417.900 477.600 ;
        RECT 431.400 471.000 433.200 483.600 ;
        RECT 436.500 482.100 438.900 483.600 ;
        RECT 436.500 471.600 438.300 482.100 ;
        RECT 439.200 479.100 441.000 480.900 ;
        RECT 458.100 477.600 459.300 490.950 ;
        RECT 476.100 483.600 477.300 490.950 ;
        RECT 479.100 486.300 480.000 497.700 ;
        RECT 504.000 497.700 505.800 498.600 ;
        RECT 481.500 490.950 483.600 493.050 ;
        RECT 481.800 489.150 483.600 490.950 ;
        RECT 500.400 490.950 502.500 493.050 ;
        RECT 500.400 489.150 502.200 490.950 ;
        RECT 478.200 485.400 480.000 486.300 ;
        RECT 504.000 486.300 504.900 497.700 ;
        RECT 506.700 493.050 507.900 500.400 ;
        RECT 524.700 499.500 525.900 500.400 ;
        RECT 530.700 499.500 531.900 500.400 ;
        RECT 524.700 498.300 531.900 499.500 ;
        RECT 524.700 493.050 525.900 498.300 ;
        RECT 551.700 493.050 552.900 503.400 ;
        RECT 557.550 500.400 559.350 506.400 ;
        RECT 560.850 500.400 562.650 507.000 ;
        RECT 565.950 503.400 567.750 506.400 ;
        RECT 570.450 503.400 572.250 507.000 ;
        RECT 573.450 503.400 575.250 506.400 ;
        RECT 576.750 503.400 578.550 507.000 ;
        RECT 581.250 504.300 583.050 506.400 ;
        RECT 581.250 503.400 584.850 504.300 ;
        RECT 565.350 501.300 567.750 503.400 ;
        RECT 574.200 502.500 575.250 503.400 ;
        RECT 581.250 502.800 585.150 503.400 ;
        RECT 574.200 501.450 579.150 502.500 ;
        RECT 577.350 500.700 579.150 501.450 ;
        RECT 557.550 493.050 558.750 500.400 ;
        RECT 580.350 499.800 582.150 501.600 ;
        RECT 583.050 501.300 585.150 502.800 ;
        RECT 586.050 500.400 587.850 507.000 ;
        RECT 589.050 502.200 590.850 506.400 ;
        RECT 589.050 500.400 591.450 502.200 ;
        RECT 608.100 500.400 609.900 506.400 ;
        RECT 570.150 498.000 571.950 498.600 ;
        RECT 581.100 498.000 582.150 499.800 ;
        RECT 570.150 496.800 582.150 498.000 ;
        RECT 505.800 490.950 507.900 493.050 ;
        RECT 523.800 490.950 525.900 493.050 ;
        RECT 529.800 490.950 531.900 493.050 ;
        RECT 550.950 490.950 553.050 493.050 ;
        RECT 553.950 490.950 556.050 493.050 ;
        RECT 557.550 491.250 563.850 493.050 ;
        RECT 557.550 490.950 562.050 491.250 ;
        RECT 504.000 485.400 505.800 486.300 ;
        RECT 478.200 484.500 483.900 485.400 ;
        RECT 439.500 471.000 441.300 477.600 ;
        RECT 455.100 471.000 456.900 477.600 ;
        RECT 458.100 471.600 459.900 477.600 ;
        RECT 461.100 471.000 462.900 477.600 ;
        RECT 476.100 471.600 477.900 483.600 ;
        RECT 479.100 471.000 480.900 481.800 ;
        RECT 482.700 477.600 483.900 484.500 ;
        RECT 482.100 471.600 483.900 477.600 ;
        RECT 500.100 484.500 505.800 485.400 ;
        RECT 500.100 477.600 501.300 484.500 ;
        RECT 506.700 483.600 507.900 490.950 ;
        RECT 524.700 485.400 525.900 490.950 ;
        RECT 530.100 489.150 531.900 490.950 ;
        RECT 524.700 484.500 531.900 485.400 ;
        RECT 524.700 483.600 525.900 484.500 ;
        RECT 500.100 471.600 501.900 477.600 ;
        RECT 503.100 471.000 504.900 481.800 ;
        RECT 506.100 471.600 507.900 483.600 ;
        RECT 521.100 471.000 522.900 483.600 ;
        RECT 524.100 471.600 525.900 483.600 ;
        RECT 527.100 471.000 528.900 483.600 ;
        RECT 530.100 471.600 531.900 484.500 ;
        RECT 533.100 471.000 534.900 483.600 ;
        RECT 551.700 477.600 552.900 490.950 ;
        RECT 554.100 489.150 555.900 490.950 ;
        RECT 557.550 483.600 558.750 490.950 ;
        RECT 559.650 488.100 561.450 488.250 ;
        RECT 565.350 488.100 567.450 488.400 ;
        RECT 559.650 486.900 567.450 488.100 ;
        RECT 559.650 486.450 561.450 486.900 ;
        RECT 565.350 486.300 567.450 486.900 ;
        RECT 570.150 484.200 571.050 496.800 ;
        RECT 581.100 495.600 589.050 496.800 ;
        RECT 581.100 495.000 582.900 495.600 ;
        RECT 584.100 493.800 585.900 494.400 ;
        RECT 577.800 492.600 585.900 493.800 ;
        RECT 587.250 493.050 589.050 495.600 ;
        RECT 577.800 490.950 579.900 492.600 ;
        RECT 586.950 490.950 589.050 493.050 ;
        RECT 579.750 485.700 581.550 486.000 ;
        RECT 590.550 485.700 591.450 500.400 ;
        RECT 608.700 498.300 609.900 500.400 ;
        RECT 611.100 501.300 612.900 506.400 ;
        RECT 614.100 502.200 615.900 507.000 ;
        RECT 617.100 501.300 618.900 506.400 ;
        RECT 632.100 503.400 633.900 506.400 ;
        RECT 635.100 503.400 636.900 507.000 ;
        RECT 650.100 503.400 651.900 507.000 ;
        RECT 653.100 503.400 654.900 506.400 ;
        RECT 656.100 503.400 657.900 507.000 ;
        RECT 611.100 499.950 618.900 501.300 ;
        RECT 608.700 497.400 612.300 498.300 ;
        RECT 608.100 493.050 609.900 494.850 ;
        RECT 611.100 493.050 612.300 497.400 ;
        RECT 614.100 493.050 615.900 494.850 ;
        RECT 632.700 493.050 633.900 503.400 ;
        RECT 653.400 493.050 654.300 503.400 ;
        RECT 671.400 500.400 673.200 507.000 ;
        RECT 676.500 499.200 678.300 506.400 ;
        RECT 674.100 498.300 678.300 499.200 ;
        RECT 695.100 498.600 696.900 506.400 ;
        RECT 699.600 500.400 701.400 507.000 ;
        RECT 702.600 502.200 704.400 506.400 ;
        RECT 723.600 502.200 725.400 506.400 ;
        RECT 702.600 500.400 705.300 502.200 ;
        RECT 701.700 498.600 703.500 499.500 ;
        RECT 671.250 493.050 673.050 494.850 ;
        RECT 674.100 493.050 675.300 498.300 ;
        RECT 695.100 497.700 703.500 498.600 ;
        RECT 677.100 493.050 678.900 494.850 ;
        RECT 695.250 493.050 697.050 494.850 ;
        RECT 607.950 490.950 610.050 493.050 ;
        RECT 610.950 490.950 613.050 493.050 ;
        RECT 613.950 490.950 616.050 493.050 ;
        RECT 616.950 490.950 619.050 493.050 ;
        RECT 631.950 490.950 634.050 493.050 ;
        RECT 634.950 490.950 637.050 493.050 ;
        RECT 649.950 490.950 652.050 493.050 ;
        RECT 652.950 490.950 655.050 493.050 ;
        RECT 655.950 490.950 658.050 493.050 ;
        RECT 670.950 490.950 673.050 493.050 ;
        RECT 673.950 490.950 676.050 493.050 ;
        RECT 676.950 490.950 679.050 493.050 ;
        RECT 695.100 490.950 697.200 493.050 ;
        RECT 579.750 485.100 591.450 485.700 ;
        RECT 551.100 471.600 552.900 477.600 ;
        RECT 554.100 471.000 555.900 477.600 ;
        RECT 557.550 471.600 559.350 483.600 ;
        RECT 560.550 471.000 562.350 483.600 ;
        RECT 566.250 483.300 571.050 484.200 ;
        RECT 573.150 484.500 591.450 485.100 ;
        RECT 573.150 484.200 581.550 484.500 ;
        RECT 566.250 482.400 567.450 483.300 ;
        RECT 564.450 480.600 567.450 482.400 ;
        RECT 568.350 482.100 570.150 482.400 ;
        RECT 573.150 482.100 574.050 484.200 ;
        RECT 590.550 483.600 591.450 484.500 ;
        RECT 568.350 481.200 574.050 482.100 ;
        RECT 574.950 482.700 576.750 483.300 ;
        RECT 574.950 481.500 582.750 482.700 ;
        RECT 568.350 480.600 570.150 481.200 ;
        RECT 580.650 480.600 582.750 481.500 ;
        RECT 565.350 477.600 567.450 479.700 ;
        RECT 571.950 479.550 573.750 480.300 ;
        RECT 576.750 479.550 578.550 480.300 ;
        RECT 571.950 478.500 578.550 479.550 ;
        RECT 565.350 471.600 567.150 477.600 ;
        RECT 569.850 471.000 571.650 477.600 ;
        RECT 572.850 471.600 574.650 478.500 ;
        RECT 575.850 471.000 577.650 477.600 ;
        RECT 580.650 471.600 582.450 480.600 ;
        RECT 586.050 471.000 587.850 483.600 ;
        RECT 589.050 481.800 591.450 483.600 ;
        RECT 611.100 483.600 612.300 490.950 ;
        RECT 617.100 489.150 618.900 490.950 ;
        RECT 611.100 482.100 613.500 483.600 ;
        RECT 589.050 471.600 590.850 481.800 ;
        RECT 609.000 479.100 610.800 480.900 ;
        RECT 608.700 471.000 610.500 477.600 ;
        RECT 611.700 471.600 613.500 482.100 ;
        RECT 616.800 471.000 618.600 483.600 ;
        RECT 632.700 477.600 633.900 490.950 ;
        RECT 635.100 489.150 636.900 490.950 ;
        RECT 650.250 489.150 652.050 490.950 ;
        RECT 653.400 483.600 654.300 490.950 ;
        RECT 656.100 489.150 657.900 490.950 ;
        RECT 632.100 471.600 633.900 477.600 ;
        RECT 635.100 471.000 636.900 477.600 ;
        RECT 650.100 471.000 651.900 483.600 ;
        RECT 653.400 482.400 657.000 483.600 ;
        RECT 655.200 471.600 657.000 482.400 ;
        RECT 674.100 477.600 675.300 490.950 ;
        RECT 688.950 486.450 691.050 487.050 ;
        RECT 694.950 486.450 697.050 487.050 ;
        RECT 688.950 485.550 697.050 486.450 ;
        RECT 688.950 484.950 691.050 485.550 ;
        RECT 694.950 484.950 697.050 485.550 ;
        RECT 698.100 477.600 699.000 497.700 ;
        RECT 704.400 493.050 705.300 500.400 ;
        RECT 722.700 500.400 725.400 502.200 ;
        RECT 726.600 500.400 728.400 507.000 ;
        RECT 722.700 493.050 723.600 500.400 ;
        RECT 724.500 498.600 726.300 499.500 ;
        RECT 731.100 498.600 732.900 506.400 ;
        RECT 749.400 500.400 751.200 507.000 ;
        RECT 754.500 499.200 756.300 506.400 ;
        RECT 770.100 503.400 771.900 507.000 ;
        RECT 773.100 503.400 774.900 506.400 ;
        RECT 724.500 497.700 732.900 498.600 ;
        RECT 752.100 498.300 756.300 499.200 ;
        RECT 700.500 490.950 702.600 493.050 ;
        RECT 703.800 490.950 705.900 493.050 ;
        RECT 722.100 490.950 724.200 493.050 ;
        RECT 725.400 490.950 727.500 493.050 ;
        RECT 700.200 489.150 702.000 490.950 ;
        RECT 704.400 483.600 705.300 490.950 ;
        RECT 722.700 483.600 723.600 490.950 ;
        RECT 726.000 489.150 727.800 490.950 ;
        RECT 671.100 471.000 672.900 477.600 ;
        RECT 674.100 471.600 675.900 477.600 ;
        RECT 677.100 471.000 678.900 477.600 ;
        RECT 695.100 471.000 696.900 477.600 ;
        RECT 698.100 471.600 699.900 477.600 ;
        RECT 701.100 471.000 702.900 483.000 ;
        RECT 704.100 471.600 705.900 483.600 ;
        RECT 722.100 471.600 723.900 483.600 ;
        RECT 725.100 471.000 726.900 483.000 ;
        RECT 729.000 477.600 729.900 497.700 ;
        RECT 730.950 493.050 732.750 494.850 ;
        RECT 749.250 493.050 751.050 494.850 ;
        RECT 752.100 493.050 753.300 498.300 ;
        RECT 755.100 493.050 756.900 494.850 ;
        RECT 773.100 493.050 774.300 503.400 ;
        RECT 788.100 501.300 789.900 506.400 ;
        RECT 791.100 502.200 792.900 507.000 ;
        RECT 794.100 501.300 795.900 506.400 ;
        RECT 788.100 499.950 795.900 501.300 ;
        RECT 797.100 500.400 798.900 506.400 ;
        RECT 797.100 498.300 798.300 500.400 ;
        RECT 794.700 497.400 798.300 498.300 ;
        RECT 812.100 497.400 813.900 507.000 ;
        RECT 818.700 498.000 820.500 506.400 ;
        RECT 839.400 500.400 841.200 507.000 ;
        RECT 844.500 499.200 846.300 506.400 ;
        RECT 842.100 498.300 846.300 499.200 ;
        RECT 863.100 498.600 864.900 506.400 ;
        RECT 867.600 500.400 869.400 507.000 ;
        RECT 870.600 502.200 872.400 506.400 ;
        RECT 870.600 500.400 873.300 502.200 ;
        RECT 869.700 498.600 871.500 499.500 ;
        RECT 791.100 493.050 792.900 494.850 ;
        RECT 794.700 493.050 795.900 497.400 ;
        RECT 818.700 496.800 822.000 498.000 ;
        RECT 797.100 493.050 798.900 494.850 ;
        RECT 812.100 493.050 813.900 494.850 ;
        RECT 818.100 493.050 819.900 494.850 ;
        RECT 821.100 493.050 822.000 496.800 ;
        RECT 839.250 493.050 841.050 494.850 ;
        RECT 842.100 493.050 843.300 498.300 ;
        RECT 863.100 497.700 871.500 498.600 ;
        RECT 845.100 493.050 846.900 494.850 ;
        RECT 863.250 493.050 865.050 494.850 ;
        RECT 730.800 490.950 732.900 493.050 ;
        RECT 748.950 490.950 751.050 493.050 ;
        RECT 751.950 490.950 754.050 493.050 ;
        RECT 754.950 490.950 757.050 493.050 ;
        RECT 769.950 490.950 772.050 493.050 ;
        RECT 772.950 490.950 775.050 493.050 ;
        RECT 787.950 490.950 790.050 493.050 ;
        RECT 790.950 490.950 793.050 493.050 ;
        RECT 793.950 490.950 796.050 493.050 ;
        RECT 796.950 490.950 799.050 493.050 ;
        RECT 811.950 490.950 814.050 493.050 ;
        RECT 814.950 490.950 817.050 493.050 ;
        RECT 817.950 490.950 820.050 493.050 ;
        RECT 820.950 490.950 823.050 493.050 ;
        RECT 838.950 490.950 841.050 493.050 ;
        RECT 841.950 490.950 844.050 493.050 ;
        RECT 844.950 490.950 847.050 493.050 ;
        RECT 863.100 490.950 865.200 493.050 ;
        RECT 733.950 480.450 736.050 481.050 ;
        RECT 748.950 480.450 751.050 481.050 ;
        RECT 733.950 479.550 751.050 480.450 ;
        RECT 733.950 478.950 736.050 479.550 ;
        RECT 748.950 478.950 751.050 479.550 ;
        RECT 752.100 477.600 753.300 490.950 ;
        RECT 770.100 489.150 771.900 490.950 ;
        RECT 773.100 477.600 774.300 490.950 ;
        RECT 788.100 489.150 789.900 490.950 ;
        RECT 794.700 483.600 795.900 490.950 ;
        RECT 815.100 489.150 816.900 490.950 ;
        RECT 796.950 486.450 799.050 487.050 ;
        RECT 817.950 486.450 820.050 487.050 ;
        RECT 796.950 485.550 820.050 486.450 ;
        RECT 796.950 484.950 799.050 485.550 ;
        RECT 817.950 484.950 820.050 485.550 ;
        RECT 728.100 471.600 729.900 477.600 ;
        RECT 731.100 471.000 732.900 477.600 ;
        RECT 749.100 471.000 750.900 477.600 ;
        RECT 752.100 471.600 753.900 477.600 ;
        RECT 755.100 471.000 756.900 477.600 ;
        RECT 770.100 471.000 771.900 477.600 ;
        RECT 773.100 471.600 774.900 477.600 ;
        RECT 788.400 471.000 790.200 483.600 ;
        RECT 793.500 482.100 795.900 483.600 ;
        RECT 793.500 471.600 795.300 482.100 ;
        RECT 796.200 479.100 798.000 480.900 ;
        RECT 821.100 478.800 822.000 490.950 ;
        RECT 815.400 477.900 822.000 478.800 ;
        RECT 815.400 477.600 816.900 477.900 ;
        RECT 796.500 471.000 798.300 477.600 ;
        RECT 812.100 471.000 813.900 477.600 ;
        RECT 815.100 471.600 816.900 477.600 ;
        RECT 821.100 477.600 822.000 477.900 ;
        RECT 842.100 477.600 843.300 490.950 ;
        RECT 850.950 486.450 853.050 487.050 ;
        RECT 859.950 486.450 862.050 486.900 ;
        RECT 850.950 485.550 862.050 486.450 ;
        RECT 850.950 484.950 853.050 485.550 ;
        RECT 859.950 484.800 862.050 485.550 ;
        RECT 866.100 477.600 867.000 497.700 ;
        RECT 872.400 493.050 873.300 500.400 ;
        RECT 874.950 498.450 877.050 502.050 ;
        RECT 888.000 500.400 889.800 507.000 ;
        RECT 892.500 501.600 894.300 506.400 ;
        RECT 895.500 503.400 897.300 507.000 ;
        RECT 892.500 500.400 897.600 501.600 ;
        RECT 874.950 498.000 879.450 498.450 ;
        RECT 875.550 497.550 879.450 498.000 ;
        RECT 868.500 490.950 870.600 493.050 ;
        RECT 871.800 490.950 873.900 493.050 ;
        RECT 868.200 489.150 870.000 490.950 ;
        RECT 872.400 483.600 873.300 490.950 ;
        RECT 878.550 486.900 879.450 497.550 ;
        RECT 887.100 493.050 888.900 494.850 ;
        RECT 893.250 493.050 895.050 494.850 ;
        RECT 896.700 493.050 897.600 500.400 ;
        RECT 911.100 501.300 912.900 506.400 ;
        RECT 914.100 502.200 915.900 507.000 ;
        RECT 917.100 501.300 918.900 506.400 ;
        RECT 911.100 499.950 918.900 501.300 ;
        RECT 920.100 500.400 921.900 506.400 ;
        RECT 920.100 498.300 921.300 500.400 ;
        RECT 917.700 497.400 921.300 498.300 ;
        RECT 935.100 497.400 936.900 507.000 ;
        RECT 941.700 498.000 943.500 506.400 ;
        RECT 959.700 503.400 961.500 507.000 ;
        RECT 962.700 501.600 964.500 506.400 ;
        RECT 959.400 500.400 964.500 501.600 ;
        RECT 967.200 500.400 969.000 507.000 ;
        RECT 906.000 495.450 910.050 496.050 ;
        RECT 905.550 493.950 910.050 495.450 ;
        RECT 886.950 490.950 889.050 493.050 ;
        RECT 889.950 490.950 892.050 493.050 ;
        RECT 892.950 490.950 895.050 493.050 ;
        RECT 895.950 490.950 898.050 493.050 ;
        RECT 890.250 489.150 892.050 490.950 ;
        RECT 877.950 484.800 880.050 486.900 ;
        RECT 896.700 483.600 897.600 490.950 ;
        RECT 905.550 490.050 906.450 493.950 ;
        RECT 914.100 493.050 915.900 494.850 ;
        RECT 917.700 493.050 918.900 497.400 ;
        RECT 941.700 496.800 945.000 498.000 ;
        RECT 922.950 495.450 927.000 496.050 ;
        RECT 920.100 493.050 921.900 494.850 ;
        RECT 922.950 493.950 927.450 495.450 ;
        RECT 910.950 490.950 913.050 493.050 ;
        RECT 913.950 490.950 916.050 493.050 ;
        RECT 916.950 490.950 919.050 493.050 ;
        RECT 919.950 490.950 922.050 493.050 ;
        RECT 903.000 489.900 906.450 490.050 ;
        RECT 901.950 488.550 906.450 489.900 ;
        RECT 911.100 489.150 912.900 490.950 ;
        RECT 901.950 487.950 906.000 488.550 ;
        RECT 901.950 487.800 904.050 487.950 ;
        RECT 917.700 483.600 918.900 490.950 ;
        RECT 926.550 486.900 927.450 493.950 ;
        RECT 935.100 493.050 936.900 494.850 ;
        RECT 941.100 493.050 942.900 494.850 ;
        RECT 944.100 493.050 945.000 496.800 ;
        RECT 954.000 495.450 958.050 496.050 ;
        RECT 953.550 493.950 958.050 495.450 ;
        RECT 934.950 490.950 937.050 493.050 ;
        RECT 937.950 490.950 940.050 493.050 ;
        RECT 940.950 490.950 943.050 493.050 ;
        RECT 943.950 490.950 946.050 493.050 ;
        RECT 938.100 489.150 939.900 490.950 ;
        RECT 925.950 484.800 928.050 486.900 ;
        RECT 818.100 471.000 819.900 477.000 ;
        RECT 821.100 471.600 822.900 477.600 ;
        RECT 839.100 471.000 840.900 477.600 ;
        RECT 842.100 471.600 843.900 477.600 ;
        RECT 845.100 471.000 846.900 477.600 ;
        RECT 863.100 471.000 864.900 477.600 ;
        RECT 866.100 471.600 867.900 477.600 ;
        RECT 869.100 471.000 870.900 483.000 ;
        RECT 872.100 471.600 873.900 483.600 ;
        RECT 887.100 482.700 894.900 483.600 ;
        RECT 887.100 471.600 888.900 482.700 ;
        RECT 890.100 471.000 891.900 481.800 ;
        RECT 893.100 471.600 894.900 482.700 ;
        RECT 896.100 471.600 897.900 483.600 ;
        RECT 911.400 471.000 913.200 483.600 ;
        RECT 916.500 482.100 918.900 483.600 ;
        RECT 916.500 471.600 918.300 482.100 ;
        RECT 919.200 479.100 921.000 480.900 ;
        RECT 944.100 478.800 945.000 490.950 ;
        RECT 946.950 489.450 949.050 490.050 ;
        RECT 953.550 489.450 954.450 493.950 ;
        RECT 959.400 493.050 960.300 500.400 ;
        RECT 986.100 497.400 987.900 507.000 ;
        RECT 992.700 498.000 994.500 506.400 ;
        RECT 997.950 504.450 1000.050 505.050 ;
        RECT 1009.950 504.450 1012.050 504.900 ;
        RECT 997.950 503.550 1012.050 504.450 ;
        RECT 997.950 502.950 1000.050 503.550 ;
        RECT 1009.950 502.800 1012.050 503.550 ;
        RECT 992.700 496.800 996.000 498.000 ;
        RECT 981.000 495.450 985.050 496.050 ;
        RECT 961.950 493.050 963.750 494.850 ;
        RECT 968.100 493.050 969.900 494.850 ;
        RECT 980.550 493.950 985.050 495.450 ;
        RECT 958.950 490.950 961.050 493.050 ;
        RECT 961.950 490.950 964.050 493.050 ;
        RECT 964.950 490.950 967.050 493.050 ;
        RECT 967.950 490.950 970.050 493.050 ;
        RECT 946.950 488.550 954.450 489.450 ;
        RECT 946.950 487.950 949.050 488.550 ;
        RECT 959.400 483.600 960.300 490.950 ;
        RECT 964.950 489.150 966.750 490.950 ;
        RECT 980.550 490.050 981.450 493.950 ;
        RECT 986.100 493.050 987.900 494.850 ;
        RECT 992.100 493.050 993.900 494.850 ;
        RECT 995.100 493.050 996.000 496.800 ;
        RECT 985.950 490.950 988.050 493.050 ;
        RECT 988.950 490.950 991.050 493.050 ;
        RECT 991.950 490.950 994.050 493.050 ;
        RECT 994.950 490.950 997.050 493.050 ;
        RECT 980.550 488.550 985.050 490.050 ;
        RECT 989.100 489.150 990.900 490.950 ;
        RECT 981.000 487.950 985.050 488.550 ;
        RECT 973.950 486.450 976.050 487.050 ;
        RECT 985.950 486.450 988.050 486.750 ;
        RECT 973.950 485.550 988.050 486.450 ;
        RECT 973.950 484.950 976.050 485.550 ;
        RECT 985.950 484.650 988.050 485.550 ;
        RECT 938.400 477.900 945.000 478.800 ;
        RECT 938.400 477.600 939.900 477.900 ;
        RECT 919.500 471.000 921.300 477.600 ;
        RECT 935.100 471.000 936.900 477.600 ;
        RECT 938.100 471.600 939.900 477.600 ;
        RECT 944.100 477.600 945.000 477.900 ;
        RECT 941.100 471.000 942.900 477.000 ;
        RECT 944.100 471.600 945.900 477.600 ;
        RECT 959.100 471.600 960.900 483.600 ;
        RECT 962.100 482.700 969.900 483.600 ;
        RECT 962.100 471.600 963.900 482.700 ;
        RECT 965.100 471.000 966.900 481.800 ;
        RECT 968.100 471.600 969.900 482.700 ;
        RECT 995.100 478.800 996.000 490.950 ;
        RECT 989.400 477.900 996.000 478.800 ;
        RECT 989.400 477.600 990.900 477.900 ;
        RECT 986.100 471.000 987.900 477.600 ;
        RECT 989.100 471.600 990.900 477.600 ;
        RECT 995.100 477.600 996.000 477.900 ;
        RECT 992.100 471.000 993.900 477.000 ;
        RECT 995.100 471.600 996.900 477.600 ;
        RECT 17.100 455.400 18.900 467.400 ;
        RECT 20.100 457.200 21.900 468.000 ;
        RECT 23.100 461.400 24.900 467.400 ;
        RECT 17.100 448.050 18.300 455.400 ;
        RECT 23.700 454.500 24.900 461.400 ;
        RECT 19.200 453.600 24.900 454.500 ;
        RECT 38.100 455.400 39.900 467.400 ;
        RECT 41.100 457.200 42.900 468.000 ;
        RECT 44.100 461.400 45.900 467.400 ;
        RECT 19.200 452.700 21.000 453.600 ;
        RECT 17.100 445.950 19.200 448.050 ;
        RECT 17.100 438.600 18.300 445.950 ;
        RECT 20.100 441.300 21.000 452.700 ;
        RECT 22.800 448.050 24.600 449.850 ;
        RECT 22.500 445.950 24.600 448.050 ;
        RECT 38.100 448.050 39.300 455.400 ;
        RECT 44.700 454.500 45.900 461.400 ;
        RECT 40.200 453.600 45.900 454.500 ;
        RECT 62.100 455.400 63.900 467.400 ;
        RECT 65.100 457.200 66.900 468.000 ;
        RECT 68.100 461.400 69.900 467.400 ;
        RECT 83.100 461.400 84.900 468.000 ;
        RECT 86.100 461.400 87.900 467.400 ;
        RECT 89.100 461.400 90.900 468.000 ;
        RECT 104.700 461.400 106.500 468.000 ;
        RECT 40.200 452.700 42.000 453.600 ;
        RECT 38.100 445.950 40.200 448.050 ;
        RECT 19.200 440.400 21.000 441.300 ;
        RECT 19.200 439.500 24.900 440.400 ;
        RECT 17.100 432.600 18.900 438.600 ;
        RECT 20.100 432.000 21.900 438.600 ;
        RECT 23.700 435.600 24.900 439.500 ;
        RECT 23.100 432.600 24.900 435.600 ;
        RECT 38.100 438.600 39.300 445.950 ;
        RECT 41.100 441.300 42.000 452.700 ;
        RECT 43.800 448.050 45.600 449.850 ;
        RECT 43.500 445.950 45.600 448.050 ;
        RECT 62.100 448.050 63.300 455.400 ;
        RECT 68.700 454.500 69.900 461.400 ;
        RECT 64.200 453.600 69.900 454.500 ;
        RECT 64.200 452.700 66.000 453.600 ;
        RECT 62.100 445.950 64.200 448.050 ;
        RECT 40.200 440.400 42.000 441.300 ;
        RECT 40.200 439.500 45.900 440.400 ;
        RECT 38.100 432.600 39.900 438.600 ;
        RECT 41.100 432.000 42.900 438.600 ;
        RECT 44.700 435.600 45.900 439.500 ;
        RECT 44.100 432.600 45.900 435.600 ;
        RECT 62.100 438.600 63.300 445.950 ;
        RECT 65.100 441.300 66.000 452.700 ;
        RECT 67.800 448.050 69.600 449.850 ;
        RECT 86.100 448.050 87.300 461.400 ;
        RECT 105.000 458.100 106.800 459.900 ;
        RECT 107.700 456.900 109.500 467.400 ;
        RECT 107.100 455.400 109.500 456.900 ;
        RECT 112.800 455.400 114.600 468.000 ;
        RECT 128.100 461.400 129.900 467.400 ;
        RECT 107.100 448.050 108.300 455.400 ;
        RECT 128.100 454.500 129.300 461.400 ;
        RECT 131.100 457.200 132.900 468.000 ;
        RECT 134.100 455.400 135.900 467.400 ;
        RECT 149.400 455.400 151.200 468.000 ;
        RECT 154.500 456.900 156.300 467.400 ;
        RECT 157.500 461.400 159.300 468.000 ;
        RECT 160.950 465.450 163.050 466.050 ;
        RECT 160.950 465.000 171.450 465.450 ;
        RECT 160.950 464.550 172.050 465.000 ;
        RECT 160.950 463.950 163.050 464.550 ;
        RECT 169.950 460.950 172.050 464.550 ;
        RECT 173.100 461.400 174.900 467.400 ;
        RECT 176.100 461.400 177.900 468.000 ;
        RECT 157.200 458.100 159.000 459.900 ;
        RECT 154.500 455.400 156.900 456.900 ;
        RECT 128.100 453.600 133.800 454.500 ;
        RECT 132.000 452.700 133.800 453.600 ;
        RECT 113.100 448.050 114.900 449.850 ;
        RECT 128.400 448.050 130.200 449.850 ;
        RECT 67.500 445.950 69.600 448.050 ;
        RECT 82.950 445.950 85.050 448.050 ;
        RECT 85.950 445.950 88.050 448.050 ;
        RECT 88.950 445.950 91.050 448.050 ;
        RECT 103.950 445.950 106.050 448.050 ;
        RECT 106.950 445.950 109.050 448.050 ;
        RECT 109.950 445.950 112.050 448.050 ;
        RECT 112.950 445.950 115.050 448.050 ;
        RECT 128.400 445.950 130.500 448.050 ;
        RECT 83.250 444.150 85.050 445.950 ;
        RECT 64.200 440.400 66.000 441.300 ;
        RECT 86.100 440.700 87.300 445.950 ;
        RECT 89.100 444.150 90.900 445.950 ;
        RECT 104.100 444.150 105.900 445.950 ;
        RECT 107.100 441.600 108.300 445.950 ;
        RECT 110.100 444.150 111.900 445.950 ;
        RECT 115.950 444.450 118.050 445.050 ;
        RECT 121.950 444.450 124.050 445.050 ;
        RECT 115.950 443.550 124.050 444.450 ;
        RECT 115.950 442.950 118.050 443.550 ;
        RECT 121.950 442.950 124.050 443.550 ;
        RECT 104.700 440.700 108.300 441.600 ;
        RECT 132.000 441.300 132.900 452.700 ;
        RECT 134.700 448.050 135.900 455.400 ;
        RECT 149.100 448.050 150.900 449.850 ;
        RECT 155.700 448.050 156.900 455.400 ;
        RECT 173.700 448.050 174.900 461.400 ;
        RECT 180.150 457.200 181.950 467.400 ;
        RECT 179.550 455.400 181.950 457.200 ;
        RECT 183.150 455.400 184.950 468.000 ;
        RECT 188.550 458.400 190.350 467.400 ;
        RECT 193.350 461.400 195.150 468.000 ;
        RECT 196.350 460.500 198.150 467.400 ;
        RECT 199.350 461.400 201.150 468.000 ;
        RECT 203.850 461.400 205.650 467.400 ;
        RECT 192.450 459.450 199.050 460.500 ;
        RECT 192.450 458.700 194.250 459.450 ;
        RECT 197.250 458.700 199.050 459.450 ;
        RECT 203.550 459.300 205.650 461.400 ;
        RECT 188.250 457.500 190.350 458.400 ;
        RECT 200.850 457.800 202.650 458.400 ;
        RECT 188.250 456.300 196.050 457.500 ;
        RECT 194.250 455.700 196.050 456.300 ;
        RECT 196.950 456.900 202.650 457.800 ;
        RECT 179.550 454.500 180.450 455.400 ;
        RECT 196.950 454.800 197.850 456.900 ;
        RECT 200.850 456.600 202.650 456.900 ;
        RECT 203.550 456.600 206.550 458.400 ;
        RECT 203.550 455.700 204.750 456.600 ;
        RECT 189.450 454.500 197.850 454.800 ;
        RECT 179.550 453.900 197.850 454.500 ;
        RECT 199.950 454.800 204.750 455.700 ;
        RECT 208.650 455.400 210.450 468.000 ;
        RECT 211.650 455.400 213.450 467.400 ;
        RECT 216.150 457.200 217.950 467.400 ;
        RECT 179.550 453.300 191.250 453.900 ;
        RECT 176.100 448.050 177.900 449.850 ;
        RECT 133.800 445.950 135.900 448.050 ;
        RECT 148.950 445.950 151.050 448.050 ;
        RECT 151.950 445.950 154.050 448.050 ;
        RECT 154.950 445.950 157.050 448.050 ;
        RECT 157.950 445.950 160.050 448.050 ;
        RECT 172.950 445.950 175.050 448.050 ;
        RECT 175.950 445.950 178.050 448.050 ;
        RECT 64.200 439.500 69.900 440.400 ;
        RECT 86.100 439.800 90.300 440.700 ;
        RECT 62.100 432.600 63.900 438.600 ;
        RECT 65.100 432.000 66.900 438.600 ;
        RECT 68.700 435.600 69.900 439.500 ;
        RECT 68.100 432.600 69.900 435.600 ;
        RECT 83.400 432.000 85.200 438.600 ;
        RECT 88.500 432.600 90.300 439.800 ;
        RECT 104.700 438.600 105.900 440.700 ;
        RECT 132.000 440.400 133.800 441.300 ;
        RECT 128.100 439.500 133.800 440.400 ;
        RECT 104.100 432.600 105.900 438.600 ;
        RECT 107.100 437.700 114.900 439.050 ;
        RECT 107.100 432.600 108.900 437.700 ;
        RECT 110.100 432.000 111.900 436.800 ;
        RECT 113.100 432.600 114.900 437.700 ;
        RECT 128.100 435.600 129.300 439.500 ;
        RECT 134.700 438.600 135.900 445.950 ;
        RECT 152.100 444.150 153.900 445.950 ;
        RECT 155.700 441.600 156.900 445.950 ;
        RECT 158.100 444.150 159.900 445.950 ;
        RECT 155.700 440.700 159.300 441.600 ;
        RECT 128.100 432.600 129.900 435.600 ;
        RECT 131.100 432.000 132.900 438.600 ;
        RECT 134.100 432.600 135.900 438.600 ;
        RECT 149.100 437.700 156.900 439.050 ;
        RECT 149.100 432.600 150.900 437.700 ;
        RECT 152.100 432.000 153.900 436.800 ;
        RECT 155.100 432.600 156.900 437.700 ;
        RECT 158.100 438.600 159.300 440.700 ;
        RECT 158.100 432.600 159.900 438.600 ;
        RECT 173.700 435.600 174.900 445.950 ;
        RECT 179.550 438.600 180.450 453.300 ;
        RECT 189.450 453.000 191.250 453.300 ;
        RECT 181.950 445.950 184.050 448.050 ;
        RECT 191.100 446.400 193.200 448.050 ;
        RECT 181.950 443.400 183.750 445.950 ;
        RECT 185.100 445.200 193.200 446.400 ;
        RECT 185.100 444.600 186.900 445.200 ;
        RECT 188.100 443.400 189.900 444.000 ;
        RECT 181.950 442.200 189.900 443.400 ;
        RECT 199.950 442.200 200.850 454.800 ;
        RECT 203.550 452.100 205.650 452.700 ;
        RECT 209.550 452.100 211.350 452.550 ;
        RECT 203.550 450.900 211.350 452.100 ;
        RECT 203.550 450.600 205.650 450.900 ;
        RECT 209.550 450.750 211.350 450.900 ;
        RECT 212.250 448.050 213.450 455.400 ;
        RECT 208.950 447.750 213.450 448.050 ;
        RECT 207.150 445.950 213.450 447.750 ;
        RECT 188.850 441.000 200.850 442.200 ;
        RECT 188.850 439.200 189.900 441.000 ;
        RECT 199.050 440.400 200.850 441.000 ;
        RECT 179.550 436.800 181.950 438.600 ;
        RECT 173.100 432.600 174.900 435.600 ;
        RECT 176.100 432.000 177.900 435.600 ;
        RECT 180.150 432.600 181.950 436.800 ;
        RECT 183.150 432.000 184.950 438.600 ;
        RECT 185.850 436.200 187.950 437.700 ;
        RECT 188.850 437.400 190.650 439.200 ;
        RECT 212.250 438.600 213.450 445.950 ;
        RECT 191.850 437.550 193.650 438.300 ;
        RECT 191.850 436.500 196.800 437.550 ;
        RECT 185.850 435.600 189.750 436.200 ;
        RECT 195.750 435.600 196.800 436.500 ;
        RECT 203.250 435.600 205.650 437.700 ;
        RECT 186.150 434.700 189.750 435.600 ;
        RECT 187.950 432.600 189.750 434.700 ;
        RECT 192.450 432.000 194.250 435.600 ;
        RECT 195.750 432.600 197.550 435.600 ;
        RECT 198.750 432.000 200.550 435.600 ;
        RECT 203.250 432.600 205.050 435.600 ;
        RECT 208.350 432.000 210.150 438.600 ;
        RECT 211.650 432.600 213.450 438.600 ;
        RECT 215.550 455.400 217.950 457.200 ;
        RECT 219.150 455.400 220.950 468.000 ;
        RECT 224.550 458.400 226.350 467.400 ;
        RECT 229.350 461.400 231.150 468.000 ;
        RECT 232.350 460.500 234.150 467.400 ;
        RECT 235.350 461.400 237.150 468.000 ;
        RECT 239.850 461.400 241.650 467.400 ;
        RECT 228.450 459.450 235.050 460.500 ;
        RECT 228.450 458.700 230.250 459.450 ;
        RECT 233.250 458.700 235.050 459.450 ;
        RECT 239.550 459.300 241.650 461.400 ;
        RECT 224.250 457.500 226.350 458.400 ;
        RECT 236.850 457.800 238.650 458.400 ;
        RECT 224.250 456.300 232.050 457.500 ;
        RECT 230.250 455.700 232.050 456.300 ;
        RECT 232.950 456.900 238.650 457.800 ;
        RECT 215.550 454.500 216.450 455.400 ;
        RECT 232.950 454.800 233.850 456.900 ;
        RECT 236.850 456.600 238.650 456.900 ;
        RECT 239.550 456.600 242.550 458.400 ;
        RECT 239.550 455.700 240.750 456.600 ;
        RECT 225.450 454.500 233.850 454.800 ;
        RECT 215.550 453.900 233.850 454.500 ;
        RECT 235.950 454.800 240.750 455.700 ;
        RECT 244.650 455.400 246.450 468.000 ;
        RECT 247.650 455.400 249.450 467.400 ;
        RECT 263.400 455.400 265.200 468.000 ;
        RECT 268.500 456.900 270.300 467.400 ;
        RECT 271.500 461.400 273.300 468.000 ;
        RECT 287.100 461.400 288.900 468.000 ;
        RECT 290.100 461.400 291.900 467.400 ;
        RECT 293.100 461.400 294.900 468.000 ;
        RECT 271.200 458.100 273.000 459.900 ;
        RECT 268.500 455.400 270.900 456.900 ;
        RECT 215.550 453.300 227.250 453.900 ;
        RECT 215.550 438.600 216.450 453.300 ;
        RECT 225.450 453.000 227.250 453.300 ;
        RECT 217.950 445.950 220.050 448.050 ;
        RECT 227.100 446.400 229.200 448.050 ;
        RECT 217.950 443.400 219.750 445.950 ;
        RECT 221.100 445.200 229.200 446.400 ;
        RECT 221.100 444.600 222.900 445.200 ;
        RECT 224.100 443.400 225.900 444.000 ;
        RECT 217.950 442.200 225.900 443.400 ;
        RECT 235.950 442.200 236.850 454.800 ;
        RECT 239.550 452.100 241.650 452.700 ;
        RECT 245.550 452.100 247.350 452.550 ;
        RECT 239.550 450.900 247.350 452.100 ;
        RECT 239.550 450.600 241.650 450.900 ;
        RECT 245.550 450.750 247.350 450.900 ;
        RECT 248.250 448.050 249.450 455.400 ;
        RECT 263.100 448.050 264.900 449.850 ;
        RECT 269.700 448.050 270.900 455.400 ;
        RECT 290.100 448.050 291.300 461.400 ;
        RECT 311.400 455.400 313.200 468.000 ;
        RECT 316.500 456.900 318.300 467.400 ;
        RECT 319.500 461.400 321.300 468.000 ;
        RECT 335.100 466.500 342.900 467.400 ;
        RECT 319.200 458.100 321.000 459.900 ;
        RECT 316.500 455.400 318.900 456.900 ;
        RECT 335.100 455.400 336.900 466.500 ;
        RECT 311.100 448.050 312.900 449.850 ;
        RECT 317.700 448.050 318.900 455.400 ;
        RECT 338.100 454.500 339.900 465.600 ;
        RECT 341.100 456.600 342.900 466.500 ;
        RECT 344.100 457.500 345.900 468.000 ;
        RECT 347.100 456.600 348.900 467.400 ;
        RECT 341.100 455.700 348.900 456.600 ;
        RECT 362.100 456.600 363.900 467.400 ;
        RECT 365.100 457.500 366.900 468.000 ;
        RECT 368.100 466.500 375.900 467.400 ;
        RECT 368.100 456.600 369.900 466.500 ;
        RECT 362.100 455.700 369.900 456.600 ;
        RECT 371.100 454.500 372.900 465.600 ;
        RECT 374.100 455.400 375.900 466.500 ;
        RECT 389.400 455.400 391.200 468.000 ;
        RECT 394.500 456.900 396.300 467.400 ;
        RECT 397.500 461.400 399.300 468.000 ;
        RECT 397.200 458.100 399.000 459.900 ;
        RECT 394.500 455.400 396.900 456.900 ;
        RECT 413.400 455.400 415.200 468.000 ;
        RECT 418.500 456.900 420.300 467.400 ;
        RECT 421.500 461.400 423.300 468.000 ;
        RECT 421.200 458.100 423.000 459.900 ;
        RECT 418.500 455.400 420.900 456.900 ;
        RECT 440.100 456.600 441.900 467.400 ;
        RECT 443.100 457.500 444.900 468.000 ;
        RECT 446.100 466.500 453.900 467.400 ;
        RECT 446.100 456.600 447.900 466.500 ;
        RECT 440.100 455.700 447.900 456.600 ;
        RECT 338.100 453.600 342.900 454.500 ;
        RECT 338.100 448.050 339.900 449.850 ;
        RECT 342.000 448.050 342.900 453.600 ;
        RECT 368.100 453.600 372.900 454.500 ;
        RECT 343.950 448.050 345.750 449.850 ;
        RECT 365.250 448.050 367.050 449.850 ;
        RECT 368.100 448.050 369.000 453.600 ;
        RECT 371.100 448.050 372.900 449.850 ;
        RECT 389.100 448.050 390.900 449.850 ;
        RECT 395.700 448.050 396.900 455.400 ;
        RECT 413.100 448.050 414.900 449.850 ;
        RECT 419.700 448.050 420.900 455.400 ;
        RECT 449.100 454.500 450.900 465.600 ;
        RECT 452.100 455.400 453.900 466.500 ;
        RECT 470.100 461.400 471.900 468.000 ;
        RECT 473.100 461.400 474.900 467.400 ;
        RECT 476.100 461.400 477.900 468.000 ;
        RECT 491.700 461.400 493.500 468.000 ;
        RECT 421.950 453.450 424.050 454.050 ;
        RECT 442.950 453.450 445.050 454.050 ;
        RECT 421.950 452.550 445.050 453.450 ;
        RECT 421.950 451.950 424.050 452.550 ;
        RECT 442.950 451.950 445.050 452.550 ;
        RECT 446.100 453.600 450.900 454.500 ;
        RECT 443.250 448.050 445.050 449.850 ;
        RECT 446.100 448.050 447.000 453.600 ;
        RECT 449.100 448.050 450.900 449.850 ;
        RECT 473.700 448.050 474.900 461.400 ;
        RECT 492.000 458.100 493.800 459.900 ;
        RECT 494.700 456.900 496.500 467.400 ;
        RECT 494.100 455.400 496.500 456.900 ;
        RECT 499.800 455.400 501.600 468.000 ;
        RECT 515.100 461.400 516.900 467.400 ;
        RECT 518.100 461.400 519.900 468.000 ;
        RECT 481.950 453.450 484.050 454.050 ;
        RECT 490.950 453.450 493.050 454.050 ;
        RECT 481.950 452.550 493.050 453.450 ;
        RECT 481.950 451.950 484.050 452.550 ;
        RECT 490.950 451.950 493.050 452.550 ;
        RECT 494.100 448.050 495.300 455.400 ;
        RECT 496.950 453.450 499.050 454.050 ;
        RECT 511.950 453.450 514.050 454.050 ;
        RECT 496.950 452.550 514.050 453.450 ;
        RECT 496.950 451.950 499.050 452.550 ;
        RECT 511.950 451.950 514.050 452.550 ;
        RECT 500.100 448.050 501.900 449.850 ;
        RECT 515.700 448.050 516.900 461.400 ;
        RECT 521.550 455.400 523.350 467.400 ;
        RECT 524.550 455.400 526.350 468.000 ;
        RECT 529.350 461.400 531.150 467.400 ;
        RECT 533.850 461.400 535.650 468.000 ;
        RECT 529.350 459.300 531.450 461.400 ;
        RECT 536.850 460.500 538.650 467.400 ;
        RECT 539.850 461.400 541.650 468.000 ;
        RECT 535.950 459.450 542.550 460.500 ;
        RECT 535.950 458.700 537.750 459.450 ;
        RECT 540.750 458.700 542.550 459.450 ;
        RECT 544.650 458.400 546.450 467.400 ;
        RECT 528.450 456.600 531.450 458.400 ;
        RECT 532.350 457.800 534.150 458.400 ;
        RECT 532.350 456.900 538.050 457.800 ;
        RECT 544.650 457.500 546.750 458.400 ;
        RECT 532.350 456.600 534.150 456.900 ;
        RECT 530.250 455.700 531.450 456.600 ;
        RECT 518.100 448.050 519.900 449.850 ;
        RECT 521.550 448.050 522.750 455.400 ;
        RECT 530.250 454.800 535.050 455.700 ;
        RECT 523.650 452.100 525.450 452.550 ;
        RECT 529.350 452.100 531.450 452.700 ;
        RECT 523.650 450.900 531.450 452.100 ;
        RECT 523.650 450.750 525.450 450.900 ;
        RECT 529.350 450.600 531.450 450.900 ;
        RECT 244.950 447.750 249.450 448.050 ;
        RECT 243.150 445.950 249.450 447.750 ;
        RECT 262.950 445.950 265.050 448.050 ;
        RECT 265.950 445.950 268.050 448.050 ;
        RECT 268.950 445.950 271.050 448.050 ;
        RECT 271.950 445.950 274.050 448.050 ;
        RECT 286.950 445.950 289.050 448.050 ;
        RECT 289.950 445.950 292.050 448.050 ;
        RECT 292.950 445.950 295.050 448.050 ;
        RECT 310.950 445.950 313.050 448.050 ;
        RECT 313.950 445.950 316.050 448.050 ;
        RECT 316.950 445.950 319.050 448.050 ;
        RECT 319.950 445.950 322.050 448.050 ;
        RECT 334.950 445.950 337.050 448.050 ;
        RECT 337.950 445.950 340.050 448.050 ;
        RECT 340.950 445.950 343.050 448.050 ;
        RECT 343.950 445.950 346.050 448.050 ;
        RECT 346.950 445.950 349.050 448.050 ;
        RECT 361.950 445.950 364.050 448.050 ;
        RECT 364.950 445.950 367.050 448.050 ;
        RECT 367.950 445.950 370.050 448.050 ;
        RECT 370.950 445.950 373.050 448.050 ;
        RECT 373.950 445.950 376.050 448.050 ;
        RECT 388.950 445.950 391.050 448.050 ;
        RECT 391.950 445.950 394.050 448.050 ;
        RECT 394.950 445.950 397.050 448.050 ;
        RECT 397.950 445.950 400.050 448.050 ;
        RECT 412.950 445.950 415.050 448.050 ;
        RECT 415.950 445.950 418.050 448.050 ;
        RECT 418.950 445.950 421.050 448.050 ;
        RECT 421.950 445.950 424.050 448.050 ;
        RECT 439.950 445.950 442.050 448.050 ;
        RECT 442.950 445.950 445.050 448.050 ;
        RECT 445.950 445.950 448.050 448.050 ;
        RECT 448.950 445.950 451.050 448.050 ;
        RECT 451.950 445.950 454.050 448.050 ;
        RECT 469.950 445.950 472.050 448.050 ;
        RECT 472.950 445.950 475.050 448.050 ;
        RECT 475.950 445.950 478.050 448.050 ;
        RECT 490.950 445.950 493.050 448.050 ;
        RECT 493.950 445.950 496.050 448.050 ;
        RECT 496.950 445.950 499.050 448.050 ;
        RECT 499.950 445.950 502.050 448.050 ;
        RECT 514.950 445.950 517.050 448.050 ;
        RECT 517.950 445.950 520.050 448.050 ;
        RECT 521.550 447.750 526.050 448.050 ;
        RECT 521.550 445.950 527.850 447.750 ;
        RECT 224.850 441.000 236.850 442.200 ;
        RECT 224.850 439.200 225.900 441.000 ;
        RECT 235.050 440.400 236.850 441.000 ;
        RECT 215.550 436.800 217.950 438.600 ;
        RECT 216.150 432.600 217.950 436.800 ;
        RECT 219.150 432.000 220.950 438.600 ;
        RECT 221.850 436.200 223.950 437.700 ;
        RECT 224.850 437.400 226.650 439.200 ;
        RECT 248.250 438.600 249.450 445.950 ;
        RECT 266.100 444.150 267.900 445.950 ;
        RECT 269.700 441.600 270.900 445.950 ;
        RECT 272.100 444.150 273.900 445.950 ;
        RECT 287.250 444.150 289.050 445.950 ;
        RECT 269.700 440.700 273.300 441.600 ;
        RECT 227.850 437.550 229.650 438.300 ;
        RECT 227.850 436.500 232.800 437.550 ;
        RECT 221.850 435.600 225.750 436.200 ;
        RECT 231.750 435.600 232.800 436.500 ;
        RECT 239.250 435.600 241.650 437.700 ;
        RECT 222.150 434.700 225.750 435.600 ;
        RECT 223.950 432.600 225.750 434.700 ;
        RECT 228.450 432.000 230.250 435.600 ;
        RECT 231.750 432.600 233.550 435.600 ;
        RECT 234.750 432.000 236.550 435.600 ;
        RECT 239.250 432.600 241.050 435.600 ;
        RECT 244.350 432.000 246.150 438.600 ;
        RECT 247.650 432.600 249.450 438.600 ;
        RECT 263.100 437.700 270.900 439.050 ;
        RECT 263.100 432.600 264.900 437.700 ;
        RECT 266.100 432.000 267.900 436.800 ;
        RECT 269.100 432.600 270.900 437.700 ;
        RECT 272.100 438.600 273.300 440.700 ;
        RECT 290.100 440.700 291.300 445.950 ;
        RECT 293.100 444.150 294.900 445.950 ;
        RECT 314.100 444.150 315.900 445.950 ;
        RECT 317.700 441.600 318.900 445.950 ;
        RECT 320.100 444.150 321.900 445.950 ;
        RECT 335.100 444.150 336.900 445.950 ;
        RECT 317.700 440.700 321.300 441.600 ;
        RECT 290.100 439.800 294.300 440.700 ;
        RECT 272.100 432.600 273.900 438.600 ;
        RECT 287.400 432.000 289.200 438.600 ;
        RECT 292.500 432.600 294.300 439.800 ;
        RECT 311.100 437.700 318.900 439.050 ;
        RECT 311.100 432.600 312.900 437.700 ;
        RECT 314.100 432.000 315.900 436.800 ;
        RECT 317.100 432.600 318.900 437.700 ;
        RECT 320.100 438.600 321.300 440.700 ;
        RECT 341.700 438.600 342.900 445.950 ;
        RECT 346.950 444.150 348.750 445.950 ;
        RECT 362.250 444.150 364.050 445.950 ;
        RECT 368.100 438.600 369.300 445.950 ;
        RECT 374.100 444.150 375.900 445.950 ;
        RECT 392.100 444.150 393.900 445.950 ;
        RECT 395.700 441.600 396.900 445.950 ;
        RECT 398.100 444.150 399.900 445.950 ;
        RECT 416.100 444.150 417.900 445.950 ;
        RECT 419.700 441.600 420.900 445.950 ;
        RECT 422.100 444.150 423.900 445.950 ;
        RECT 440.250 444.150 442.050 445.950 ;
        RECT 395.700 440.700 399.300 441.600 ;
        RECT 419.700 440.700 423.300 441.600 ;
        RECT 320.100 432.600 321.900 438.600 ;
        RECT 337.500 432.000 339.300 438.600 ;
        RECT 342.000 432.600 343.800 438.600 ;
        RECT 346.500 432.000 348.300 438.600 ;
        RECT 362.700 432.000 364.500 438.600 ;
        RECT 367.200 432.600 369.000 438.600 ;
        RECT 371.700 432.000 373.500 438.600 ;
        RECT 389.100 437.700 396.900 439.050 ;
        RECT 389.100 432.600 390.900 437.700 ;
        RECT 392.100 432.000 393.900 436.800 ;
        RECT 395.100 432.600 396.900 437.700 ;
        RECT 398.100 438.600 399.300 440.700 ;
        RECT 398.100 432.600 399.900 438.600 ;
        RECT 413.100 437.700 420.900 439.050 ;
        RECT 413.100 432.600 414.900 437.700 ;
        RECT 416.100 432.000 417.900 436.800 ;
        RECT 419.100 432.600 420.900 437.700 ;
        RECT 422.100 438.600 423.300 440.700 ;
        RECT 446.100 438.600 447.300 445.950 ;
        RECT 452.100 444.150 453.900 445.950 ;
        RECT 470.100 444.150 471.900 445.950 ;
        RECT 448.950 441.450 451.050 442.050 ;
        RECT 466.950 441.450 469.050 442.050 ;
        RECT 448.950 440.550 469.050 441.450 ;
        RECT 473.700 440.700 474.900 445.950 ;
        RECT 475.950 444.150 477.750 445.950 ;
        RECT 491.100 444.150 492.900 445.950 ;
        RECT 494.100 441.600 495.300 445.950 ;
        RECT 497.100 444.150 498.900 445.950 ;
        RECT 448.950 439.950 451.050 440.550 ;
        RECT 466.950 439.950 469.050 440.550 ;
        RECT 470.700 439.800 474.900 440.700 ;
        RECT 491.700 440.700 495.300 441.600 ;
        RECT 422.100 432.600 423.900 438.600 ;
        RECT 440.700 432.000 442.500 438.600 ;
        RECT 445.200 432.600 447.000 438.600 ;
        RECT 449.700 432.000 451.500 438.600 ;
        RECT 470.700 432.600 472.500 439.800 ;
        RECT 491.700 438.600 492.900 440.700 ;
        RECT 475.800 432.000 477.600 438.600 ;
        RECT 491.100 432.600 492.900 438.600 ;
        RECT 494.100 437.700 501.900 439.050 ;
        RECT 494.100 432.600 495.900 437.700 ;
        RECT 497.100 432.000 498.900 436.800 ;
        RECT 500.100 432.600 501.900 437.700 ;
        RECT 515.700 435.600 516.900 445.950 ;
        RECT 521.550 438.600 522.750 445.950 ;
        RECT 534.150 442.200 535.050 454.800 ;
        RECT 537.150 454.800 538.050 456.900 ;
        RECT 538.950 456.300 546.750 457.500 ;
        RECT 538.950 455.700 540.750 456.300 ;
        RECT 550.050 455.400 551.850 468.000 ;
        RECT 553.050 457.200 554.850 467.400 ;
        RECT 553.050 455.400 555.450 457.200 ;
        RECT 537.150 454.500 545.550 454.800 ;
        RECT 554.550 454.500 555.450 455.400 ;
        RECT 537.150 453.900 555.450 454.500 ;
        RECT 543.750 453.300 555.450 453.900 ;
        RECT 543.750 453.000 545.550 453.300 ;
        RECT 541.800 446.400 543.900 448.050 ;
        RECT 541.800 445.200 549.900 446.400 ;
        RECT 550.950 445.950 553.050 448.050 ;
        RECT 548.100 444.600 549.900 445.200 ;
        RECT 545.100 443.400 546.900 444.000 ;
        RECT 551.250 443.400 553.050 445.950 ;
        RECT 545.100 442.200 553.050 443.400 ;
        RECT 534.150 441.000 546.150 442.200 ;
        RECT 534.150 440.400 535.950 441.000 ;
        RECT 545.100 439.200 546.150 441.000 ;
        RECT 515.100 432.600 516.900 435.600 ;
        RECT 518.100 432.000 519.900 435.600 ;
        RECT 521.550 432.600 523.350 438.600 ;
        RECT 524.850 432.000 526.650 438.600 ;
        RECT 529.350 435.600 531.750 437.700 ;
        RECT 541.350 437.550 543.150 438.300 ;
        RECT 538.200 436.500 543.150 437.550 ;
        RECT 544.350 437.400 546.150 439.200 ;
        RECT 554.550 438.600 555.450 453.300 ;
        RECT 538.200 435.600 539.250 436.500 ;
        RECT 547.050 436.200 549.150 437.700 ;
        RECT 545.250 435.600 549.150 436.200 ;
        RECT 529.950 432.600 531.750 435.600 ;
        RECT 534.450 432.000 536.250 435.600 ;
        RECT 537.450 432.600 539.250 435.600 ;
        RECT 540.750 432.000 542.550 435.600 ;
        RECT 545.250 434.700 548.850 435.600 ;
        RECT 545.250 432.600 547.050 434.700 ;
        RECT 550.050 432.000 551.850 438.600 ;
        RECT 553.050 436.800 555.450 438.600 ;
        RECT 557.550 455.400 559.350 467.400 ;
        RECT 560.550 455.400 562.350 468.000 ;
        RECT 565.350 461.400 567.150 467.400 ;
        RECT 569.850 461.400 571.650 468.000 ;
        RECT 565.350 459.300 567.450 461.400 ;
        RECT 572.850 460.500 574.650 467.400 ;
        RECT 575.850 461.400 577.650 468.000 ;
        RECT 571.950 459.450 578.550 460.500 ;
        RECT 571.950 458.700 573.750 459.450 ;
        RECT 576.750 458.700 578.550 459.450 ;
        RECT 580.650 458.400 582.450 467.400 ;
        RECT 564.450 456.600 567.450 458.400 ;
        RECT 568.350 457.800 570.150 458.400 ;
        RECT 568.350 456.900 574.050 457.800 ;
        RECT 580.650 457.500 582.750 458.400 ;
        RECT 568.350 456.600 570.150 456.900 ;
        RECT 566.250 455.700 567.450 456.600 ;
        RECT 557.550 448.050 558.750 455.400 ;
        RECT 566.250 454.800 571.050 455.700 ;
        RECT 559.650 452.100 561.450 452.550 ;
        RECT 565.350 452.100 567.450 452.700 ;
        RECT 559.650 450.900 567.450 452.100 ;
        RECT 559.650 450.750 561.450 450.900 ;
        RECT 565.350 450.600 567.450 450.900 ;
        RECT 557.550 447.750 562.050 448.050 ;
        RECT 557.550 445.950 563.850 447.750 ;
        RECT 557.550 438.600 558.750 445.950 ;
        RECT 570.150 442.200 571.050 454.800 ;
        RECT 573.150 454.800 574.050 456.900 ;
        RECT 574.950 456.300 582.750 457.500 ;
        RECT 574.950 455.700 576.750 456.300 ;
        RECT 586.050 455.400 587.850 468.000 ;
        RECT 589.050 457.200 590.850 467.400 ;
        RECT 589.050 455.400 591.450 457.200 ;
        RECT 605.400 455.400 607.200 468.000 ;
        RECT 610.500 456.900 612.300 467.400 ;
        RECT 613.500 461.400 615.300 468.000 ;
        RECT 632.100 461.400 633.900 468.000 ;
        RECT 635.100 461.400 636.900 467.400 ;
        RECT 638.100 462.000 639.900 468.000 ;
        RECT 635.400 461.100 636.900 461.400 ;
        RECT 641.100 461.400 642.900 467.400 ;
        RECT 656.100 461.400 657.900 468.000 ;
        RECT 659.100 461.400 660.900 467.400 ;
        RECT 662.100 461.400 663.900 468.000 ;
        RECT 677.100 461.400 678.900 468.000 ;
        RECT 680.100 461.400 681.900 467.400 ;
        RECT 683.100 461.400 684.900 468.000 ;
        RECT 701.100 461.400 702.900 468.000 ;
        RECT 704.100 461.400 705.900 467.400 ;
        RECT 707.100 462.000 708.900 468.000 ;
        RECT 641.100 461.100 642.000 461.400 ;
        RECT 635.400 460.200 642.000 461.100 ;
        RECT 613.200 458.100 615.000 459.900 ;
        RECT 610.500 455.400 612.900 456.900 ;
        RECT 573.150 454.500 581.550 454.800 ;
        RECT 590.550 454.500 591.450 455.400 ;
        RECT 573.150 453.900 591.450 454.500 ;
        RECT 579.750 453.300 591.450 453.900 ;
        RECT 579.750 453.000 581.550 453.300 ;
        RECT 577.800 446.400 579.900 448.050 ;
        RECT 577.800 445.200 585.900 446.400 ;
        RECT 586.950 445.950 589.050 448.050 ;
        RECT 584.100 444.600 585.900 445.200 ;
        RECT 581.100 443.400 582.900 444.000 ;
        RECT 587.250 443.400 589.050 445.950 ;
        RECT 581.100 442.200 589.050 443.400 ;
        RECT 570.150 441.000 582.150 442.200 ;
        RECT 570.150 440.400 571.950 441.000 ;
        RECT 581.100 439.200 582.150 441.000 ;
        RECT 553.050 432.600 554.850 436.800 ;
        RECT 557.550 432.600 559.350 438.600 ;
        RECT 560.850 432.000 562.650 438.600 ;
        RECT 565.350 435.600 567.750 437.700 ;
        RECT 577.350 437.550 579.150 438.300 ;
        RECT 574.200 436.500 579.150 437.550 ;
        RECT 580.350 437.400 582.150 439.200 ;
        RECT 590.550 438.600 591.450 453.300 ;
        RECT 595.950 453.450 598.050 453.900 ;
        RECT 601.950 453.450 604.050 454.050 ;
        RECT 607.950 453.450 610.050 454.050 ;
        RECT 595.950 452.550 610.050 453.450 ;
        RECT 595.950 451.800 598.050 452.550 ;
        RECT 601.950 451.950 604.050 452.550 ;
        RECT 607.950 451.950 610.050 452.550 ;
        RECT 605.100 448.050 606.900 449.850 ;
        RECT 611.700 448.050 612.900 455.400 ;
        RECT 613.950 453.450 616.050 454.050 ;
        RECT 637.950 453.450 640.050 454.050 ;
        RECT 613.950 452.550 640.050 453.450 ;
        RECT 613.950 451.950 616.050 452.550 ;
        RECT 637.950 451.950 640.050 452.550 ;
        RECT 635.100 448.050 636.900 449.850 ;
        RECT 641.100 448.050 642.000 460.200 ;
        RECT 659.700 448.050 660.900 461.400 ;
        RECT 680.100 448.050 681.300 461.400 ;
        RECT 704.400 461.100 705.900 461.400 ;
        RECT 710.100 461.400 711.900 467.400 ;
        RECT 725.700 461.400 727.500 468.000 ;
        RECT 710.100 461.100 711.000 461.400 ;
        RECT 704.400 460.200 711.000 461.100 ;
        RECT 704.100 448.050 705.900 449.850 ;
        RECT 710.100 448.050 711.000 460.200 ;
        RECT 726.000 458.100 727.800 459.900 ;
        RECT 728.700 456.900 730.500 467.400 ;
        RECT 728.100 455.400 730.500 456.900 ;
        RECT 733.800 455.400 735.600 468.000 ;
        RECT 749.100 461.400 750.900 468.000 ;
        RECT 752.100 461.400 753.900 467.400 ;
        RECT 755.100 461.400 756.900 468.000 ;
        RECT 770.100 461.400 771.900 468.000 ;
        RECT 773.100 461.400 774.900 467.400 ;
        RECT 776.100 461.400 777.900 468.000 ;
        RECT 794.100 461.400 795.900 468.000 ;
        RECT 797.100 461.400 798.900 467.400 ;
        RECT 728.100 448.050 729.300 455.400 ;
        RECT 736.950 453.450 739.050 454.050 ;
        RECT 748.950 453.450 751.050 454.050 ;
        RECT 736.950 452.550 751.050 453.450 ;
        RECT 736.950 451.950 739.050 452.550 ;
        RECT 748.950 451.950 751.050 452.550 ;
        RECT 737.550 450.450 738.450 451.950 ;
        RECT 734.100 448.050 735.900 449.850 ;
        RECT 737.550 449.550 741.450 450.450 ;
        RECT 604.950 445.950 607.050 448.050 ;
        RECT 607.950 445.950 610.050 448.050 ;
        RECT 610.950 445.950 613.050 448.050 ;
        RECT 613.950 445.950 616.050 448.050 ;
        RECT 631.950 445.950 634.050 448.050 ;
        RECT 634.950 445.950 637.050 448.050 ;
        RECT 637.950 445.950 640.050 448.050 ;
        RECT 640.950 445.950 643.050 448.050 ;
        RECT 655.950 445.950 658.050 448.050 ;
        RECT 658.950 445.950 661.050 448.050 ;
        RECT 661.950 445.950 664.050 448.050 ;
        RECT 676.950 445.950 679.050 448.050 ;
        RECT 679.950 445.950 682.050 448.050 ;
        RECT 682.950 445.950 685.050 448.050 ;
        RECT 700.950 445.950 703.050 448.050 ;
        RECT 703.950 445.950 706.050 448.050 ;
        RECT 706.950 445.950 709.050 448.050 ;
        RECT 709.950 445.950 712.050 448.050 ;
        RECT 724.950 445.950 727.050 448.050 ;
        RECT 727.950 445.950 730.050 448.050 ;
        RECT 730.950 445.950 733.050 448.050 ;
        RECT 733.950 445.950 736.050 448.050 ;
        RECT 608.100 444.150 609.900 445.950 ;
        RECT 611.700 441.600 612.900 445.950 ;
        RECT 614.100 444.150 615.900 445.950 ;
        RECT 616.950 444.450 619.050 445.050 ;
        RECT 625.950 444.450 628.050 445.050 ;
        RECT 616.950 443.550 628.050 444.450 ;
        RECT 632.100 444.150 633.900 445.950 ;
        RECT 638.100 444.150 639.900 445.950 ;
        RECT 616.950 442.950 619.050 443.550 ;
        RECT 625.950 442.950 628.050 443.550 ;
        RECT 641.100 442.200 642.000 445.950 ;
        RECT 656.100 444.150 657.900 445.950 ;
        RECT 611.700 440.700 615.300 441.600 ;
        RECT 574.200 435.600 575.250 436.500 ;
        RECT 583.050 436.200 585.150 437.700 ;
        RECT 581.250 435.600 585.150 436.200 ;
        RECT 565.950 432.600 567.750 435.600 ;
        RECT 570.450 432.000 572.250 435.600 ;
        RECT 573.450 432.600 575.250 435.600 ;
        RECT 576.750 432.000 578.550 435.600 ;
        RECT 581.250 434.700 584.850 435.600 ;
        RECT 581.250 432.600 583.050 434.700 ;
        RECT 586.050 432.000 587.850 438.600 ;
        RECT 589.050 436.800 591.450 438.600 ;
        RECT 605.100 437.700 612.900 439.050 ;
        RECT 589.050 432.600 590.850 436.800 ;
        RECT 605.100 432.600 606.900 437.700 ;
        RECT 608.100 432.000 609.900 436.800 ;
        RECT 611.100 432.600 612.900 437.700 ;
        RECT 614.100 438.600 615.300 440.700 ;
        RECT 614.100 432.600 615.900 438.600 ;
        RECT 632.100 432.000 633.900 441.600 ;
        RECT 638.700 441.000 642.000 442.200 ;
        RECT 638.700 432.600 640.500 441.000 ;
        RECT 659.700 440.700 660.900 445.950 ;
        RECT 661.950 444.150 663.750 445.950 ;
        RECT 677.250 444.150 679.050 445.950 ;
        RECT 656.700 439.800 660.900 440.700 ;
        RECT 670.950 441.450 673.050 442.050 ;
        RECT 676.950 441.450 679.050 442.050 ;
        RECT 670.950 440.550 679.050 441.450 ;
        RECT 670.950 439.950 673.050 440.550 ;
        RECT 676.950 439.950 679.050 440.550 ;
        RECT 680.100 440.700 681.300 445.950 ;
        RECT 683.100 444.150 684.900 445.950 ;
        RECT 701.100 444.150 702.900 445.950 ;
        RECT 707.100 444.150 708.900 445.950 ;
        RECT 710.100 442.200 711.000 445.950 ;
        RECT 725.100 444.150 726.900 445.950 ;
        RECT 680.100 439.800 684.300 440.700 ;
        RECT 656.700 432.600 658.500 439.800 ;
        RECT 661.800 432.000 663.600 438.600 ;
        RECT 677.400 432.000 679.200 438.600 ;
        RECT 682.500 432.600 684.300 439.800 ;
        RECT 701.100 432.000 702.900 441.600 ;
        RECT 707.700 441.000 711.000 442.200 ;
        RECT 728.100 441.600 729.300 445.950 ;
        RECT 731.100 444.150 732.900 445.950 ;
        RECT 740.550 445.050 741.450 449.550 ;
        RECT 752.100 448.050 753.300 461.400 ;
        RECT 773.100 448.050 774.300 461.400 ;
        RECT 794.100 448.050 795.900 449.850 ;
        RECT 797.100 448.050 798.300 461.400 ;
        RECT 815.400 455.400 817.200 468.000 ;
        RECT 820.500 456.900 822.300 467.400 ;
        RECT 823.500 461.400 825.300 468.000 ;
        RECT 823.200 458.100 825.000 459.900 ;
        RECT 820.500 455.400 822.900 456.900 ;
        RECT 839.400 455.400 841.200 468.000 ;
        RECT 844.500 456.900 846.300 467.400 ;
        RECT 847.500 461.400 849.300 468.000 ;
        RECT 847.200 458.100 849.000 459.900 ;
        RECT 844.500 455.400 846.900 456.900 ;
        RECT 866.100 455.400 867.900 467.400 ;
        RECT 869.100 456.000 870.900 468.000 ;
        RECT 872.100 461.400 873.900 467.400 ;
        RECT 875.100 461.400 876.900 468.000 ;
        RECT 815.100 448.050 816.900 449.850 ;
        RECT 821.700 448.050 822.900 455.400 ;
        RECT 839.100 448.050 840.900 449.850 ;
        RECT 845.700 448.050 846.900 455.400 ;
        RECT 866.700 448.050 867.600 455.400 ;
        RECT 870.000 448.050 871.800 449.850 ;
        RECT 748.950 445.950 751.050 448.050 ;
        RECT 751.950 445.950 754.050 448.050 ;
        RECT 754.950 445.950 757.050 448.050 ;
        RECT 769.950 445.950 772.050 448.050 ;
        RECT 772.950 445.950 775.050 448.050 ;
        RECT 775.950 445.950 778.050 448.050 ;
        RECT 793.950 445.950 796.050 448.050 ;
        RECT 796.950 445.950 799.050 448.050 ;
        RECT 814.950 445.950 817.050 448.050 ;
        RECT 817.950 445.950 820.050 448.050 ;
        RECT 820.950 445.950 823.050 448.050 ;
        RECT 823.950 445.950 826.050 448.050 ;
        RECT 838.950 445.950 841.050 448.050 ;
        RECT 841.950 445.950 844.050 448.050 ;
        RECT 844.950 445.950 847.050 448.050 ;
        RECT 847.950 445.950 850.050 448.050 ;
        RECT 866.100 445.950 868.200 448.050 ;
        RECT 869.400 445.950 871.500 448.050 ;
        RECT 736.950 443.550 741.450 445.050 ;
        RECT 749.250 444.150 751.050 445.950 ;
        RECT 736.950 442.950 741.000 443.550 ;
        RECT 707.700 432.600 709.500 441.000 ;
        RECT 725.700 440.700 729.300 441.600 ;
        RECT 752.100 440.700 753.300 445.950 ;
        RECT 755.100 444.150 756.900 445.950 ;
        RECT 770.250 444.150 772.050 445.950 ;
        RECT 773.100 440.700 774.300 445.950 ;
        RECT 776.100 444.150 777.900 445.950 ;
        RECT 725.700 438.600 726.900 440.700 ;
        RECT 752.100 439.800 756.300 440.700 ;
        RECT 773.100 439.800 777.300 440.700 ;
        RECT 725.100 432.600 726.900 438.600 ;
        RECT 728.100 437.700 735.900 439.050 ;
        RECT 728.100 432.600 729.900 437.700 ;
        RECT 731.100 432.000 732.900 436.800 ;
        RECT 734.100 432.600 735.900 437.700 ;
        RECT 749.400 432.000 751.200 438.600 ;
        RECT 754.500 432.600 756.300 439.800 ;
        RECT 770.400 432.000 772.200 438.600 ;
        RECT 775.500 432.600 777.300 439.800 ;
        RECT 797.100 435.600 798.300 445.950 ;
        RECT 818.100 444.150 819.900 445.950 ;
        RECT 821.700 441.600 822.900 445.950 ;
        RECT 824.100 444.150 825.900 445.950 ;
        RECT 842.100 444.150 843.900 445.950 ;
        RECT 845.700 441.600 846.900 445.950 ;
        RECT 848.100 444.150 849.900 445.950 ;
        RECT 821.700 440.700 825.300 441.600 ;
        RECT 845.700 440.700 849.300 441.600 ;
        RECT 815.100 437.700 822.900 439.050 ;
        RECT 794.100 432.000 795.900 435.600 ;
        RECT 797.100 432.600 798.900 435.600 ;
        RECT 815.100 432.600 816.900 437.700 ;
        RECT 818.100 432.000 819.900 436.800 ;
        RECT 821.100 432.600 822.900 437.700 ;
        RECT 824.100 438.600 825.300 440.700 ;
        RECT 824.100 432.600 825.900 438.600 ;
        RECT 839.100 437.700 846.900 439.050 ;
        RECT 839.100 432.600 840.900 437.700 ;
        RECT 842.100 432.000 843.900 436.800 ;
        RECT 845.100 432.600 846.900 437.700 ;
        RECT 848.100 438.600 849.300 440.700 ;
        RECT 866.700 438.600 867.600 445.950 ;
        RECT 873.000 441.300 873.900 461.400 ;
        RECT 890.100 456.300 891.900 467.400 ;
        RECT 893.100 457.200 894.900 468.000 ;
        RECT 896.100 456.300 897.900 467.400 ;
        RECT 890.100 455.400 897.900 456.300 ;
        RECT 899.100 455.400 900.900 467.400 ;
        RECT 914.100 461.400 915.900 468.000 ;
        RECT 917.100 461.400 918.900 467.400 ;
        RECT 920.100 462.000 921.900 468.000 ;
        RECT 917.400 461.100 918.900 461.400 ;
        RECT 923.100 461.400 924.900 467.400 ;
        RECT 941.100 461.400 942.900 468.000 ;
        RECT 944.100 461.400 945.900 467.400 ;
        RECT 947.100 462.000 948.900 468.000 ;
        RECT 923.100 461.100 924.000 461.400 ;
        RECT 917.400 460.200 924.000 461.100 ;
        RECT 944.400 461.100 945.900 461.400 ;
        RECT 950.100 461.400 951.900 467.400 ;
        RECT 950.100 461.100 951.000 461.400 ;
        RECT 944.400 460.200 951.000 461.100 ;
        RECT 893.250 448.050 895.050 449.850 ;
        RECT 899.700 448.050 900.600 455.400 ;
        RECT 917.100 448.050 918.900 449.850 ;
        RECT 923.100 448.050 924.000 460.200 ;
        RECT 931.950 456.450 934.050 457.050 ;
        RECT 940.950 456.450 943.050 457.050 ;
        RECT 931.950 455.550 943.050 456.450 ;
        RECT 931.950 454.950 934.050 455.550 ;
        RECT 940.950 454.950 943.050 455.550 ;
        RECT 934.950 453.450 937.050 454.050 ;
        RECT 946.950 453.450 949.050 453.900 ;
        RECT 934.950 452.550 949.050 453.450 ;
        RECT 934.950 451.950 937.050 452.550 ;
        RECT 946.950 451.800 949.050 452.550 ;
        RECT 925.950 450.450 930.000 451.050 ;
        RECT 925.950 448.950 930.450 450.450 ;
        RECT 874.800 445.950 876.900 448.050 ;
        RECT 889.950 445.950 892.050 448.050 ;
        RECT 892.950 445.950 895.050 448.050 ;
        RECT 895.950 445.950 898.050 448.050 ;
        RECT 898.950 445.950 901.050 448.050 ;
        RECT 913.950 445.950 916.050 448.050 ;
        RECT 916.950 445.950 919.050 448.050 ;
        RECT 919.950 445.950 922.050 448.050 ;
        RECT 922.950 445.950 925.050 448.050 ;
        RECT 874.950 444.150 876.750 445.950 ;
        RECT 890.100 444.150 891.900 445.950 ;
        RECT 896.250 444.150 898.050 445.950 ;
        RECT 877.950 441.450 880.050 442.050 ;
        RECT 889.950 441.450 892.050 442.050 ;
        RECT 868.500 440.400 876.900 441.300 ;
        RECT 868.500 439.500 870.300 440.400 ;
        RECT 848.100 432.600 849.900 438.600 ;
        RECT 866.700 436.800 869.400 438.600 ;
        RECT 867.600 432.600 869.400 436.800 ;
        RECT 870.600 432.000 872.400 438.600 ;
        RECT 875.100 432.600 876.900 440.400 ;
        RECT 877.950 440.550 892.050 441.450 ;
        RECT 877.950 439.950 880.050 440.550 ;
        RECT 889.950 439.950 892.050 440.550 ;
        RECT 899.700 438.600 900.600 445.950 ;
        RECT 914.100 444.150 915.900 445.950 ;
        RECT 920.100 444.150 921.900 445.950 ;
        RECT 923.100 442.200 924.000 445.950 ;
        RECT 929.550 444.450 930.450 448.950 ;
        RECT 944.100 448.050 945.900 449.850 ;
        RECT 950.100 448.050 951.000 460.200 ;
        RECT 965.100 456.300 966.900 467.400 ;
        RECT 968.100 457.200 969.900 468.000 ;
        RECT 971.100 456.300 972.900 467.400 ;
        RECT 965.100 455.400 972.900 456.300 ;
        RECT 974.100 455.400 975.900 467.400 ;
        RECT 992.700 461.400 994.500 468.000 ;
        RECT 993.000 458.100 994.800 459.900 ;
        RECT 995.700 456.900 997.500 467.400 ;
        RECT 995.100 455.400 997.500 456.900 ;
        RECT 1000.800 455.400 1002.600 468.000 ;
        RECT 970.950 453.450 973.050 454.200 ;
        RECT 959.550 452.550 973.050 453.450 ;
        RECT 940.950 445.950 943.050 448.050 ;
        RECT 943.950 445.950 946.050 448.050 ;
        RECT 946.950 445.950 949.050 448.050 ;
        RECT 949.950 445.950 952.050 448.050 ;
        RECT 937.950 444.450 940.050 445.050 ;
        RECT 929.550 443.550 940.050 444.450 ;
        RECT 941.100 444.150 942.900 445.950 ;
        RECT 947.100 444.150 948.900 445.950 ;
        RECT 937.950 442.950 940.050 443.550 ;
        RECT 950.100 442.200 951.000 445.950 ;
        RECT 959.550 445.050 960.450 452.550 ;
        RECT 970.950 452.100 973.050 452.550 ;
        RECT 968.250 448.050 970.050 449.850 ;
        RECT 974.700 448.050 975.600 455.400 ;
        RECT 995.100 448.050 996.300 455.400 ;
        RECT 1001.100 448.050 1002.900 449.850 ;
        RECT 964.950 445.950 967.050 448.050 ;
        RECT 967.950 445.950 970.050 448.050 ;
        RECT 970.950 445.950 973.050 448.050 ;
        RECT 973.950 445.950 976.050 448.050 ;
        RECT 991.950 445.950 994.050 448.050 ;
        RECT 994.950 445.950 997.050 448.050 ;
        RECT 997.950 445.950 1000.050 448.050 ;
        RECT 1000.950 445.950 1003.050 448.050 ;
        RECT 959.550 443.550 964.050 445.050 ;
        RECT 965.100 444.150 966.900 445.950 ;
        RECT 971.250 444.150 973.050 445.950 ;
        RECT 960.000 442.950 964.050 443.550 ;
        RECT 891.000 432.000 892.800 438.600 ;
        RECT 895.500 437.400 900.600 438.600 ;
        RECT 895.500 432.600 897.300 437.400 ;
        RECT 898.500 432.000 900.300 435.600 ;
        RECT 914.100 432.000 915.900 441.600 ;
        RECT 920.700 441.000 924.000 442.200 ;
        RECT 920.700 432.600 922.500 441.000 ;
        RECT 941.100 432.000 942.900 441.600 ;
        RECT 947.700 441.000 951.000 442.200 ;
        RECT 947.700 432.600 949.500 441.000 ;
        RECT 974.700 438.600 975.600 445.950 ;
        RECT 992.100 444.150 993.900 445.950 ;
        RECT 995.100 441.600 996.300 445.950 ;
        RECT 998.100 444.150 999.900 445.950 ;
        RECT 992.700 440.700 996.300 441.600 ;
        RECT 992.700 438.600 993.900 440.700 ;
        RECT 966.000 432.000 967.800 438.600 ;
        RECT 970.500 437.400 975.600 438.600 ;
        RECT 970.500 432.600 972.300 437.400 ;
        RECT 973.500 432.000 975.300 435.600 ;
        RECT 992.100 432.600 993.900 438.600 ;
        RECT 995.100 437.700 1002.900 439.050 ;
        RECT 995.100 432.600 996.900 437.700 ;
        RECT 998.100 432.000 999.900 436.800 ;
        RECT 1001.100 432.600 1002.900 437.700 ;
        RECT 3.150 424.200 4.950 428.400 ;
        RECT 2.550 422.400 4.950 424.200 ;
        RECT 6.150 422.400 7.950 429.000 ;
        RECT 10.950 426.300 12.750 428.400 ;
        RECT 9.150 425.400 12.750 426.300 ;
        RECT 15.450 425.400 17.250 429.000 ;
        RECT 18.750 425.400 20.550 428.400 ;
        RECT 21.750 425.400 23.550 429.000 ;
        RECT 26.250 425.400 28.050 428.400 ;
        RECT 8.850 424.800 12.750 425.400 ;
        RECT 8.850 423.300 10.950 424.800 ;
        RECT 18.750 424.500 19.800 425.400 ;
        RECT 2.550 407.700 3.450 422.400 ;
        RECT 11.850 421.800 13.650 423.600 ;
        RECT 14.850 423.450 19.800 424.500 ;
        RECT 14.850 422.700 16.650 423.450 ;
        RECT 26.250 423.300 28.650 425.400 ;
        RECT 31.350 422.400 33.150 429.000 ;
        RECT 34.650 422.400 36.450 428.400 ;
        RECT 39.150 424.200 40.950 428.400 ;
        RECT 11.850 420.000 12.900 421.800 ;
        RECT 22.050 420.000 23.850 420.600 ;
        RECT 11.850 418.800 23.850 420.000 ;
        RECT 4.950 417.600 12.900 418.800 ;
        RECT 4.950 415.050 6.750 417.600 ;
        RECT 11.100 417.000 12.900 417.600 ;
        RECT 8.100 415.800 9.900 416.400 ;
        RECT 4.950 412.950 7.050 415.050 ;
        RECT 8.100 414.600 16.200 415.800 ;
        RECT 14.100 412.950 16.200 414.600 ;
        RECT 12.450 407.700 14.250 408.000 ;
        RECT 2.550 407.100 14.250 407.700 ;
        RECT 2.550 406.500 20.850 407.100 ;
        RECT 2.550 405.600 3.450 406.500 ;
        RECT 12.450 406.200 20.850 406.500 ;
        RECT 2.550 403.800 4.950 405.600 ;
        RECT 3.150 393.600 4.950 403.800 ;
        RECT 6.150 393.000 7.950 405.600 ;
        RECT 17.250 404.700 19.050 405.300 ;
        RECT 11.250 403.500 19.050 404.700 ;
        RECT 19.950 404.100 20.850 406.200 ;
        RECT 22.950 406.200 23.850 418.800 ;
        RECT 35.250 415.050 36.450 422.400 ;
        RECT 30.150 413.250 36.450 415.050 ;
        RECT 31.950 412.950 36.450 413.250 ;
        RECT 26.550 410.100 28.650 410.400 ;
        RECT 32.550 410.100 34.350 410.250 ;
        RECT 26.550 408.900 34.350 410.100 ;
        RECT 26.550 408.300 28.650 408.900 ;
        RECT 32.550 408.450 34.350 408.900 ;
        RECT 22.950 405.300 27.750 406.200 ;
        RECT 35.250 405.600 36.450 412.950 ;
        RECT 26.550 404.400 27.750 405.300 ;
        RECT 23.850 404.100 25.650 404.400 ;
        RECT 11.250 402.600 13.350 403.500 ;
        RECT 19.950 403.200 25.650 404.100 ;
        RECT 23.850 402.600 25.650 403.200 ;
        RECT 26.550 402.600 29.550 404.400 ;
        RECT 11.550 393.600 13.350 402.600 ;
        RECT 15.450 401.550 17.250 402.300 ;
        RECT 20.250 401.550 22.050 402.300 ;
        RECT 15.450 400.500 22.050 401.550 ;
        RECT 16.350 393.000 18.150 399.600 ;
        RECT 19.350 393.600 21.150 400.500 ;
        RECT 26.550 399.600 28.650 401.700 ;
        RECT 22.350 393.000 24.150 399.600 ;
        RECT 26.850 393.600 28.650 399.600 ;
        RECT 31.650 393.000 33.450 405.600 ;
        RECT 34.650 393.600 36.450 405.600 ;
        RECT 38.550 422.400 40.950 424.200 ;
        RECT 42.150 422.400 43.950 429.000 ;
        RECT 46.950 426.300 48.750 428.400 ;
        RECT 45.150 425.400 48.750 426.300 ;
        RECT 51.450 425.400 53.250 429.000 ;
        RECT 54.750 425.400 56.550 428.400 ;
        RECT 57.750 425.400 59.550 429.000 ;
        RECT 62.250 425.400 64.050 428.400 ;
        RECT 44.850 424.800 48.750 425.400 ;
        RECT 44.850 423.300 46.950 424.800 ;
        RECT 54.750 424.500 55.800 425.400 ;
        RECT 38.550 407.700 39.450 422.400 ;
        RECT 47.850 421.800 49.650 423.600 ;
        RECT 50.850 423.450 55.800 424.500 ;
        RECT 50.850 422.700 52.650 423.450 ;
        RECT 62.250 423.300 64.650 425.400 ;
        RECT 67.350 422.400 69.150 429.000 ;
        RECT 70.650 422.400 72.450 428.400 ;
        RECT 47.850 420.000 48.900 421.800 ;
        RECT 58.050 420.000 59.850 420.600 ;
        RECT 47.850 418.800 59.850 420.000 ;
        RECT 40.950 417.600 48.900 418.800 ;
        RECT 40.950 415.050 42.750 417.600 ;
        RECT 47.100 417.000 48.900 417.600 ;
        RECT 44.100 415.800 45.900 416.400 ;
        RECT 40.950 412.950 43.050 415.050 ;
        RECT 44.100 414.600 52.200 415.800 ;
        RECT 50.100 412.950 52.200 414.600 ;
        RECT 48.450 407.700 50.250 408.000 ;
        RECT 38.550 407.100 50.250 407.700 ;
        RECT 38.550 406.500 56.850 407.100 ;
        RECT 38.550 405.600 39.450 406.500 ;
        RECT 48.450 406.200 56.850 406.500 ;
        RECT 38.550 403.800 40.950 405.600 ;
        RECT 39.150 393.600 40.950 403.800 ;
        RECT 42.150 393.000 43.950 405.600 ;
        RECT 53.250 404.700 55.050 405.300 ;
        RECT 47.250 403.500 55.050 404.700 ;
        RECT 55.950 404.100 56.850 406.200 ;
        RECT 58.950 406.200 59.850 418.800 ;
        RECT 71.250 415.050 72.450 422.400 ;
        RECT 86.100 423.300 87.900 428.400 ;
        RECT 89.100 424.200 90.900 429.000 ;
        RECT 92.100 423.300 93.900 428.400 ;
        RECT 86.100 421.950 93.900 423.300 ;
        RECT 95.100 422.400 96.900 428.400 ;
        RECT 99.150 424.200 100.950 428.400 ;
        RECT 98.550 422.400 100.950 424.200 ;
        RECT 102.150 422.400 103.950 429.000 ;
        RECT 106.950 426.300 108.750 428.400 ;
        RECT 105.150 425.400 108.750 426.300 ;
        RECT 111.450 425.400 113.250 429.000 ;
        RECT 114.750 425.400 116.550 428.400 ;
        RECT 117.750 425.400 119.550 429.000 ;
        RECT 122.250 425.400 124.050 428.400 ;
        RECT 104.850 424.800 108.750 425.400 ;
        RECT 104.850 423.300 106.950 424.800 ;
        RECT 114.750 424.500 115.800 425.400 ;
        RECT 95.100 420.300 96.300 422.400 ;
        RECT 92.700 419.400 96.300 420.300 ;
        RECT 89.100 415.050 90.900 416.850 ;
        RECT 92.700 415.050 93.900 419.400 ;
        RECT 95.100 415.050 96.900 416.850 ;
        RECT 66.150 413.250 72.450 415.050 ;
        RECT 67.950 412.950 72.450 413.250 ;
        RECT 85.950 412.950 88.050 415.050 ;
        RECT 88.950 412.950 91.050 415.050 ;
        RECT 91.950 412.950 94.050 415.050 ;
        RECT 94.950 412.950 97.050 415.050 ;
        RECT 62.550 410.100 64.650 410.400 ;
        RECT 68.550 410.100 70.350 410.250 ;
        RECT 62.550 408.900 70.350 410.100 ;
        RECT 62.550 408.300 64.650 408.900 ;
        RECT 68.550 408.450 70.350 408.900 ;
        RECT 58.950 405.300 63.750 406.200 ;
        RECT 71.250 405.600 72.450 412.950 ;
        RECT 86.100 411.150 87.900 412.950 ;
        RECT 92.700 405.600 93.900 412.950 ;
        RECT 62.550 404.400 63.750 405.300 ;
        RECT 59.850 404.100 61.650 404.400 ;
        RECT 47.250 402.600 49.350 403.500 ;
        RECT 55.950 403.200 61.650 404.100 ;
        RECT 59.850 402.600 61.650 403.200 ;
        RECT 62.550 402.600 65.550 404.400 ;
        RECT 47.550 393.600 49.350 402.600 ;
        RECT 51.450 401.550 53.250 402.300 ;
        RECT 56.250 401.550 58.050 402.300 ;
        RECT 51.450 400.500 58.050 401.550 ;
        RECT 52.350 393.000 54.150 399.600 ;
        RECT 55.350 393.600 57.150 400.500 ;
        RECT 62.550 399.600 64.650 401.700 ;
        RECT 58.350 393.000 60.150 399.600 ;
        RECT 62.850 393.600 64.650 399.600 ;
        RECT 67.650 393.000 69.450 405.600 ;
        RECT 70.650 393.600 72.450 405.600 ;
        RECT 86.400 393.000 88.200 405.600 ;
        RECT 91.500 404.100 93.900 405.600 ;
        RECT 98.550 407.700 99.450 422.400 ;
        RECT 107.850 421.800 109.650 423.600 ;
        RECT 110.850 423.450 115.800 424.500 ;
        RECT 110.850 422.700 112.650 423.450 ;
        RECT 122.250 423.300 124.650 425.400 ;
        RECT 127.350 422.400 129.150 429.000 ;
        RECT 130.650 422.400 132.450 428.400 ;
        RECT 149.100 422.400 150.900 428.400 ;
        RECT 107.850 420.000 108.900 421.800 ;
        RECT 118.050 420.000 119.850 420.600 ;
        RECT 107.850 418.800 119.850 420.000 ;
        RECT 100.950 417.600 108.900 418.800 ;
        RECT 100.950 415.050 102.750 417.600 ;
        RECT 107.100 417.000 108.900 417.600 ;
        RECT 104.100 415.800 105.900 416.400 ;
        RECT 100.950 412.950 103.050 415.050 ;
        RECT 104.100 414.600 112.200 415.800 ;
        RECT 110.100 412.950 112.200 414.600 ;
        RECT 108.450 407.700 110.250 408.000 ;
        RECT 98.550 407.100 110.250 407.700 ;
        RECT 98.550 406.500 116.850 407.100 ;
        RECT 98.550 405.600 99.450 406.500 ;
        RECT 108.450 406.200 116.850 406.500 ;
        RECT 91.500 393.600 93.300 404.100 ;
        RECT 98.550 403.800 100.950 405.600 ;
        RECT 94.200 401.100 96.000 402.900 ;
        RECT 94.500 393.000 96.300 399.600 ;
        RECT 99.150 393.600 100.950 403.800 ;
        RECT 102.150 393.000 103.950 405.600 ;
        RECT 113.250 404.700 115.050 405.300 ;
        RECT 107.250 403.500 115.050 404.700 ;
        RECT 115.950 404.100 116.850 406.200 ;
        RECT 118.950 406.200 119.850 418.800 ;
        RECT 131.250 415.050 132.450 422.400 ;
        RECT 149.700 420.300 150.900 422.400 ;
        RECT 152.100 423.300 153.900 428.400 ;
        RECT 155.100 424.200 156.900 429.000 ;
        RECT 158.100 423.300 159.900 428.400 ;
        RECT 152.100 421.950 159.900 423.300 ;
        RECT 176.100 425.400 177.900 428.400 ;
        RECT 176.100 421.500 177.300 425.400 ;
        RECT 179.100 422.400 180.900 429.000 ;
        RECT 182.100 422.400 183.900 428.400 ;
        RECT 200.400 422.400 202.200 429.000 ;
        RECT 176.100 420.600 181.800 421.500 ;
        RECT 149.700 419.400 153.300 420.300 ;
        RECT 149.100 415.050 150.900 416.850 ;
        RECT 152.100 415.050 153.300 419.400 ;
        RECT 180.000 419.700 181.800 420.600 ;
        RECT 155.100 415.050 156.900 416.850 ;
        RECT 126.150 413.250 132.450 415.050 ;
        RECT 127.950 412.950 132.450 413.250 ;
        RECT 148.950 412.950 151.050 415.050 ;
        RECT 151.950 412.950 154.050 415.050 ;
        RECT 154.950 412.950 157.050 415.050 ;
        RECT 157.950 412.950 160.050 415.050 ;
        RECT 176.400 412.950 178.500 415.050 ;
        RECT 122.550 410.100 124.650 410.400 ;
        RECT 128.550 410.100 130.350 410.250 ;
        RECT 122.550 408.900 130.350 410.100 ;
        RECT 122.550 408.300 124.650 408.900 ;
        RECT 128.550 408.450 130.350 408.900 ;
        RECT 118.950 405.300 123.750 406.200 ;
        RECT 131.250 405.600 132.450 412.950 ;
        RECT 122.550 404.400 123.750 405.300 ;
        RECT 119.850 404.100 121.650 404.400 ;
        RECT 107.250 402.600 109.350 403.500 ;
        RECT 115.950 403.200 121.650 404.100 ;
        RECT 119.850 402.600 121.650 403.200 ;
        RECT 122.550 402.600 125.550 404.400 ;
        RECT 107.550 393.600 109.350 402.600 ;
        RECT 111.450 401.550 113.250 402.300 ;
        RECT 116.250 401.550 118.050 402.300 ;
        RECT 111.450 400.500 118.050 401.550 ;
        RECT 112.350 393.000 114.150 399.600 ;
        RECT 115.350 393.600 117.150 400.500 ;
        RECT 122.550 399.600 124.650 401.700 ;
        RECT 118.350 393.000 120.150 399.600 ;
        RECT 122.850 393.600 124.650 399.600 ;
        RECT 127.650 393.000 129.450 405.600 ;
        RECT 130.650 393.600 132.450 405.600 ;
        RECT 152.100 405.600 153.300 412.950 ;
        RECT 158.100 411.150 159.900 412.950 ;
        RECT 176.400 411.150 178.200 412.950 ;
        RECT 154.950 408.450 157.050 409.050 ;
        RECT 166.950 408.450 169.050 409.050 ;
        RECT 154.950 407.550 169.050 408.450 ;
        RECT 154.950 406.950 157.050 407.550 ;
        RECT 166.950 406.950 169.050 407.550 ;
        RECT 180.000 408.300 180.900 419.700 ;
        RECT 182.700 415.050 183.900 422.400 ;
        RECT 205.500 421.200 207.300 428.400 ;
        RECT 221.100 422.400 222.900 428.400 ;
        RECT 203.100 420.300 207.300 421.200 ;
        RECT 221.700 420.300 222.900 422.400 ;
        RECT 224.100 423.300 225.900 428.400 ;
        RECT 227.100 424.200 228.900 429.000 ;
        RECT 230.100 423.300 231.900 428.400 ;
        RECT 224.100 421.950 231.900 423.300 ;
        RECT 248.100 423.300 249.900 428.400 ;
        RECT 251.100 424.200 252.900 429.000 ;
        RECT 254.100 423.300 255.900 428.400 ;
        RECT 248.100 421.950 255.900 423.300 ;
        RECT 257.100 422.400 258.900 428.400 ;
        RECT 272.100 423.300 273.900 428.400 ;
        RECT 275.100 424.200 276.900 429.000 ;
        RECT 278.100 423.300 279.900 428.400 ;
        RECT 257.100 420.300 258.300 422.400 ;
        RECT 272.100 421.950 279.900 423.300 ;
        RECT 281.100 422.400 282.900 428.400 ;
        RECT 299.100 425.400 300.900 429.000 ;
        RECT 302.100 425.400 303.900 428.400 ;
        RECT 305.100 425.400 306.900 429.000 ;
        RECT 281.100 420.300 282.300 422.400 ;
        RECT 200.250 415.050 202.050 416.850 ;
        RECT 203.100 415.050 204.300 420.300 ;
        RECT 221.700 419.400 225.300 420.300 ;
        RECT 206.100 415.050 207.900 416.850 ;
        RECT 221.100 415.050 222.900 416.850 ;
        RECT 224.100 415.050 225.300 419.400 ;
        RECT 254.700 419.400 258.300 420.300 ;
        RECT 278.700 419.400 282.300 420.300 ;
        RECT 227.100 415.050 228.900 416.850 ;
        RECT 251.100 415.050 252.900 416.850 ;
        RECT 254.700 415.050 255.900 419.400 ;
        RECT 257.100 415.050 258.900 416.850 ;
        RECT 275.100 415.050 276.900 416.850 ;
        RECT 278.700 415.050 279.900 419.400 ;
        RECT 281.100 415.050 282.900 416.850 ;
        RECT 302.700 415.050 303.600 425.400 ;
        RECT 309.150 424.200 310.950 428.400 ;
        RECT 308.550 422.400 310.950 424.200 ;
        RECT 312.150 422.400 313.950 429.000 ;
        RECT 316.950 426.300 318.750 428.400 ;
        RECT 315.150 425.400 318.750 426.300 ;
        RECT 321.450 425.400 323.250 429.000 ;
        RECT 324.750 425.400 326.550 428.400 ;
        RECT 327.750 425.400 329.550 429.000 ;
        RECT 332.250 425.400 334.050 428.400 ;
        RECT 314.850 424.800 318.750 425.400 ;
        RECT 314.850 423.300 316.950 424.800 ;
        RECT 324.750 424.500 325.800 425.400 ;
        RECT 181.800 412.950 183.900 415.050 ;
        RECT 199.950 412.950 202.050 415.050 ;
        RECT 202.950 412.950 205.050 415.050 ;
        RECT 205.950 412.950 208.050 415.050 ;
        RECT 220.950 412.950 223.050 415.050 ;
        RECT 223.950 412.950 226.050 415.050 ;
        RECT 226.950 412.950 229.050 415.050 ;
        RECT 229.950 412.950 232.050 415.050 ;
        RECT 247.950 412.950 250.050 415.050 ;
        RECT 250.950 412.950 253.050 415.050 ;
        RECT 253.950 412.950 256.050 415.050 ;
        RECT 256.950 412.950 259.050 415.050 ;
        RECT 271.950 412.950 274.050 415.050 ;
        RECT 274.950 412.950 277.050 415.050 ;
        RECT 277.950 412.950 280.050 415.050 ;
        RECT 280.950 412.950 283.050 415.050 ;
        RECT 298.950 412.950 301.050 415.050 ;
        RECT 301.950 412.950 304.050 415.050 ;
        RECT 304.950 412.950 307.050 415.050 ;
        RECT 180.000 407.400 181.800 408.300 ;
        RECT 176.100 406.500 181.800 407.400 ;
        RECT 152.100 404.100 154.500 405.600 ;
        RECT 150.000 401.100 151.800 402.900 ;
        RECT 149.700 393.000 151.500 399.600 ;
        RECT 152.700 393.600 154.500 404.100 ;
        RECT 157.800 393.000 159.600 405.600 ;
        RECT 176.100 399.600 177.300 406.500 ;
        RECT 182.700 405.600 183.900 412.950 ;
        RECT 176.100 393.600 177.900 399.600 ;
        RECT 179.100 393.000 180.900 403.800 ;
        RECT 182.100 393.600 183.900 405.600 ;
        RECT 203.100 399.600 204.300 412.950 ;
        RECT 224.100 405.600 225.300 412.950 ;
        RECT 230.100 411.150 231.900 412.950 ;
        RECT 248.100 411.150 249.900 412.950 ;
        RECT 254.700 405.600 255.900 412.950 ;
        RECT 272.100 411.150 273.900 412.950 ;
        RECT 262.950 408.450 265.050 409.050 ;
        RECT 274.950 408.450 277.050 408.750 ;
        RECT 262.950 407.550 277.050 408.450 ;
        RECT 262.950 406.950 265.050 407.550 ;
        RECT 274.950 406.650 277.050 407.550 ;
        RECT 278.700 405.600 279.900 412.950 ;
        RECT 299.100 411.150 300.900 412.950 ;
        RECT 289.950 408.450 292.050 409.050 ;
        RECT 295.950 408.450 300.000 409.050 ;
        RECT 289.950 407.550 300.450 408.450 ;
        RECT 289.950 406.950 292.050 407.550 ;
        RECT 295.950 406.950 300.000 407.550 ;
        RECT 224.100 404.100 226.500 405.600 ;
        RECT 222.000 401.100 223.800 402.900 ;
        RECT 200.100 393.000 201.900 399.600 ;
        RECT 203.100 393.600 204.900 399.600 ;
        RECT 206.100 393.000 207.900 399.600 ;
        RECT 221.700 393.000 223.500 399.600 ;
        RECT 224.700 393.600 226.500 404.100 ;
        RECT 229.800 393.000 231.600 405.600 ;
        RECT 248.400 393.000 250.200 405.600 ;
        RECT 253.500 404.100 255.900 405.600 ;
        RECT 253.500 393.600 255.300 404.100 ;
        RECT 256.200 401.100 258.000 402.900 ;
        RECT 256.500 393.000 258.300 399.600 ;
        RECT 272.400 393.000 274.200 405.600 ;
        RECT 277.500 404.100 279.900 405.600 ;
        RECT 280.950 405.450 283.050 406.050 ;
        RECT 292.950 405.450 295.050 405.900 ;
        RECT 302.700 405.600 303.600 412.950 ;
        RECT 304.950 411.150 306.750 412.950 ;
        RECT 308.550 407.700 309.450 422.400 ;
        RECT 317.850 421.800 319.650 423.600 ;
        RECT 320.850 423.450 325.800 424.500 ;
        RECT 320.850 422.700 322.650 423.450 ;
        RECT 332.250 423.300 334.650 425.400 ;
        RECT 337.350 422.400 339.150 429.000 ;
        RECT 340.650 422.400 342.450 428.400 ;
        RECT 345.150 424.200 346.950 428.400 ;
        RECT 317.850 420.000 318.900 421.800 ;
        RECT 328.050 420.000 329.850 420.600 ;
        RECT 317.850 418.800 329.850 420.000 ;
        RECT 310.950 417.600 318.900 418.800 ;
        RECT 310.950 415.050 312.750 417.600 ;
        RECT 317.100 417.000 318.900 417.600 ;
        RECT 314.100 415.800 315.900 416.400 ;
        RECT 310.950 412.950 313.050 415.050 ;
        RECT 314.100 414.600 322.200 415.800 ;
        RECT 320.100 412.950 322.200 414.600 ;
        RECT 318.450 407.700 320.250 408.000 ;
        RECT 308.550 407.100 320.250 407.700 ;
        RECT 308.550 406.500 326.850 407.100 ;
        RECT 308.550 405.600 309.450 406.500 ;
        RECT 318.450 406.200 326.850 406.500 ;
        RECT 280.950 404.550 295.050 405.450 ;
        RECT 277.500 393.600 279.300 404.100 ;
        RECT 280.950 403.950 283.050 404.550 ;
        RECT 292.950 403.800 295.050 404.550 ;
        RECT 300.000 404.400 303.600 405.600 ;
        RECT 280.200 401.100 282.000 402.900 ;
        RECT 280.500 393.000 282.300 399.600 ;
        RECT 300.000 393.600 301.800 404.400 ;
        RECT 305.100 393.000 306.900 405.600 ;
        RECT 308.550 403.800 310.950 405.600 ;
        RECT 309.150 393.600 310.950 403.800 ;
        RECT 312.150 393.000 313.950 405.600 ;
        RECT 323.250 404.700 325.050 405.300 ;
        RECT 317.250 403.500 325.050 404.700 ;
        RECT 325.950 404.100 326.850 406.200 ;
        RECT 328.950 406.200 329.850 418.800 ;
        RECT 341.250 415.050 342.450 422.400 ;
        RECT 336.150 413.250 342.450 415.050 ;
        RECT 337.950 412.950 342.450 413.250 ;
        RECT 332.550 410.100 334.650 410.400 ;
        RECT 338.550 410.100 340.350 410.250 ;
        RECT 332.550 408.900 340.350 410.100 ;
        RECT 332.550 408.300 334.650 408.900 ;
        RECT 338.550 408.450 340.350 408.900 ;
        RECT 328.950 405.300 333.750 406.200 ;
        RECT 341.250 405.600 342.450 412.950 ;
        RECT 332.550 404.400 333.750 405.300 ;
        RECT 329.850 404.100 331.650 404.400 ;
        RECT 317.250 402.600 319.350 403.500 ;
        RECT 325.950 403.200 331.650 404.100 ;
        RECT 329.850 402.600 331.650 403.200 ;
        RECT 332.550 402.600 335.550 404.400 ;
        RECT 317.550 393.600 319.350 402.600 ;
        RECT 321.450 401.550 323.250 402.300 ;
        RECT 326.250 401.550 328.050 402.300 ;
        RECT 321.450 400.500 328.050 401.550 ;
        RECT 322.350 393.000 324.150 399.600 ;
        RECT 325.350 393.600 327.150 400.500 ;
        RECT 332.550 399.600 334.650 401.700 ;
        RECT 328.350 393.000 330.150 399.600 ;
        RECT 332.850 393.600 334.650 399.600 ;
        RECT 337.650 393.000 339.450 405.600 ;
        RECT 340.650 393.600 342.450 405.600 ;
        RECT 344.550 422.400 346.950 424.200 ;
        RECT 348.150 422.400 349.950 429.000 ;
        RECT 352.950 426.300 354.750 428.400 ;
        RECT 351.150 425.400 354.750 426.300 ;
        RECT 357.450 425.400 359.250 429.000 ;
        RECT 360.750 425.400 362.550 428.400 ;
        RECT 363.750 425.400 365.550 429.000 ;
        RECT 368.250 425.400 370.050 428.400 ;
        RECT 350.850 424.800 354.750 425.400 ;
        RECT 350.850 423.300 352.950 424.800 ;
        RECT 360.750 424.500 361.800 425.400 ;
        RECT 344.550 407.700 345.450 422.400 ;
        RECT 353.850 421.800 355.650 423.600 ;
        RECT 356.850 423.450 361.800 424.500 ;
        RECT 356.850 422.700 358.650 423.450 ;
        RECT 368.250 423.300 370.650 425.400 ;
        RECT 373.350 422.400 375.150 429.000 ;
        RECT 376.650 422.400 378.450 428.400 ;
        RECT 392.100 425.400 393.900 428.400 ;
        RECT 395.100 425.400 396.900 429.000 ;
        RECT 353.850 420.000 354.900 421.800 ;
        RECT 364.050 420.000 365.850 420.600 ;
        RECT 353.850 418.800 365.850 420.000 ;
        RECT 346.950 417.600 354.900 418.800 ;
        RECT 346.950 415.050 348.750 417.600 ;
        RECT 353.100 417.000 354.900 417.600 ;
        RECT 350.100 415.800 351.900 416.400 ;
        RECT 346.950 412.950 349.050 415.050 ;
        RECT 350.100 414.600 358.200 415.800 ;
        RECT 356.100 412.950 358.200 414.600 ;
        RECT 354.450 407.700 356.250 408.000 ;
        RECT 344.550 407.100 356.250 407.700 ;
        RECT 344.550 406.500 362.850 407.100 ;
        RECT 344.550 405.600 345.450 406.500 ;
        RECT 354.450 406.200 362.850 406.500 ;
        RECT 344.550 403.800 346.950 405.600 ;
        RECT 345.150 393.600 346.950 403.800 ;
        RECT 348.150 393.000 349.950 405.600 ;
        RECT 359.250 404.700 361.050 405.300 ;
        RECT 353.250 403.500 361.050 404.700 ;
        RECT 361.950 404.100 362.850 406.200 ;
        RECT 364.950 406.200 365.850 418.800 ;
        RECT 377.250 415.050 378.450 422.400 ;
        RECT 392.700 415.050 393.900 425.400 ;
        RECT 410.100 422.400 411.900 429.000 ;
        RECT 413.100 421.500 414.900 428.400 ;
        RECT 416.100 422.400 417.900 429.000 ;
        RECT 419.100 421.500 420.900 428.400 ;
        RECT 422.100 422.400 423.900 429.000 ;
        RECT 425.100 421.500 426.900 428.400 ;
        RECT 428.100 422.400 429.900 429.000 ;
        RECT 431.100 421.500 432.900 428.400 ;
        RECT 434.100 422.400 435.900 429.000 ;
        RECT 449.700 422.400 451.500 429.000 ;
        RECT 454.200 422.400 456.000 428.400 ;
        RECT 458.700 422.400 460.500 429.000 ;
        RECT 476.100 422.400 477.900 428.400 ;
        RECT 479.100 422.400 480.900 429.000 ;
        RECT 482.100 425.400 483.900 428.400 ;
        RECT 413.100 420.300 417.000 421.500 ;
        RECT 419.100 420.300 423.000 421.500 ;
        RECT 425.100 420.300 429.000 421.500 ;
        RECT 431.100 420.300 433.950 421.500 ;
        RECT 415.800 419.400 417.000 420.300 ;
        RECT 421.800 419.400 423.000 420.300 ;
        RECT 427.800 419.400 429.000 420.300 ;
        RECT 415.800 418.200 420.000 419.400 ;
        RECT 412.800 415.050 414.600 416.850 ;
        RECT 372.150 413.250 378.450 415.050 ;
        RECT 373.950 412.950 378.450 413.250 ;
        RECT 391.950 412.950 394.050 415.050 ;
        RECT 394.950 412.950 397.050 415.050 ;
        RECT 412.800 412.950 414.900 415.050 ;
        RECT 368.550 410.100 370.650 410.400 ;
        RECT 374.550 410.100 376.350 410.250 ;
        RECT 368.550 408.900 376.350 410.100 ;
        RECT 368.550 408.300 370.650 408.900 ;
        RECT 374.550 408.450 376.350 408.900 ;
        RECT 364.950 405.300 369.750 406.200 ;
        RECT 377.250 405.600 378.450 412.950 ;
        RECT 368.550 404.400 369.750 405.300 ;
        RECT 365.850 404.100 367.650 404.400 ;
        RECT 353.250 402.600 355.350 403.500 ;
        RECT 361.950 403.200 367.650 404.100 ;
        RECT 365.850 402.600 367.650 403.200 ;
        RECT 368.550 402.600 371.550 404.400 ;
        RECT 353.550 393.600 355.350 402.600 ;
        RECT 357.450 401.550 359.250 402.300 ;
        RECT 362.250 401.550 364.050 402.300 ;
        RECT 357.450 400.500 364.050 401.550 ;
        RECT 358.350 393.000 360.150 399.600 ;
        RECT 361.350 393.600 363.150 400.500 ;
        RECT 368.550 399.600 370.650 401.700 ;
        RECT 364.350 393.000 366.150 399.600 ;
        RECT 368.850 393.600 370.650 399.600 ;
        RECT 373.650 393.000 375.450 405.600 ;
        RECT 376.650 393.600 378.450 405.600 ;
        RECT 392.700 399.600 393.900 412.950 ;
        RECT 395.100 411.150 396.900 412.950 ;
        RECT 415.800 407.700 417.000 418.200 ;
        RECT 418.200 417.600 420.000 418.200 ;
        RECT 421.800 418.200 426.000 419.400 ;
        RECT 421.800 407.700 423.000 418.200 ;
        RECT 424.200 417.600 426.000 418.200 ;
        RECT 427.800 418.200 432.000 419.400 ;
        RECT 427.800 407.700 429.000 418.200 ;
        RECT 430.200 417.600 432.000 418.200 ;
        RECT 432.900 415.050 433.950 420.300 ;
        RECT 442.950 420.450 445.050 421.050 ;
        RECT 451.950 420.450 454.050 421.050 ;
        RECT 442.950 419.550 454.050 420.450 ;
        RECT 442.950 418.950 445.050 419.550 ;
        RECT 451.950 418.950 454.050 419.550 ;
        RECT 449.250 415.050 451.050 416.850 ;
        RECT 455.100 415.050 456.300 422.400 ;
        RECT 461.100 415.050 462.900 416.850 ;
        RECT 476.100 415.050 477.300 422.400 ;
        RECT 482.700 421.500 483.900 425.400 ;
        RECT 478.200 420.600 483.900 421.500 ;
        RECT 497.100 425.400 498.900 428.400 ;
        RECT 497.100 421.500 498.300 425.400 ;
        RECT 500.100 422.400 501.900 429.000 ;
        RECT 503.100 422.400 504.900 428.400 ;
        RECT 497.100 420.600 502.800 421.500 ;
        RECT 478.200 419.700 480.000 420.600 ;
        RECT 430.800 412.950 433.950 415.050 ;
        RECT 448.950 412.950 451.050 415.050 ;
        RECT 451.950 412.950 454.050 415.050 ;
        RECT 454.950 412.950 457.050 415.050 ;
        RECT 457.950 412.950 460.050 415.050 ;
        RECT 460.950 412.950 463.050 415.050 ;
        RECT 476.100 412.950 478.200 415.050 ;
        RECT 432.900 407.700 433.950 412.950 ;
        RECT 452.250 411.150 454.050 412.950 ;
        RECT 413.100 406.500 417.000 407.700 ;
        RECT 419.100 406.500 423.000 407.700 ;
        RECT 425.100 406.500 429.000 407.700 ;
        RECT 431.100 406.500 433.950 407.700 ;
        RECT 455.100 407.400 456.000 412.950 ;
        RECT 458.100 411.150 459.900 412.950 ;
        RECT 455.100 406.500 459.900 407.400 ;
        RECT 392.100 393.600 393.900 399.600 ;
        RECT 395.100 393.000 396.900 399.600 ;
        RECT 410.100 393.000 411.900 405.600 ;
        RECT 413.100 393.600 414.900 406.500 ;
        RECT 416.100 393.000 417.900 405.600 ;
        RECT 419.100 393.600 420.900 406.500 ;
        RECT 422.100 393.000 423.900 405.600 ;
        RECT 425.100 393.600 426.900 406.500 ;
        RECT 428.100 393.000 429.900 405.600 ;
        RECT 431.100 393.600 432.900 406.500 ;
        RECT 434.100 393.000 435.900 405.600 ;
        RECT 449.100 404.400 456.900 405.300 ;
        RECT 449.100 393.600 450.900 404.400 ;
        RECT 452.100 393.000 453.900 403.500 ;
        RECT 455.100 394.500 456.900 404.400 ;
        RECT 458.100 395.400 459.900 406.500 ;
        RECT 476.100 405.600 477.300 412.950 ;
        RECT 479.100 408.300 480.000 419.700 ;
        RECT 501.000 419.700 502.800 420.600 ;
        RECT 481.500 412.950 483.600 415.050 ;
        RECT 481.800 411.150 483.600 412.950 ;
        RECT 497.400 412.950 499.500 415.050 ;
        RECT 497.400 411.150 499.200 412.950 ;
        RECT 478.200 407.400 480.000 408.300 ;
        RECT 501.000 408.300 501.900 419.700 ;
        RECT 503.700 415.050 504.900 422.400 ;
        RECT 518.100 425.400 519.900 428.400 ;
        RECT 518.100 421.500 519.300 425.400 ;
        RECT 521.100 422.400 522.900 429.000 ;
        RECT 524.100 422.400 525.900 428.400 ;
        RECT 539.100 422.400 540.900 428.400 ;
        RECT 518.100 420.600 523.800 421.500 ;
        RECT 522.000 419.700 523.800 420.600 ;
        RECT 502.800 412.950 504.900 415.050 ;
        RECT 501.000 407.400 502.800 408.300 ;
        RECT 478.200 406.500 483.900 407.400 ;
        RECT 461.100 394.500 462.900 405.600 ;
        RECT 455.100 393.600 462.900 394.500 ;
        RECT 476.100 393.600 477.900 405.600 ;
        RECT 479.100 393.000 480.900 403.800 ;
        RECT 482.700 399.600 483.900 406.500 ;
        RECT 482.100 393.600 483.900 399.600 ;
        RECT 497.100 406.500 502.800 407.400 ;
        RECT 497.100 399.600 498.300 406.500 ;
        RECT 503.700 405.600 504.900 412.950 ;
        RECT 518.400 412.950 520.500 415.050 ;
        RECT 518.400 411.150 520.200 412.950 ;
        RECT 522.000 408.300 522.900 419.700 ;
        RECT 524.700 415.050 525.900 422.400 ;
        RECT 539.700 420.300 540.900 422.400 ;
        RECT 542.100 423.300 543.900 428.400 ;
        RECT 545.100 424.200 546.900 429.000 ;
        RECT 548.100 423.300 549.900 428.400 ;
        RECT 563.100 425.400 564.900 428.400 ;
        RECT 566.100 425.400 567.900 429.000 ;
        RECT 542.100 421.950 549.900 423.300 ;
        RECT 539.700 419.400 543.300 420.300 ;
        RECT 539.100 415.050 540.900 416.850 ;
        RECT 542.100 415.050 543.300 419.400 ;
        RECT 550.950 417.450 555.000 418.050 ;
        RECT 545.100 415.050 546.900 416.850 ;
        RECT 550.950 415.950 555.450 417.450 ;
        RECT 556.950 415.950 559.050 418.050 ;
        RECT 523.800 412.950 525.900 415.050 ;
        RECT 538.950 412.950 541.050 415.050 ;
        RECT 541.950 412.950 544.050 415.050 ;
        RECT 544.950 412.950 547.050 415.050 ;
        RECT 547.950 412.950 550.050 415.050 ;
        RECT 522.000 407.400 523.800 408.300 ;
        RECT 497.100 393.600 498.900 399.600 ;
        RECT 500.100 393.000 501.900 403.800 ;
        RECT 503.100 393.600 504.900 405.600 ;
        RECT 518.100 406.500 523.800 407.400 ;
        RECT 518.100 399.600 519.300 406.500 ;
        RECT 524.700 405.600 525.900 412.950 ;
        RECT 529.950 408.450 532.050 409.050 ;
        RECT 538.950 408.450 541.050 409.050 ;
        RECT 529.950 407.550 541.050 408.450 ;
        RECT 529.950 406.950 532.050 407.550 ;
        RECT 538.950 406.950 541.050 407.550 ;
        RECT 518.100 393.600 519.900 399.600 ;
        RECT 521.100 393.000 522.900 403.800 ;
        RECT 524.100 393.600 525.900 405.600 ;
        RECT 542.100 405.600 543.300 412.950 ;
        RECT 548.100 411.150 549.900 412.950 ;
        RECT 554.550 412.050 555.450 415.950 ;
        RECT 550.950 410.550 555.450 412.050 ;
        RECT 557.550 412.050 558.450 415.950 ;
        RECT 563.700 415.050 564.900 425.400 ;
        RECT 569.550 422.400 571.350 428.400 ;
        RECT 572.850 422.400 574.650 429.000 ;
        RECT 577.950 425.400 579.750 428.400 ;
        RECT 582.450 425.400 584.250 429.000 ;
        RECT 585.450 425.400 587.250 428.400 ;
        RECT 588.750 425.400 590.550 429.000 ;
        RECT 593.250 426.300 595.050 428.400 ;
        RECT 593.250 425.400 596.850 426.300 ;
        RECT 577.350 423.300 579.750 425.400 ;
        RECT 586.200 424.500 587.250 425.400 ;
        RECT 593.250 424.800 597.150 425.400 ;
        RECT 586.200 423.450 591.150 424.500 ;
        RECT 589.350 422.700 591.150 423.450 ;
        RECT 569.550 415.050 570.750 422.400 ;
        RECT 592.350 421.800 594.150 423.600 ;
        RECT 595.050 423.300 597.150 424.800 ;
        RECT 598.050 422.400 599.850 429.000 ;
        RECT 601.050 424.200 602.850 428.400 ;
        RECT 601.050 422.400 603.450 424.200 ;
        RECT 617.400 422.400 619.200 429.000 ;
        RECT 582.150 420.000 583.950 420.600 ;
        RECT 593.100 420.000 594.150 421.800 ;
        RECT 582.150 418.800 594.150 420.000 ;
        RECT 562.950 412.950 565.050 415.050 ;
        RECT 565.950 412.950 568.050 415.050 ;
        RECT 569.550 413.250 575.850 415.050 ;
        RECT 569.550 412.950 574.050 413.250 ;
        RECT 557.550 410.550 562.050 412.050 ;
        RECT 550.950 409.950 555.000 410.550 ;
        RECT 558.000 409.950 562.050 410.550 ;
        RECT 542.100 404.100 544.500 405.600 ;
        RECT 540.000 401.100 541.800 402.900 ;
        RECT 539.700 393.000 541.500 399.600 ;
        RECT 542.700 393.600 544.500 404.100 ;
        RECT 547.800 393.000 549.600 405.600 ;
        RECT 563.700 399.600 564.900 412.950 ;
        RECT 566.100 411.150 567.900 412.950 ;
        RECT 569.550 405.600 570.750 412.950 ;
        RECT 571.650 410.100 573.450 410.250 ;
        RECT 577.350 410.100 579.450 410.400 ;
        RECT 571.650 408.900 579.450 410.100 ;
        RECT 571.650 408.450 573.450 408.900 ;
        RECT 577.350 408.300 579.450 408.900 ;
        RECT 582.150 406.200 583.050 418.800 ;
        RECT 593.100 417.600 601.050 418.800 ;
        RECT 593.100 417.000 594.900 417.600 ;
        RECT 596.100 415.800 597.900 416.400 ;
        RECT 589.800 414.600 597.900 415.800 ;
        RECT 599.250 415.050 601.050 417.600 ;
        RECT 589.800 412.950 591.900 414.600 ;
        RECT 598.950 412.950 601.050 415.050 ;
        RECT 591.750 407.700 593.550 408.000 ;
        RECT 602.550 407.700 603.450 422.400 ;
        RECT 622.500 421.200 624.300 428.400 ;
        RECT 638.100 422.400 639.900 428.400 ;
        RECT 620.100 420.300 624.300 421.200 ;
        RECT 638.700 420.300 639.900 422.400 ;
        RECT 641.100 423.300 642.900 428.400 ;
        RECT 644.100 424.200 645.900 429.000 ;
        RECT 647.100 423.300 648.900 428.400 ;
        RECT 641.100 421.950 648.900 423.300 ;
        RECT 662.700 421.200 664.500 428.400 ;
        RECT 667.800 422.400 669.600 429.000 ;
        RECT 683.700 422.400 685.500 429.000 ;
        RECT 688.200 422.400 690.000 428.400 ;
        RECT 692.700 422.400 694.500 429.000 ;
        RECT 713.100 425.400 714.900 429.000 ;
        RECT 716.100 425.400 717.900 428.400 ;
        RECT 662.700 420.300 666.900 421.200 ;
        RECT 617.250 415.050 619.050 416.850 ;
        RECT 620.100 415.050 621.300 420.300 ;
        RECT 638.700 419.400 642.300 420.300 ;
        RECT 623.100 415.050 624.900 416.850 ;
        RECT 638.100 415.050 639.900 416.850 ;
        RECT 641.100 415.050 642.300 419.400 ;
        RECT 649.950 417.450 652.050 418.050 ;
        RECT 655.950 417.450 658.050 418.050 ;
        RECT 644.100 415.050 645.900 416.850 ;
        RECT 649.950 416.550 658.050 417.450 ;
        RECT 649.950 415.950 652.050 416.550 ;
        RECT 655.950 415.950 658.050 416.550 ;
        RECT 662.100 415.050 663.900 416.850 ;
        RECT 665.700 415.050 666.900 420.300 ;
        RECT 667.950 415.050 669.750 416.850 ;
        RECT 683.250 415.050 685.050 416.850 ;
        RECT 689.100 415.050 690.300 422.400 ;
        RECT 695.100 415.050 696.900 416.850 ;
        RECT 716.100 415.050 717.300 425.400 ;
        RECT 735.600 424.200 737.400 428.400 ;
        RECT 734.700 422.400 737.400 424.200 ;
        RECT 738.600 422.400 740.400 429.000 ;
        RECT 734.700 415.050 735.600 422.400 ;
        RECT 736.500 420.600 738.300 421.500 ;
        RECT 743.100 420.600 744.900 428.400 ;
        RECT 736.500 419.700 744.900 420.600 ;
        RECT 758.100 420.600 759.900 428.400 ;
        RECT 762.600 422.400 764.400 429.000 ;
        RECT 765.600 424.200 767.400 428.400 ;
        RECT 765.600 422.400 768.300 424.200 ;
        RECT 782.400 422.400 784.200 429.000 ;
        RECT 764.700 420.600 766.500 421.500 ;
        RECT 758.100 419.700 766.500 420.600 ;
        RECT 616.950 412.950 619.050 415.050 ;
        RECT 619.950 412.950 622.050 415.050 ;
        RECT 622.950 412.950 625.050 415.050 ;
        RECT 637.950 412.950 640.050 415.050 ;
        RECT 640.950 412.950 643.050 415.050 ;
        RECT 643.950 412.950 646.050 415.050 ;
        RECT 646.950 412.950 649.050 415.050 ;
        RECT 661.950 412.950 664.050 415.050 ;
        RECT 664.950 412.950 667.050 415.050 ;
        RECT 667.950 412.950 670.050 415.050 ;
        RECT 682.950 412.950 685.050 415.050 ;
        RECT 685.950 412.950 688.050 415.050 ;
        RECT 688.950 412.950 691.050 415.050 ;
        RECT 691.950 412.950 694.050 415.050 ;
        RECT 694.950 412.950 697.050 415.050 ;
        RECT 712.950 412.950 715.050 415.050 ;
        RECT 715.950 412.950 718.050 415.050 ;
        RECT 734.100 412.950 736.200 415.050 ;
        RECT 737.400 412.950 739.500 415.050 ;
        RECT 591.750 407.100 603.450 407.700 ;
        RECT 563.100 393.600 564.900 399.600 ;
        RECT 566.100 393.000 567.900 399.600 ;
        RECT 569.550 393.600 571.350 405.600 ;
        RECT 572.550 393.000 574.350 405.600 ;
        RECT 578.250 405.300 583.050 406.200 ;
        RECT 585.150 406.500 603.450 407.100 ;
        RECT 585.150 406.200 593.550 406.500 ;
        RECT 578.250 404.400 579.450 405.300 ;
        RECT 576.450 402.600 579.450 404.400 ;
        RECT 580.350 404.100 582.150 404.400 ;
        RECT 585.150 404.100 586.050 406.200 ;
        RECT 602.550 405.600 603.450 406.500 ;
        RECT 580.350 403.200 586.050 404.100 ;
        RECT 586.950 404.700 588.750 405.300 ;
        RECT 586.950 403.500 594.750 404.700 ;
        RECT 580.350 402.600 582.150 403.200 ;
        RECT 592.650 402.600 594.750 403.500 ;
        RECT 577.350 399.600 579.450 401.700 ;
        RECT 583.950 401.550 585.750 402.300 ;
        RECT 588.750 401.550 590.550 402.300 ;
        RECT 583.950 400.500 590.550 401.550 ;
        RECT 577.350 393.600 579.150 399.600 ;
        RECT 581.850 393.000 583.650 399.600 ;
        RECT 584.850 393.600 586.650 400.500 ;
        RECT 587.850 393.000 589.650 399.600 ;
        RECT 592.650 393.600 594.450 402.600 ;
        RECT 598.050 393.000 599.850 405.600 ;
        RECT 601.050 403.800 603.450 405.600 ;
        RECT 601.050 393.600 602.850 403.800 ;
        RECT 620.100 399.600 621.300 412.950 ;
        RECT 641.100 405.600 642.300 412.950 ;
        RECT 647.100 411.150 648.900 412.950 ;
        RECT 641.100 404.100 643.500 405.600 ;
        RECT 639.000 401.100 640.800 402.900 ;
        RECT 617.100 393.000 618.900 399.600 ;
        RECT 620.100 393.600 621.900 399.600 ;
        RECT 623.100 393.000 624.900 399.600 ;
        RECT 638.700 393.000 640.500 399.600 ;
        RECT 641.700 393.600 643.500 404.100 ;
        RECT 646.800 393.000 648.600 405.600 ;
        RECT 665.700 399.600 666.900 412.950 ;
        RECT 686.250 411.150 688.050 412.950 ;
        RECT 676.950 408.450 679.050 409.050 ;
        RECT 685.950 408.450 688.050 409.050 ;
        RECT 676.950 407.550 688.050 408.450 ;
        RECT 676.950 406.950 679.050 407.550 ;
        RECT 685.950 406.950 688.050 407.550 ;
        RECT 689.100 407.400 690.000 412.950 ;
        RECT 692.100 411.150 693.900 412.950 ;
        RECT 713.100 411.150 714.900 412.950 ;
        RECT 689.100 406.500 693.900 407.400 ;
        RECT 683.100 404.400 690.900 405.300 ;
        RECT 662.100 393.000 663.900 399.600 ;
        RECT 665.100 393.600 666.900 399.600 ;
        RECT 668.100 393.000 669.900 399.600 ;
        RECT 683.100 393.600 684.900 404.400 ;
        RECT 686.100 393.000 687.900 403.500 ;
        RECT 689.100 394.500 690.900 404.400 ;
        RECT 692.100 395.400 693.900 406.500 ;
        RECT 695.100 394.500 696.900 405.600 ;
        RECT 716.100 399.600 717.300 412.950 ;
        RECT 734.700 405.600 735.600 412.950 ;
        RECT 738.000 411.150 739.800 412.950 ;
        RECT 689.100 393.600 696.900 394.500 ;
        RECT 713.100 393.000 714.900 399.600 ;
        RECT 716.100 393.600 717.900 399.600 ;
        RECT 734.100 393.600 735.900 405.600 ;
        RECT 737.100 393.000 738.900 405.000 ;
        RECT 741.000 399.600 741.900 419.700 ;
        RECT 742.950 415.050 744.750 416.850 ;
        RECT 758.250 415.050 760.050 416.850 ;
        RECT 742.800 412.950 744.900 415.050 ;
        RECT 758.100 412.950 760.200 415.050 ;
        RECT 761.100 399.600 762.000 419.700 ;
        RECT 767.400 415.050 768.300 422.400 ;
        RECT 787.500 421.200 789.300 428.400 ;
        RECT 803.100 422.400 804.900 428.400 ;
        RECT 785.100 420.300 789.300 421.200 ;
        RECT 803.700 420.300 804.900 422.400 ;
        RECT 806.100 423.300 807.900 428.400 ;
        RECT 809.100 424.200 810.900 429.000 ;
        RECT 812.100 423.300 813.900 428.400 ;
        RECT 827.100 425.400 828.900 429.000 ;
        RECT 830.100 425.400 831.900 428.400 ;
        RECT 806.100 421.950 813.900 423.300 ;
        RECT 782.250 415.050 784.050 416.850 ;
        RECT 785.100 415.050 786.300 420.300 ;
        RECT 803.700 419.400 807.300 420.300 ;
        RECT 788.100 415.050 789.900 416.850 ;
        RECT 803.100 415.050 804.900 416.850 ;
        RECT 806.100 415.050 807.300 419.400 ;
        RECT 809.100 415.050 810.900 416.850 ;
        RECT 830.100 415.050 831.300 425.400 ;
        RECT 850.500 420.000 852.300 428.400 ;
        RECT 849.000 418.800 852.300 420.000 ;
        RECT 857.100 419.400 858.900 429.000 ;
        RECT 873.000 422.400 874.800 429.000 ;
        RECT 877.500 423.600 879.300 428.400 ;
        RECT 880.500 425.400 882.300 429.000 ;
        RECT 877.500 422.400 882.600 423.600 ;
        RECT 849.000 415.050 849.900 418.800 ;
        RECT 851.100 415.050 852.900 416.850 ;
        RECT 857.100 415.050 858.900 416.850 ;
        RECT 872.100 415.050 873.900 416.850 ;
        RECT 878.250 415.050 880.050 416.850 ;
        RECT 881.700 415.050 882.600 422.400 ;
        RECT 899.100 423.300 900.900 428.400 ;
        RECT 902.100 424.200 903.900 429.000 ;
        RECT 905.100 423.300 906.900 428.400 ;
        RECT 899.100 421.950 906.900 423.300 ;
        RECT 908.100 422.400 909.900 428.400 ;
        RECT 923.100 423.300 924.900 428.400 ;
        RECT 926.100 424.200 927.900 429.000 ;
        RECT 929.100 423.300 930.900 428.400 ;
        RECT 908.100 420.300 909.300 422.400 ;
        RECT 923.100 421.950 930.900 423.300 ;
        RECT 932.100 422.400 933.900 428.400 ;
        RECT 932.100 420.300 933.300 422.400 ;
        RECT 905.700 419.400 909.300 420.300 ;
        RECT 929.700 419.400 933.300 420.300 ;
        RECT 949.500 420.000 951.300 428.400 ;
        RECT 902.100 415.050 903.900 416.850 ;
        RECT 905.700 415.050 906.900 419.400 ;
        RECT 910.950 417.450 915.000 418.050 ;
        RECT 918.000 417.450 922.050 418.050 ;
        RECT 908.100 415.050 909.900 416.850 ;
        RECT 910.950 415.950 915.450 417.450 ;
        RECT 763.500 412.950 765.600 415.050 ;
        RECT 766.800 412.950 768.900 415.050 ;
        RECT 781.950 412.950 784.050 415.050 ;
        RECT 784.950 412.950 787.050 415.050 ;
        RECT 787.950 412.950 790.050 415.050 ;
        RECT 802.950 412.950 805.050 415.050 ;
        RECT 805.950 412.950 808.050 415.050 ;
        RECT 808.950 412.950 811.050 415.050 ;
        RECT 811.950 412.950 814.050 415.050 ;
        RECT 826.950 412.950 829.050 415.050 ;
        RECT 829.950 412.950 832.050 415.050 ;
        RECT 847.950 412.950 850.050 415.050 ;
        RECT 850.950 412.950 853.050 415.050 ;
        RECT 853.950 412.950 856.050 415.050 ;
        RECT 856.950 412.950 859.050 415.050 ;
        RECT 871.950 412.950 874.050 415.050 ;
        RECT 874.950 412.950 877.050 415.050 ;
        RECT 877.950 412.950 880.050 415.050 ;
        RECT 880.950 412.950 883.050 415.050 ;
        RECT 898.950 412.950 901.050 415.050 ;
        RECT 901.950 412.950 904.050 415.050 ;
        RECT 904.950 412.950 907.050 415.050 ;
        RECT 907.950 412.950 910.050 415.050 ;
        RECT 763.200 411.150 765.000 412.950 ;
        RECT 767.400 405.600 768.300 412.950 ;
        RECT 740.100 393.600 741.900 399.600 ;
        RECT 743.100 393.000 744.900 399.600 ;
        RECT 758.100 393.000 759.900 399.600 ;
        RECT 761.100 393.600 762.900 399.600 ;
        RECT 764.100 393.000 765.900 405.000 ;
        RECT 767.100 393.600 768.900 405.600 ;
        RECT 785.100 399.600 786.300 412.950 ;
        RECT 806.100 405.600 807.300 412.950 ;
        RECT 812.100 411.150 813.900 412.950 ;
        RECT 827.100 411.150 828.900 412.950 ;
        RECT 806.100 404.100 808.500 405.600 ;
        RECT 804.000 401.100 805.800 402.900 ;
        RECT 782.100 393.000 783.900 399.600 ;
        RECT 785.100 393.600 786.900 399.600 ;
        RECT 788.100 393.000 789.900 399.600 ;
        RECT 803.700 393.000 805.500 399.600 ;
        RECT 806.700 393.600 808.500 404.100 ;
        RECT 811.800 393.000 813.600 405.600 ;
        RECT 830.100 399.600 831.300 412.950 ;
        RECT 849.000 400.800 849.900 412.950 ;
        RECT 854.100 411.150 855.900 412.950 ;
        RECT 875.250 411.150 877.050 412.950 ;
        RECT 850.950 408.450 853.050 409.050 ;
        RECT 871.950 408.450 874.050 409.050 ;
        RECT 850.950 407.550 874.050 408.450 ;
        RECT 850.950 406.950 853.050 407.550 ;
        RECT 871.950 406.950 874.050 407.550 ;
        RECT 881.700 405.600 882.600 412.950 ;
        RECT 899.100 411.150 900.900 412.950 ;
        RECT 905.700 405.600 906.900 412.950 ;
        RECT 914.550 412.050 915.450 415.950 ;
        RECT 910.950 410.550 915.450 412.050 ;
        RECT 917.550 415.950 922.050 417.450 ;
        RECT 917.550 412.050 918.450 415.950 ;
        RECT 926.100 415.050 927.900 416.850 ;
        RECT 929.700 415.050 930.900 419.400 ;
        RECT 948.000 418.800 951.300 420.000 ;
        RECT 956.100 419.400 957.900 429.000 ;
        RECT 971.100 425.400 972.900 428.400 ;
        RECT 974.100 425.400 975.900 429.000 ;
        RECT 989.700 425.400 991.500 429.000 ;
        RECT 942.000 417.450 946.050 418.050 ;
        RECT 932.100 415.050 933.900 416.850 ;
        RECT 941.550 415.950 946.050 417.450 ;
        RECT 922.950 412.950 925.050 415.050 ;
        RECT 925.950 412.950 928.050 415.050 ;
        RECT 928.950 412.950 931.050 415.050 ;
        RECT 931.950 412.950 934.050 415.050 ;
        RECT 917.550 410.550 922.050 412.050 ;
        RECT 923.100 411.150 924.900 412.950 ;
        RECT 910.950 409.950 915.000 410.550 ;
        RECT 918.000 409.950 922.050 410.550 ;
        RECT 929.700 405.600 930.900 412.950 ;
        RECT 941.550 412.050 942.450 415.950 ;
        RECT 948.000 415.050 948.900 418.800 ;
        RECT 967.950 417.450 970.050 418.050 ;
        RECT 950.100 415.050 951.900 416.850 ;
        RECT 956.100 415.050 957.900 416.850 ;
        RECT 962.550 416.550 970.050 417.450 ;
        RECT 946.950 412.950 949.050 415.050 ;
        RECT 949.950 412.950 952.050 415.050 ;
        RECT 952.950 412.950 955.050 415.050 ;
        RECT 955.950 412.950 958.050 415.050 ;
        RECT 941.550 410.550 946.050 412.050 ;
        RECT 942.000 409.950 946.050 410.550 ;
        RECT 931.950 408.450 934.050 409.050 ;
        RECT 937.950 408.450 940.050 409.050 ;
        RECT 931.950 407.550 940.050 408.450 ;
        RECT 931.950 406.950 934.050 407.550 ;
        RECT 937.950 406.950 940.050 407.550 ;
        RECT 872.100 404.700 879.900 405.600 ;
        RECT 849.000 399.900 855.600 400.800 ;
        RECT 849.000 399.600 849.900 399.900 ;
        RECT 827.100 393.000 828.900 399.600 ;
        RECT 830.100 393.600 831.900 399.600 ;
        RECT 848.100 393.600 849.900 399.600 ;
        RECT 854.100 399.600 855.600 399.900 ;
        RECT 851.100 393.000 852.900 399.000 ;
        RECT 854.100 393.600 855.900 399.600 ;
        RECT 857.100 393.000 858.900 399.600 ;
        RECT 872.100 393.600 873.900 404.700 ;
        RECT 875.100 393.000 876.900 403.800 ;
        RECT 878.100 393.600 879.900 404.700 ;
        RECT 881.100 393.600 882.900 405.600 ;
        RECT 899.400 393.000 901.200 405.600 ;
        RECT 904.500 404.100 906.900 405.600 ;
        RECT 904.500 393.600 906.300 404.100 ;
        RECT 907.200 401.100 909.000 402.900 ;
        RECT 907.500 393.000 909.300 399.600 ;
        RECT 923.400 393.000 925.200 405.600 ;
        RECT 928.500 404.100 930.900 405.600 ;
        RECT 928.500 393.600 930.300 404.100 ;
        RECT 931.200 401.100 933.000 402.900 ;
        RECT 948.000 400.800 948.900 412.950 ;
        RECT 953.100 411.150 954.900 412.950 ;
        RECT 962.550 411.450 963.450 416.550 ;
        RECT 967.950 415.950 970.050 416.550 ;
        RECT 971.700 415.050 972.900 425.400 ;
        RECT 992.700 423.600 994.500 428.400 ;
        RECT 989.400 422.400 994.500 423.600 ;
        RECT 997.200 422.400 999.000 429.000 ;
        RECT 989.400 415.050 990.300 422.400 ;
        RECT 991.950 420.450 994.050 421.050 ;
        RECT 1003.950 420.450 1006.050 421.050 ;
        RECT 991.950 419.550 1006.050 420.450 ;
        RECT 991.950 418.950 994.050 419.550 ;
        RECT 1003.950 418.950 1006.050 419.550 ;
        RECT 991.950 415.050 993.750 416.850 ;
        RECT 998.100 415.050 999.900 416.850 ;
        RECT 970.950 412.950 973.050 415.050 ;
        RECT 973.950 412.950 976.050 415.050 ;
        RECT 988.950 412.950 991.050 415.050 ;
        RECT 991.950 412.950 994.050 415.050 ;
        RECT 994.950 412.950 997.050 415.050 ;
        RECT 997.950 412.950 1000.050 415.050 ;
        RECT 959.550 410.550 963.450 411.450 ;
        RECT 959.550 409.050 960.450 410.550 ;
        RECT 955.950 407.550 960.450 409.050 ;
        RECT 955.950 406.950 960.000 407.550 ;
        RECT 955.950 405.450 958.050 405.900 ;
        RECT 964.950 405.450 967.050 406.050 ;
        RECT 955.950 404.550 967.050 405.450 ;
        RECT 955.950 403.800 958.050 404.550 ;
        RECT 964.950 403.950 967.050 404.550 ;
        RECT 948.000 399.900 954.600 400.800 ;
        RECT 948.000 399.600 948.900 399.900 ;
        RECT 931.500 393.000 933.300 399.600 ;
        RECT 947.100 393.600 948.900 399.600 ;
        RECT 953.100 399.600 954.600 399.900 ;
        RECT 971.700 399.600 972.900 412.950 ;
        RECT 974.100 411.150 975.900 412.950 ;
        RECT 989.400 405.600 990.300 412.950 ;
        RECT 994.950 411.150 996.750 412.950 ;
        RECT 950.100 393.000 951.900 399.000 ;
        RECT 953.100 393.600 954.900 399.600 ;
        RECT 956.100 393.000 957.900 399.600 ;
        RECT 971.100 393.600 972.900 399.600 ;
        RECT 974.100 393.000 975.900 399.600 ;
        RECT 989.100 393.600 990.900 405.600 ;
        RECT 992.100 404.700 999.900 405.600 ;
        RECT 992.100 393.600 993.900 404.700 ;
        RECT 995.100 393.000 996.900 403.800 ;
        RECT 998.100 393.600 999.900 404.700 ;
        RECT 17.100 383.400 18.900 390.000 ;
        RECT 20.100 383.400 21.900 389.400 ;
        RECT 17.100 370.050 18.900 371.850 ;
        RECT 20.100 370.050 21.300 383.400 ;
        RECT 35.400 377.400 37.200 390.000 ;
        RECT 40.500 378.900 42.300 389.400 ;
        RECT 43.500 383.400 45.300 390.000 ;
        RECT 59.100 383.400 60.900 390.000 ;
        RECT 62.100 383.400 63.900 389.400 ;
        RECT 65.100 383.400 66.900 390.000 ;
        RECT 43.200 380.100 45.000 381.900 ;
        RECT 40.500 377.400 42.900 378.900 ;
        RECT 35.100 370.050 36.900 371.850 ;
        RECT 41.700 370.050 42.900 377.400 ;
        RECT 62.700 370.050 63.900 383.400 ;
        RECT 69.150 379.200 70.950 389.400 ;
        RECT 68.550 377.400 70.950 379.200 ;
        RECT 72.150 377.400 73.950 390.000 ;
        RECT 77.550 380.400 79.350 389.400 ;
        RECT 82.350 383.400 84.150 390.000 ;
        RECT 85.350 382.500 87.150 389.400 ;
        RECT 88.350 383.400 90.150 390.000 ;
        RECT 92.850 383.400 94.650 389.400 ;
        RECT 81.450 381.450 88.050 382.500 ;
        RECT 81.450 380.700 83.250 381.450 ;
        RECT 86.250 380.700 88.050 381.450 ;
        RECT 92.550 381.300 94.650 383.400 ;
        RECT 77.250 379.500 79.350 380.400 ;
        RECT 89.850 379.800 91.650 380.400 ;
        RECT 77.250 378.300 85.050 379.500 ;
        RECT 83.250 377.700 85.050 378.300 ;
        RECT 85.950 378.900 91.650 379.800 ;
        RECT 68.550 376.500 69.450 377.400 ;
        RECT 85.950 376.800 86.850 378.900 ;
        RECT 89.850 378.600 91.650 378.900 ;
        RECT 92.550 378.600 95.550 380.400 ;
        RECT 92.550 377.700 93.750 378.600 ;
        RECT 78.450 376.500 86.850 376.800 ;
        RECT 68.550 375.900 86.850 376.500 ;
        RECT 88.950 376.800 93.750 377.700 ;
        RECT 97.650 377.400 99.450 390.000 ;
        RECT 100.650 377.400 102.450 389.400 ;
        RECT 116.100 377.400 117.900 389.400 ;
        RECT 119.100 378.300 120.900 389.400 ;
        RECT 122.100 379.200 123.900 390.000 ;
        RECT 125.100 378.300 126.900 389.400 ;
        RECT 119.100 377.400 126.900 378.300 ;
        RECT 140.100 377.400 141.900 390.000 ;
        RECT 145.200 378.600 147.000 389.400 ;
        RECT 143.400 377.400 147.000 378.600 ;
        RECT 161.100 377.400 162.900 390.000 ;
        RECT 68.550 375.300 80.250 375.900 ;
        RECT 16.950 367.950 19.050 370.050 ;
        RECT 19.950 367.950 22.050 370.050 ;
        RECT 34.950 367.950 37.050 370.050 ;
        RECT 37.950 367.950 40.050 370.050 ;
        RECT 40.950 367.950 43.050 370.050 ;
        RECT 43.950 367.950 46.050 370.050 ;
        RECT 58.950 367.950 61.050 370.050 ;
        RECT 61.950 367.950 64.050 370.050 ;
        RECT 64.950 367.950 67.050 370.050 ;
        RECT 20.100 357.600 21.300 367.950 ;
        RECT 38.100 366.150 39.900 367.950 ;
        RECT 41.700 363.600 42.900 367.950 ;
        RECT 44.100 366.150 45.900 367.950 ;
        RECT 59.100 366.150 60.900 367.950 ;
        RECT 41.700 362.700 45.300 363.600 ;
        RECT 62.700 362.700 63.900 367.950 ;
        RECT 64.950 366.150 66.750 367.950 ;
        RECT 35.100 359.700 42.900 361.050 ;
        RECT 17.100 354.000 18.900 357.600 ;
        RECT 20.100 354.600 21.900 357.600 ;
        RECT 35.100 354.600 36.900 359.700 ;
        RECT 38.100 354.000 39.900 358.800 ;
        RECT 41.100 354.600 42.900 359.700 ;
        RECT 44.100 360.600 45.300 362.700 ;
        RECT 59.700 361.800 63.900 362.700 ;
        RECT 44.100 354.600 45.900 360.600 ;
        RECT 59.700 354.600 61.500 361.800 ;
        RECT 68.550 360.600 69.450 375.300 ;
        RECT 78.450 375.000 80.250 375.300 ;
        RECT 70.950 367.950 73.050 370.050 ;
        RECT 80.100 368.400 82.200 370.050 ;
        RECT 70.950 365.400 72.750 367.950 ;
        RECT 74.100 367.200 82.200 368.400 ;
        RECT 74.100 366.600 75.900 367.200 ;
        RECT 77.100 365.400 78.900 366.000 ;
        RECT 70.950 364.200 78.900 365.400 ;
        RECT 88.950 364.200 89.850 376.800 ;
        RECT 92.550 374.100 94.650 374.700 ;
        RECT 98.550 374.100 100.350 374.550 ;
        RECT 92.550 372.900 100.350 374.100 ;
        RECT 92.550 372.600 94.650 372.900 ;
        RECT 98.550 372.750 100.350 372.900 ;
        RECT 101.250 370.050 102.450 377.400 ;
        RECT 116.400 370.050 117.300 377.400 ;
        RECT 118.950 375.450 121.050 376.050 ;
        RECT 139.950 375.450 142.050 376.050 ;
        RECT 118.950 374.550 142.050 375.450 ;
        RECT 118.950 373.950 121.050 374.550 ;
        RECT 139.950 373.950 142.050 374.550 ;
        RECT 130.950 372.450 133.050 373.050 ;
        RECT 136.950 372.450 139.050 373.050 ;
        RECT 121.950 370.050 123.750 371.850 ;
        RECT 130.950 371.550 139.050 372.450 ;
        RECT 130.950 370.950 133.050 371.550 ;
        RECT 136.950 370.950 139.050 371.550 ;
        RECT 140.250 370.050 142.050 371.850 ;
        RECT 143.400 370.050 144.300 377.400 ;
        RECT 164.100 376.500 165.900 389.400 ;
        RECT 167.100 377.400 168.900 390.000 ;
        RECT 170.100 376.500 171.900 389.400 ;
        RECT 173.100 377.400 174.900 390.000 ;
        RECT 176.100 376.500 177.900 389.400 ;
        RECT 179.100 377.400 180.900 390.000 ;
        RECT 182.100 376.500 183.900 389.400 ;
        RECT 185.100 377.400 186.900 390.000 ;
        RECT 189.150 379.200 190.950 389.400 ;
        RECT 188.550 377.400 190.950 379.200 ;
        RECT 192.150 377.400 193.950 390.000 ;
        RECT 197.550 380.400 199.350 389.400 ;
        RECT 202.350 383.400 204.150 390.000 ;
        RECT 205.350 382.500 207.150 389.400 ;
        RECT 208.350 383.400 210.150 390.000 ;
        RECT 212.850 383.400 214.650 389.400 ;
        RECT 201.450 381.450 208.050 382.500 ;
        RECT 201.450 380.700 203.250 381.450 ;
        RECT 206.250 380.700 208.050 381.450 ;
        RECT 212.550 381.300 214.650 383.400 ;
        RECT 197.250 379.500 199.350 380.400 ;
        RECT 209.850 379.800 211.650 380.400 ;
        RECT 197.250 378.300 205.050 379.500 ;
        RECT 203.250 377.700 205.050 378.300 ;
        RECT 205.950 378.900 211.650 379.800 ;
        RECT 188.550 376.500 189.450 377.400 ;
        RECT 205.950 376.800 206.850 378.900 ;
        RECT 209.850 378.600 211.650 378.900 ;
        RECT 212.550 378.600 215.550 380.400 ;
        RECT 212.550 377.700 213.750 378.600 ;
        RECT 198.450 376.500 206.850 376.800 ;
        RECT 164.100 375.300 168.000 376.500 ;
        RECT 170.100 375.300 174.000 376.500 ;
        RECT 176.100 375.300 180.000 376.500 ;
        RECT 182.100 375.300 184.950 376.500 ;
        RECT 146.100 370.050 147.900 371.850 ;
        RECT 97.950 369.750 102.450 370.050 ;
        RECT 96.150 367.950 102.450 369.750 ;
        RECT 115.950 367.950 118.050 370.050 ;
        RECT 118.950 367.950 121.050 370.050 ;
        RECT 121.950 367.950 124.050 370.050 ;
        RECT 124.950 367.950 127.050 370.050 ;
        RECT 139.950 367.950 142.050 370.050 ;
        RECT 142.950 367.950 145.050 370.050 ;
        RECT 145.950 367.950 148.050 370.050 ;
        RECT 163.800 367.950 165.900 370.050 ;
        RECT 77.850 363.000 89.850 364.200 ;
        RECT 77.850 361.200 78.900 363.000 ;
        RECT 88.050 362.400 89.850 363.000 ;
        RECT 64.800 354.000 66.600 360.600 ;
        RECT 68.550 358.800 70.950 360.600 ;
        RECT 69.150 354.600 70.950 358.800 ;
        RECT 72.150 354.000 73.950 360.600 ;
        RECT 74.850 358.200 76.950 359.700 ;
        RECT 77.850 359.400 79.650 361.200 ;
        RECT 101.250 360.600 102.450 367.950 ;
        RECT 80.850 359.550 82.650 360.300 ;
        RECT 80.850 358.500 85.800 359.550 ;
        RECT 74.850 357.600 78.750 358.200 ;
        RECT 84.750 357.600 85.800 358.500 ;
        RECT 92.250 357.600 94.650 359.700 ;
        RECT 75.150 356.700 78.750 357.600 ;
        RECT 76.950 354.600 78.750 356.700 ;
        RECT 81.450 354.000 83.250 357.600 ;
        RECT 84.750 354.600 86.550 357.600 ;
        RECT 87.750 354.000 89.550 357.600 ;
        RECT 92.250 354.600 94.050 357.600 ;
        RECT 97.350 354.000 99.150 360.600 ;
        RECT 100.650 354.600 102.450 360.600 ;
        RECT 116.400 360.600 117.300 367.950 ;
        RECT 118.950 366.150 120.750 367.950 ;
        RECT 125.100 366.150 126.900 367.950 ;
        RECT 121.950 363.450 124.050 364.050 ;
        RECT 130.950 363.450 133.050 364.050 ;
        RECT 121.950 362.550 133.050 363.450 ;
        RECT 121.950 361.950 124.050 362.550 ;
        RECT 130.950 361.950 133.050 362.550 ;
        RECT 116.400 359.400 121.500 360.600 ;
        RECT 116.700 354.000 118.500 357.600 ;
        RECT 119.700 354.600 121.500 359.400 ;
        RECT 124.200 354.000 126.000 360.600 ;
        RECT 143.400 357.600 144.300 367.950 ;
        RECT 163.800 366.150 165.600 367.950 ;
        RECT 166.800 364.800 168.000 375.300 ;
        RECT 169.200 364.800 171.000 365.400 ;
        RECT 166.800 363.600 171.000 364.800 ;
        RECT 172.800 364.800 174.000 375.300 ;
        RECT 175.200 364.800 177.000 365.400 ;
        RECT 172.800 363.600 177.000 364.800 ;
        RECT 178.800 364.800 180.000 375.300 ;
        RECT 183.900 370.050 184.950 375.300 ;
        RECT 181.800 367.950 184.950 370.050 ;
        RECT 181.200 364.800 183.000 365.400 ;
        RECT 178.800 363.600 183.000 364.800 ;
        RECT 166.800 362.700 168.000 363.600 ;
        RECT 172.800 362.700 174.000 363.600 ;
        RECT 178.800 362.700 180.000 363.600 ;
        RECT 183.900 362.700 184.950 367.950 ;
        RECT 164.100 361.500 168.000 362.700 ;
        RECT 170.100 361.500 174.000 362.700 ;
        RECT 176.100 361.500 180.000 362.700 ;
        RECT 182.100 361.500 184.950 362.700 ;
        RECT 188.550 375.900 206.850 376.500 ;
        RECT 208.950 376.800 213.750 377.700 ;
        RECT 217.650 377.400 219.450 390.000 ;
        RECT 220.650 377.400 222.450 389.400 ;
        RECT 239.100 383.400 240.900 390.000 ;
        RECT 242.100 383.400 243.900 389.400 ;
        RECT 245.100 383.400 246.900 390.000 ;
        RECT 188.550 375.300 200.250 375.900 ;
        RECT 140.100 354.000 141.900 357.600 ;
        RECT 143.100 354.600 144.900 357.600 ;
        RECT 146.100 354.000 147.900 357.600 ;
        RECT 161.100 354.000 162.900 360.600 ;
        RECT 164.100 354.600 165.900 361.500 ;
        RECT 167.100 354.000 168.900 360.600 ;
        RECT 170.100 354.600 171.900 361.500 ;
        RECT 173.100 354.000 174.900 360.600 ;
        RECT 176.100 354.600 177.900 361.500 ;
        RECT 179.100 354.000 180.900 360.600 ;
        RECT 182.100 354.600 183.900 361.500 ;
        RECT 188.550 360.600 189.450 375.300 ;
        RECT 198.450 375.000 200.250 375.300 ;
        RECT 190.950 367.950 193.050 370.050 ;
        RECT 200.100 368.400 202.200 370.050 ;
        RECT 190.950 365.400 192.750 367.950 ;
        RECT 194.100 367.200 202.200 368.400 ;
        RECT 194.100 366.600 195.900 367.200 ;
        RECT 197.100 365.400 198.900 366.000 ;
        RECT 190.950 364.200 198.900 365.400 ;
        RECT 208.950 364.200 209.850 376.800 ;
        RECT 212.550 374.100 214.650 374.700 ;
        RECT 218.550 374.100 220.350 374.550 ;
        RECT 212.550 372.900 220.350 374.100 ;
        RECT 212.550 372.600 214.650 372.900 ;
        RECT 218.550 372.750 220.350 372.900 ;
        RECT 221.250 370.050 222.450 377.400 ;
        RECT 242.700 370.050 243.900 383.400 ;
        RECT 263.100 377.400 264.900 390.000 ;
        RECT 266.100 376.500 267.900 389.400 ;
        RECT 269.100 377.400 270.900 390.000 ;
        RECT 272.100 376.500 273.900 389.400 ;
        RECT 275.100 377.400 276.900 390.000 ;
        RECT 278.100 376.500 279.900 389.400 ;
        RECT 281.100 377.400 282.900 390.000 ;
        RECT 284.100 376.500 285.900 389.400 ;
        RECT 287.100 377.400 288.900 390.000 ;
        RECT 291.150 379.200 292.950 389.400 ;
        RECT 290.550 377.400 292.950 379.200 ;
        RECT 294.150 377.400 295.950 390.000 ;
        RECT 299.550 380.400 301.350 389.400 ;
        RECT 304.350 383.400 306.150 390.000 ;
        RECT 307.350 382.500 309.150 389.400 ;
        RECT 310.350 383.400 312.150 390.000 ;
        RECT 314.850 383.400 316.650 389.400 ;
        RECT 303.450 381.450 310.050 382.500 ;
        RECT 303.450 380.700 305.250 381.450 ;
        RECT 308.250 380.700 310.050 381.450 ;
        RECT 314.550 381.300 316.650 383.400 ;
        RECT 299.250 379.500 301.350 380.400 ;
        RECT 311.850 379.800 313.650 380.400 ;
        RECT 299.250 378.300 307.050 379.500 ;
        RECT 305.250 377.700 307.050 378.300 ;
        RECT 307.950 378.900 313.650 379.800 ;
        RECT 290.550 376.500 291.450 377.400 ;
        RECT 307.950 376.800 308.850 378.900 ;
        RECT 311.850 378.600 313.650 378.900 ;
        RECT 314.550 378.600 317.550 380.400 ;
        RECT 314.550 377.700 315.750 378.600 ;
        RECT 300.450 376.500 308.850 376.800 ;
        RECT 266.100 375.300 270.000 376.500 ;
        RECT 272.100 375.300 276.000 376.500 ;
        RECT 278.100 375.300 282.000 376.500 ;
        RECT 284.100 375.300 286.950 376.500 ;
        RECT 217.950 369.750 222.450 370.050 ;
        RECT 216.150 367.950 222.450 369.750 ;
        RECT 238.950 367.950 241.050 370.050 ;
        RECT 241.950 367.950 244.050 370.050 ;
        RECT 244.950 367.950 247.050 370.050 ;
        RECT 265.800 367.950 267.900 370.050 ;
        RECT 197.850 363.000 209.850 364.200 ;
        RECT 197.850 361.200 198.900 363.000 ;
        RECT 208.050 362.400 209.850 363.000 ;
        RECT 185.100 354.000 186.900 360.600 ;
        RECT 188.550 358.800 190.950 360.600 ;
        RECT 189.150 354.600 190.950 358.800 ;
        RECT 192.150 354.000 193.950 360.600 ;
        RECT 194.850 358.200 196.950 359.700 ;
        RECT 197.850 359.400 199.650 361.200 ;
        RECT 221.250 360.600 222.450 367.950 ;
        RECT 239.100 366.150 240.900 367.950 ;
        RECT 242.700 362.700 243.900 367.950 ;
        RECT 244.950 366.150 246.750 367.950 ;
        RECT 265.800 366.150 267.600 367.950 ;
        RECT 268.800 364.800 270.000 375.300 ;
        RECT 271.200 364.800 273.000 365.400 ;
        RECT 268.800 363.600 273.000 364.800 ;
        RECT 274.800 364.800 276.000 375.300 ;
        RECT 277.200 364.800 279.000 365.400 ;
        RECT 274.800 363.600 279.000 364.800 ;
        RECT 280.800 364.800 282.000 375.300 ;
        RECT 285.900 370.050 286.950 375.300 ;
        RECT 283.800 367.950 286.950 370.050 ;
        RECT 283.200 364.800 285.000 365.400 ;
        RECT 280.800 363.600 285.000 364.800 ;
        RECT 268.800 362.700 270.000 363.600 ;
        RECT 274.800 362.700 276.000 363.600 ;
        RECT 280.800 362.700 282.000 363.600 ;
        RECT 285.900 362.700 286.950 367.950 ;
        RECT 200.850 359.550 202.650 360.300 ;
        RECT 200.850 358.500 205.800 359.550 ;
        RECT 194.850 357.600 198.750 358.200 ;
        RECT 204.750 357.600 205.800 358.500 ;
        RECT 212.250 357.600 214.650 359.700 ;
        RECT 195.150 356.700 198.750 357.600 ;
        RECT 196.950 354.600 198.750 356.700 ;
        RECT 201.450 354.000 203.250 357.600 ;
        RECT 204.750 354.600 206.550 357.600 ;
        RECT 207.750 354.000 209.550 357.600 ;
        RECT 212.250 354.600 214.050 357.600 ;
        RECT 217.350 354.000 219.150 360.600 ;
        RECT 220.650 354.600 222.450 360.600 ;
        RECT 239.700 361.800 243.900 362.700 ;
        RECT 239.700 354.600 241.500 361.800 ;
        RECT 266.100 361.500 270.000 362.700 ;
        RECT 272.100 361.500 276.000 362.700 ;
        RECT 278.100 361.500 282.000 362.700 ;
        RECT 284.100 361.500 286.950 362.700 ;
        RECT 290.550 375.900 308.850 376.500 ;
        RECT 310.950 376.800 315.750 377.700 ;
        RECT 319.650 377.400 321.450 390.000 ;
        RECT 322.650 377.400 324.450 389.400 ;
        RECT 341.100 383.400 342.900 390.000 ;
        RECT 344.100 383.400 345.900 389.400 ;
        RECT 347.100 383.400 348.900 390.000 ;
        RECT 362.700 383.400 364.500 390.000 ;
        RECT 290.550 375.300 302.250 375.900 ;
        RECT 244.800 354.000 246.600 360.600 ;
        RECT 263.100 354.000 264.900 360.600 ;
        RECT 266.100 354.600 267.900 361.500 ;
        RECT 269.100 354.000 270.900 360.600 ;
        RECT 272.100 354.600 273.900 361.500 ;
        RECT 275.100 354.000 276.900 360.600 ;
        RECT 278.100 354.600 279.900 361.500 ;
        RECT 281.100 354.000 282.900 360.600 ;
        RECT 284.100 354.600 285.900 361.500 ;
        RECT 290.550 360.600 291.450 375.300 ;
        RECT 300.450 375.000 302.250 375.300 ;
        RECT 292.950 367.950 295.050 370.050 ;
        RECT 302.100 368.400 304.200 370.050 ;
        RECT 292.950 365.400 294.750 367.950 ;
        RECT 296.100 367.200 304.200 368.400 ;
        RECT 296.100 366.600 297.900 367.200 ;
        RECT 299.100 365.400 300.900 366.000 ;
        RECT 292.950 364.200 300.900 365.400 ;
        RECT 310.950 364.200 311.850 376.800 ;
        RECT 314.550 374.100 316.650 374.700 ;
        RECT 320.550 374.100 322.350 374.550 ;
        RECT 314.550 372.900 322.350 374.100 ;
        RECT 314.550 372.600 316.650 372.900 ;
        RECT 320.550 372.750 322.350 372.900 ;
        RECT 323.250 370.050 324.450 377.400 ;
        RECT 344.100 370.050 345.300 383.400 ;
        RECT 363.000 380.100 364.800 381.900 ;
        RECT 365.700 378.900 367.500 389.400 ;
        RECT 365.100 377.400 367.500 378.900 ;
        RECT 370.800 377.400 372.600 390.000 ;
        RECT 386.100 383.400 387.900 390.000 ;
        RECT 389.100 383.400 390.900 389.400 ;
        RECT 392.100 383.400 393.900 390.000 ;
        RECT 407.700 383.400 409.500 390.000 ;
        RECT 361.950 375.450 364.050 376.050 ;
        RECT 353.550 374.550 364.050 375.450 ;
        RECT 319.950 369.750 324.450 370.050 ;
        RECT 318.150 367.950 324.450 369.750 ;
        RECT 340.950 367.950 343.050 370.050 ;
        RECT 343.950 367.950 346.050 370.050 ;
        RECT 346.950 367.950 349.050 370.050 ;
        RECT 299.850 363.000 311.850 364.200 ;
        RECT 299.850 361.200 300.900 363.000 ;
        RECT 310.050 362.400 311.850 363.000 ;
        RECT 287.100 354.000 288.900 360.600 ;
        RECT 290.550 358.800 292.950 360.600 ;
        RECT 291.150 354.600 292.950 358.800 ;
        RECT 294.150 354.000 295.950 360.600 ;
        RECT 296.850 358.200 298.950 359.700 ;
        RECT 299.850 359.400 301.650 361.200 ;
        RECT 323.250 360.600 324.450 367.950 ;
        RECT 341.250 366.150 343.050 367.950 ;
        RECT 344.100 362.700 345.300 367.950 ;
        RECT 347.100 366.150 348.900 367.950 ;
        RECT 353.550 367.050 354.450 374.550 ;
        RECT 361.950 373.950 364.050 374.550 ;
        RECT 357.000 372.450 361.050 373.050 ;
        RECT 349.950 365.550 354.450 367.050 ;
        RECT 356.550 370.950 361.050 372.450 ;
        RECT 356.550 367.050 357.450 370.950 ;
        RECT 365.100 370.050 366.300 377.400 ;
        RECT 371.100 370.050 372.900 371.850 ;
        RECT 389.100 370.050 390.300 383.400 ;
        RECT 408.000 380.100 409.800 381.900 ;
        RECT 410.700 378.900 412.500 389.400 ;
        RECT 410.100 377.400 412.500 378.900 ;
        RECT 415.800 377.400 417.600 390.000 ;
        RECT 431.700 383.400 433.500 390.000 ;
        RECT 432.000 380.100 433.800 381.900 ;
        RECT 434.700 378.900 436.500 389.400 ;
        RECT 434.100 377.400 436.500 378.900 ;
        RECT 439.800 377.400 441.600 390.000 ;
        RECT 455.100 383.400 456.900 389.400 ;
        RECT 458.100 383.400 459.900 390.000 ;
        RECT 410.100 370.050 411.300 377.400 ;
        RECT 416.100 370.050 417.900 371.850 ;
        RECT 434.100 370.050 435.300 377.400 ;
        RECT 436.950 375.450 439.050 376.050 ;
        RECT 451.950 375.450 454.050 376.050 ;
        RECT 436.950 374.550 454.050 375.450 ;
        RECT 436.950 373.950 439.050 374.550 ;
        RECT 451.950 373.950 454.050 374.550 ;
        RECT 440.100 370.050 441.900 371.850 ;
        RECT 455.700 370.050 456.900 383.400 ;
        RECT 461.550 377.400 463.350 389.400 ;
        RECT 464.550 377.400 466.350 390.000 ;
        RECT 469.350 383.400 471.150 389.400 ;
        RECT 473.850 383.400 475.650 390.000 ;
        RECT 469.350 381.300 471.450 383.400 ;
        RECT 476.850 382.500 478.650 389.400 ;
        RECT 479.850 383.400 481.650 390.000 ;
        RECT 475.950 381.450 482.550 382.500 ;
        RECT 475.950 380.700 477.750 381.450 ;
        RECT 480.750 380.700 482.550 381.450 ;
        RECT 484.650 380.400 486.450 389.400 ;
        RECT 468.450 378.600 471.450 380.400 ;
        RECT 472.350 379.800 474.150 380.400 ;
        RECT 472.350 378.900 478.050 379.800 ;
        RECT 484.650 379.500 486.750 380.400 ;
        RECT 472.350 378.600 474.150 378.900 ;
        RECT 470.250 377.700 471.450 378.600 ;
        RECT 458.100 370.050 459.900 371.850 ;
        RECT 461.550 370.050 462.750 377.400 ;
        RECT 470.250 376.800 475.050 377.700 ;
        RECT 463.650 374.100 465.450 374.550 ;
        RECT 469.350 374.100 471.450 374.700 ;
        RECT 463.650 372.900 471.450 374.100 ;
        RECT 463.650 372.750 465.450 372.900 ;
        RECT 469.350 372.600 471.450 372.900 ;
        RECT 361.950 367.950 364.050 370.050 ;
        RECT 364.950 367.950 367.050 370.050 ;
        RECT 367.950 367.950 370.050 370.050 ;
        RECT 370.950 367.950 373.050 370.050 ;
        RECT 385.950 367.950 388.050 370.050 ;
        RECT 388.950 367.950 391.050 370.050 ;
        RECT 391.950 367.950 394.050 370.050 ;
        RECT 406.950 367.950 409.050 370.050 ;
        RECT 409.950 367.950 412.050 370.050 ;
        RECT 412.950 367.950 415.050 370.050 ;
        RECT 415.950 367.950 418.050 370.050 ;
        RECT 430.950 367.950 433.050 370.050 ;
        RECT 433.950 367.950 436.050 370.050 ;
        RECT 436.950 367.950 439.050 370.050 ;
        RECT 439.950 367.950 442.050 370.050 ;
        RECT 454.950 367.950 457.050 370.050 ;
        RECT 457.950 367.950 460.050 370.050 ;
        RECT 461.550 369.750 466.050 370.050 ;
        RECT 461.550 367.950 467.850 369.750 ;
        RECT 356.550 365.550 361.050 367.050 ;
        RECT 362.100 366.150 363.900 367.950 ;
        RECT 349.950 364.950 354.000 365.550 ;
        RECT 357.000 364.950 361.050 365.550 ;
        RECT 365.100 363.600 366.300 367.950 ;
        RECT 368.100 366.150 369.900 367.950 ;
        RECT 386.250 366.150 388.050 367.950 ;
        RECT 362.700 362.700 366.300 363.600 ;
        RECT 389.100 362.700 390.300 367.950 ;
        RECT 392.100 366.150 393.900 367.950 ;
        RECT 407.100 366.150 408.900 367.950 ;
        RECT 410.100 363.600 411.300 367.950 ;
        RECT 413.100 366.150 414.900 367.950 ;
        RECT 431.100 366.150 432.900 367.950 ;
        RECT 434.100 363.600 435.300 367.950 ;
        RECT 437.100 366.150 438.900 367.950 ;
        RECT 407.700 362.700 411.300 363.600 ;
        RECT 431.700 362.700 435.300 363.600 ;
        RECT 344.100 361.800 348.300 362.700 ;
        RECT 302.850 359.550 304.650 360.300 ;
        RECT 302.850 358.500 307.800 359.550 ;
        RECT 296.850 357.600 300.750 358.200 ;
        RECT 306.750 357.600 307.800 358.500 ;
        RECT 314.250 357.600 316.650 359.700 ;
        RECT 297.150 356.700 300.750 357.600 ;
        RECT 298.950 354.600 300.750 356.700 ;
        RECT 303.450 354.000 305.250 357.600 ;
        RECT 306.750 354.600 308.550 357.600 ;
        RECT 309.750 354.000 311.550 357.600 ;
        RECT 314.250 354.600 316.050 357.600 ;
        RECT 319.350 354.000 321.150 360.600 ;
        RECT 322.650 354.600 324.450 360.600 ;
        RECT 341.400 354.000 343.200 360.600 ;
        RECT 346.500 354.600 348.300 361.800 ;
        RECT 362.700 360.600 363.900 362.700 ;
        RECT 389.100 361.800 393.300 362.700 ;
        RECT 362.100 354.600 363.900 360.600 ;
        RECT 365.100 359.700 372.900 361.050 ;
        RECT 365.100 354.600 366.900 359.700 ;
        RECT 368.100 354.000 369.900 358.800 ;
        RECT 371.100 354.600 372.900 359.700 ;
        RECT 386.400 354.000 388.200 360.600 ;
        RECT 391.500 354.600 393.300 361.800 ;
        RECT 407.700 360.600 408.900 362.700 ;
        RECT 407.100 354.600 408.900 360.600 ;
        RECT 410.100 359.700 417.900 361.050 ;
        RECT 431.700 360.600 432.900 362.700 ;
        RECT 410.100 354.600 411.900 359.700 ;
        RECT 413.100 354.000 414.900 358.800 ;
        RECT 416.100 354.600 417.900 359.700 ;
        RECT 431.100 354.600 432.900 360.600 ;
        RECT 434.100 359.700 441.900 361.050 ;
        RECT 434.100 354.600 435.900 359.700 ;
        RECT 437.100 354.000 438.900 358.800 ;
        RECT 440.100 354.600 441.900 359.700 ;
        RECT 455.700 357.600 456.900 367.950 ;
        RECT 461.550 360.600 462.750 367.950 ;
        RECT 474.150 364.200 475.050 376.800 ;
        RECT 477.150 376.800 478.050 378.900 ;
        RECT 478.950 378.300 486.750 379.500 ;
        RECT 478.950 377.700 480.750 378.300 ;
        RECT 490.050 377.400 491.850 390.000 ;
        RECT 493.050 379.200 494.850 389.400 ;
        RECT 498.150 379.200 499.950 389.400 ;
        RECT 493.050 377.400 495.450 379.200 ;
        RECT 477.150 376.500 485.550 376.800 ;
        RECT 494.550 376.500 495.450 377.400 ;
        RECT 477.150 375.900 495.450 376.500 ;
        RECT 483.750 375.300 495.450 375.900 ;
        RECT 483.750 375.000 485.550 375.300 ;
        RECT 481.800 368.400 483.900 370.050 ;
        RECT 481.800 367.200 489.900 368.400 ;
        RECT 490.950 367.950 493.050 370.050 ;
        RECT 488.100 366.600 489.900 367.200 ;
        RECT 485.100 365.400 486.900 366.000 ;
        RECT 491.250 365.400 493.050 367.950 ;
        RECT 485.100 364.200 493.050 365.400 ;
        RECT 474.150 363.000 486.150 364.200 ;
        RECT 474.150 362.400 475.950 363.000 ;
        RECT 485.100 361.200 486.150 363.000 ;
        RECT 455.100 354.600 456.900 357.600 ;
        RECT 458.100 354.000 459.900 357.600 ;
        RECT 461.550 354.600 463.350 360.600 ;
        RECT 464.850 354.000 466.650 360.600 ;
        RECT 469.350 357.600 471.750 359.700 ;
        RECT 481.350 359.550 483.150 360.300 ;
        RECT 478.200 358.500 483.150 359.550 ;
        RECT 484.350 359.400 486.150 361.200 ;
        RECT 494.550 360.600 495.450 375.300 ;
        RECT 478.200 357.600 479.250 358.500 ;
        RECT 487.050 358.200 489.150 359.700 ;
        RECT 485.250 357.600 489.150 358.200 ;
        RECT 469.950 354.600 471.750 357.600 ;
        RECT 474.450 354.000 476.250 357.600 ;
        RECT 477.450 354.600 479.250 357.600 ;
        RECT 480.750 354.000 482.550 357.600 ;
        RECT 485.250 356.700 488.850 357.600 ;
        RECT 485.250 354.600 487.050 356.700 ;
        RECT 490.050 354.000 491.850 360.600 ;
        RECT 493.050 358.800 495.450 360.600 ;
        RECT 497.550 377.400 499.950 379.200 ;
        RECT 501.150 377.400 502.950 390.000 ;
        RECT 506.550 380.400 508.350 389.400 ;
        RECT 511.350 383.400 513.150 390.000 ;
        RECT 514.350 382.500 516.150 389.400 ;
        RECT 517.350 383.400 519.150 390.000 ;
        RECT 521.850 383.400 523.650 389.400 ;
        RECT 510.450 381.450 517.050 382.500 ;
        RECT 510.450 380.700 512.250 381.450 ;
        RECT 515.250 380.700 517.050 381.450 ;
        RECT 521.550 381.300 523.650 383.400 ;
        RECT 506.250 379.500 508.350 380.400 ;
        RECT 518.850 379.800 520.650 380.400 ;
        RECT 506.250 378.300 514.050 379.500 ;
        RECT 512.250 377.700 514.050 378.300 ;
        RECT 514.950 378.900 520.650 379.800 ;
        RECT 497.550 376.500 498.450 377.400 ;
        RECT 514.950 376.800 515.850 378.900 ;
        RECT 518.850 378.600 520.650 378.900 ;
        RECT 521.550 378.600 524.550 380.400 ;
        RECT 521.550 377.700 522.750 378.600 ;
        RECT 507.450 376.500 515.850 376.800 ;
        RECT 497.550 375.900 515.850 376.500 ;
        RECT 517.950 376.800 522.750 377.700 ;
        RECT 526.650 377.400 528.450 390.000 ;
        RECT 529.650 377.400 531.450 389.400 ;
        RECT 497.550 375.300 509.250 375.900 ;
        RECT 497.550 360.600 498.450 375.300 ;
        RECT 507.450 375.000 509.250 375.300 ;
        RECT 499.950 367.950 502.050 370.050 ;
        RECT 509.100 368.400 511.200 370.050 ;
        RECT 499.950 365.400 501.750 367.950 ;
        RECT 503.100 367.200 511.200 368.400 ;
        RECT 503.100 366.600 504.900 367.200 ;
        RECT 506.100 365.400 507.900 366.000 ;
        RECT 499.950 364.200 507.900 365.400 ;
        RECT 517.950 364.200 518.850 376.800 ;
        RECT 521.550 374.100 523.650 374.700 ;
        RECT 527.550 374.100 529.350 374.550 ;
        RECT 521.550 372.900 529.350 374.100 ;
        RECT 521.550 372.600 523.650 372.900 ;
        RECT 527.550 372.750 529.350 372.900 ;
        RECT 530.250 370.050 531.450 377.400 ;
        RECT 545.100 383.400 546.900 389.400 ;
        RECT 545.100 376.500 546.300 383.400 ;
        RECT 548.100 379.200 549.900 390.000 ;
        RECT 551.100 377.400 552.900 389.400 ;
        RECT 569.100 383.400 570.900 390.000 ;
        RECT 572.100 383.400 573.900 389.400 ;
        RECT 545.100 375.600 550.800 376.500 ;
        RECT 549.000 374.700 550.800 375.600 ;
        RECT 526.950 369.750 531.450 370.050 ;
        RECT 525.150 367.950 531.450 369.750 ;
        RECT 545.400 370.050 547.200 371.850 ;
        RECT 545.400 367.950 547.500 370.050 ;
        RECT 506.850 363.000 518.850 364.200 ;
        RECT 506.850 361.200 507.900 363.000 ;
        RECT 517.050 362.400 518.850 363.000 ;
        RECT 497.550 358.800 499.950 360.600 ;
        RECT 493.050 354.600 494.850 358.800 ;
        RECT 498.150 354.600 499.950 358.800 ;
        RECT 501.150 354.000 502.950 360.600 ;
        RECT 503.850 358.200 505.950 359.700 ;
        RECT 506.850 359.400 508.650 361.200 ;
        RECT 530.250 360.600 531.450 367.950 ;
        RECT 549.000 363.300 549.900 374.700 ;
        RECT 551.700 370.050 552.900 377.400 ;
        RECT 569.100 370.050 570.900 371.850 ;
        RECT 572.100 370.050 573.300 383.400 ;
        RECT 587.100 377.400 588.900 390.000 ;
        RECT 590.100 377.400 591.900 389.400 ;
        RECT 593.100 377.400 594.900 390.000 ;
        RECT 608.100 383.400 609.900 389.400 ;
        RECT 611.100 383.400 612.900 390.000 ;
        RECT 626.100 383.400 627.900 390.000 ;
        RECT 629.100 383.400 630.900 389.400 ;
        RECT 632.100 384.000 633.900 390.000 ;
        RECT 590.400 370.050 591.450 377.400 ;
        RECT 608.700 370.050 609.900 383.400 ;
        RECT 629.400 383.100 630.900 383.400 ;
        RECT 635.100 383.400 636.900 389.400 ;
        RECT 635.100 383.100 636.000 383.400 ;
        RECT 629.400 382.200 636.000 383.100 ;
        RECT 611.100 370.050 612.900 371.850 ;
        RECT 629.100 370.050 630.900 371.850 ;
        RECT 635.100 370.050 636.000 382.200 ;
        RECT 653.100 378.300 654.900 389.400 ;
        RECT 656.100 379.200 657.900 390.000 ;
        RECT 659.100 378.300 660.900 389.400 ;
        RECT 653.100 377.400 660.900 378.300 ;
        RECT 662.100 377.400 663.900 389.400 ;
        RECT 677.100 383.400 678.900 390.000 ;
        RECT 680.100 383.400 681.900 389.400 ;
        RECT 683.100 384.000 684.900 390.000 ;
        RECT 680.400 383.100 681.900 383.400 ;
        RECT 686.100 383.400 687.900 389.400 ;
        RECT 686.100 383.100 687.000 383.400 ;
        RECT 680.400 382.200 687.000 383.100 ;
        RECT 656.250 370.050 658.050 371.850 ;
        RECT 662.700 370.050 663.600 377.400 ;
        RECT 680.100 370.050 681.900 371.850 ;
        RECT 686.100 370.050 687.000 382.200 ;
        RECT 701.100 377.400 702.900 390.000 ;
        RECT 706.200 378.600 708.000 389.400 ;
        RECT 704.400 377.400 708.000 378.600 ;
        RECT 725.400 377.400 727.200 390.000 ;
        RECT 730.500 378.900 732.300 389.400 ;
        RECT 733.500 383.400 735.300 390.000 ;
        RECT 733.200 380.100 735.000 381.900 ;
        RECT 730.500 377.400 732.900 378.900 ;
        RECT 749.400 377.400 751.200 390.000 ;
        RECT 754.500 378.900 756.300 389.400 ;
        RECT 757.500 383.400 759.300 390.000 ;
        RECT 776.100 383.400 777.900 390.000 ;
        RECT 779.100 383.400 780.900 389.400 ;
        RECT 782.100 383.400 783.900 390.000 ;
        RECT 797.100 383.400 798.900 390.000 ;
        RECT 800.100 383.400 801.900 389.400 ;
        RECT 803.100 384.000 804.900 390.000 ;
        RECT 757.200 380.100 759.000 381.900 ;
        RECT 754.500 377.400 756.900 378.900 ;
        RECT 701.250 370.050 703.050 371.850 ;
        RECT 704.400 370.050 705.300 377.400 ;
        RECT 707.100 370.050 708.900 371.850 ;
        RECT 725.100 370.050 726.900 371.850 ;
        RECT 731.700 370.050 732.900 377.400 ;
        RECT 749.100 370.050 750.900 371.850 ;
        RECT 755.700 370.050 756.900 377.400 ;
        RECT 779.700 370.050 780.900 383.400 ;
        RECT 800.400 383.100 801.900 383.400 ;
        RECT 806.100 383.400 807.900 389.400 ;
        RECT 806.100 383.100 807.000 383.400 ;
        RECT 800.400 382.200 807.000 383.100 ;
        RECT 800.100 370.050 801.900 371.850 ;
        RECT 806.100 370.050 807.000 382.200 ;
        RECT 821.100 378.300 822.900 389.400 ;
        RECT 824.100 379.200 825.900 390.000 ;
        RECT 827.100 378.300 828.900 389.400 ;
        RECT 821.100 377.400 828.900 378.300 ;
        RECT 830.100 377.400 831.900 389.400 ;
        RECT 845.100 383.400 846.900 390.000 ;
        RECT 848.100 383.400 849.900 389.400 ;
        RECT 851.100 384.000 852.900 390.000 ;
        RECT 848.400 383.100 849.900 383.400 ;
        RECT 854.100 383.400 855.900 389.400 ;
        RECT 869.100 383.400 870.900 390.000 ;
        RECT 872.100 383.400 873.900 389.400 ;
        RECT 875.100 384.000 876.900 390.000 ;
        RECT 854.100 383.100 855.000 383.400 ;
        RECT 848.400 382.200 855.000 383.100 ;
        RECT 872.400 383.100 873.900 383.400 ;
        RECT 878.100 383.400 879.900 389.400 ;
        RECT 893.700 383.400 895.500 390.000 ;
        RECT 878.100 383.100 879.000 383.400 ;
        RECT 872.400 382.200 879.000 383.100 ;
        RECT 838.950 378.450 841.050 379.050 ;
        RECT 844.950 378.450 847.050 379.050 ;
        RECT 838.950 377.550 847.050 378.450 ;
        RECT 824.250 370.050 826.050 371.850 ;
        RECT 830.700 370.050 831.600 377.400 ;
        RECT 838.950 376.950 841.050 377.550 ;
        RECT 844.950 376.950 847.050 377.550 ;
        RECT 848.100 370.050 849.900 371.850 ;
        RECT 854.100 370.050 855.000 382.200 ;
        RECT 859.950 375.450 862.050 376.050 ;
        RECT 871.950 375.450 874.050 379.050 ;
        RECT 859.950 375.000 874.050 375.450 ;
        RECT 859.950 374.550 873.450 375.000 ;
        RECT 859.950 373.950 862.050 374.550 ;
        RECT 872.100 370.050 873.900 371.850 ;
        RECT 878.100 370.050 879.000 382.200 ;
        RECT 894.000 380.100 895.800 381.900 ;
        RECT 896.700 378.900 898.500 389.400 ;
        RECT 896.100 377.400 898.500 378.900 ;
        RECT 901.800 377.400 903.600 390.000 ;
        RECT 917.400 377.400 919.200 390.000 ;
        RECT 922.500 378.900 924.300 389.400 ;
        RECT 925.500 383.400 927.300 390.000 ;
        RECT 944.100 383.400 945.900 390.000 ;
        RECT 947.100 383.400 948.900 389.400 ;
        RECT 950.100 384.000 951.900 390.000 ;
        RECT 947.400 383.100 948.900 383.400 ;
        RECT 953.100 383.400 954.900 389.400 ;
        RECT 968.100 383.400 969.900 389.400 ;
        RECT 971.100 384.000 972.900 390.000 ;
        RECT 953.100 383.100 954.000 383.400 ;
        RECT 947.400 382.200 954.000 383.100 ;
        RECT 925.200 380.100 927.000 381.900 ;
        RECT 922.500 377.400 924.900 378.900 ;
        RECT 888.000 372.450 892.050 373.050 ;
        RECT 887.550 370.950 892.050 372.450 ;
        RECT 550.800 367.950 552.900 370.050 ;
        RECT 568.950 367.950 571.050 370.050 ;
        RECT 571.950 367.950 574.050 370.050 ;
        RECT 587.400 367.950 589.500 370.050 ;
        RECT 590.400 367.950 594.600 370.050 ;
        RECT 607.950 367.950 610.050 370.050 ;
        RECT 610.950 367.950 613.050 370.050 ;
        RECT 625.950 367.950 628.050 370.050 ;
        RECT 628.950 367.950 631.050 370.050 ;
        RECT 631.950 367.950 634.050 370.050 ;
        RECT 634.950 367.950 637.050 370.050 ;
        RECT 652.950 367.950 655.050 370.050 ;
        RECT 655.950 367.950 658.050 370.050 ;
        RECT 658.950 367.950 661.050 370.050 ;
        RECT 661.950 367.950 664.050 370.050 ;
        RECT 676.950 367.950 679.050 370.050 ;
        RECT 679.950 367.950 682.050 370.050 ;
        RECT 682.950 367.950 685.050 370.050 ;
        RECT 685.950 367.950 688.050 370.050 ;
        RECT 700.950 367.950 703.050 370.050 ;
        RECT 703.950 367.950 706.050 370.050 ;
        RECT 706.950 367.950 709.050 370.050 ;
        RECT 724.950 367.950 727.050 370.050 ;
        RECT 727.950 367.950 730.050 370.050 ;
        RECT 730.950 367.950 733.050 370.050 ;
        RECT 733.950 367.950 736.050 370.050 ;
        RECT 748.950 367.950 751.050 370.050 ;
        RECT 751.950 367.950 754.050 370.050 ;
        RECT 754.950 367.950 757.050 370.050 ;
        RECT 757.950 367.950 760.050 370.050 ;
        RECT 775.950 367.950 778.050 370.050 ;
        RECT 778.950 367.950 781.050 370.050 ;
        RECT 781.950 367.950 784.050 370.050 ;
        RECT 796.950 367.950 799.050 370.050 ;
        RECT 799.950 367.950 802.050 370.050 ;
        RECT 802.950 367.950 805.050 370.050 ;
        RECT 805.950 367.950 808.050 370.050 ;
        RECT 820.950 367.950 823.050 370.050 ;
        RECT 823.950 367.950 826.050 370.050 ;
        RECT 826.950 367.950 829.050 370.050 ;
        RECT 829.950 367.950 832.050 370.050 ;
        RECT 844.950 367.950 847.050 370.050 ;
        RECT 847.950 367.950 850.050 370.050 ;
        RECT 850.950 367.950 853.050 370.050 ;
        RECT 853.950 367.950 856.050 370.050 ;
        RECT 868.950 367.950 871.050 370.050 ;
        RECT 871.950 367.950 874.050 370.050 ;
        RECT 874.950 367.950 877.050 370.050 ;
        RECT 877.950 367.950 880.050 370.050 ;
        RECT 549.000 362.400 550.800 363.300 ;
        RECT 509.850 359.550 511.650 360.300 ;
        RECT 509.850 358.500 514.800 359.550 ;
        RECT 503.850 357.600 507.750 358.200 ;
        RECT 513.750 357.600 514.800 358.500 ;
        RECT 521.250 357.600 523.650 359.700 ;
        RECT 504.150 356.700 507.750 357.600 ;
        RECT 505.950 354.600 507.750 356.700 ;
        RECT 510.450 354.000 512.250 357.600 ;
        RECT 513.750 354.600 515.550 357.600 ;
        RECT 516.750 354.000 518.550 357.600 ;
        RECT 521.250 354.600 523.050 357.600 ;
        RECT 526.350 354.000 528.150 360.600 ;
        RECT 529.650 354.600 531.450 360.600 ;
        RECT 545.100 361.500 550.800 362.400 ;
        RECT 545.100 357.600 546.300 361.500 ;
        RECT 551.700 360.600 552.900 367.950 ;
        RECT 545.100 354.600 546.900 357.600 ;
        RECT 548.100 354.000 549.900 360.600 ;
        RECT 551.100 354.600 552.900 360.600 ;
        RECT 572.100 357.600 573.300 367.950 ;
        RECT 587.400 366.150 589.200 367.950 ;
        RECT 590.400 360.600 591.450 367.950 ;
        RECT 569.100 354.000 570.900 357.600 ;
        RECT 572.100 354.600 573.900 357.600 ;
        RECT 587.100 354.000 588.900 360.600 ;
        RECT 590.100 354.600 591.900 360.600 ;
        RECT 593.100 354.000 594.900 360.600 ;
        RECT 608.700 357.600 609.900 367.950 ;
        RECT 626.100 366.150 627.900 367.950 ;
        RECT 632.100 366.150 633.900 367.950 ;
        RECT 635.100 364.200 636.000 367.950 ;
        RECT 653.100 366.150 654.900 367.950 ;
        RECT 659.250 366.150 661.050 367.950 ;
        RECT 608.100 354.600 609.900 357.600 ;
        RECT 611.100 354.000 612.900 357.600 ;
        RECT 626.100 354.000 627.900 363.600 ;
        RECT 632.700 363.000 636.000 364.200 ;
        RECT 632.700 354.600 634.500 363.000 ;
        RECT 662.700 360.600 663.600 367.950 ;
        RECT 677.100 366.150 678.900 367.950 ;
        RECT 683.100 366.150 684.900 367.950 ;
        RECT 686.100 364.200 687.000 367.950 ;
        RECT 654.000 354.000 655.800 360.600 ;
        RECT 658.500 359.400 663.600 360.600 ;
        RECT 658.500 354.600 660.300 359.400 ;
        RECT 661.500 354.000 663.300 357.600 ;
        RECT 677.100 354.000 678.900 363.600 ;
        RECT 683.700 363.000 687.000 364.200 ;
        RECT 683.700 354.600 685.500 363.000 ;
        RECT 704.400 357.600 705.300 367.950 ;
        RECT 728.100 366.150 729.900 367.950 ;
        RECT 731.700 363.600 732.900 367.950 ;
        RECT 734.100 366.150 735.900 367.950 ;
        RECT 752.100 366.150 753.900 367.950 ;
        RECT 755.700 363.600 756.900 367.950 ;
        RECT 758.100 366.150 759.900 367.950 ;
        RECT 776.100 366.150 777.900 367.950 ;
        RECT 731.700 362.700 735.300 363.600 ;
        RECT 755.700 362.700 759.300 363.600 ;
        RECT 779.700 362.700 780.900 367.950 ;
        RECT 781.950 366.150 783.750 367.950 ;
        RECT 787.950 366.450 790.050 367.050 ;
        RECT 793.950 366.450 796.050 367.050 ;
        RECT 787.950 365.550 796.050 366.450 ;
        RECT 797.100 366.150 798.900 367.950 ;
        RECT 803.100 366.150 804.900 367.950 ;
        RECT 787.950 364.950 790.050 365.550 ;
        RECT 793.950 364.950 796.050 365.550 ;
        RECT 806.100 364.200 807.000 367.950 ;
        RECT 821.100 366.150 822.900 367.950 ;
        RECT 827.250 366.150 829.050 367.950 ;
        RECT 725.100 359.700 732.900 361.050 ;
        RECT 701.100 354.000 702.900 357.600 ;
        RECT 704.100 354.600 705.900 357.600 ;
        RECT 707.100 354.000 708.900 357.600 ;
        RECT 725.100 354.600 726.900 359.700 ;
        RECT 728.100 354.000 729.900 358.800 ;
        RECT 731.100 354.600 732.900 359.700 ;
        RECT 734.100 360.600 735.300 362.700 ;
        RECT 734.100 354.600 735.900 360.600 ;
        RECT 749.100 359.700 756.900 361.050 ;
        RECT 749.100 354.600 750.900 359.700 ;
        RECT 752.100 354.000 753.900 358.800 ;
        RECT 755.100 354.600 756.900 359.700 ;
        RECT 758.100 360.600 759.300 362.700 ;
        RECT 776.700 361.800 780.900 362.700 ;
        RECT 758.100 354.600 759.900 360.600 ;
        RECT 776.700 354.600 778.500 361.800 ;
        RECT 781.800 354.000 783.600 360.600 ;
        RECT 797.100 354.000 798.900 363.600 ;
        RECT 803.700 363.000 807.000 364.200 ;
        RECT 803.700 354.600 805.500 363.000 ;
        RECT 830.700 360.600 831.600 367.950 ;
        RECT 845.100 366.150 846.900 367.950 ;
        RECT 851.100 366.150 852.900 367.950 ;
        RECT 854.100 364.200 855.000 367.950 ;
        RECT 869.100 366.150 870.900 367.950 ;
        RECT 875.100 366.150 876.900 367.950 ;
        RECT 878.100 364.200 879.000 367.950 ;
        RECT 880.950 366.450 883.050 367.050 ;
        RECT 887.550 366.450 888.450 370.950 ;
        RECT 896.100 370.050 897.300 377.400 ;
        RECT 898.950 375.450 901.050 376.050 ;
        RECT 919.950 375.450 922.050 376.050 ;
        RECT 898.950 374.550 922.050 375.450 ;
        RECT 898.950 373.950 901.050 374.550 ;
        RECT 919.950 373.950 922.050 374.550 ;
        RECT 912.000 372.450 916.050 373.050 ;
        RECT 902.100 370.050 903.900 371.850 ;
        RECT 911.550 370.950 916.050 372.450 ;
        RECT 892.950 367.950 895.050 370.050 ;
        RECT 895.950 367.950 898.050 370.050 ;
        RECT 898.950 367.950 901.050 370.050 ;
        RECT 901.950 367.950 904.050 370.050 ;
        RECT 880.950 365.550 888.450 366.450 ;
        RECT 893.100 366.150 894.900 367.950 ;
        RECT 880.950 364.950 883.050 365.550 ;
        RECT 822.000 354.000 823.800 360.600 ;
        RECT 826.500 359.400 831.600 360.600 ;
        RECT 826.500 354.600 828.300 359.400 ;
        RECT 829.500 354.000 831.300 357.600 ;
        RECT 845.100 354.000 846.900 363.600 ;
        RECT 851.700 363.000 855.000 364.200 ;
        RECT 851.700 354.600 853.500 363.000 ;
        RECT 869.100 354.000 870.900 363.600 ;
        RECT 875.700 363.000 879.000 364.200 ;
        RECT 896.100 363.600 897.300 367.950 ;
        RECT 899.100 366.150 900.900 367.950 ;
        RECT 911.550 367.050 912.450 370.950 ;
        RECT 917.100 370.050 918.900 371.850 ;
        RECT 923.700 370.050 924.900 377.400 ;
        RECT 947.100 370.050 948.900 371.850 ;
        RECT 953.100 370.050 954.000 382.200 ;
        RECT 969.000 383.100 969.900 383.400 ;
        RECT 974.100 383.400 975.900 389.400 ;
        RECT 977.100 383.400 978.900 390.000 ;
        RECT 992.100 383.400 993.900 390.000 ;
        RECT 995.100 383.400 996.900 389.400 ;
        RECT 998.100 383.400 999.900 390.000 ;
        RECT 974.100 383.100 975.600 383.400 ;
        RECT 969.000 382.200 975.600 383.100 ;
        RECT 969.000 370.050 969.900 382.200 ;
        RECT 976.950 375.450 979.050 376.050 ;
        RECT 985.950 375.450 988.050 376.050 ;
        RECT 976.950 374.550 988.050 375.450 ;
        RECT 976.950 373.950 979.050 374.550 ;
        RECT 985.950 373.950 988.050 374.550 ;
        RECT 987.000 372.450 991.050 373.050 ;
        RECT 974.100 370.050 975.900 371.850 ;
        RECT 986.550 370.950 991.050 372.450 ;
        RECT 916.950 367.950 919.050 370.050 ;
        RECT 919.950 367.950 922.050 370.050 ;
        RECT 922.950 367.950 925.050 370.050 ;
        RECT 925.950 367.950 928.050 370.050 ;
        RECT 943.950 367.950 946.050 370.050 ;
        RECT 946.950 367.950 949.050 370.050 ;
        RECT 949.950 367.950 952.050 370.050 ;
        RECT 952.950 367.950 955.050 370.050 ;
        RECT 967.950 367.950 970.050 370.050 ;
        RECT 970.950 367.950 973.050 370.050 ;
        RECT 973.950 367.950 976.050 370.050 ;
        RECT 976.950 367.950 979.050 370.050 ;
        RECT 911.550 365.550 916.050 367.050 ;
        RECT 920.100 366.150 921.900 367.950 ;
        RECT 912.000 364.950 916.050 365.550 ;
        RECT 875.700 354.600 877.500 363.000 ;
        RECT 893.700 362.700 897.300 363.600 ;
        RECT 923.700 363.600 924.900 367.950 ;
        RECT 926.100 366.150 927.900 367.950 ;
        RECT 944.100 366.150 945.900 367.950 ;
        RECT 950.100 366.150 951.900 367.950 ;
        RECT 953.100 364.200 954.000 367.950 ;
        RECT 923.700 362.700 927.300 363.600 ;
        RECT 893.700 360.600 894.900 362.700 ;
        RECT 893.100 354.600 894.900 360.600 ;
        RECT 896.100 359.700 903.900 361.050 ;
        RECT 896.100 354.600 897.900 359.700 ;
        RECT 899.100 354.000 900.900 358.800 ;
        RECT 902.100 354.600 903.900 359.700 ;
        RECT 917.100 359.700 924.900 361.050 ;
        RECT 917.100 354.600 918.900 359.700 ;
        RECT 920.100 354.000 921.900 358.800 ;
        RECT 923.100 354.600 924.900 359.700 ;
        RECT 926.100 360.600 927.300 362.700 ;
        RECT 926.100 354.600 927.900 360.600 ;
        RECT 931.950 360.450 934.050 360.900 ;
        RECT 937.950 360.450 940.050 361.050 ;
        RECT 931.950 359.550 940.050 360.450 ;
        RECT 931.950 358.800 934.050 359.550 ;
        RECT 937.950 358.950 940.050 359.550 ;
        RECT 944.100 354.000 945.900 363.600 ;
        RECT 950.700 363.000 954.000 364.200 ;
        RECT 969.000 364.200 969.900 367.950 ;
        RECT 971.100 366.150 972.900 367.950 ;
        RECT 977.100 366.150 978.900 367.950 ;
        RECT 986.550 367.050 987.450 370.950 ;
        RECT 995.700 370.050 996.900 383.400 ;
        RECT 991.950 367.950 994.050 370.050 ;
        RECT 994.950 367.950 997.050 370.050 ;
        RECT 997.950 367.950 1000.050 370.050 ;
        RECT 986.550 365.550 991.050 367.050 ;
        RECT 992.100 366.150 993.900 367.950 ;
        RECT 987.000 364.950 991.050 365.550 ;
        RECT 969.000 363.000 972.300 364.200 ;
        RECT 950.700 354.600 952.500 363.000 ;
        RECT 970.500 354.600 972.300 363.000 ;
        RECT 977.100 354.000 978.900 363.600 ;
        RECT 995.700 362.700 996.900 367.950 ;
        RECT 997.950 366.150 999.750 367.950 ;
        RECT 992.700 361.800 996.900 362.700 ;
        RECT 992.700 354.600 994.500 361.800 ;
        RECT 997.800 354.000 999.600 360.600 ;
        RECT 14.700 343.200 16.500 350.400 ;
        RECT 19.800 344.400 21.600 351.000 ;
        RECT 35.100 344.400 36.900 350.400 ;
        RECT 38.100 344.400 39.900 351.000 ;
        RECT 41.100 347.400 42.900 350.400 ;
        RECT 56.700 347.400 58.500 351.000 ;
        RECT 14.700 342.300 18.900 343.200 ;
        RECT 14.100 337.050 15.900 338.850 ;
        RECT 17.700 337.050 18.900 342.300 ;
        RECT 19.950 337.050 21.750 338.850 ;
        RECT 35.100 337.050 36.300 344.400 ;
        RECT 41.700 343.500 42.900 347.400 ;
        RECT 59.700 345.600 61.500 350.400 ;
        RECT 37.200 342.600 42.900 343.500 ;
        RECT 56.400 344.400 61.500 345.600 ;
        RECT 64.200 344.400 66.000 351.000 ;
        RECT 83.100 344.400 84.900 350.400 ;
        RECT 37.200 341.700 39.000 342.600 ;
        RECT 13.950 334.950 16.050 337.050 ;
        RECT 16.950 334.950 19.050 337.050 ;
        RECT 19.950 334.950 22.050 337.050 ;
        RECT 35.100 334.950 37.200 337.050 ;
        RECT 17.700 321.600 18.900 334.950 ;
        RECT 35.100 327.600 36.300 334.950 ;
        RECT 38.100 330.300 39.000 341.700 ;
        RECT 56.400 337.050 57.300 344.400 ;
        RECT 83.700 342.300 84.900 344.400 ;
        RECT 86.100 345.300 87.900 350.400 ;
        RECT 89.100 346.200 90.900 351.000 ;
        RECT 92.100 345.300 93.900 350.400 ;
        RECT 96.150 346.200 97.950 350.400 ;
        RECT 86.100 343.950 93.900 345.300 ;
        RECT 95.550 344.400 97.950 346.200 ;
        RECT 99.150 344.400 100.950 351.000 ;
        RECT 103.950 348.300 105.750 350.400 ;
        RECT 102.150 347.400 105.750 348.300 ;
        RECT 108.450 347.400 110.250 351.000 ;
        RECT 111.750 347.400 113.550 350.400 ;
        RECT 114.750 347.400 116.550 351.000 ;
        RECT 119.250 347.400 121.050 350.400 ;
        RECT 101.850 346.800 105.750 347.400 ;
        RECT 101.850 345.300 103.950 346.800 ;
        RECT 111.750 346.500 112.800 347.400 ;
        RECT 83.700 341.400 87.300 342.300 ;
        RECT 58.950 337.050 60.750 338.850 ;
        RECT 65.100 337.050 66.900 338.850 ;
        RECT 83.100 337.050 84.900 338.850 ;
        RECT 86.100 337.050 87.300 341.400 ;
        RECT 89.100 337.050 90.900 338.850 ;
        RECT 40.500 334.950 42.600 337.050 ;
        RECT 55.950 334.950 58.050 337.050 ;
        RECT 58.950 334.950 61.050 337.050 ;
        RECT 61.950 334.950 64.050 337.050 ;
        RECT 64.950 334.950 67.050 337.050 ;
        RECT 82.950 334.950 85.050 337.050 ;
        RECT 85.950 334.950 88.050 337.050 ;
        RECT 88.950 334.950 91.050 337.050 ;
        RECT 91.950 334.950 94.050 337.050 ;
        RECT 40.800 333.150 42.600 334.950 ;
        RECT 37.200 329.400 39.000 330.300 ;
        RECT 37.200 328.500 42.900 329.400 ;
        RECT 14.100 315.000 15.900 321.600 ;
        RECT 17.100 315.600 18.900 321.600 ;
        RECT 20.100 315.000 21.900 321.600 ;
        RECT 35.100 315.600 36.900 327.600 ;
        RECT 38.100 315.000 39.900 325.800 ;
        RECT 41.700 321.600 42.900 328.500 ;
        RECT 56.400 327.600 57.300 334.950 ;
        RECT 61.950 333.150 63.750 334.950 ;
        RECT 58.950 330.450 61.050 331.050 ;
        RECT 76.950 330.450 79.050 331.050 ;
        RECT 58.950 329.550 79.050 330.450 ;
        RECT 58.950 328.950 61.050 329.550 ;
        RECT 76.950 328.950 79.050 329.550 ;
        RECT 86.100 327.600 87.300 334.950 ;
        RECT 92.100 333.150 93.900 334.950 ;
        RECT 95.550 329.700 96.450 344.400 ;
        RECT 104.850 343.800 106.650 345.600 ;
        RECT 107.850 345.450 112.800 346.500 ;
        RECT 107.850 344.700 109.650 345.450 ;
        RECT 119.250 345.300 121.650 347.400 ;
        RECT 124.350 344.400 126.150 351.000 ;
        RECT 127.650 344.400 129.450 350.400 ;
        RECT 143.100 347.400 144.900 351.000 ;
        RECT 146.100 347.400 147.900 350.400 ;
        RECT 104.850 342.000 105.900 343.800 ;
        RECT 115.050 342.000 116.850 342.600 ;
        RECT 104.850 340.800 116.850 342.000 ;
        RECT 97.950 339.600 105.900 340.800 ;
        RECT 97.950 337.050 99.750 339.600 ;
        RECT 104.100 339.000 105.900 339.600 ;
        RECT 101.100 337.800 102.900 338.400 ;
        RECT 97.950 334.950 100.050 337.050 ;
        RECT 101.100 336.600 109.200 337.800 ;
        RECT 107.100 334.950 109.200 336.600 ;
        RECT 105.450 329.700 107.250 330.000 ;
        RECT 95.550 329.100 107.250 329.700 ;
        RECT 95.550 328.500 113.850 329.100 ;
        RECT 95.550 327.600 96.450 328.500 ;
        RECT 105.450 328.200 113.850 328.500 ;
        RECT 41.100 315.600 42.900 321.600 ;
        RECT 56.100 315.600 57.900 327.600 ;
        RECT 59.100 326.700 66.900 327.600 ;
        RECT 59.100 315.600 60.900 326.700 ;
        RECT 62.100 315.000 63.900 325.800 ;
        RECT 65.100 315.600 66.900 326.700 ;
        RECT 86.100 326.100 88.500 327.600 ;
        RECT 84.000 323.100 85.800 324.900 ;
        RECT 83.700 315.000 85.500 321.600 ;
        RECT 86.700 315.600 88.500 326.100 ;
        RECT 91.800 315.000 93.600 327.600 ;
        RECT 95.550 325.800 97.950 327.600 ;
        RECT 96.150 315.600 97.950 325.800 ;
        RECT 99.150 315.000 100.950 327.600 ;
        RECT 110.250 326.700 112.050 327.300 ;
        RECT 104.250 325.500 112.050 326.700 ;
        RECT 112.950 326.100 113.850 328.200 ;
        RECT 115.950 328.200 116.850 340.800 ;
        RECT 128.250 337.050 129.450 344.400 ;
        RECT 146.100 337.050 147.300 347.400 ;
        RECT 161.100 341.400 162.900 351.000 ;
        RECT 167.700 342.000 169.500 350.400 ;
        RECT 185.700 343.200 187.500 350.400 ;
        RECT 190.800 344.400 192.600 351.000 ;
        RECT 206.100 344.400 207.900 350.400 ;
        RECT 185.700 342.300 189.900 343.200 ;
        RECT 167.700 340.800 171.000 342.000 ;
        RECT 161.100 337.050 162.900 338.850 ;
        RECT 167.100 337.050 168.900 338.850 ;
        RECT 170.100 337.050 171.000 340.800 ;
        RECT 185.100 337.050 186.900 338.850 ;
        RECT 188.700 337.050 189.900 342.300 ;
        RECT 206.700 342.300 207.900 344.400 ;
        RECT 209.100 345.300 210.900 350.400 ;
        RECT 212.100 346.200 213.900 351.000 ;
        RECT 215.100 345.300 216.900 350.400 ;
        RECT 209.100 343.950 216.900 345.300 ;
        RECT 230.100 344.400 231.900 350.400 ;
        RECT 233.100 345.000 234.900 351.000 ;
        RECT 239.700 350.400 240.900 351.000 ;
        RECT 236.100 347.400 237.900 350.400 ;
        RECT 239.100 347.400 240.900 350.400 ;
        RECT 206.700 341.400 210.300 342.300 ;
        RECT 190.950 337.050 192.750 338.850 ;
        RECT 206.100 337.050 207.900 338.850 ;
        RECT 209.100 337.050 210.300 341.400 ;
        RECT 212.100 337.050 213.900 338.850 ;
        RECT 230.100 337.050 231.000 344.400 ;
        RECT 236.700 343.200 237.600 347.400 ;
        RECT 232.200 342.300 237.600 343.200 ;
        RECT 254.700 343.200 256.500 350.400 ;
        RECT 259.800 344.400 261.600 351.000 ;
        RECT 278.100 344.400 279.900 350.400 ;
        RECT 254.700 342.300 258.900 343.200 ;
        RECT 232.200 341.400 234.300 342.300 ;
        RECT 123.150 335.250 129.450 337.050 ;
        RECT 124.950 334.950 129.450 335.250 ;
        RECT 142.950 334.950 145.050 337.050 ;
        RECT 145.950 334.950 148.050 337.050 ;
        RECT 160.950 334.950 163.050 337.050 ;
        RECT 163.950 334.950 166.050 337.050 ;
        RECT 166.950 334.950 169.050 337.050 ;
        RECT 169.950 334.950 172.050 337.050 ;
        RECT 184.950 334.950 187.050 337.050 ;
        RECT 187.950 334.950 190.050 337.050 ;
        RECT 190.950 334.950 193.050 337.050 ;
        RECT 205.950 334.950 208.050 337.050 ;
        RECT 208.950 334.950 211.050 337.050 ;
        RECT 211.950 334.950 214.050 337.050 ;
        RECT 214.950 334.950 217.050 337.050 ;
        RECT 230.100 334.950 232.200 337.050 ;
        RECT 119.550 332.100 121.650 332.400 ;
        RECT 125.550 332.100 127.350 332.250 ;
        RECT 119.550 330.900 127.350 332.100 ;
        RECT 119.550 330.300 121.650 330.900 ;
        RECT 125.550 330.450 127.350 330.900 ;
        RECT 115.950 327.300 120.750 328.200 ;
        RECT 128.250 327.600 129.450 334.950 ;
        RECT 143.100 333.150 144.900 334.950 ;
        RECT 119.550 326.400 120.750 327.300 ;
        RECT 116.850 326.100 118.650 326.400 ;
        RECT 104.250 324.600 106.350 325.500 ;
        RECT 112.950 325.200 118.650 326.100 ;
        RECT 116.850 324.600 118.650 325.200 ;
        RECT 119.550 324.600 122.550 326.400 ;
        RECT 104.550 315.600 106.350 324.600 ;
        RECT 108.450 323.550 110.250 324.300 ;
        RECT 113.250 323.550 115.050 324.300 ;
        RECT 108.450 322.500 115.050 323.550 ;
        RECT 109.350 315.000 111.150 321.600 ;
        RECT 112.350 315.600 114.150 322.500 ;
        RECT 119.550 321.600 121.650 323.700 ;
        RECT 115.350 315.000 117.150 321.600 ;
        RECT 119.850 315.600 121.650 321.600 ;
        RECT 124.650 315.000 126.450 327.600 ;
        RECT 127.650 315.600 129.450 327.600 ;
        RECT 146.100 321.600 147.300 334.950 ;
        RECT 164.100 333.150 165.900 334.950 ;
        RECT 170.100 322.800 171.000 334.950 ;
        RECT 164.400 321.900 171.000 322.800 ;
        RECT 164.400 321.600 165.900 321.900 ;
        RECT 143.100 315.000 144.900 321.600 ;
        RECT 146.100 315.600 147.900 321.600 ;
        RECT 161.100 315.000 162.900 321.600 ;
        RECT 164.100 315.600 165.900 321.600 ;
        RECT 170.100 321.600 171.000 321.900 ;
        RECT 188.700 321.600 189.900 334.950 ;
        RECT 209.100 327.600 210.300 334.950 ;
        RECT 215.100 333.150 216.900 334.950 ;
        RECT 231.000 327.600 232.200 334.950 ;
        RECT 233.400 330.900 234.300 341.400 ;
        RECT 238.800 337.050 240.600 338.850 ;
        RECT 254.100 337.050 255.900 338.850 ;
        RECT 257.700 337.050 258.900 342.300 ;
        RECT 278.700 342.300 279.900 344.400 ;
        RECT 281.100 345.300 282.900 350.400 ;
        RECT 284.100 346.200 285.900 351.000 ;
        RECT 287.100 345.300 288.900 350.400 ;
        RECT 281.100 343.950 288.900 345.300 ;
        RECT 302.400 344.400 304.200 351.000 ;
        RECT 307.500 343.200 309.300 350.400 ;
        RECT 326.100 345.300 327.900 350.400 ;
        RECT 329.100 346.200 330.900 351.000 ;
        RECT 332.100 345.300 333.900 350.400 ;
        RECT 326.100 343.950 333.900 345.300 ;
        RECT 335.100 344.400 336.900 350.400 ;
        RECT 339.150 346.200 340.950 350.400 ;
        RECT 338.550 344.400 340.950 346.200 ;
        RECT 342.150 344.400 343.950 351.000 ;
        RECT 346.950 348.300 348.750 350.400 ;
        RECT 345.150 347.400 348.750 348.300 ;
        RECT 351.450 347.400 353.250 351.000 ;
        RECT 354.750 347.400 356.550 350.400 ;
        RECT 357.750 347.400 359.550 351.000 ;
        RECT 362.250 347.400 364.050 350.400 ;
        RECT 344.850 346.800 348.750 347.400 ;
        RECT 344.850 345.300 346.950 346.800 ;
        RECT 354.750 346.500 355.800 347.400 ;
        RECT 305.100 342.300 309.300 343.200 ;
        RECT 335.100 342.300 336.300 344.400 ;
        RECT 278.700 341.400 282.300 342.300 ;
        RECT 259.950 337.050 261.750 338.850 ;
        RECT 278.100 337.050 279.900 338.850 ;
        RECT 281.100 337.050 282.300 341.400 ;
        RECT 284.100 337.050 285.900 338.850 ;
        RECT 302.250 337.050 304.050 338.850 ;
        RECT 305.100 337.050 306.300 342.300 ;
        RECT 332.700 341.400 336.300 342.300 ;
        RECT 308.100 337.050 309.900 338.850 ;
        RECT 329.100 337.050 330.900 338.850 ;
        RECT 332.700 337.050 333.900 341.400 ;
        RECT 335.100 337.050 336.900 338.850 ;
        RECT 235.500 334.950 237.600 337.050 ;
        RECT 238.800 334.950 240.900 337.050 ;
        RECT 253.950 334.950 256.050 337.050 ;
        RECT 256.950 334.950 259.050 337.050 ;
        RECT 259.950 334.950 262.050 337.050 ;
        RECT 277.950 334.950 280.050 337.050 ;
        RECT 280.950 334.950 283.050 337.050 ;
        RECT 283.950 334.950 286.050 337.050 ;
        RECT 286.950 334.950 289.050 337.050 ;
        RECT 301.950 334.950 304.050 337.050 ;
        RECT 304.950 334.950 307.050 337.050 ;
        RECT 307.950 334.950 310.050 337.050 ;
        RECT 325.950 334.950 328.050 337.050 ;
        RECT 328.950 334.950 331.050 337.050 ;
        RECT 331.950 334.950 334.050 337.050 ;
        RECT 334.950 334.950 337.050 337.050 ;
        RECT 235.200 333.150 237.000 334.950 ;
        RECT 233.100 330.300 234.900 330.900 ;
        RECT 233.100 329.100 240.900 330.300 ;
        RECT 239.700 327.600 240.900 329.100 ;
        RECT 209.100 326.100 211.500 327.600 ;
        RECT 207.000 323.100 208.800 324.900 ;
        RECT 167.100 315.000 168.900 321.000 ;
        RECT 170.100 315.600 171.900 321.600 ;
        RECT 185.100 315.000 186.900 321.600 ;
        RECT 188.100 315.600 189.900 321.600 ;
        RECT 191.100 315.000 192.900 321.600 ;
        RECT 206.700 315.000 208.500 321.600 ;
        RECT 209.700 315.600 211.500 326.100 ;
        RECT 214.800 315.000 216.600 327.600 ;
        RECT 231.000 326.100 233.400 327.600 ;
        RECT 231.600 315.600 233.400 326.100 ;
        RECT 234.600 315.000 236.400 327.600 ;
        RECT 239.100 315.600 240.900 327.600 ;
        RECT 257.700 321.600 258.900 334.950 ;
        RECT 281.100 327.600 282.300 334.950 ;
        RECT 287.100 333.150 288.900 334.950 ;
        RECT 281.100 326.100 283.500 327.600 ;
        RECT 279.000 323.100 280.800 324.900 ;
        RECT 254.100 315.000 255.900 321.600 ;
        RECT 257.100 315.600 258.900 321.600 ;
        RECT 260.100 315.000 261.900 321.600 ;
        RECT 278.700 315.000 280.500 321.600 ;
        RECT 281.700 315.600 283.500 326.100 ;
        RECT 286.800 315.000 288.600 327.600 ;
        RECT 305.100 321.600 306.300 334.950 ;
        RECT 326.100 333.150 327.900 334.950 ;
        RECT 332.700 327.600 333.900 334.950 ;
        RECT 302.100 315.000 303.900 321.600 ;
        RECT 305.100 315.600 306.900 321.600 ;
        RECT 308.100 315.000 309.900 321.600 ;
        RECT 326.400 315.000 328.200 327.600 ;
        RECT 331.500 326.100 333.900 327.600 ;
        RECT 338.550 329.700 339.450 344.400 ;
        RECT 347.850 343.800 349.650 345.600 ;
        RECT 350.850 345.450 355.800 346.500 ;
        RECT 350.850 344.700 352.650 345.450 ;
        RECT 362.250 345.300 364.650 347.400 ;
        RECT 367.350 344.400 369.150 351.000 ;
        RECT 370.650 344.400 372.450 350.400 ;
        RECT 386.400 344.400 388.200 351.000 ;
        RECT 347.850 342.000 348.900 343.800 ;
        RECT 358.050 342.000 359.850 342.600 ;
        RECT 347.850 340.800 359.850 342.000 ;
        RECT 340.950 339.600 348.900 340.800 ;
        RECT 340.950 337.050 342.750 339.600 ;
        RECT 347.100 339.000 348.900 339.600 ;
        RECT 344.100 337.800 345.900 338.400 ;
        RECT 340.950 334.950 343.050 337.050 ;
        RECT 344.100 336.600 352.200 337.800 ;
        RECT 350.100 334.950 352.200 336.600 ;
        RECT 348.450 329.700 350.250 330.000 ;
        RECT 338.550 329.100 350.250 329.700 ;
        RECT 338.550 328.500 356.850 329.100 ;
        RECT 338.550 327.600 339.450 328.500 ;
        RECT 348.450 328.200 356.850 328.500 ;
        RECT 331.500 315.600 333.300 326.100 ;
        RECT 338.550 325.800 340.950 327.600 ;
        RECT 334.200 323.100 336.000 324.900 ;
        RECT 334.500 315.000 336.300 321.600 ;
        RECT 339.150 315.600 340.950 325.800 ;
        RECT 342.150 315.000 343.950 327.600 ;
        RECT 353.250 326.700 355.050 327.300 ;
        RECT 347.250 325.500 355.050 326.700 ;
        RECT 355.950 326.100 356.850 328.200 ;
        RECT 358.950 328.200 359.850 340.800 ;
        RECT 371.250 337.050 372.450 344.400 ;
        RECT 391.500 343.200 393.300 350.400 ;
        RECT 410.400 344.400 412.200 351.000 ;
        RECT 415.500 343.200 417.300 350.400 ;
        RECT 389.100 342.300 393.300 343.200 ;
        RECT 413.100 342.300 417.300 343.200 ;
        RECT 431.100 347.400 432.900 350.400 ;
        RECT 431.100 343.500 432.300 347.400 ;
        RECT 434.100 344.400 435.900 351.000 ;
        RECT 437.100 344.400 438.900 350.400 ;
        RECT 452.100 344.400 453.900 350.400 ;
        RECT 431.100 342.600 436.800 343.500 ;
        RECT 386.250 337.050 388.050 338.850 ;
        RECT 389.100 337.050 390.300 342.300 ;
        RECT 392.100 337.050 393.900 338.850 ;
        RECT 410.250 337.050 412.050 338.850 ;
        RECT 413.100 337.050 414.300 342.300 ;
        RECT 435.000 341.700 436.800 342.600 ;
        RECT 416.100 337.050 417.900 338.850 ;
        RECT 366.150 335.250 372.450 337.050 ;
        RECT 367.950 334.950 372.450 335.250 ;
        RECT 385.950 334.950 388.050 337.050 ;
        RECT 388.950 334.950 391.050 337.050 ;
        RECT 391.950 334.950 394.050 337.050 ;
        RECT 409.950 334.950 412.050 337.050 ;
        RECT 412.950 334.950 415.050 337.050 ;
        RECT 415.950 334.950 418.050 337.050 ;
        RECT 431.400 334.950 433.500 337.050 ;
        RECT 362.550 332.100 364.650 332.400 ;
        RECT 368.550 332.100 370.350 332.250 ;
        RECT 362.550 330.900 370.350 332.100 ;
        RECT 362.550 330.300 364.650 330.900 ;
        RECT 368.550 330.450 370.350 330.900 ;
        RECT 358.950 327.300 363.750 328.200 ;
        RECT 371.250 327.600 372.450 334.950 ;
        RECT 362.550 326.400 363.750 327.300 ;
        RECT 359.850 326.100 361.650 326.400 ;
        RECT 347.250 324.600 349.350 325.500 ;
        RECT 355.950 325.200 361.650 326.100 ;
        RECT 359.850 324.600 361.650 325.200 ;
        RECT 362.550 324.600 365.550 326.400 ;
        RECT 347.550 315.600 349.350 324.600 ;
        RECT 351.450 323.550 353.250 324.300 ;
        RECT 356.250 323.550 358.050 324.300 ;
        RECT 351.450 322.500 358.050 323.550 ;
        RECT 352.350 315.000 354.150 321.600 ;
        RECT 355.350 315.600 357.150 322.500 ;
        RECT 362.550 321.600 364.650 323.700 ;
        RECT 358.350 315.000 360.150 321.600 ;
        RECT 362.850 315.600 364.650 321.600 ;
        RECT 367.650 315.000 369.450 327.600 ;
        RECT 370.650 315.600 372.450 327.600 ;
        RECT 389.100 321.600 390.300 334.950 ;
        RECT 400.950 324.450 403.050 325.050 ;
        RECT 409.950 324.450 412.050 324.900 ;
        RECT 400.950 323.550 412.050 324.450 ;
        RECT 400.950 322.950 403.050 323.550 ;
        RECT 409.950 322.800 412.050 323.550 ;
        RECT 413.100 321.600 414.300 334.950 ;
        RECT 431.400 333.150 433.200 334.950 ;
        RECT 435.000 330.300 435.900 341.700 ;
        RECT 437.700 337.050 438.900 344.400 ;
        RECT 452.700 342.300 453.900 344.400 ;
        RECT 455.100 345.300 456.900 350.400 ;
        RECT 458.100 346.200 459.900 351.000 ;
        RECT 461.100 345.300 462.900 350.400 ;
        RECT 455.100 343.950 462.900 345.300 ;
        RECT 476.100 347.400 477.900 350.400 ;
        RECT 476.100 343.500 477.300 347.400 ;
        RECT 479.100 344.400 480.900 351.000 ;
        RECT 482.100 344.400 483.900 350.400 ;
        RECT 500.400 344.400 502.200 351.000 ;
        RECT 476.100 342.600 481.800 343.500 ;
        RECT 452.700 341.400 456.300 342.300 ;
        RECT 452.100 337.050 453.900 338.850 ;
        RECT 455.100 337.050 456.300 341.400 ;
        RECT 480.000 341.700 481.800 342.600 ;
        RECT 458.100 337.050 459.900 338.850 ;
        RECT 436.800 334.950 438.900 337.050 ;
        RECT 451.950 334.950 454.050 337.050 ;
        RECT 454.950 334.950 457.050 337.050 ;
        RECT 457.950 334.950 460.050 337.050 ;
        RECT 460.950 334.950 463.050 337.050 ;
        RECT 476.400 334.950 478.500 337.050 ;
        RECT 435.000 329.400 436.800 330.300 ;
        RECT 431.100 328.500 436.800 329.400 ;
        RECT 431.100 321.600 432.300 328.500 ;
        RECT 437.700 327.600 438.900 334.950 ;
        RECT 386.100 315.000 387.900 321.600 ;
        RECT 389.100 315.600 390.900 321.600 ;
        RECT 392.100 315.000 393.900 321.600 ;
        RECT 410.100 315.000 411.900 321.600 ;
        RECT 413.100 315.600 414.900 321.600 ;
        RECT 416.100 315.000 417.900 321.600 ;
        RECT 431.100 315.600 432.900 321.600 ;
        RECT 434.100 315.000 435.900 325.800 ;
        RECT 437.100 315.600 438.900 327.600 ;
        RECT 455.100 327.600 456.300 334.950 ;
        RECT 461.100 333.150 462.900 334.950 ;
        RECT 476.400 333.150 478.200 334.950 ;
        RECT 480.000 330.300 480.900 341.700 ;
        RECT 482.700 337.050 483.900 344.400 ;
        RECT 505.500 343.200 507.300 350.400 ;
        RECT 521.100 347.400 522.900 350.400 ;
        RECT 524.100 347.400 525.900 351.000 ;
        RECT 539.100 347.400 540.900 350.400 ;
        RECT 503.100 342.300 507.300 343.200 ;
        RECT 500.250 337.050 502.050 338.850 ;
        RECT 503.100 337.050 504.300 342.300 ;
        RECT 506.100 337.050 507.900 338.850 ;
        RECT 521.700 337.050 522.900 347.400 ;
        RECT 539.100 343.500 540.300 347.400 ;
        RECT 542.100 344.400 543.900 351.000 ;
        RECT 545.100 344.400 546.900 350.400 ;
        RECT 539.100 342.600 544.800 343.500 ;
        RECT 543.000 341.700 544.800 342.600 ;
        RECT 481.800 334.950 483.900 337.050 ;
        RECT 499.950 334.950 502.050 337.050 ;
        RECT 502.950 334.950 505.050 337.050 ;
        RECT 505.950 334.950 508.050 337.050 ;
        RECT 520.950 334.950 523.050 337.050 ;
        RECT 523.950 334.950 526.050 337.050 ;
        RECT 539.400 334.950 541.500 337.050 ;
        RECT 480.000 329.400 481.800 330.300 ;
        RECT 476.100 328.500 481.800 329.400 ;
        RECT 455.100 326.100 457.500 327.600 ;
        RECT 453.000 323.100 454.800 324.900 ;
        RECT 452.700 315.000 454.500 321.600 ;
        RECT 455.700 315.600 457.500 326.100 ;
        RECT 460.800 315.000 462.600 327.600 ;
        RECT 476.100 321.600 477.300 328.500 ;
        RECT 482.700 327.600 483.900 334.950 ;
        RECT 476.100 315.600 477.900 321.600 ;
        RECT 479.100 315.000 480.900 325.800 ;
        RECT 482.100 315.600 483.900 327.600 ;
        RECT 503.100 321.600 504.300 334.950 ;
        RECT 521.700 321.600 522.900 334.950 ;
        RECT 524.100 333.150 525.900 334.950 ;
        RECT 539.400 333.150 541.200 334.950 ;
        RECT 543.000 330.300 543.900 341.700 ;
        RECT 545.700 337.050 546.900 344.400 ;
        RECT 563.100 345.300 564.900 350.400 ;
        RECT 566.100 346.200 567.900 351.000 ;
        RECT 569.100 345.300 570.900 350.400 ;
        RECT 563.100 343.950 570.900 345.300 ;
        RECT 572.100 344.400 573.900 350.400 ;
        RECT 576.150 346.200 577.950 350.400 ;
        RECT 575.550 344.400 577.950 346.200 ;
        RECT 579.150 344.400 580.950 351.000 ;
        RECT 583.950 348.300 585.750 350.400 ;
        RECT 582.150 347.400 585.750 348.300 ;
        RECT 588.450 347.400 590.250 351.000 ;
        RECT 591.750 347.400 593.550 350.400 ;
        RECT 594.750 347.400 596.550 351.000 ;
        RECT 599.250 347.400 601.050 350.400 ;
        RECT 581.850 346.800 585.750 347.400 ;
        RECT 581.850 345.300 583.950 346.800 ;
        RECT 591.750 346.500 592.800 347.400 ;
        RECT 572.100 342.300 573.300 344.400 ;
        RECT 569.700 341.400 573.300 342.300 ;
        RECT 566.100 337.050 567.900 338.850 ;
        RECT 569.700 337.050 570.900 341.400 ;
        RECT 572.100 337.050 573.900 338.850 ;
        RECT 544.800 334.950 546.900 337.050 ;
        RECT 562.950 334.950 565.050 337.050 ;
        RECT 565.950 334.950 568.050 337.050 ;
        RECT 568.950 334.950 571.050 337.050 ;
        RECT 571.950 334.950 574.050 337.050 ;
        RECT 543.000 329.400 544.800 330.300 ;
        RECT 539.100 328.500 544.800 329.400 ;
        RECT 539.100 321.600 540.300 328.500 ;
        RECT 545.700 327.600 546.900 334.950 ;
        RECT 563.100 333.150 564.900 334.950 ;
        RECT 569.700 327.600 570.900 334.950 ;
        RECT 500.100 315.000 501.900 321.600 ;
        RECT 503.100 315.600 504.900 321.600 ;
        RECT 506.100 315.000 507.900 321.600 ;
        RECT 521.100 315.600 522.900 321.600 ;
        RECT 524.100 315.000 525.900 321.600 ;
        RECT 539.100 315.600 540.900 321.600 ;
        RECT 542.100 315.000 543.900 325.800 ;
        RECT 545.100 315.600 546.900 327.600 ;
        RECT 563.400 315.000 565.200 327.600 ;
        RECT 568.500 326.100 570.900 327.600 ;
        RECT 575.550 329.700 576.450 344.400 ;
        RECT 584.850 343.800 586.650 345.600 ;
        RECT 587.850 345.450 592.800 346.500 ;
        RECT 587.850 344.700 589.650 345.450 ;
        RECT 599.250 345.300 601.650 347.400 ;
        RECT 604.350 344.400 606.150 351.000 ;
        RECT 607.650 344.400 609.450 350.400 ;
        RECT 626.100 347.400 627.900 351.000 ;
        RECT 629.100 347.400 630.900 350.400 ;
        RECT 584.850 342.000 585.900 343.800 ;
        RECT 595.050 342.000 596.850 342.600 ;
        RECT 584.850 340.800 596.850 342.000 ;
        RECT 577.950 339.600 585.900 340.800 ;
        RECT 577.950 337.050 579.750 339.600 ;
        RECT 584.100 339.000 585.900 339.600 ;
        RECT 581.100 337.800 582.900 338.400 ;
        RECT 577.950 334.950 580.050 337.050 ;
        RECT 581.100 336.600 589.200 337.800 ;
        RECT 587.100 334.950 589.200 336.600 ;
        RECT 585.450 329.700 587.250 330.000 ;
        RECT 575.550 329.100 587.250 329.700 ;
        RECT 575.550 328.500 593.850 329.100 ;
        RECT 575.550 327.600 576.450 328.500 ;
        RECT 585.450 328.200 593.850 328.500 ;
        RECT 568.500 315.600 570.300 326.100 ;
        RECT 575.550 325.800 577.950 327.600 ;
        RECT 571.200 323.100 573.000 324.900 ;
        RECT 571.500 315.000 573.300 321.600 ;
        RECT 576.150 315.600 577.950 325.800 ;
        RECT 579.150 315.000 580.950 327.600 ;
        RECT 590.250 326.700 592.050 327.300 ;
        RECT 584.250 325.500 592.050 326.700 ;
        RECT 592.950 326.100 593.850 328.200 ;
        RECT 595.950 328.200 596.850 340.800 ;
        RECT 608.250 337.050 609.450 344.400 ;
        RECT 629.100 337.050 630.300 347.400 ;
        RECT 645.000 344.400 646.800 351.000 ;
        RECT 649.500 345.600 651.300 350.400 ;
        RECT 652.500 347.400 654.300 351.000 ;
        RECT 649.500 344.400 654.600 345.600 ;
        RECT 668.100 344.400 669.900 350.400 ;
        RECT 671.100 344.400 672.900 351.000 ;
        RECT 634.950 342.450 637.050 343.050 ;
        RECT 646.950 342.450 649.050 343.050 ;
        RECT 634.950 341.550 649.050 342.450 ;
        RECT 634.950 340.950 637.050 341.550 ;
        RECT 646.950 340.950 649.050 341.550 ;
        RECT 644.100 337.050 645.900 338.850 ;
        RECT 650.250 337.050 652.050 338.850 ;
        RECT 653.700 337.050 654.600 344.400 ;
        RECT 668.700 337.050 669.900 344.400 ;
        RECT 686.100 342.600 687.900 350.400 ;
        RECT 690.600 344.400 692.400 351.000 ;
        RECT 693.600 346.200 695.400 350.400 ;
        RECT 693.600 344.400 696.300 346.200 ;
        RECT 692.700 342.600 694.500 343.500 ;
        RECT 686.100 341.700 694.500 342.600 ;
        RECT 671.100 337.050 672.900 338.850 ;
        RECT 686.250 337.050 688.050 338.850 ;
        RECT 603.150 335.250 609.450 337.050 ;
        RECT 604.950 334.950 609.450 335.250 ;
        RECT 625.950 334.950 628.050 337.050 ;
        RECT 628.950 334.950 631.050 337.050 ;
        RECT 643.950 334.950 646.050 337.050 ;
        RECT 646.950 334.950 649.050 337.050 ;
        RECT 649.950 334.950 652.050 337.050 ;
        RECT 652.950 334.950 655.050 337.050 ;
        RECT 667.950 334.950 670.050 337.050 ;
        RECT 670.950 334.950 673.050 337.050 ;
        RECT 686.100 334.950 688.200 337.050 ;
        RECT 599.550 332.100 601.650 332.400 ;
        RECT 605.550 332.100 607.350 332.250 ;
        RECT 599.550 330.900 607.350 332.100 ;
        RECT 599.550 330.300 601.650 330.900 ;
        RECT 605.550 330.450 607.350 330.900 ;
        RECT 595.950 327.300 600.750 328.200 ;
        RECT 608.250 327.600 609.450 334.950 ;
        RECT 626.100 333.150 627.900 334.950 ;
        RECT 599.550 326.400 600.750 327.300 ;
        RECT 596.850 326.100 598.650 326.400 ;
        RECT 584.250 324.600 586.350 325.500 ;
        RECT 592.950 325.200 598.650 326.100 ;
        RECT 596.850 324.600 598.650 325.200 ;
        RECT 599.550 324.600 602.550 326.400 ;
        RECT 584.550 315.600 586.350 324.600 ;
        RECT 588.450 323.550 590.250 324.300 ;
        RECT 593.250 323.550 595.050 324.300 ;
        RECT 588.450 322.500 595.050 323.550 ;
        RECT 589.350 315.000 591.150 321.600 ;
        RECT 592.350 315.600 594.150 322.500 ;
        RECT 599.550 321.600 601.650 323.700 ;
        RECT 595.350 315.000 597.150 321.600 ;
        RECT 599.850 315.600 601.650 321.600 ;
        RECT 604.650 315.000 606.450 327.600 ;
        RECT 607.650 315.600 609.450 327.600 ;
        RECT 629.100 321.600 630.300 334.950 ;
        RECT 647.250 333.150 649.050 334.950 ;
        RECT 634.950 330.450 637.050 331.050 ;
        RECT 649.950 330.450 652.050 331.050 ;
        RECT 634.950 329.550 652.050 330.450 ;
        RECT 634.950 328.950 637.050 329.550 ;
        RECT 649.950 328.950 652.050 329.550 ;
        RECT 653.700 327.600 654.600 334.950 ;
        RECT 668.700 327.600 669.900 334.950 ;
        RECT 644.100 326.700 651.900 327.600 ;
        RECT 626.100 315.000 627.900 321.600 ;
        RECT 629.100 315.600 630.900 321.600 ;
        RECT 644.100 315.600 645.900 326.700 ;
        RECT 647.100 315.000 648.900 325.800 ;
        RECT 650.100 315.600 651.900 326.700 ;
        RECT 653.100 315.600 654.900 327.600 ;
        RECT 668.100 315.600 669.900 327.600 ;
        RECT 671.100 315.000 672.900 327.600 ;
        RECT 689.100 321.600 690.000 341.700 ;
        RECT 695.400 337.050 696.300 344.400 ;
        RECT 713.700 343.200 715.500 350.400 ;
        RECT 718.800 344.400 720.600 351.000 ;
        RECT 734.400 344.400 736.200 351.000 ;
        RECT 739.500 343.200 741.300 350.400 ;
        RECT 755.100 347.400 756.900 351.000 ;
        RECT 758.100 347.400 759.900 350.400 ;
        RECT 713.700 342.300 717.900 343.200 ;
        RECT 713.100 337.050 714.900 338.850 ;
        RECT 716.700 337.050 717.900 342.300 ;
        RECT 737.100 342.300 741.300 343.200 ;
        RECT 718.950 337.050 720.750 338.850 ;
        RECT 734.250 337.050 736.050 338.850 ;
        RECT 737.100 337.050 738.300 342.300 ;
        RECT 740.100 337.050 741.900 338.850 ;
        RECT 758.100 337.050 759.300 347.400 ;
        RECT 776.100 344.400 777.900 350.400 ;
        RECT 776.700 342.300 777.900 344.400 ;
        RECT 779.100 345.300 780.900 350.400 ;
        RECT 782.100 346.200 783.900 351.000 ;
        RECT 785.100 345.300 786.900 350.400 ;
        RECT 779.100 343.950 786.900 345.300 ;
        RECT 776.700 341.400 780.300 342.300 ;
        RECT 800.100 341.400 801.900 351.000 ;
        RECT 806.700 342.000 808.500 350.400 ;
        RECT 827.100 344.400 828.900 350.400 ;
        RECT 827.700 342.300 828.900 344.400 ;
        RECT 830.100 345.300 831.900 350.400 ;
        RECT 833.100 346.200 834.900 351.000 ;
        RECT 836.100 345.300 837.900 350.400 ;
        RECT 830.100 343.950 837.900 345.300 ;
        RECT 852.000 344.400 853.800 351.000 ;
        RECT 856.500 345.600 858.300 350.400 ;
        RECT 859.500 347.400 861.300 351.000 ;
        RECT 856.500 344.400 861.600 345.600 ;
        RECT 760.950 339.450 763.050 340.050 ;
        RECT 760.950 338.550 771.450 339.450 ;
        RECT 760.950 337.950 763.050 338.550 ;
        RECT 691.500 334.950 693.600 337.050 ;
        RECT 694.800 334.950 696.900 337.050 ;
        RECT 712.950 334.950 715.050 337.050 ;
        RECT 715.950 334.950 718.050 337.050 ;
        RECT 718.950 334.950 721.050 337.050 ;
        RECT 733.950 334.950 736.050 337.050 ;
        RECT 736.950 334.950 739.050 337.050 ;
        RECT 739.950 334.950 742.050 337.050 ;
        RECT 754.950 334.950 757.050 337.050 ;
        RECT 757.950 334.950 760.050 337.050 ;
        RECT 691.200 333.150 693.000 334.950 ;
        RECT 695.400 327.600 696.300 334.950 ;
        RECT 686.100 315.000 687.900 321.600 ;
        RECT 689.100 315.600 690.900 321.600 ;
        RECT 692.100 315.000 693.900 327.000 ;
        RECT 695.100 315.600 696.900 327.600 ;
        RECT 716.700 321.600 717.900 334.950 ;
        RECT 718.950 330.450 721.050 330.750 ;
        RECT 733.950 330.450 736.050 331.050 ;
        RECT 718.950 329.550 736.050 330.450 ;
        RECT 718.950 328.650 721.050 329.550 ;
        RECT 733.950 328.950 736.050 329.550 ;
        RECT 737.100 321.600 738.300 334.950 ;
        RECT 755.100 333.150 756.900 334.950 ;
        RECT 758.100 321.600 759.300 334.950 ;
        RECT 770.550 334.050 771.450 338.550 ;
        RECT 776.100 337.050 777.900 338.850 ;
        RECT 779.100 337.050 780.300 341.400 ;
        RECT 806.700 340.800 810.000 342.000 ;
        RECT 827.700 341.400 831.300 342.300 ;
        RECT 782.100 337.050 783.900 338.850 ;
        RECT 800.100 337.050 801.900 338.850 ;
        RECT 806.100 337.050 807.900 338.850 ;
        RECT 809.100 337.050 810.000 340.800 ;
        RECT 827.100 337.050 828.900 338.850 ;
        RECT 830.100 337.050 831.300 341.400 ;
        RECT 838.950 339.450 841.050 340.050 ;
        RECT 844.950 339.450 847.050 340.050 ;
        RECT 833.100 337.050 834.900 338.850 ;
        RECT 838.950 338.550 847.050 339.450 ;
        RECT 838.950 337.950 841.050 338.550 ;
        RECT 844.950 337.950 847.050 338.550 ;
        RECT 851.100 337.050 852.900 338.850 ;
        RECT 857.250 337.050 859.050 338.850 ;
        RECT 860.700 337.050 861.600 344.400 ;
        RECT 868.950 345.450 871.050 346.050 ;
        RECT 874.950 345.450 877.050 349.050 ;
        RECT 868.950 345.000 877.050 345.450 ;
        RECT 868.950 344.550 876.450 345.000 ;
        RECT 868.950 343.950 871.050 344.550 ;
        RECT 878.100 341.400 879.900 351.000 ;
        RECT 884.700 342.000 886.500 350.400 ;
        RECT 902.100 347.400 903.900 351.000 ;
        RECT 905.100 347.400 906.900 350.400 ;
        RECT 908.100 347.400 909.900 351.000 ;
        RECT 923.100 347.400 924.900 351.000 ;
        RECT 926.100 347.400 927.900 350.400 ;
        RECT 884.700 340.800 888.000 342.000 ;
        RECT 878.100 337.050 879.900 338.850 ;
        RECT 884.100 337.050 885.900 338.850 ;
        RECT 887.100 337.050 888.000 340.800 ;
        RECT 897.000 339.450 901.050 340.050 ;
        RECT 896.550 337.950 901.050 339.450 ;
        RECT 775.950 334.950 778.050 337.050 ;
        RECT 778.950 334.950 781.050 337.050 ;
        RECT 781.950 334.950 784.050 337.050 ;
        RECT 784.950 334.950 787.050 337.050 ;
        RECT 799.950 334.950 802.050 337.050 ;
        RECT 802.950 334.950 805.050 337.050 ;
        RECT 805.950 334.950 808.050 337.050 ;
        RECT 808.950 334.950 811.050 337.050 ;
        RECT 826.950 334.950 829.050 337.050 ;
        RECT 829.950 334.950 832.050 337.050 ;
        RECT 832.950 334.950 835.050 337.050 ;
        RECT 835.950 334.950 838.050 337.050 ;
        RECT 850.950 334.950 853.050 337.050 ;
        RECT 853.950 334.950 856.050 337.050 ;
        RECT 856.950 334.950 859.050 337.050 ;
        RECT 859.950 334.950 862.050 337.050 ;
        RECT 877.950 334.950 880.050 337.050 ;
        RECT 880.950 334.950 883.050 337.050 ;
        RECT 883.950 334.950 886.050 337.050 ;
        RECT 886.950 334.950 889.050 337.050 ;
        RECT 770.550 332.550 775.050 334.050 ;
        RECT 771.000 331.950 775.050 332.550 ;
        RECT 779.100 327.600 780.300 334.950 ;
        RECT 785.100 333.150 786.900 334.950 ;
        RECT 803.100 333.150 804.900 334.950 ;
        RECT 779.100 326.100 781.500 327.600 ;
        RECT 777.000 323.100 778.800 324.900 ;
        RECT 713.100 315.000 714.900 321.600 ;
        RECT 716.100 315.600 717.900 321.600 ;
        RECT 719.100 315.000 720.900 321.600 ;
        RECT 734.100 315.000 735.900 321.600 ;
        RECT 737.100 315.600 738.900 321.600 ;
        RECT 740.100 315.000 741.900 321.600 ;
        RECT 755.100 315.000 756.900 321.600 ;
        RECT 758.100 315.600 759.900 321.600 ;
        RECT 776.700 315.000 778.500 321.600 ;
        RECT 779.700 315.600 781.500 326.100 ;
        RECT 784.800 315.000 786.600 327.600 ;
        RECT 809.100 322.800 810.000 334.950 ;
        RECT 830.100 327.600 831.300 334.950 ;
        RECT 836.100 333.150 837.900 334.950 ;
        RECT 854.250 333.150 856.050 334.950 ;
        RECT 835.950 330.450 838.050 331.050 ;
        RECT 850.950 330.450 853.050 331.050 ;
        RECT 835.950 329.550 853.050 330.450 ;
        RECT 835.950 328.950 838.050 329.550 ;
        RECT 850.950 328.950 853.050 329.550 ;
        RECT 860.700 327.600 861.600 334.950 ;
        RECT 881.100 333.150 882.900 334.950 ;
        RECT 830.100 326.100 832.500 327.600 ;
        RECT 828.000 323.100 829.800 324.900 ;
        RECT 803.400 321.900 810.000 322.800 ;
        RECT 803.400 321.600 804.900 321.900 ;
        RECT 800.100 315.000 801.900 321.600 ;
        RECT 803.100 315.600 804.900 321.600 ;
        RECT 809.100 321.600 810.000 321.900 ;
        RECT 806.100 315.000 807.900 321.000 ;
        RECT 809.100 315.600 810.900 321.600 ;
        RECT 827.700 315.000 829.500 321.600 ;
        RECT 830.700 315.600 832.500 326.100 ;
        RECT 835.800 315.000 837.600 327.600 ;
        RECT 851.100 326.700 858.900 327.600 ;
        RECT 851.100 315.600 852.900 326.700 ;
        RECT 854.100 315.000 855.900 325.800 ;
        RECT 857.100 315.600 858.900 326.700 ;
        RECT 860.100 315.600 861.900 327.600 ;
        RECT 887.100 322.800 888.000 334.950 ;
        RECT 889.950 333.450 892.050 334.050 ;
        RECT 896.550 333.450 897.450 337.950 ;
        RECT 905.400 337.050 906.300 347.400 ;
        RECT 910.950 339.450 913.050 340.050 ;
        RECT 910.950 338.550 918.450 339.450 ;
        RECT 910.950 337.950 913.050 338.550 ;
        RECT 901.950 334.950 904.050 337.050 ;
        RECT 904.950 334.950 907.050 337.050 ;
        RECT 907.950 334.950 910.050 337.050 ;
        RECT 889.950 332.550 897.450 333.450 ;
        RECT 902.250 333.150 904.050 334.950 ;
        RECT 889.950 331.950 892.050 332.550 ;
        RECT 905.400 327.600 906.300 334.950 ;
        RECT 908.100 333.150 909.900 334.950 ;
        RECT 917.550 334.050 918.450 338.550 ;
        RECT 926.100 337.050 927.300 347.400 ;
        RECT 941.400 344.400 943.200 351.000 ;
        RECT 946.500 343.200 948.300 350.400 ;
        RECT 962.700 347.400 964.500 351.000 ;
        RECT 965.700 345.600 967.500 350.400 ;
        RECT 944.100 342.300 948.300 343.200 ;
        RECT 962.400 344.400 967.500 345.600 ;
        RECT 970.200 344.400 972.000 351.000 ;
        RECT 941.250 337.050 943.050 338.850 ;
        RECT 944.100 337.050 945.300 342.300 ;
        RECT 947.100 337.050 948.900 338.850 ;
        RECT 962.400 337.050 963.300 344.400 ;
        RECT 967.950 342.450 970.050 343.200 ;
        RECT 979.950 342.450 982.050 343.050 ;
        RECT 967.950 341.550 982.050 342.450 ;
        RECT 986.100 342.600 987.900 350.400 ;
        RECT 990.600 344.400 992.400 351.000 ;
        RECT 993.600 346.200 995.400 350.400 ;
        RECT 993.600 344.400 996.300 346.200 ;
        RECT 992.700 342.600 994.500 343.500 ;
        RECT 986.100 341.700 994.500 342.600 ;
        RECT 967.950 341.100 970.050 341.550 ;
        RECT 979.950 340.950 982.050 341.550 ;
        RECT 964.950 337.050 966.750 338.850 ;
        RECT 971.100 337.050 972.900 338.850 ;
        RECT 986.250 337.050 988.050 338.850 ;
        RECT 922.950 334.950 925.050 337.050 ;
        RECT 925.950 334.950 928.050 337.050 ;
        RECT 940.950 334.950 943.050 337.050 ;
        RECT 943.950 334.950 946.050 337.050 ;
        RECT 946.950 334.950 949.050 337.050 ;
        RECT 961.950 334.950 964.050 337.050 ;
        RECT 964.950 334.950 967.050 337.050 ;
        RECT 967.950 334.950 970.050 337.050 ;
        RECT 970.950 334.950 973.050 337.050 ;
        RECT 986.100 334.950 988.200 337.050 ;
        RECT 917.550 332.550 922.050 334.050 ;
        RECT 923.100 333.150 924.900 334.950 ;
        RECT 918.000 331.950 922.050 332.550 ;
        RECT 881.400 321.900 888.000 322.800 ;
        RECT 881.400 321.600 882.900 321.900 ;
        RECT 878.100 315.000 879.900 321.600 ;
        RECT 881.100 315.600 882.900 321.600 ;
        RECT 887.100 321.600 888.000 321.900 ;
        RECT 884.100 315.000 885.900 321.000 ;
        RECT 887.100 315.600 888.900 321.600 ;
        RECT 902.100 315.000 903.900 327.600 ;
        RECT 905.400 326.400 909.000 327.600 ;
        RECT 907.200 315.600 909.000 326.400 ;
        RECT 926.100 321.600 927.300 334.950 ;
        RECT 931.950 330.450 934.050 330.900 ;
        RECT 940.950 330.450 943.050 331.050 ;
        RECT 931.950 329.550 943.050 330.450 ;
        RECT 931.950 328.800 934.050 329.550 ;
        RECT 940.950 328.950 943.050 329.550 ;
        RECT 944.100 321.600 945.300 334.950 ;
        RECT 962.400 327.600 963.300 334.950 ;
        RECT 967.950 333.150 969.750 334.950 ;
        RECT 923.100 315.000 924.900 321.600 ;
        RECT 926.100 315.600 927.900 321.600 ;
        RECT 941.100 315.000 942.900 321.600 ;
        RECT 944.100 315.600 945.900 321.600 ;
        RECT 947.100 315.000 948.900 321.600 ;
        RECT 962.100 315.600 963.900 327.600 ;
        RECT 965.100 326.700 972.900 327.600 ;
        RECT 965.100 315.600 966.900 326.700 ;
        RECT 968.100 315.000 969.900 325.800 ;
        RECT 971.100 315.600 972.900 326.700 ;
        RECT 989.100 321.600 990.000 341.700 ;
        RECT 995.400 337.050 996.300 344.400 ;
        RECT 991.500 334.950 993.600 337.050 ;
        RECT 994.800 334.950 996.900 337.050 ;
        RECT 991.200 333.150 993.000 334.950 ;
        RECT 995.400 327.600 996.300 334.950 ;
        RECT 986.100 315.000 987.900 321.600 ;
        RECT 989.100 315.600 990.900 321.600 ;
        RECT 992.100 315.000 993.900 327.000 ;
        RECT 995.100 315.600 996.900 327.600 ;
        RECT 14.100 305.400 15.900 312.000 ;
        RECT 17.100 305.400 18.900 311.400 ;
        RECT 20.100 305.400 21.900 312.000 ;
        RECT 17.700 292.050 18.900 305.400 ;
        RECT 24.150 301.200 25.950 311.400 ;
        RECT 23.550 299.400 25.950 301.200 ;
        RECT 27.150 299.400 28.950 312.000 ;
        RECT 32.550 302.400 34.350 311.400 ;
        RECT 37.350 305.400 39.150 312.000 ;
        RECT 40.350 304.500 42.150 311.400 ;
        RECT 43.350 305.400 45.150 312.000 ;
        RECT 47.850 305.400 49.650 311.400 ;
        RECT 36.450 303.450 43.050 304.500 ;
        RECT 36.450 302.700 38.250 303.450 ;
        RECT 41.250 302.700 43.050 303.450 ;
        RECT 47.550 303.300 49.650 305.400 ;
        RECT 32.250 301.500 34.350 302.400 ;
        RECT 44.850 301.800 46.650 302.400 ;
        RECT 32.250 300.300 40.050 301.500 ;
        RECT 38.250 299.700 40.050 300.300 ;
        RECT 40.950 300.900 46.650 301.800 ;
        RECT 23.550 298.500 24.450 299.400 ;
        RECT 40.950 298.800 41.850 300.900 ;
        RECT 44.850 300.600 46.650 300.900 ;
        RECT 47.550 300.600 50.550 302.400 ;
        RECT 47.550 299.700 48.750 300.600 ;
        RECT 33.450 298.500 41.850 298.800 ;
        RECT 23.550 297.900 41.850 298.500 ;
        RECT 43.950 298.800 48.750 299.700 ;
        RECT 52.650 299.400 54.450 312.000 ;
        RECT 55.650 299.400 57.450 311.400 ;
        RECT 74.100 299.400 75.900 312.000 ;
        RECT 79.200 300.600 81.000 311.400 ;
        RECT 77.400 299.400 81.000 300.600 ;
        RECT 98.100 305.400 99.900 311.400 ;
        RECT 23.550 297.300 35.250 297.900 ;
        RECT 13.950 289.950 16.050 292.050 ;
        RECT 16.950 289.950 19.050 292.050 ;
        RECT 19.950 289.950 22.050 292.050 ;
        RECT 14.100 288.150 15.900 289.950 ;
        RECT 17.700 284.700 18.900 289.950 ;
        RECT 19.950 288.150 21.750 289.950 ;
        RECT 14.700 283.800 18.900 284.700 ;
        RECT 14.700 276.600 16.500 283.800 ;
        RECT 23.550 282.600 24.450 297.300 ;
        RECT 33.450 297.000 35.250 297.300 ;
        RECT 25.950 289.950 28.050 292.050 ;
        RECT 35.100 290.400 37.200 292.050 ;
        RECT 25.950 287.400 27.750 289.950 ;
        RECT 29.100 289.200 37.200 290.400 ;
        RECT 29.100 288.600 30.900 289.200 ;
        RECT 32.100 287.400 33.900 288.000 ;
        RECT 25.950 286.200 33.900 287.400 ;
        RECT 43.950 286.200 44.850 298.800 ;
        RECT 47.550 296.100 49.650 296.700 ;
        RECT 53.550 296.100 55.350 296.550 ;
        RECT 47.550 294.900 55.350 296.100 ;
        RECT 47.550 294.600 49.650 294.900 ;
        RECT 53.550 294.750 55.350 294.900 ;
        RECT 56.250 292.050 57.450 299.400 ;
        RECT 74.250 292.050 76.050 293.850 ;
        RECT 77.400 292.050 78.300 299.400 ;
        RECT 98.100 298.500 99.300 305.400 ;
        RECT 101.100 301.200 102.900 312.000 ;
        RECT 104.100 299.400 105.900 311.400 ;
        RECT 119.100 299.400 120.900 311.400 ;
        RECT 122.100 300.300 123.900 311.400 ;
        RECT 125.100 301.200 126.900 312.000 ;
        RECT 128.100 300.300 129.900 311.400 ;
        RECT 143.100 305.400 144.900 312.000 ;
        RECT 146.100 305.400 147.900 311.400 ;
        RECT 149.100 306.000 150.900 312.000 ;
        RECT 146.400 305.100 147.900 305.400 ;
        RECT 152.100 305.400 153.900 311.400 ;
        RECT 170.100 305.400 171.900 312.000 ;
        RECT 173.100 305.400 174.900 311.400 ;
        RECT 176.100 305.400 177.900 312.000 ;
        RECT 194.100 305.400 195.900 312.000 ;
        RECT 197.100 305.400 198.900 311.400 ;
        RECT 212.100 305.400 213.900 312.000 ;
        RECT 215.100 305.400 216.900 311.400 ;
        RECT 218.100 306.000 219.900 312.000 ;
        RECT 152.100 305.100 153.000 305.400 ;
        RECT 146.400 304.200 153.000 305.100 ;
        RECT 122.100 299.400 129.900 300.300 ;
        RECT 98.100 297.600 103.800 298.500 ;
        RECT 102.000 296.700 103.800 297.600 ;
        RECT 80.100 292.050 81.900 293.850 ;
        RECT 98.400 292.050 100.200 293.850 ;
        RECT 52.950 291.750 57.450 292.050 ;
        RECT 51.150 289.950 57.450 291.750 ;
        RECT 73.950 289.950 76.050 292.050 ;
        RECT 76.950 289.950 79.050 292.050 ;
        RECT 79.950 289.950 82.050 292.050 ;
        RECT 98.400 289.950 100.500 292.050 ;
        RECT 32.850 285.000 44.850 286.200 ;
        RECT 32.850 283.200 33.900 285.000 ;
        RECT 43.050 284.400 44.850 285.000 ;
        RECT 19.800 276.000 21.600 282.600 ;
        RECT 23.550 280.800 25.950 282.600 ;
        RECT 24.150 276.600 25.950 280.800 ;
        RECT 27.150 276.000 28.950 282.600 ;
        RECT 29.850 280.200 31.950 281.700 ;
        RECT 32.850 281.400 34.650 283.200 ;
        RECT 56.250 282.600 57.450 289.950 ;
        RECT 58.950 288.450 61.050 289.050 ;
        RECT 70.950 288.450 73.050 289.050 ;
        RECT 58.950 287.550 73.050 288.450 ;
        RECT 58.950 286.950 61.050 287.550 ;
        RECT 70.950 286.950 73.050 287.550 ;
        RECT 35.850 281.550 37.650 282.300 ;
        RECT 35.850 280.500 40.800 281.550 ;
        RECT 29.850 279.600 33.750 280.200 ;
        RECT 39.750 279.600 40.800 280.500 ;
        RECT 47.250 279.600 49.650 281.700 ;
        RECT 30.150 278.700 33.750 279.600 ;
        RECT 31.950 276.600 33.750 278.700 ;
        RECT 36.450 276.000 38.250 279.600 ;
        RECT 39.750 276.600 41.550 279.600 ;
        RECT 42.750 276.000 44.550 279.600 ;
        RECT 47.250 276.600 49.050 279.600 ;
        RECT 52.350 276.000 54.150 282.600 ;
        RECT 55.650 276.600 57.450 282.600 ;
        RECT 77.400 279.600 78.300 289.950 ;
        RECT 102.000 285.300 102.900 296.700 ;
        RECT 104.700 292.050 105.900 299.400 ;
        RECT 119.400 292.050 120.300 299.400 ;
        RECT 121.950 297.450 124.050 298.050 ;
        RECT 136.950 297.450 139.050 298.050 ;
        RECT 148.950 297.450 151.050 298.050 ;
        RECT 121.950 296.550 151.050 297.450 ;
        RECT 121.950 295.950 124.050 296.550 ;
        RECT 136.950 295.950 139.050 296.550 ;
        RECT 148.950 295.950 151.050 296.550 ;
        RECT 124.950 292.050 126.750 293.850 ;
        RECT 146.100 292.050 147.900 293.850 ;
        RECT 152.100 292.050 153.000 304.200 ;
        RECT 173.100 292.050 174.300 305.400 ;
        RECT 194.100 292.050 195.900 293.850 ;
        RECT 197.100 292.050 198.300 305.400 ;
        RECT 215.400 305.100 216.900 305.400 ;
        RECT 221.100 305.400 222.900 311.400 ;
        RECT 239.100 305.400 240.900 312.000 ;
        RECT 242.100 305.400 243.900 311.400 ;
        RECT 245.100 305.400 246.900 312.000 ;
        RECT 260.700 305.400 262.500 312.000 ;
        RECT 221.100 305.100 222.000 305.400 ;
        RECT 215.400 304.200 222.000 305.100 ;
        RECT 199.950 300.450 202.050 301.050 ;
        RECT 217.950 300.450 220.050 301.050 ;
        RECT 199.950 299.550 220.050 300.450 ;
        RECT 199.950 298.950 202.050 299.550 ;
        RECT 217.950 298.950 220.050 299.550 ;
        RECT 202.950 297.450 205.050 298.050 ;
        RECT 211.950 297.450 214.050 298.050 ;
        RECT 202.950 296.550 214.050 297.450 ;
        RECT 202.950 295.950 205.050 296.550 ;
        RECT 211.950 295.950 214.050 296.550 ;
        RECT 215.100 292.050 216.900 293.850 ;
        RECT 221.100 292.050 222.000 304.200 ;
        RECT 242.100 292.050 243.300 305.400 ;
        RECT 261.000 302.100 262.800 303.900 ;
        RECT 263.700 300.900 265.500 311.400 ;
        RECT 263.100 299.400 265.500 300.900 ;
        RECT 268.800 299.400 270.600 312.000 ;
        RECT 273.150 301.200 274.950 311.400 ;
        RECT 272.550 299.400 274.950 301.200 ;
        RECT 276.150 299.400 277.950 312.000 ;
        RECT 281.550 302.400 283.350 311.400 ;
        RECT 286.350 305.400 288.150 312.000 ;
        RECT 289.350 304.500 291.150 311.400 ;
        RECT 292.350 305.400 294.150 312.000 ;
        RECT 296.850 305.400 298.650 311.400 ;
        RECT 285.450 303.450 292.050 304.500 ;
        RECT 285.450 302.700 287.250 303.450 ;
        RECT 290.250 302.700 292.050 303.450 ;
        RECT 296.550 303.300 298.650 305.400 ;
        RECT 281.250 301.500 283.350 302.400 ;
        RECT 293.850 301.800 295.650 302.400 ;
        RECT 281.250 300.300 289.050 301.500 ;
        RECT 287.250 299.700 289.050 300.300 ;
        RECT 289.950 300.900 295.650 301.800 ;
        RECT 263.100 292.050 264.300 299.400 ;
        RECT 272.550 298.500 273.450 299.400 ;
        RECT 289.950 298.800 290.850 300.900 ;
        RECT 293.850 300.600 295.650 300.900 ;
        RECT 296.550 300.600 299.550 302.400 ;
        RECT 296.550 299.700 297.750 300.600 ;
        RECT 282.450 298.500 290.850 298.800 ;
        RECT 272.550 297.900 290.850 298.500 ;
        RECT 292.950 298.800 297.750 299.700 ;
        RECT 301.650 299.400 303.450 312.000 ;
        RECT 304.650 299.400 306.450 311.400 ;
        RECT 320.400 299.400 322.200 312.000 ;
        RECT 325.500 300.900 327.300 311.400 ;
        RECT 328.500 305.400 330.300 312.000 ;
        RECT 344.100 305.400 345.900 312.000 ;
        RECT 347.100 305.400 348.900 311.400 ;
        RECT 350.100 305.400 351.900 312.000 ;
        RECT 328.200 302.100 330.000 303.900 ;
        RECT 325.500 299.400 327.900 300.900 ;
        RECT 272.550 297.300 284.250 297.900 ;
        RECT 269.100 292.050 270.900 293.850 ;
        RECT 103.800 289.950 105.900 292.050 ;
        RECT 118.950 289.950 121.050 292.050 ;
        RECT 121.950 289.950 124.050 292.050 ;
        RECT 124.950 289.950 127.050 292.050 ;
        RECT 127.950 289.950 130.050 292.050 ;
        RECT 142.950 289.950 145.050 292.050 ;
        RECT 145.950 289.950 148.050 292.050 ;
        RECT 148.950 289.950 151.050 292.050 ;
        RECT 151.950 289.950 154.050 292.050 ;
        RECT 169.950 289.950 172.050 292.050 ;
        RECT 172.950 289.950 175.050 292.050 ;
        RECT 175.950 289.950 178.050 292.050 ;
        RECT 193.950 289.950 196.050 292.050 ;
        RECT 196.950 289.950 199.050 292.050 ;
        RECT 211.950 289.950 214.050 292.050 ;
        RECT 214.950 289.950 217.050 292.050 ;
        RECT 217.950 289.950 220.050 292.050 ;
        RECT 220.950 289.950 223.050 292.050 ;
        RECT 238.950 289.950 241.050 292.050 ;
        RECT 241.950 289.950 244.050 292.050 ;
        RECT 244.950 289.950 247.050 292.050 ;
        RECT 259.950 289.950 262.050 292.050 ;
        RECT 262.950 289.950 265.050 292.050 ;
        RECT 265.950 289.950 268.050 292.050 ;
        RECT 268.950 289.950 271.050 292.050 ;
        RECT 102.000 284.400 103.800 285.300 ;
        RECT 98.100 283.500 103.800 284.400 ;
        RECT 98.100 279.600 99.300 283.500 ;
        RECT 104.700 282.600 105.900 289.950 ;
        RECT 74.100 276.000 75.900 279.600 ;
        RECT 77.100 276.600 78.900 279.600 ;
        RECT 80.100 276.000 81.900 279.600 ;
        RECT 98.100 276.600 99.900 279.600 ;
        RECT 101.100 276.000 102.900 282.600 ;
        RECT 104.100 276.600 105.900 282.600 ;
        RECT 119.400 282.600 120.300 289.950 ;
        RECT 121.950 288.150 123.750 289.950 ;
        RECT 128.100 288.150 129.900 289.950 ;
        RECT 143.100 288.150 144.900 289.950 ;
        RECT 149.100 288.150 150.900 289.950 ;
        RECT 152.100 286.200 153.000 289.950 ;
        RECT 170.250 288.150 172.050 289.950 ;
        RECT 119.400 281.400 124.500 282.600 ;
        RECT 119.700 276.000 121.500 279.600 ;
        RECT 122.700 276.600 124.500 281.400 ;
        RECT 127.200 276.000 129.000 282.600 ;
        RECT 143.100 276.000 144.900 285.600 ;
        RECT 149.700 285.000 153.000 286.200 ;
        RECT 149.700 276.600 151.500 285.000 ;
        RECT 173.100 284.700 174.300 289.950 ;
        RECT 176.100 288.150 177.900 289.950 ;
        RECT 173.100 283.800 177.300 284.700 ;
        RECT 170.400 276.000 172.200 282.600 ;
        RECT 175.500 276.600 177.300 283.800 ;
        RECT 197.100 279.600 198.300 289.950 ;
        RECT 212.100 288.150 213.900 289.950 ;
        RECT 218.100 288.150 219.900 289.950 ;
        RECT 221.100 286.200 222.000 289.950 ;
        RECT 239.250 288.150 241.050 289.950 ;
        RECT 194.100 276.000 195.900 279.600 ;
        RECT 197.100 276.600 198.900 279.600 ;
        RECT 212.100 276.000 213.900 285.600 ;
        RECT 218.700 285.000 222.000 286.200 ;
        RECT 218.700 276.600 220.500 285.000 ;
        RECT 242.100 284.700 243.300 289.950 ;
        RECT 245.100 288.150 246.900 289.950 ;
        RECT 260.100 288.150 261.900 289.950 ;
        RECT 263.100 285.600 264.300 289.950 ;
        RECT 266.100 288.150 267.900 289.950 ;
        RECT 260.700 284.700 264.300 285.600 ;
        RECT 242.100 283.800 246.300 284.700 ;
        RECT 239.400 276.000 241.200 282.600 ;
        RECT 244.500 276.600 246.300 283.800 ;
        RECT 260.700 282.600 261.900 284.700 ;
        RECT 260.100 276.600 261.900 282.600 ;
        RECT 263.100 281.700 270.900 283.050 ;
        RECT 263.100 276.600 264.900 281.700 ;
        RECT 266.100 276.000 267.900 280.800 ;
        RECT 269.100 276.600 270.900 281.700 ;
        RECT 272.550 282.600 273.450 297.300 ;
        RECT 282.450 297.000 284.250 297.300 ;
        RECT 274.950 289.950 277.050 292.050 ;
        RECT 284.100 290.400 286.200 292.050 ;
        RECT 274.950 287.400 276.750 289.950 ;
        RECT 278.100 289.200 286.200 290.400 ;
        RECT 278.100 288.600 279.900 289.200 ;
        RECT 281.100 287.400 282.900 288.000 ;
        RECT 274.950 286.200 282.900 287.400 ;
        RECT 292.950 286.200 293.850 298.800 ;
        RECT 296.550 296.100 298.650 296.700 ;
        RECT 302.550 296.100 304.350 296.550 ;
        RECT 296.550 294.900 304.350 296.100 ;
        RECT 296.550 294.600 298.650 294.900 ;
        RECT 302.550 294.750 304.350 294.900 ;
        RECT 305.250 292.050 306.450 299.400 ;
        RECT 320.100 292.050 321.900 293.850 ;
        RECT 326.700 292.050 327.900 299.400 ;
        RECT 331.950 294.450 334.050 295.050 ;
        RECT 337.950 294.450 340.050 295.050 ;
        RECT 331.950 293.550 340.050 294.450 ;
        RECT 331.950 292.950 334.050 293.550 ;
        RECT 337.950 292.950 340.050 293.550 ;
        RECT 347.700 292.050 348.900 305.400 ;
        RECT 353.550 299.400 355.350 311.400 ;
        RECT 356.550 299.400 358.350 312.000 ;
        RECT 361.350 305.400 363.150 311.400 ;
        RECT 365.850 305.400 367.650 312.000 ;
        RECT 361.350 303.300 363.450 305.400 ;
        RECT 368.850 304.500 370.650 311.400 ;
        RECT 371.850 305.400 373.650 312.000 ;
        RECT 367.950 303.450 374.550 304.500 ;
        RECT 367.950 302.700 369.750 303.450 ;
        RECT 372.750 302.700 374.550 303.450 ;
        RECT 376.650 302.400 378.450 311.400 ;
        RECT 360.450 300.600 363.450 302.400 ;
        RECT 364.350 301.800 366.150 302.400 ;
        RECT 364.350 300.900 370.050 301.800 ;
        RECT 376.650 301.500 378.750 302.400 ;
        RECT 364.350 300.600 366.150 300.900 ;
        RECT 362.250 299.700 363.450 300.600 ;
        RECT 353.550 292.050 354.750 299.400 ;
        RECT 362.250 298.800 367.050 299.700 ;
        RECT 355.650 296.100 357.450 296.550 ;
        RECT 361.350 296.100 363.450 296.700 ;
        RECT 355.650 294.900 363.450 296.100 ;
        RECT 355.650 294.750 357.450 294.900 ;
        RECT 361.350 294.600 363.450 294.900 ;
        RECT 301.950 291.750 306.450 292.050 ;
        RECT 300.150 289.950 306.450 291.750 ;
        RECT 319.950 289.950 322.050 292.050 ;
        RECT 322.950 289.950 325.050 292.050 ;
        RECT 325.950 289.950 328.050 292.050 ;
        RECT 328.950 289.950 331.050 292.050 ;
        RECT 343.950 289.950 346.050 292.050 ;
        RECT 346.950 289.950 349.050 292.050 ;
        RECT 349.950 289.950 352.050 292.050 ;
        RECT 353.550 291.750 358.050 292.050 ;
        RECT 353.550 289.950 359.850 291.750 ;
        RECT 281.850 285.000 293.850 286.200 ;
        RECT 281.850 283.200 282.900 285.000 ;
        RECT 292.050 284.400 293.850 285.000 ;
        RECT 272.550 280.800 274.950 282.600 ;
        RECT 273.150 276.600 274.950 280.800 ;
        RECT 276.150 276.000 277.950 282.600 ;
        RECT 278.850 280.200 280.950 281.700 ;
        RECT 281.850 281.400 283.650 283.200 ;
        RECT 305.250 282.600 306.450 289.950 ;
        RECT 323.100 288.150 324.900 289.950 ;
        RECT 326.700 285.600 327.900 289.950 ;
        RECT 329.100 288.150 330.900 289.950 ;
        RECT 344.100 288.150 345.900 289.950 ;
        RECT 326.700 284.700 330.300 285.600 ;
        RECT 347.700 284.700 348.900 289.950 ;
        RECT 349.950 288.150 351.750 289.950 ;
        RECT 284.850 281.550 286.650 282.300 ;
        RECT 284.850 280.500 289.800 281.550 ;
        RECT 278.850 279.600 282.750 280.200 ;
        RECT 288.750 279.600 289.800 280.500 ;
        RECT 296.250 279.600 298.650 281.700 ;
        RECT 279.150 278.700 282.750 279.600 ;
        RECT 280.950 276.600 282.750 278.700 ;
        RECT 285.450 276.000 287.250 279.600 ;
        RECT 288.750 276.600 290.550 279.600 ;
        RECT 291.750 276.000 293.550 279.600 ;
        RECT 296.250 276.600 298.050 279.600 ;
        RECT 301.350 276.000 303.150 282.600 ;
        RECT 304.650 276.600 306.450 282.600 ;
        RECT 320.100 281.700 327.900 283.050 ;
        RECT 320.100 276.600 321.900 281.700 ;
        RECT 323.100 276.000 324.900 280.800 ;
        RECT 326.100 276.600 327.900 281.700 ;
        RECT 329.100 282.600 330.300 284.700 ;
        RECT 344.700 283.800 348.900 284.700 ;
        RECT 329.100 276.600 330.900 282.600 ;
        RECT 344.700 276.600 346.500 283.800 ;
        RECT 353.550 282.600 354.750 289.950 ;
        RECT 366.150 286.200 367.050 298.800 ;
        RECT 369.150 298.800 370.050 300.900 ;
        RECT 370.950 300.300 378.750 301.500 ;
        RECT 370.950 299.700 372.750 300.300 ;
        RECT 382.050 299.400 383.850 312.000 ;
        RECT 385.050 301.200 386.850 311.400 ;
        RECT 390.150 301.200 391.950 311.400 ;
        RECT 385.050 299.400 387.450 301.200 ;
        RECT 369.150 298.500 377.550 298.800 ;
        RECT 386.550 298.500 387.450 299.400 ;
        RECT 369.150 297.900 387.450 298.500 ;
        RECT 375.750 297.300 387.450 297.900 ;
        RECT 375.750 297.000 377.550 297.300 ;
        RECT 373.800 290.400 375.900 292.050 ;
        RECT 373.800 289.200 381.900 290.400 ;
        RECT 382.950 289.950 385.050 292.050 ;
        RECT 380.100 288.600 381.900 289.200 ;
        RECT 377.100 287.400 378.900 288.000 ;
        RECT 383.250 287.400 385.050 289.950 ;
        RECT 377.100 286.200 385.050 287.400 ;
        RECT 366.150 285.000 378.150 286.200 ;
        RECT 366.150 284.400 367.950 285.000 ;
        RECT 377.100 283.200 378.150 285.000 ;
        RECT 349.800 276.000 351.600 282.600 ;
        RECT 353.550 276.600 355.350 282.600 ;
        RECT 356.850 276.000 358.650 282.600 ;
        RECT 361.350 279.600 363.750 281.700 ;
        RECT 373.350 281.550 375.150 282.300 ;
        RECT 370.200 280.500 375.150 281.550 ;
        RECT 376.350 281.400 378.150 283.200 ;
        RECT 386.550 282.600 387.450 297.300 ;
        RECT 370.200 279.600 371.250 280.500 ;
        RECT 379.050 280.200 381.150 281.700 ;
        RECT 377.250 279.600 381.150 280.200 ;
        RECT 361.950 276.600 363.750 279.600 ;
        RECT 366.450 276.000 368.250 279.600 ;
        RECT 369.450 276.600 371.250 279.600 ;
        RECT 372.750 276.000 374.550 279.600 ;
        RECT 377.250 278.700 380.850 279.600 ;
        RECT 377.250 276.600 379.050 278.700 ;
        RECT 382.050 276.000 383.850 282.600 ;
        RECT 385.050 280.800 387.450 282.600 ;
        RECT 389.550 299.400 391.950 301.200 ;
        RECT 393.150 299.400 394.950 312.000 ;
        RECT 398.550 302.400 400.350 311.400 ;
        RECT 403.350 305.400 405.150 312.000 ;
        RECT 406.350 304.500 408.150 311.400 ;
        RECT 409.350 305.400 411.150 312.000 ;
        RECT 413.850 305.400 415.650 311.400 ;
        RECT 402.450 303.450 409.050 304.500 ;
        RECT 402.450 302.700 404.250 303.450 ;
        RECT 407.250 302.700 409.050 303.450 ;
        RECT 413.550 303.300 415.650 305.400 ;
        RECT 398.250 301.500 400.350 302.400 ;
        RECT 410.850 301.800 412.650 302.400 ;
        RECT 398.250 300.300 406.050 301.500 ;
        RECT 404.250 299.700 406.050 300.300 ;
        RECT 406.950 300.900 412.650 301.800 ;
        RECT 389.550 298.500 390.450 299.400 ;
        RECT 406.950 298.800 407.850 300.900 ;
        RECT 410.850 300.600 412.650 300.900 ;
        RECT 413.550 300.600 416.550 302.400 ;
        RECT 413.550 299.700 414.750 300.600 ;
        RECT 399.450 298.500 407.850 298.800 ;
        RECT 389.550 297.900 407.850 298.500 ;
        RECT 409.950 298.800 414.750 299.700 ;
        RECT 418.650 299.400 420.450 312.000 ;
        RECT 421.650 299.400 423.450 311.400 ;
        RECT 437.700 305.400 439.500 312.000 ;
        RECT 438.000 302.100 439.800 303.900 ;
        RECT 440.700 300.900 442.500 311.400 ;
        RECT 389.550 297.300 401.250 297.900 ;
        RECT 389.550 282.600 390.450 297.300 ;
        RECT 399.450 297.000 401.250 297.300 ;
        RECT 391.950 289.950 394.050 292.050 ;
        RECT 401.100 290.400 403.200 292.050 ;
        RECT 391.950 287.400 393.750 289.950 ;
        RECT 395.100 289.200 403.200 290.400 ;
        RECT 395.100 288.600 396.900 289.200 ;
        RECT 398.100 287.400 399.900 288.000 ;
        RECT 391.950 286.200 399.900 287.400 ;
        RECT 409.950 286.200 410.850 298.800 ;
        RECT 413.550 296.100 415.650 296.700 ;
        RECT 419.550 296.100 421.350 296.550 ;
        RECT 413.550 294.900 421.350 296.100 ;
        RECT 413.550 294.600 415.650 294.900 ;
        RECT 419.550 294.750 421.350 294.900 ;
        RECT 422.250 292.050 423.450 299.400 ;
        RECT 440.100 299.400 442.500 300.900 ;
        RECT 445.800 299.400 447.600 312.000 ;
        RECT 461.100 305.400 462.900 311.400 ;
        RECT 464.100 305.400 465.900 312.000 ;
        RECT 479.700 305.400 481.500 312.000 ;
        RECT 440.100 292.050 441.300 299.400 ;
        RECT 446.100 292.050 447.900 293.850 ;
        RECT 461.700 292.050 462.900 305.400 ;
        RECT 480.000 302.100 481.800 303.900 ;
        RECT 482.700 300.900 484.500 311.400 ;
        RECT 482.100 299.400 484.500 300.900 ;
        RECT 487.800 299.400 489.600 312.000 ;
        RECT 503.100 305.400 504.900 311.400 ;
        RECT 506.100 305.400 507.900 312.000 ;
        RECT 474.000 294.450 478.050 295.050 ;
        RECT 464.100 292.050 465.900 293.850 ;
        RECT 473.550 292.950 478.050 294.450 ;
        RECT 418.950 291.750 423.450 292.050 ;
        RECT 417.150 289.950 423.450 291.750 ;
        RECT 436.950 289.950 439.050 292.050 ;
        RECT 439.950 289.950 442.050 292.050 ;
        RECT 442.950 289.950 445.050 292.050 ;
        RECT 445.950 289.950 448.050 292.050 ;
        RECT 460.950 289.950 463.050 292.050 ;
        RECT 463.950 289.950 466.050 292.050 ;
        RECT 398.850 285.000 410.850 286.200 ;
        RECT 398.850 283.200 399.900 285.000 ;
        RECT 409.050 284.400 410.850 285.000 ;
        RECT 389.550 280.800 391.950 282.600 ;
        RECT 385.050 276.600 386.850 280.800 ;
        RECT 390.150 276.600 391.950 280.800 ;
        RECT 393.150 276.000 394.950 282.600 ;
        RECT 395.850 280.200 397.950 281.700 ;
        RECT 398.850 281.400 400.650 283.200 ;
        RECT 422.250 282.600 423.450 289.950 ;
        RECT 437.100 288.150 438.900 289.950 ;
        RECT 440.100 285.600 441.300 289.950 ;
        RECT 443.100 288.150 444.900 289.950 ;
        RECT 437.700 284.700 441.300 285.600 ;
        RECT 437.700 282.600 438.900 284.700 ;
        RECT 401.850 281.550 403.650 282.300 ;
        RECT 401.850 280.500 406.800 281.550 ;
        RECT 395.850 279.600 399.750 280.200 ;
        RECT 405.750 279.600 406.800 280.500 ;
        RECT 413.250 279.600 415.650 281.700 ;
        RECT 396.150 278.700 399.750 279.600 ;
        RECT 397.950 276.600 399.750 278.700 ;
        RECT 402.450 276.000 404.250 279.600 ;
        RECT 405.750 276.600 407.550 279.600 ;
        RECT 408.750 276.000 410.550 279.600 ;
        RECT 413.250 276.600 415.050 279.600 ;
        RECT 418.350 276.000 420.150 282.600 ;
        RECT 421.650 276.600 423.450 282.600 ;
        RECT 437.100 276.600 438.900 282.600 ;
        RECT 440.100 281.700 447.900 283.050 ;
        RECT 440.100 276.600 441.900 281.700 ;
        RECT 443.100 276.000 444.900 280.800 ;
        RECT 446.100 276.600 447.900 281.700 ;
        RECT 461.700 279.600 462.900 289.950 ;
        RECT 466.950 288.450 469.050 289.050 ;
        RECT 473.550 288.450 474.450 292.950 ;
        RECT 482.100 292.050 483.300 299.400 ;
        RECT 488.100 292.050 489.900 293.850 ;
        RECT 503.700 292.050 504.900 305.400 ;
        RECT 509.550 299.400 511.350 311.400 ;
        RECT 512.550 299.400 514.350 312.000 ;
        RECT 517.350 305.400 519.150 311.400 ;
        RECT 521.850 305.400 523.650 312.000 ;
        RECT 517.350 303.300 519.450 305.400 ;
        RECT 524.850 304.500 526.650 311.400 ;
        RECT 527.850 305.400 529.650 312.000 ;
        RECT 523.950 303.450 530.550 304.500 ;
        RECT 523.950 302.700 525.750 303.450 ;
        RECT 528.750 302.700 530.550 303.450 ;
        RECT 532.650 302.400 534.450 311.400 ;
        RECT 516.450 300.600 519.450 302.400 ;
        RECT 520.350 301.800 522.150 302.400 ;
        RECT 520.350 300.900 526.050 301.800 ;
        RECT 532.650 301.500 534.750 302.400 ;
        RECT 520.350 300.600 522.150 300.900 ;
        RECT 518.250 299.700 519.450 300.600 ;
        RECT 506.100 292.050 507.900 293.850 ;
        RECT 509.550 292.050 510.750 299.400 ;
        RECT 518.250 298.800 523.050 299.700 ;
        RECT 511.650 296.100 513.450 296.550 ;
        RECT 517.350 296.100 519.450 296.700 ;
        RECT 511.650 294.900 519.450 296.100 ;
        RECT 511.650 294.750 513.450 294.900 ;
        RECT 517.350 294.600 519.450 294.900 ;
        RECT 478.950 289.950 481.050 292.050 ;
        RECT 481.950 289.950 484.050 292.050 ;
        RECT 484.950 289.950 487.050 292.050 ;
        RECT 487.950 289.950 490.050 292.050 ;
        RECT 502.950 289.950 505.050 292.050 ;
        RECT 505.950 289.950 508.050 292.050 ;
        RECT 509.550 291.750 514.050 292.050 ;
        RECT 509.550 289.950 515.850 291.750 ;
        RECT 466.950 287.550 474.450 288.450 ;
        RECT 479.100 288.150 480.900 289.950 ;
        RECT 466.950 286.950 469.050 287.550 ;
        RECT 482.100 285.600 483.300 289.950 ;
        RECT 485.100 288.150 486.900 289.950 ;
        RECT 479.700 284.700 483.300 285.600 ;
        RECT 479.700 282.600 480.900 284.700 ;
        RECT 461.100 276.600 462.900 279.600 ;
        RECT 464.100 276.000 465.900 279.600 ;
        RECT 479.100 276.600 480.900 282.600 ;
        RECT 482.100 281.700 489.900 283.050 ;
        RECT 482.100 276.600 483.900 281.700 ;
        RECT 485.100 276.000 486.900 280.800 ;
        RECT 488.100 276.600 489.900 281.700 ;
        RECT 503.700 279.600 504.900 289.950 ;
        RECT 509.550 282.600 510.750 289.950 ;
        RECT 522.150 286.200 523.050 298.800 ;
        RECT 525.150 298.800 526.050 300.900 ;
        RECT 526.950 300.300 534.750 301.500 ;
        RECT 526.950 299.700 528.750 300.300 ;
        RECT 538.050 299.400 539.850 312.000 ;
        RECT 541.050 301.200 542.850 311.400 ;
        RECT 560.100 305.400 561.900 312.000 ;
        RECT 563.100 305.400 564.900 311.400 ;
        RECT 541.050 299.400 543.450 301.200 ;
        RECT 525.150 298.500 533.550 298.800 ;
        RECT 542.550 298.500 543.450 299.400 ;
        RECT 525.150 297.900 543.450 298.500 ;
        RECT 531.750 297.300 543.450 297.900 ;
        RECT 531.750 297.000 533.550 297.300 ;
        RECT 529.800 290.400 531.900 292.050 ;
        RECT 529.800 289.200 537.900 290.400 ;
        RECT 538.950 289.950 541.050 292.050 ;
        RECT 536.100 288.600 537.900 289.200 ;
        RECT 533.100 287.400 534.900 288.000 ;
        RECT 539.250 287.400 541.050 289.950 ;
        RECT 533.100 286.200 541.050 287.400 ;
        RECT 522.150 285.000 534.150 286.200 ;
        RECT 522.150 284.400 523.950 285.000 ;
        RECT 533.100 283.200 534.150 285.000 ;
        RECT 503.100 276.600 504.900 279.600 ;
        RECT 506.100 276.000 507.900 279.600 ;
        RECT 509.550 276.600 511.350 282.600 ;
        RECT 512.850 276.000 514.650 282.600 ;
        RECT 517.350 279.600 519.750 281.700 ;
        RECT 529.350 281.550 531.150 282.300 ;
        RECT 526.200 280.500 531.150 281.550 ;
        RECT 532.350 281.400 534.150 283.200 ;
        RECT 542.550 282.600 543.450 297.300 ;
        RECT 560.100 292.050 561.900 293.850 ;
        RECT 563.100 292.050 564.300 305.400 ;
        RECT 566.550 299.400 568.350 311.400 ;
        RECT 569.550 299.400 571.350 312.000 ;
        RECT 574.350 305.400 576.150 311.400 ;
        RECT 578.850 305.400 580.650 312.000 ;
        RECT 574.350 303.300 576.450 305.400 ;
        RECT 581.850 304.500 583.650 311.400 ;
        RECT 584.850 305.400 586.650 312.000 ;
        RECT 580.950 303.450 587.550 304.500 ;
        RECT 580.950 302.700 582.750 303.450 ;
        RECT 585.750 302.700 587.550 303.450 ;
        RECT 589.650 302.400 591.450 311.400 ;
        RECT 573.450 300.600 576.450 302.400 ;
        RECT 577.350 301.800 579.150 302.400 ;
        RECT 577.350 300.900 583.050 301.800 ;
        RECT 589.650 301.500 591.750 302.400 ;
        RECT 577.350 300.600 579.150 300.900 ;
        RECT 575.250 299.700 576.450 300.600 ;
        RECT 566.550 292.050 567.750 299.400 ;
        RECT 575.250 298.800 580.050 299.700 ;
        RECT 568.650 296.100 570.450 296.550 ;
        RECT 574.350 296.100 576.450 296.700 ;
        RECT 568.650 294.900 576.450 296.100 ;
        RECT 568.650 294.750 570.450 294.900 ;
        RECT 574.350 294.600 576.450 294.900 ;
        RECT 559.950 289.950 562.050 292.050 ;
        RECT 562.950 289.950 565.050 292.050 ;
        RECT 566.550 291.750 571.050 292.050 ;
        RECT 566.550 289.950 572.850 291.750 ;
        RECT 544.950 285.450 547.050 286.050 ;
        RECT 559.950 285.450 562.050 285.750 ;
        RECT 544.950 284.550 562.050 285.450 ;
        RECT 544.950 283.950 547.050 284.550 ;
        RECT 559.950 283.650 562.050 284.550 ;
        RECT 526.200 279.600 527.250 280.500 ;
        RECT 535.050 280.200 537.150 281.700 ;
        RECT 533.250 279.600 537.150 280.200 ;
        RECT 517.950 276.600 519.750 279.600 ;
        RECT 522.450 276.000 524.250 279.600 ;
        RECT 525.450 276.600 527.250 279.600 ;
        RECT 528.750 276.000 530.550 279.600 ;
        RECT 533.250 278.700 536.850 279.600 ;
        RECT 533.250 276.600 535.050 278.700 ;
        RECT 538.050 276.000 539.850 282.600 ;
        RECT 541.050 280.800 543.450 282.600 ;
        RECT 541.050 276.600 542.850 280.800 ;
        RECT 563.100 279.600 564.300 289.950 ;
        RECT 566.550 282.600 567.750 289.950 ;
        RECT 579.150 286.200 580.050 298.800 ;
        RECT 582.150 298.800 583.050 300.900 ;
        RECT 583.950 300.300 591.750 301.500 ;
        RECT 583.950 299.700 585.750 300.300 ;
        RECT 595.050 299.400 596.850 312.000 ;
        RECT 598.050 301.200 599.850 311.400 ;
        RECT 598.050 299.400 600.450 301.200 ;
        RECT 614.100 300.600 615.900 311.400 ;
        RECT 617.100 301.500 618.900 312.000 ;
        RECT 620.100 310.500 627.900 311.400 ;
        RECT 620.100 300.600 621.900 310.500 ;
        RECT 614.100 299.700 621.900 300.600 ;
        RECT 582.150 298.500 590.550 298.800 ;
        RECT 599.550 298.500 600.450 299.400 ;
        RECT 623.100 298.500 624.900 309.600 ;
        RECT 626.100 299.400 627.900 310.500 ;
        RECT 641.100 299.400 642.900 312.000 ;
        RECT 645.600 299.400 648.900 311.400 ;
        RECT 651.600 299.400 653.400 312.000 ;
        RECT 671.100 300.300 672.900 311.400 ;
        RECT 674.100 301.200 675.900 312.000 ;
        RECT 677.100 300.300 678.900 311.400 ;
        RECT 671.100 299.400 678.900 300.300 ;
        RECT 680.100 299.400 681.900 311.400 ;
        RECT 696.000 300.600 697.800 311.400 ;
        RECT 696.000 299.400 699.600 300.600 ;
        RECT 701.100 299.400 702.900 312.000 ;
        RECT 719.400 299.400 721.200 312.000 ;
        RECT 724.500 300.900 726.300 311.400 ;
        RECT 727.500 305.400 729.300 312.000 ;
        RECT 727.200 302.100 729.000 303.900 ;
        RECT 724.500 299.400 726.900 300.900 ;
        RECT 582.150 297.900 600.450 298.500 ;
        RECT 588.750 297.300 600.450 297.900 ;
        RECT 616.950 297.450 619.050 298.050 ;
        RECT 588.750 297.000 590.550 297.300 ;
        RECT 586.800 290.400 588.900 292.050 ;
        RECT 586.800 289.200 594.900 290.400 ;
        RECT 595.950 289.950 598.050 292.050 ;
        RECT 593.100 288.600 594.900 289.200 ;
        RECT 590.100 287.400 591.900 288.000 ;
        RECT 596.250 287.400 598.050 289.950 ;
        RECT 590.100 286.200 598.050 287.400 ;
        RECT 579.150 285.000 591.150 286.200 ;
        RECT 579.150 284.400 580.950 285.000 ;
        RECT 590.100 283.200 591.150 285.000 ;
        RECT 560.100 276.000 561.900 279.600 ;
        RECT 563.100 276.600 564.900 279.600 ;
        RECT 566.550 276.600 568.350 282.600 ;
        RECT 569.850 276.000 571.650 282.600 ;
        RECT 574.350 279.600 576.750 281.700 ;
        RECT 586.350 281.550 588.150 282.300 ;
        RECT 583.200 280.500 588.150 281.550 ;
        RECT 589.350 281.400 591.150 283.200 ;
        RECT 599.550 282.600 600.450 297.300 ;
        RECT 611.550 296.550 619.050 297.450 ;
        RECT 611.550 294.450 612.450 296.550 ;
        RECT 616.950 295.950 619.050 296.550 ;
        RECT 620.100 297.600 624.900 298.500 ;
        RECT 608.550 293.550 612.450 294.450 ;
        RECT 608.550 285.450 609.450 293.550 ;
        RECT 617.250 292.050 619.050 293.850 ;
        RECT 620.100 292.050 621.000 297.600 ;
        RECT 625.950 297.450 628.050 298.050 ;
        RECT 631.950 297.450 634.050 298.050 ;
        RECT 625.950 296.550 634.050 297.450 ;
        RECT 625.950 295.950 628.050 296.550 ;
        RECT 631.950 295.950 634.050 296.550 ;
        RECT 623.100 292.050 624.900 293.850 ;
        RECT 641.100 292.050 642.900 293.850 ;
        RECT 646.950 292.050 648.000 299.400 ;
        RECT 649.950 297.450 652.050 298.050 ;
        RECT 658.950 297.450 661.050 298.050 ;
        RECT 649.950 296.550 661.050 297.450 ;
        RECT 649.950 295.950 652.050 296.550 ;
        RECT 658.950 295.950 661.050 296.550 ;
        RECT 652.950 292.050 654.750 293.850 ;
        RECT 674.250 292.050 676.050 293.850 ;
        RECT 680.700 292.050 681.600 299.400 ;
        RECT 685.950 295.950 688.050 298.050 ;
        RECT 613.950 289.950 616.050 292.050 ;
        RECT 616.950 289.950 619.050 292.050 ;
        RECT 619.950 289.950 622.050 292.050 ;
        RECT 622.950 289.950 625.050 292.050 ;
        RECT 625.950 289.950 628.050 292.050 ;
        RECT 640.950 289.950 643.050 292.050 ;
        RECT 643.950 289.950 646.050 292.050 ;
        RECT 614.250 288.150 616.050 289.950 ;
        RECT 616.950 285.450 619.050 286.050 ;
        RECT 608.550 284.550 619.050 285.450 ;
        RECT 616.950 283.950 619.050 284.550 ;
        RECT 620.100 282.600 621.300 289.950 ;
        RECT 626.100 288.150 627.900 289.950 ;
        RECT 644.250 288.150 646.050 289.950 ;
        RECT 646.950 289.950 649.050 292.050 ;
        RECT 649.950 289.950 652.050 292.050 ;
        RECT 652.950 289.950 655.050 292.050 ;
        RECT 670.950 289.950 673.050 292.050 ;
        RECT 673.950 289.950 676.050 292.050 ;
        RECT 676.950 289.950 679.050 292.050 ;
        RECT 679.950 289.950 682.050 292.050 ;
        RECT 646.950 285.300 648.000 289.950 ;
        RECT 649.950 288.150 651.750 289.950 ;
        RECT 671.100 288.150 672.900 289.950 ;
        RECT 677.250 288.150 679.050 289.950 ;
        RECT 646.950 284.100 651.300 285.300 ;
        RECT 583.200 279.600 584.250 280.500 ;
        RECT 592.050 280.200 594.150 281.700 ;
        RECT 590.250 279.600 594.150 280.200 ;
        RECT 574.950 276.600 576.750 279.600 ;
        RECT 579.450 276.000 581.250 279.600 ;
        RECT 582.450 276.600 584.250 279.600 ;
        RECT 585.750 276.000 587.550 279.600 ;
        RECT 590.250 278.700 593.850 279.600 ;
        RECT 590.250 276.600 592.050 278.700 ;
        RECT 595.050 276.000 596.850 282.600 ;
        RECT 598.050 280.800 600.450 282.600 ;
        RECT 598.050 276.600 599.850 280.800 ;
        RECT 614.700 276.000 616.500 282.600 ;
        RECT 619.200 276.600 621.000 282.600 ;
        RECT 623.700 276.000 625.500 282.600 ;
        RECT 641.100 282.000 648.900 282.900 ;
        RECT 650.400 282.600 651.300 284.100 ;
        RECT 680.700 282.600 681.600 289.950 ;
        RECT 686.550 286.050 687.450 295.950 ;
        RECT 695.100 292.050 696.900 293.850 ;
        RECT 698.700 292.050 699.600 299.400 ;
        RECT 703.950 294.450 708.000 295.050 ;
        RECT 700.950 292.050 702.750 293.850 ;
        RECT 703.950 292.950 708.450 294.450 ;
        RECT 694.950 289.950 697.050 292.050 ;
        RECT 697.950 289.950 700.050 292.050 ;
        RECT 700.950 289.950 703.050 292.050 ;
        RECT 684.000 285.900 687.450 286.050 ;
        RECT 682.950 284.550 687.450 285.900 ;
        RECT 682.950 283.950 687.000 284.550 ;
        RECT 682.950 283.800 685.050 283.950 ;
        RECT 641.100 276.600 642.900 282.000 ;
        RECT 644.100 276.000 645.900 281.100 ;
        RECT 647.100 277.500 648.900 282.000 ;
        RECT 650.100 278.400 651.900 282.600 ;
        RECT 653.100 277.500 654.900 282.600 ;
        RECT 647.100 276.600 654.900 277.500 ;
        RECT 672.000 276.000 673.800 282.600 ;
        RECT 676.500 281.400 681.600 282.600 ;
        RECT 676.500 276.600 678.300 281.400 ;
        RECT 698.700 279.600 699.600 289.950 ;
        RECT 707.550 289.050 708.450 292.950 ;
        RECT 719.100 292.050 720.900 293.850 ;
        RECT 725.700 292.050 726.900 299.400 ;
        RECT 727.950 300.450 730.050 301.050 ;
        RECT 736.950 300.450 739.050 301.050 ;
        RECT 727.950 299.550 739.050 300.450 ;
        RECT 727.950 298.950 730.050 299.550 ;
        RECT 736.950 298.950 739.050 299.550 ;
        RECT 743.100 299.400 744.900 311.400 ;
        RECT 746.100 299.400 747.900 312.000 ;
        RECT 761.100 305.400 762.900 311.400 ;
        RECT 764.100 305.400 765.900 312.000 ;
        RECT 782.100 305.400 783.900 312.000 ;
        RECT 785.100 305.400 786.900 311.400 ;
        RECT 788.100 305.400 789.900 312.000 ;
        RECT 730.950 294.450 733.050 295.050 ;
        RECT 736.950 294.450 739.050 294.900 ;
        RECT 730.950 293.550 739.050 294.450 ;
        RECT 730.950 292.950 733.050 293.550 ;
        RECT 736.950 292.800 739.050 293.550 ;
        RECT 743.700 292.050 744.900 299.400 ;
        RECT 745.950 297.450 748.050 298.050 ;
        RECT 745.950 296.550 756.450 297.450 ;
        RECT 745.950 295.950 748.050 296.550 ;
        RECT 748.950 294.450 753.000 295.050 ;
        RECT 748.950 292.950 753.450 294.450 ;
        RECT 718.950 289.950 721.050 292.050 ;
        RECT 721.950 289.950 724.050 292.050 ;
        RECT 724.950 289.950 727.050 292.050 ;
        RECT 727.950 289.950 730.050 292.050 ;
        RECT 742.950 289.950 745.050 292.050 ;
        RECT 745.950 289.950 748.050 292.050 ;
        RECT 703.950 287.550 708.450 289.050 ;
        RECT 722.100 288.150 723.900 289.950 ;
        RECT 703.950 286.950 708.000 287.550 ;
        RECT 725.700 285.600 726.900 289.950 ;
        RECT 728.100 288.150 729.900 289.950 ;
        RECT 725.700 284.700 729.300 285.600 ;
        RECT 719.100 281.700 726.900 283.050 ;
        RECT 679.500 276.000 681.300 279.600 ;
        RECT 695.100 276.000 696.900 279.600 ;
        RECT 698.100 276.600 699.900 279.600 ;
        RECT 701.100 276.000 702.900 279.600 ;
        RECT 719.100 276.600 720.900 281.700 ;
        RECT 722.100 276.000 723.900 280.800 ;
        RECT 725.100 276.600 726.900 281.700 ;
        RECT 728.100 282.600 729.300 284.700 ;
        RECT 743.700 282.600 744.900 289.950 ;
        RECT 746.100 288.150 747.900 289.950 ;
        RECT 752.550 289.050 753.450 292.950 ;
        RECT 748.950 287.550 753.450 289.050 ;
        RECT 748.950 286.950 753.000 287.550 ;
        RECT 745.950 285.450 748.050 286.050 ;
        RECT 755.550 285.450 756.450 296.550 ;
        RECT 761.700 292.050 762.900 305.400 ;
        RECT 764.100 292.050 765.900 293.850 ;
        RECT 785.700 292.050 786.900 305.400 ;
        RECT 803.400 299.400 805.200 312.000 ;
        RECT 808.500 300.900 810.300 311.400 ;
        RECT 811.500 305.400 813.300 312.000 ;
        RECT 811.200 302.100 813.000 303.900 ;
        RECT 808.500 299.400 810.900 300.900 ;
        RECT 827.100 299.400 828.900 311.400 ;
        RECT 830.100 300.000 831.900 312.000 ;
        RECT 833.100 305.400 834.900 311.400 ;
        RECT 836.100 305.400 837.900 312.000 ;
        RECT 803.100 292.050 804.900 293.850 ;
        RECT 809.700 292.050 810.900 299.400 ;
        RECT 827.700 292.050 828.600 299.400 ;
        RECT 831.000 292.050 832.800 293.850 ;
        RECT 760.950 289.950 763.050 292.050 ;
        RECT 763.950 289.950 766.050 292.050 ;
        RECT 781.950 289.950 784.050 292.050 ;
        RECT 784.950 289.950 787.050 292.050 ;
        RECT 787.950 289.950 790.050 292.050 ;
        RECT 802.950 289.950 805.050 292.050 ;
        RECT 805.950 289.950 808.050 292.050 ;
        RECT 808.950 289.950 811.050 292.050 ;
        RECT 811.950 289.950 814.050 292.050 ;
        RECT 827.100 289.950 829.200 292.050 ;
        RECT 830.400 289.950 832.500 292.050 ;
        RECT 745.950 284.550 756.450 285.450 ;
        RECT 745.950 283.950 748.050 284.550 ;
        RECT 728.100 276.600 729.900 282.600 ;
        RECT 743.100 276.600 744.900 282.600 ;
        RECT 746.100 276.000 747.900 282.600 ;
        RECT 761.700 279.600 762.900 289.950 ;
        RECT 782.100 288.150 783.900 289.950 ;
        RECT 785.700 284.700 786.900 289.950 ;
        RECT 787.950 288.150 789.750 289.950 ;
        RECT 806.100 288.150 807.900 289.950 ;
        RECT 809.700 285.600 810.900 289.950 ;
        RECT 812.100 288.150 813.900 289.950 ;
        RECT 809.700 284.700 813.300 285.600 ;
        RECT 782.700 283.800 786.900 284.700 ;
        RECT 761.100 276.600 762.900 279.600 ;
        RECT 764.100 276.000 765.900 279.600 ;
        RECT 782.700 276.600 784.500 283.800 ;
        RECT 787.800 276.000 789.600 282.600 ;
        RECT 803.100 281.700 810.900 283.050 ;
        RECT 803.100 276.600 804.900 281.700 ;
        RECT 806.100 276.000 807.900 280.800 ;
        RECT 809.100 276.600 810.900 281.700 ;
        RECT 812.100 282.600 813.300 284.700 ;
        RECT 827.700 282.600 828.600 289.950 ;
        RECT 834.000 285.300 834.900 305.400 ;
        RECT 851.100 299.400 852.900 312.000 ;
        RECT 856.200 300.600 858.000 311.400 ;
        RECT 875.100 305.400 876.900 312.000 ;
        RECT 878.100 305.400 879.900 311.400 ;
        RECT 881.100 305.400 882.900 312.000 ;
        RECT 896.100 305.400 897.900 312.000 ;
        RECT 899.100 305.400 900.900 311.400 ;
        RECT 854.400 299.400 858.000 300.600 ;
        RECT 851.250 292.050 853.050 293.850 ;
        RECT 854.400 292.050 855.300 299.400 ;
        RECT 857.100 292.050 858.900 293.850 ;
        RECT 878.100 292.050 879.300 305.400 ;
        RECT 835.800 289.950 837.900 292.050 ;
        RECT 850.950 289.950 853.050 292.050 ;
        RECT 853.950 289.950 856.050 292.050 ;
        RECT 856.950 289.950 859.050 292.050 ;
        RECT 874.950 289.950 877.050 292.050 ;
        RECT 877.950 289.950 880.050 292.050 ;
        RECT 880.950 289.950 883.050 292.050 ;
        RECT 896.100 289.950 898.200 292.050 ;
        RECT 835.950 288.150 837.750 289.950 ;
        RECT 838.950 285.450 841.050 286.050 ;
        RECT 850.950 285.450 853.050 286.050 ;
        RECT 829.500 284.400 837.900 285.300 ;
        RECT 829.500 283.500 831.300 284.400 ;
        RECT 812.100 276.600 813.900 282.600 ;
        RECT 827.700 280.800 830.400 282.600 ;
        RECT 828.600 276.600 830.400 280.800 ;
        RECT 831.600 276.000 833.400 282.600 ;
        RECT 836.100 276.600 837.900 284.400 ;
        RECT 838.950 284.550 853.050 285.450 ;
        RECT 838.950 283.950 841.050 284.550 ;
        RECT 850.950 283.950 853.050 284.550 ;
        RECT 854.400 279.600 855.300 289.950 ;
        RECT 875.250 288.150 877.050 289.950 ;
        RECT 856.950 285.450 859.050 285.750 ;
        RECT 865.950 285.450 868.050 286.050 ;
        RECT 856.950 284.550 868.050 285.450 ;
        RECT 856.950 283.650 859.050 284.550 ;
        RECT 865.950 283.950 868.050 284.550 ;
        RECT 878.100 284.700 879.300 289.950 ;
        RECT 881.100 288.150 882.900 289.950 ;
        RECT 896.250 288.150 898.050 289.950 ;
        RECT 899.100 285.300 900.000 305.400 ;
        RECT 902.100 300.000 903.900 312.000 ;
        RECT 905.100 299.400 906.900 311.400 ;
        RECT 923.400 299.400 925.200 312.000 ;
        RECT 928.500 300.900 930.300 311.400 ;
        RECT 931.500 305.400 933.300 312.000 ;
        RECT 931.200 302.100 933.000 303.900 ;
        RECT 928.500 299.400 930.900 300.900 ;
        RECT 950.100 300.300 951.900 311.400 ;
        RECT 953.100 301.200 954.900 312.000 ;
        RECT 956.100 300.300 957.900 311.400 ;
        RECT 950.100 299.400 957.900 300.300 ;
        RECT 959.100 299.400 960.900 311.400 ;
        RECT 974.100 305.400 975.900 311.400 ;
        RECT 977.100 305.400 978.900 312.000 ;
        RECT 979.950 309.450 982.050 310.050 ;
        RECT 985.950 309.450 988.050 310.050 ;
        RECT 979.950 308.550 988.050 309.450 ;
        RECT 979.950 307.950 982.050 308.550 ;
        RECT 985.950 307.950 988.050 308.550 ;
        RECT 992.100 305.400 993.900 312.000 ;
        RECT 995.100 305.400 996.900 311.400 ;
        RECT 998.100 306.000 999.900 312.000 ;
        RECT 901.200 292.050 903.000 293.850 ;
        RECT 905.400 292.050 906.300 299.400 ;
        RECT 923.100 292.050 924.900 293.850 ;
        RECT 929.700 292.050 930.900 299.400 ;
        RECT 953.250 292.050 955.050 293.850 ;
        RECT 959.700 292.050 960.600 299.400 ;
        RECT 974.700 292.050 975.900 305.400 ;
        RECT 995.400 305.100 996.900 305.400 ;
        RECT 1001.100 305.400 1002.900 311.400 ;
        RECT 1001.100 305.100 1002.000 305.400 ;
        RECT 995.400 304.200 1002.000 305.100 ;
        RECT 982.950 300.450 985.050 301.050 ;
        RECT 997.950 300.450 1000.050 301.050 ;
        RECT 982.950 299.550 1000.050 300.450 ;
        RECT 982.950 298.950 985.050 299.550 ;
        RECT 997.950 298.950 1000.050 299.550 ;
        RECT 977.100 292.050 978.900 293.850 ;
        RECT 995.100 292.050 996.900 293.850 ;
        RECT 1001.100 292.050 1002.000 304.200 ;
        RECT 1003.950 294.450 1008.000 295.050 ;
        RECT 1003.950 292.950 1008.450 294.450 ;
        RECT 901.500 289.950 903.600 292.050 ;
        RECT 904.800 289.950 906.900 292.050 ;
        RECT 922.950 289.950 925.050 292.050 ;
        RECT 925.950 289.950 928.050 292.050 ;
        RECT 928.950 289.950 931.050 292.050 ;
        RECT 931.950 289.950 934.050 292.050 ;
        RECT 949.950 289.950 952.050 292.050 ;
        RECT 952.950 289.950 955.050 292.050 ;
        RECT 955.950 289.950 958.050 292.050 ;
        RECT 958.950 289.950 961.050 292.050 ;
        RECT 973.950 289.950 976.050 292.050 ;
        RECT 976.950 289.950 979.050 292.050 ;
        RECT 991.950 289.950 994.050 292.050 ;
        RECT 994.950 289.950 997.050 292.050 ;
        RECT 997.950 289.950 1000.050 292.050 ;
        RECT 1000.950 289.950 1003.050 292.050 ;
        RECT 878.100 283.800 882.300 284.700 ;
        RECT 851.100 276.000 852.900 279.600 ;
        RECT 854.100 276.600 855.900 279.600 ;
        RECT 857.100 276.000 858.900 279.600 ;
        RECT 875.400 276.000 877.200 282.600 ;
        RECT 880.500 276.600 882.300 283.800 ;
        RECT 896.100 284.400 904.500 285.300 ;
        RECT 896.100 276.600 897.900 284.400 ;
        RECT 902.700 283.500 904.500 284.400 ;
        RECT 905.400 282.600 906.300 289.950 ;
        RECT 926.100 288.150 927.900 289.950 ;
        RECT 929.700 285.600 930.900 289.950 ;
        RECT 932.100 288.150 933.900 289.950 ;
        RECT 950.100 288.150 951.900 289.950 ;
        RECT 956.250 288.150 958.050 289.950 ;
        RECT 929.700 284.700 933.300 285.600 ;
        RECT 900.600 276.000 902.400 282.600 ;
        RECT 903.600 280.800 906.300 282.600 ;
        RECT 923.100 281.700 930.900 283.050 ;
        RECT 903.600 276.600 905.400 280.800 ;
        RECT 923.100 276.600 924.900 281.700 ;
        RECT 926.100 276.000 927.900 280.800 ;
        RECT 929.100 276.600 930.900 281.700 ;
        RECT 932.100 282.600 933.300 284.700 ;
        RECT 937.950 285.450 940.050 286.050 ;
        RECT 955.950 285.450 958.050 286.050 ;
        RECT 937.950 284.550 958.050 285.450 ;
        RECT 937.950 283.950 940.050 284.550 ;
        RECT 955.950 283.950 958.050 284.550 ;
        RECT 959.700 282.600 960.600 289.950 ;
        RECT 932.100 276.600 933.900 282.600 ;
        RECT 951.000 276.000 952.800 282.600 ;
        RECT 955.500 281.400 960.600 282.600 ;
        RECT 955.500 276.600 957.300 281.400 ;
        RECT 974.700 279.600 975.900 289.950 ;
        RECT 992.100 288.150 993.900 289.950 ;
        RECT 998.100 288.150 999.900 289.950 ;
        RECT 1001.100 286.200 1002.000 289.950 ;
        RECT 1007.550 289.050 1008.450 292.950 ;
        RECT 1003.950 287.550 1008.450 289.050 ;
        RECT 1003.950 286.950 1008.000 287.550 ;
        RECT 958.500 276.000 960.300 279.600 ;
        RECT 974.100 276.600 975.900 279.600 ;
        RECT 977.100 276.000 978.900 279.600 ;
        RECT 992.100 276.000 993.900 285.600 ;
        RECT 998.700 285.000 1002.000 286.200 ;
        RECT 998.700 276.600 1000.500 285.000 ;
        RECT 14.100 266.400 15.900 272.400 ;
        RECT 17.100 266.400 18.900 273.000 ;
        RECT 20.100 269.400 21.900 272.400 ;
        RECT 14.100 259.050 15.300 266.400 ;
        RECT 20.700 265.500 21.900 269.400 ;
        RECT 38.100 266.400 39.900 272.400 ;
        RECT 16.200 264.600 21.900 265.500 ;
        RECT 16.200 263.700 18.000 264.600 ;
        RECT 14.100 256.950 16.200 259.050 ;
        RECT 14.100 249.600 15.300 256.950 ;
        RECT 17.100 252.300 18.000 263.700 ;
        RECT 38.700 264.300 39.900 266.400 ;
        RECT 41.100 267.300 42.900 272.400 ;
        RECT 44.100 268.200 45.900 273.000 ;
        RECT 47.100 267.300 48.900 272.400 ;
        RECT 51.150 268.200 52.950 272.400 ;
        RECT 41.100 265.950 48.900 267.300 ;
        RECT 50.550 266.400 52.950 268.200 ;
        RECT 54.150 266.400 55.950 273.000 ;
        RECT 58.950 270.300 60.750 272.400 ;
        RECT 57.150 269.400 60.750 270.300 ;
        RECT 63.450 269.400 65.250 273.000 ;
        RECT 66.750 269.400 68.550 272.400 ;
        RECT 69.750 269.400 71.550 273.000 ;
        RECT 74.250 269.400 76.050 272.400 ;
        RECT 56.850 268.800 60.750 269.400 ;
        RECT 56.850 267.300 58.950 268.800 ;
        RECT 66.750 268.500 67.800 269.400 ;
        RECT 38.700 263.400 42.300 264.300 ;
        RECT 38.100 259.050 39.900 260.850 ;
        RECT 41.100 259.050 42.300 263.400 ;
        RECT 44.100 259.050 45.900 260.850 ;
        RECT 19.500 256.950 21.600 259.050 ;
        RECT 37.950 256.950 40.050 259.050 ;
        RECT 40.950 256.950 43.050 259.050 ;
        RECT 43.950 256.950 46.050 259.050 ;
        RECT 46.950 256.950 49.050 259.050 ;
        RECT 19.800 255.150 21.600 256.950 ;
        RECT 16.200 251.400 18.000 252.300 ;
        RECT 16.200 250.500 21.900 251.400 ;
        RECT 14.100 237.600 15.900 249.600 ;
        RECT 17.100 237.000 18.900 247.800 ;
        RECT 20.700 243.600 21.900 250.500 ;
        RECT 41.100 249.600 42.300 256.950 ;
        RECT 47.100 255.150 48.900 256.950 ;
        RECT 50.550 251.700 51.450 266.400 ;
        RECT 59.850 265.800 61.650 267.600 ;
        RECT 62.850 267.450 67.800 268.500 ;
        RECT 62.850 266.700 64.650 267.450 ;
        RECT 74.250 267.300 76.650 269.400 ;
        RECT 79.350 266.400 81.150 273.000 ;
        RECT 82.650 266.400 84.450 272.400 ;
        RECT 59.850 264.000 60.900 265.800 ;
        RECT 70.050 264.000 71.850 264.600 ;
        RECT 59.850 262.800 71.850 264.000 ;
        RECT 52.950 261.600 60.900 262.800 ;
        RECT 52.950 259.050 54.750 261.600 ;
        RECT 59.100 261.000 60.900 261.600 ;
        RECT 56.100 259.800 57.900 260.400 ;
        RECT 52.950 256.950 55.050 259.050 ;
        RECT 56.100 258.600 64.200 259.800 ;
        RECT 62.100 256.950 64.200 258.600 ;
        RECT 60.450 251.700 62.250 252.000 ;
        RECT 50.550 251.100 62.250 251.700 ;
        RECT 50.550 250.500 68.850 251.100 ;
        RECT 50.550 249.600 51.450 250.500 ;
        RECT 60.450 250.200 68.850 250.500 ;
        RECT 41.100 248.100 43.500 249.600 ;
        RECT 39.000 245.100 40.800 246.900 ;
        RECT 20.100 237.600 21.900 243.600 ;
        RECT 38.700 237.000 40.500 243.600 ;
        RECT 41.700 237.600 43.500 248.100 ;
        RECT 46.800 237.000 48.600 249.600 ;
        RECT 50.550 247.800 52.950 249.600 ;
        RECT 51.150 237.600 52.950 247.800 ;
        RECT 54.150 237.000 55.950 249.600 ;
        RECT 65.250 248.700 67.050 249.300 ;
        RECT 59.250 247.500 67.050 248.700 ;
        RECT 67.950 248.100 68.850 250.200 ;
        RECT 70.950 250.200 71.850 262.800 ;
        RECT 83.250 259.050 84.450 266.400 ;
        RECT 98.100 267.300 99.900 272.400 ;
        RECT 101.100 268.200 102.900 273.000 ;
        RECT 104.100 267.300 105.900 272.400 ;
        RECT 98.100 265.950 105.900 267.300 ;
        RECT 107.100 266.400 108.900 272.400 ;
        RECT 107.100 264.300 108.300 266.400 ;
        RECT 104.700 263.400 108.300 264.300 ;
        RECT 124.500 264.000 126.300 272.400 ;
        RECT 101.100 259.050 102.900 260.850 ;
        RECT 104.700 259.050 105.900 263.400 ;
        RECT 123.000 262.800 126.300 264.000 ;
        RECT 131.100 263.400 132.900 273.000 ;
        RECT 146.700 265.200 148.500 272.400 ;
        RECT 151.800 266.400 153.600 273.000 ;
        RECT 167.100 266.400 168.900 272.400 ;
        RECT 170.100 266.400 171.900 273.000 ;
        RECT 173.100 269.400 174.900 272.400 ;
        RECT 191.100 269.400 192.900 273.000 ;
        RECT 194.100 269.400 195.900 272.400 ;
        RECT 146.700 264.300 150.900 265.200 ;
        RECT 107.100 259.050 108.900 260.850 ;
        RECT 123.000 259.050 123.900 262.800 ;
        RECT 125.100 259.050 126.900 260.850 ;
        RECT 131.100 259.050 132.900 260.850 ;
        RECT 146.100 259.050 147.900 260.850 ;
        RECT 149.700 259.050 150.900 264.300 ;
        RECT 151.950 259.050 153.750 260.850 ;
        RECT 167.100 259.050 168.300 266.400 ;
        RECT 173.700 265.500 174.900 269.400 ;
        RECT 169.200 264.600 174.900 265.500 ;
        RECT 169.200 263.700 171.000 264.600 ;
        RECT 78.150 257.250 84.450 259.050 ;
        RECT 79.950 256.950 84.450 257.250 ;
        RECT 97.950 256.950 100.050 259.050 ;
        RECT 100.950 256.950 103.050 259.050 ;
        RECT 103.950 256.950 106.050 259.050 ;
        RECT 106.950 256.950 109.050 259.050 ;
        RECT 121.950 256.950 124.050 259.050 ;
        RECT 124.950 256.950 127.050 259.050 ;
        RECT 127.950 256.950 130.050 259.050 ;
        RECT 130.950 256.950 133.050 259.050 ;
        RECT 145.950 256.950 148.050 259.050 ;
        RECT 148.950 256.950 151.050 259.050 ;
        RECT 151.950 256.950 154.050 259.050 ;
        RECT 167.100 256.950 169.200 259.050 ;
        RECT 74.550 254.100 76.650 254.400 ;
        RECT 80.550 254.100 82.350 254.250 ;
        RECT 74.550 252.900 82.350 254.100 ;
        RECT 74.550 252.300 76.650 252.900 ;
        RECT 80.550 252.450 82.350 252.900 ;
        RECT 70.950 249.300 75.750 250.200 ;
        RECT 83.250 249.600 84.450 256.950 ;
        RECT 98.100 255.150 99.900 256.950 ;
        RECT 104.700 249.600 105.900 256.950 ;
        RECT 74.550 248.400 75.750 249.300 ;
        RECT 71.850 248.100 73.650 248.400 ;
        RECT 59.250 246.600 61.350 247.500 ;
        RECT 67.950 247.200 73.650 248.100 ;
        RECT 71.850 246.600 73.650 247.200 ;
        RECT 74.550 246.600 77.550 248.400 ;
        RECT 59.550 237.600 61.350 246.600 ;
        RECT 63.450 245.550 65.250 246.300 ;
        RECT 68.250 245.550 70.050 246.300 ;
        RECT 63.450 244.500 70.050 245.550 ;
        RECT 64.350 237.000 66.150 243.600 ;
        RECT 67.350 237.600 69.150 244.500 ;
        RECT 74.550 243.600 76.650 245.700 ;
        RECT 70.350 237.000 72.150 243.600 ;
        RECT 74.850 237.600 76.650 243.600 ;
        RECT 79.650 237.000 81.450 249.600 ;
        RECT 82.650 237.600 84.450 249.600 ;
        RECT 98.400 237.000 100.200 249.600 ;
        RECT 103.500 248.100 105.900 249.600 ;
        RECT 103.500 237.600 105.300 248.100 ;
        RECT 106.200 245.100 108.000 246.900 ;
        RECT 123.000 244.800 123.900 256.950 ;
        RECT 128.100 255.150 129.900 256.950 ;
        RECT 124.950 252.450 127.050 253.050 ;
        RECT 133.950 252.450 136.050 253.050 ;
        RECT 124.950 251.550 136.050 252.450 ;
        RECT 124.950 250.950 127.050 251.550 ;
        RECT 133.950 250.950 136.050 251.550 ;
        RECT 123.000 243.900 129.600 244.800 ;
        RECT 123.000 243.600 123.900 243.900 ;
        RECT 106.500 237.000 108.300 243.600 ;
        RECT 122.100 237.600 123.900 243.600 ;
        RECT 128.100 243.600 129.600 243.900 ;
        RECT 149.700 243.600 150.900 256.950 ;
        RECT 167.100 249.600 168.300 256.950 ;
        RECT 170.100 252.300 171.000 263.700 ;
        RECT 194.100 259.050 195.300 269.400 ;
        RECT 209.100 267.300 210.900 272.400 ;
        RECT 212.100 268.200 213.900 273.000 ;
        RECT 215.100 267.300 216.900 272.400 ;
        RECT 209.100 265.950 216.900 267.300 ;
        RECT 218.100 266.400 219.900 272.400 ;
        RECT 233.100 269.400 234.900 272.400 ;
        RECT 236.100 269.400 237.900 273.000 ;
        RECT 251.100 269.400 252.900 273.000 ;
        RECT 254.100 269.400 255.900 272.400 ;
        RECT 218.100 264.300 219.300 266.400 ;
        RECT 215.700 263.400 219.300 264.300 ;
        RECT 212.100 259.050 213.900 260.850 ;
        RECT 215.700 259.050 216.900 263.400 ;
        RECT 218.100 259.050 219.900 260.850 ;
        RECT 233.700 259.050 234.900 269.400 ;
        RECT 254.100 259.050 255.300 269.400 ;
        RECT 269.700 265.200 271.500 272.400 ;
        RECT 274.800 266.400 276.600 273.000 ;
        RECT 293.100 267.300 294.900 272.400 ;
        RECT 296.100 268.200 297.900 273.000 ;
        RECT 299.100 267.300 300.900 272.400 ;
        RECT 293.100 265.950 300.900 267.300 ;
        RECT 302.100 266.400 303.900 272.400 ;
        RECT 306.150 268.200 307.950 272.400 ;
        RECT 305.550 266.400 307.950 268.200 ;
        RECT 309.150 266.400 310.950 273.000 ;
        RECT 313.950 270.300 315.750 272.400 ;
        RECT 312.150 269.400 315.750 270.300 ;
        RECT 318.450 269.400 320.250 273.000 ;
        RECT 321.750 269.400 323.550 272.400 ;
        RECT 324.750 269.400 326.550 273.000 ;
        RECT 329.250 269.400 331.050 272.400 ;
        RECT 311.850 268.800 315.750 269.400 ;
        RECT 311.850 267.300 313.950 268.800 ;
        RECT 321.750 268.500 322.800 269.400 ;
        RECT 269.700 264.300 273.900 265.200 ;
        RECT 302.100 264.300 303.300 266.400 ;
        RECT 269.100 259.050 270.900 260.850 ;
        RECT 272.700 259.050 273.900 264.300 ;
        RECT 299.700 263.400 303.300 264.300 ;
        RECT 274.950 259.050 276.750 260.850 ;
        RECT 296.100 259.050 297.900 260.850 ;
        RECT 299.700 259.050 300.900 263.400 ;
        RECT 302.100 259.050 303.900 260.850 ;
        RECT 172.500 256.950 174.600 259.050 ;
        RECT 190.950 256.950 193.050 259.050 ;
        RECT 193.950 256.950 196.050 259.050 ;
        RECT 208.950 256.950 211.050 259.050 ;
        RECT 211.950 256.950 214.050 259.050 ;
        RECT 214.950 256.950 217.050 259.050 ;
        RECT 217.950 256.950 220.050 259.050 ;
        RECT 232.950 256.950 235.050 259.050 ;
        RECT 235.950 256.950 238.050 259.050 ;
        RECT 250.950 256.950 253.050 259.050 ;
        RECT 253.950 256.950 256.050 259.050 ;
        RECT 268.950 256.950 271.050 259.050 ;
        RECT 271.950 256.950 274.050 259.050 ;
        RECT 274.950 256.950 277.050 259.050 ;
        RECT 292.950 256.950 295.050 259.050 ;
        RECT 295.950 256.950 298.050 259.050 ;
        RECT 298.950 256.950 301.050 259.050 ;
        RECT 301.950 256.950 304.050 259.050 ;
        RECT 172.800 255.150 174.600 256.950 ;
        RECT 191.100 255.150 192.900 256.950 ;
        RECT 169.200 251.400 171.000 252.300 ;
        RECT 169.200 250.500 174.900 251.400 ;
        RECT 125.100 237.000 126.900 243.000 ;
        RECT 128.100 237.600 129.900 243.600 ;
        RECT 131.100 237.000 132.900 243.600 ;
        RECT 146.100 237.000 147.900 243.600 ;
        RECT 149.100 237.600 150.900 243.600 ;
        RECT 152.100 237.000 153.900 243.600 ;
        RECT 167.100 237.600 168.900 249.600 ;
        RECT 170.100 237.000 171.900 247.800 ;
        RECT 173.700 243.600 174.900 250.500 ;
        RECT 194.100 243.600 195.300 256.950 ;
        RECT 209.100 255.150 210.900 256.950 ;
        RECT 215.700 249.600 216.900 256.950 ;
        RECT 173.100 237.600 174.900 243.600 ;
        RECT 191.100 237.000 192.900 243.600 ;
        RECT 194.100 237.600 195.900 243.600 ;
        RECT 209.400 237.000 211.200 249.600 ;
        RECT 214.500 248.100 216.900 249.600 ;
        RECT 214.500 237.600 216.300 248.100 ;
        RECT 217.200 245.100 219.000 246.900 ;
        RECT 233.700 243.600 234.900 256.950 ;
        RECT 236.100 255.150 237.900 256.950 ;
        RECT 251.100 255.150 252.900 256.950 ;
        RECT 254.100 243.600 255.300 256.950 ;
        RECT 272.700 243.600 273.900 256.950 ;
        RECT 293.100 255.150 294.900 256.950 ;
        RECT 299.700 249.600 300.900 256.950 ;
        RECT 217.500 237.000 219.300 243.600 ;
        RECT 233.100 237.600 234.900 243.600 ;
        RECT 236.100 237.000 237.900 243.600 ;
        RECT 251.100 237.000 252.900 243.600 ;
        RECT 254.100 237.600 255.900 243.600 ;
        RECT 269.100 237.000 270.900 243.600 ;
        RECT 272.100 237.600 273.900 243.600 ;
        RECT 275.100 237.000 276.900 243.600 ;
        RECT 293.400 237.000 295.200 249.600 ;
        RECT 298.500 248.100 300.900 249.600 ;
        RECT 305.550 251.700 306.450 266.400 ;
        RECT 314.850 265.800 316.650 267.600 ;
        RECT 317.850 267.450 322.800 268.500 ;
        RECT 317.850 266.700 319.650 267.450 ;
        RECT 329.250 267.300 331.650 269.400 ;
        RECT 334.350 266.400 336.150 273.000 ;
        RECT 337.650 266.400 339.450 272.400 ;
        RECT 356.400 266.400 358.200 273.000 ;
        RECT 314.850 264.000 315.900 265.800 ;
        RECT 325.050 264.000 326.850 264.600 ;
        RECT 314.850 262.800 326.850 264.000 ;
        RECT 307.950 261.600 315.900 262.800 ;
        RECT 307.950 259.050 309.750 261.600 ;
        RECT 314.100 261.000 315.900 261.600 ;
        RECT 311.100 259.800 312.900 260.400 ;
        RECT 307.950 256.950 310.050 259.050 ;
        RECT 311.100 258.600 319.200 259.800 ;
        RECT 317.100 256.950 319.200 258.600 ;
        RECT 315.450 251.700 317.250 252.000 ;
        RECT 305.550 251.100 317.250 251.700 ;
        RECT 305.550 250.500 323.850 251.100 ;
        RECT 305.550 249.600 306.450 250.500 ;
        RECT 315.450 250.200 323.850 250.500 ;
        RECT 298.500 237.600 300.300 248.100 ;
        RECT 305.550 247.800 307.950 249.600 ;
        RECT 301.200 245.100 303.000 246.900 ;
        RECT 301.500 237.000 303.300 243.600 ;
        RECT 306.150 237.600 307.950 247.800 ;
        RECT 309.150 237.000 310.950 249.600 ;
        RECT 320.250 248.700 322.050 249.300 ;
        RECT 314.250 247.500 322.050 248.700 ;
        RECT 322.950 248.100 323.850 250.200 ;
        RECT 325.950 250.200 326.850 262.800 ;
        RECT 338.250 259.050 339.450 266.400 ;
        RECT 361.500 265.200 363.300 272.400 ;
        RECT 359.100 264.300 363.300 265.200 ;
        RECT 380.700 265.200 382.500 272.400 ;
        RECT 385.800 266.400 387.600 273.000 ;
        RECT 401.400 266.400 403.200 273.000 ;
        RECT 406.500 265.200 408.300 272.400 ;
        RECT 425.100 266.400 426.900 272.400 ;
        RECT 380.700 264.300 384.900 265.200 ;
        RECT 356.250 259.050 358.050 260.850 ;
        RECT 359.100 259.050 360.300 264.300 ;
        RECT 362.100 259.050 363.900 260.850 ;
        RECT 380.100 259.050 381.900 260.850 ;
        RECT 383.700 259.050 384.900 264.300 ;
        RECT 404.100 264.300 408.300 265.200 ;
        RECT 425.700 264.300 426.900 266.400 ;
        RECT 428.100 267.300 429.900 272.400 ;
        RECT 431.100 268.200 432.900 273.000 ;
        RECT 434.100 267.300 435.900 272.400 ;
        RECT 428.100 265.950 435.900 267.300 ;
        RECT 449.700 265.200 451.500 272.400 ;
        RECT 454.800 266.400 456.600 273.000 ;
        RECT 459.150 268.200 460.950 272.400 ;
        RECT 458.550 266.400 460.950 268.200 ;
        RECT 462.150 266.400 463.950 273.000 ;
        RECT 466.950 270.300 468.750 272.400 ;
        RECT 465.150 269.400 468.750 270.300 ;
        RECT 471.450 269.400 473.250 273.000 ;
        RECT 474.750 269.400 476.550 272.400 ;
        RECT 477.750 269.400 479.550 273.000 ;
        RECT 482.250 269.400 484.050 272.400 ;
        RECT 464.850 268.800 468.750 269.400 ;
        RECT 464.850 267.300 466.950 268.800 ;
        RECT 474.750 268.500 475.800 269.400 ;
        RECT 449.700 264.300 453.900 265.200 ;
        RECT 385.950 259.050 387.750 260.850 ;
        RECT 401.250 259.050 403.050 260.850 ;
        RECT 404.100 259.050 405.300 264.300 ;
        RECT 425.700 263.400 429.300 264.300 ;
        RECT 420.000 261.450 424.050 262.050 ;
        RECT 407.100 259.050 408.900 260.850 ;
        RECT 419.550 259.950 424.050 261.450 ;
        RECT 333.150 257.250 339.450 259.050 ;
        RECT 334.950 256.950 339.450 257.250 ;
        RECT 355.950 256.950 358.050 259.050 ;
        RECT 358.950 256.950 361.050 259.050 ;
        RECT 361.950 256.950 364.050 259.050 ;
        RECT 379.950 256.950 382.050 259.050 ;
        RECT 382.950 256.950 385.050 259.050 ;
        RECT 385.950 256.950 388.050 259.050 ;
        RECT 400.950 256.950 403.050 259.050 ;
        RECT 403.950 256.950 406.050 259.050 ;
        RECT 406.950 256.950 409.050 259.050 ;
        RECT 329.550 254.100 331.650 254.400 ;
        RECT 335.550 254.100 337.350 254.250 ;
        RECT 329.550 252.900 337.350 254.100 ;
        RECT 329.550 252.300 331.650 252.900 ;
        RECT 335.550 252.450 337.350 252.900 ;
        RECT 325.950 249.300 330.750 250.200 ;
        RECT 338.250 249.600 339.450 256.950 ;
        RECT 329.550 248.400 330.750 249.300 ;
        RECT 326.850 248.100 328.650 248.400 ;
        RECT 314.250 246.600 316.350 247.500 ;
        RECT 322.950 247.200 328.650 248.100 ;
        RECT 326.850 246.600 328.650 247.200 ;
        RECT 329.550 246.600 332.550 248.400 ;
        RECT 314.550 237.600 316.350 246.600 ;
        RECT 318.450 245.550 320.250 246.300 ;
        RECT 323.250 245.550 325.050 246.300 ;
        RECT 318.450 244.500 325.050 245.550 ;
        RECT 319.350 237.000 321.150 243.600 ;
        RECT 322.350 237.600 324.150 244.500 ;
        RECT 329.550 243.600 331.650 245.700 ;
        RECT 325.350 237.000 327.150 243.600 ;
        RECT 329.850 237.600 331.650 243.600 ;
        RECT 334.650 237.000 336.450 249.600 ;
        RECT 337.650 237.600 339.450 249.600 ;
        RECT 359.100 243.600 360.300 256.950 ;
        RECT 383.700 243.600 384.900 256.950 ;
        RECT 404.100 243.600 405.300 256.950 ;
        RECT 419.550 256.050 420.450 259.950 ;
        RECT 425.100 259.050 426.900 260.850 ;
        RECT 428.100 259.050 429.300 263.400 ;
        RECT 431.100 259.050 432.900 260.850 ;
        RECT 449.100 259.050 450.900 260.850 ;
        RECT 452.700 259.050 453.900 264.300 ;
        RECT 454.950 259.050 456.750 260.850 ;
        RECT 424.950 256.950 427.050 259.050 ;
        RECT 427.950 256.950 430.050 259.050 ;
        RECT 430.950 256.950 433.050 259.050 ;
        RECT 433.950 256.950 436.050 259.050 ;
        RECT 448.950 256.950 451.050 259.050 ;
        RECT 451.950 256.950 454.050 259.050 ;
        RECT 454.950 256.950 457.050 259.050 ;
        RECT 419.550 254.550 424.050 256.050 ;
        RECT 420.000 253.950 424.050 254.550 ;
        RECT 428.100 249.600 429.300 256.950 ;
        RECT 434.100 255.150 435.900 256.950 ;
        RECT 428.100 248.100 430.500 249.600 ;
        RECT 426.000 245.100 427.800 246.900 ;
        RECT 356.100 237.000 357.900 243.600 ;
        RECT 359.100 237.600 360.900 243.600 ;
        RECT 362.100 237.000 363.900 243.600 ;
        RECT 380.100 237.000 381.900 243.600 ;
        RECT 383.100 237.600 384.900 243.600 ;
        RECT 386.100 237.000 387.900 243.600 ;
        RECT 401.100 237.000 402.900 243.600 ;
        RECT 404.100 237.600 405.900 243.600 ;
        RECT 407.100 237.000 408.900 243.600 ;
        RECT 425.700 237.000 427.500 243.600 ;
        RECT 428.700 237.600 430.500 248.100 ;
        RECT 433.800 237.000 435.600 249.600 ;
        RECT 452.700 243.600 453.900 256.950 ;
        RECT 458.550 251.700 459.450 266.400 ;
        RECT 467.850 265.800 469.650 267.600 ;
        RECT 470.850 267.450 475.800 268.500 ;
        RECT 470.850 266.700 472.650 267.450 ;
        RECT 482.250 267.300 484.650 269.400 ;
        RECT 487.350 266.400 489.150 273.000 ;
        RECT 490.650 266.400 492.450 272.400 ;
        RECT 467.850 264.000 468.900 265.800 ;
        RECT 478.050 264.000 479.850 264.600 ;
        RECT 467.850 262.800 479.850 264.000 ;
        RECT 460.950 261.600 468.900 262.800 ;
        RECT 460.950 259.050 462.750 261.600 ;
        RECT 467.100 261.000 468.900 261.600 ;
        RECT 464.100 259.800 465.900 260.400 ;
        RECT 460.950 256.950 463.050 259.050 ;
        RECT 464.100 258.600 472.200 259.800 ;
        RECT 470.100 256.950 472.200 258.600 ;
        RECT 468.450 251.700 470.250 252.000 ;
        RECT 458.550 251.100 470.250 251.700 ;
        RECT 458.550 250.500 476.850 251.100 ;
        RECT 458.550 249.600 459.450 250.500 ;
        RECT 468.450 250.200 476.850 250.500 ;
        RECT 458.550 247.800 460.950 249.600 ;
        RECT 449.100 237.000 450.900 243.600 ;
        RECT 452.100 237.600 453.900 243.600 ;
        RECT 455.100 237.000 456.900 243.600 ;
        RECT 459.150 237.600 460.950 247.800 ;
        RECT 462.150 237.000 463.950 249.600 ;
        RECT 473.250 248.700 475.050 249.300 ;
        RECT 467.250 247.500 475.050 248.700 ;
        RECT 475.950 248.100 476.850 250.200 ;
        RECT 478.950 250.200 479.850 262.800 ;
        RECT 491.250 259.050 492.450 266.400 ;
        RECT 509.100 263.400 510.900 273.000 ;
        RECT 515.700 264.000 517.500 272.400 ;
        RECT 536.100 269.400 537.900 273.000 ;
        RECT 539.100 269.400 540.900 272.400 ;
        RECT 515.700 262.800 519.000 264.000 ;
        RECT 509.100 259.050 510.900 260.850 ;
        RECT 515.100 259.050 516.900 260.850 ;
        RECT 518.100 259.050 519.000 262.800 ;
        RECT 539.100 259.050 540.300 269.400 ;
        RECT 554.100 263.400 555.900 273.000 ;
        RECT 560.700 264.000 562.500 272.400 ;
        RECT 578.100 267.300 579.900 272.400 ;
        RECT 581.100 268.200 582.900 273.000 ;
        RECT 584.100 267.300 585.900 272.400 ;
        RECT 578.100 265.950 585.900 267.300 ;
        RECT 587.100 266.400 588.900 272.400 ;
        RECT 602.700 269.400 604.500 273.000 ;
        RECT 605.700 267.600 607.500 272.400 ;
        RECT 602.400 266.400 607.500 267.600 ;
        RECT 610.200 266.400 612.000 273.000 ;
        RECT 629.400 266.400 631.200 273.000 ;
        RECT 587.100 264.300 588.300 266.400 ;
        RECT 560.700 262.800 564.000 264.000 ;
        RECT 541.950 261.450 544.050 262.050 ;
        RECT 541.950 260.550 549.450 261.450 ;
        RECT 541.950 259.950 544.050 260.550 ;
        RECT 486.150 257.250 492.450 259.050 ;
        RECT 487.950 256.950 492.450 257.250 ;
        RECT 508.950 256.950 511.050 259.050 ;
        RECT 511.950 256.950 514.050 259.050 ;
        RECT 514.950 256.950 517.050 259.050 ;
        RECT 517.950 256.950 520.050 259.050 ;
        RECT 535.950 256.950 538.050 259.050 ;
        RECT 538.950 256.950 541.050 259.050 ;
        RECT 482.550 254.100 484.650 254.400 ;
        RECT 488.550 254.100 490.350 254.250 ;
        RECT 482.550 252.900 490.350 254.100 ;
        RECT 482.550 252.300 484.650 252.900 ;
        RECT 488.550 252.450 490.350 252.900 ;
        RECT 478.950 249.300 483.750 250.200 ;
        RECT 491.250 249.600 492.450 256.950 ;
        RECT 512.100 255.150 513.900 256.950 ;
        RECT 499.950 252.450 502.050 253.050 ;
        RECT 508.950 252.450 511.050 253.050 ;
        RECT 499.950 251.550 511.050 252.450 ;
        RECT 499.950 250.950 502.050 251.550 ;
        RECT 508.950 250.950 511.050 251.550 ;
        RECT 482.550 248.400 483.750 249.300 ;
        RECT 479.850 248.100 481.650 248.400 ;
        RECT 467.250 246.600 469.350 247.500 ;
        RECT 475.950 247.200 481.650 248.100 ;
        RECT 479.850 246.600 481.650 247.200 ;
        RECT 482.550 246.600 485.550 248.400 ;
        RECT 467.550 237.600 469.350 246.600 ;
        RECT 471.450 245.550 473.250 246.300 ;
        RECT 476.250 245.550 478.050 246.300 ;
        RECT 471.450 244.500 478.050 245.550 ;
        RECT 472.350 237.000 474.150 243.600 ;
        RECT 475.350 237.600 477.150 244.500 ;
        RECT 482.550 243.600 484.650 245.700 ;
        RECT 478.350 237.000 480.150 243.600 ;
        RECT 482.850 237.600 484.650 243.600 ;
        RECT 487.650 237.000 489.450 249.600 ;
        RECT 490.650 237.600 492.450 249.600 ;
        RECT 518.100 244.800 519.000 256.950 ;
        RECT 536.100 255.150 537.900 256.950 ;
        RECT 512.400 243.900 519.000 244.800 ;
        RECT 512.400 243.600 513.900 243.900 ;
        RECT 509.100 237.000 510.900 243.600 ;
        RECT 512.100 237.600 513.900 243.600 ;
        RECT 518.100 243.600 519.000 243.900 ;
        RECT 539.100 243.600 540.300 256.950 ;
        RECT 548.550 256.050 549.450 260.550 ;
        RECT 554.100 259.050 555.900 260.850 ;
        RECT 560.100 259.050 561.900 260.850 ;
        RECT 563.100 259.050 564.000 262.800 ;
        RECT 584.700 263.400 588.300 264.300 ;
        RECT 581.100 259.050 582.900 260.850 ;
        RECT 584.700 259.050 585.900 263.400 ;
        RECT 589.950 261.450 592.050 262.050 ;
        RECT 587.100 259.050 588.900 260.850 ;
        RECT 589.950 260.550 597.450 261.450 ;
        RECT 589.950 259.950 592.050 260.550 ;
        RECT 553.950 256.950 556.050 259.050 ;
        RECT 556.950 256.950 559.050 259.050 ;
        RECT 559.950 256.950 562.050 259.050 ;
        RECT 562.950 256.950 565.050 259.050 ;
        RECT 577.950 256.950 580.050 259.050 ;
        RECT 580.950 256.950 583.050 259.050 ;
        RECT 583.950 256.950 586.050 259.050 ;
        RECT 586.950 256.950 589.050 259.050 ;
        RECT 548.550 254.550 553.050 256.050 ;
        RECT 557.100 255.150 558.900 256.950 ;
        RECT 549.000 253.950 553.050 254.550 ;
        RECT 563.100 244.800 564.000 256.950 ;
        RECT 578.100 255.150 579.900 256.950 ;
        RECT 584.700 249.600 585.900 256.950 ;
        RECT 586.950 252.450 589.050 252.750 ;
        RECT 592.950 252.450 595.050 253.050 ;
        RECT 586.950 251.550 595.050 252.450 ;
        RECT 586.950 250.650 589.050 251.550 ;
        RECT 592.950 250.950 595.050 251.550 ;
        RECT 596.550 250.050 597.450 260.550 ;
        RECT 602.400 259.050 603.300 266.400 ;
        RECT 634.500 265.200 636.300 272.400 ;
        RECT 653.400 266.400 655.200 273.000 ;
        RECT 658.500 265.200 660.300 272.400 ;
        RECT 677.100 269.400 678.900 272.400 ;
        RECT 680.100 269.400 681.900 273.000 ;
        RECT 695.100 269.400 696.900 272.400 ;
        RECT 698.100 269.400 699.900 273.000 ;
        RECT 713.100 269.400 714.900 272.400 ;
        RECT 716.100 269.400 717.900 273.000 ;
        RECT 632.100 264.300 636.300 265.200 ;
        RECT 656.100 264.300 660.300 265.200 ;
        RECT 604.950 259.050 606.750 260.850 ;
        RECT 611.100 259.050 612.900 260.850 ;
        RECT 629.250 259.050 631.050 260.850 ;
        RECT 632.100 259.050 633.300 264.300 ;
        RECT 635.100 259.050 636.900 260.850 ;
        RECT 653.250 259.050 655.050 260.850 ;
        RECT 656.100 259.050 657.300 264.300 ;
        RECT 659.100 259.050 660.900 260.850 ;
        RECT 677.700 259.050 678.900 269.400 ;
        RECT 695.700 259.050 696.900 269.400 ;
        RECT 713.700 259.050 714.900 269.400 ;
        RECT 732.600 268.200 734.400 272.400 ;
        RECT 731.700 266.400 734.400 268.200 ;
        RECT 735.600 266.400 737.400 273.000 ;
        RECT 731.700 259.050 732.600 266.400 ;
        RECT 733.500 264.600 735.300 265.500 ;
        RECT 740.100 264.600 741.900 272.400 ;
        RECT 755.100 269.400 756.900 272.400 ;
        RECT 758.100 269.400 759.900 273.000 ;
        RECT 733.500 263.700 741.900 264.600 ;
        RECT 601.950 256.950 604.050 259.050 ;
        RECT 604.950 256.950 607.050 259.050 ;
        RECT 607.950 256.950 610.050 259.050 ;
        RECT 610.950 256.950 613.050 259.050 ;
        RECT 628.950 256.950 631.050 259.050 ;
        RECT 631.950 256.950 634.050 259.050 ;
        RECT 634.950 256.950 637.050 259.050 ;
        RECT 652.950 256.950 655.050 259.050 ;
        RECT 655.950 256.950 658.050 259.050 ;
        RECT 658.950 256.950 661.050 259.050 ;
        RECT 676.950 256.950 679.050 259.050 ;
        RECT 679.950 256.950 682.050 259.050 ;
        RECT 694.950 256.950 697.050 259.050 ;
        RECT 697.950 256.950 700.050 259.050 ;
        RECT 712.950 256.950 715.050 259.050 ;
        RECT 715.950 256.950 718.050 259.050 ;
        RECT 731.100 256.950 733.200 259.050 ;
        RECT 734.400 256.950 736.500 259.050 ;
        RECT 594.000 249.900 597.450 250.050 ;
        RECT 557.400 243.900 564.000 244.800 ;
        RECT 557.400 243.600 558.900 243.900 ;
        RECT 515.100 237.000 516.900 243.000 ;
        RECT 518.100 237.600 519.900 243.600 ;
        RECT 536.100 237.000 537.900 243.600 ;
        RECT 539.100 237.600 540.900 243.600 ;
        RECT 554.100 237.000 555.900 243.600 ;
        RECT 557.100 237.600 558.900 243.600 ;
        RECT 563.100 243.600 564.000 243.900 ;
        RECT 560.100 237.000 561.900 243.000 ;
        RECT 563.100 237.600 564.900 243.600 ;
        RECT 568.950 240.450 571.050 241.050 ;
        RECT 574.950 240.450 577.050 241.050 ;
        RECT 568.950 239.550 577.050 240.450 ;
        RECT 568.950 238.950 571.050 239.550 ;
        RECT 574.950 238.950 577.050 239.550 ;
        RECT 578.400 237.000 580.200 249.600 ;
        RECT 583.500 248.100 585.900 249.600 ;
        RECT 592.950 248.550 597.450 249.900 ;
        RECT 602.400 249.600 603.300 256.950 ;
        RECT 607.950 255.150 609.750 256.950 ;
        RECT 604.950 252.450 607.050 252.750 ;
        RECT 610.950 252.450 613.050 253.050 ;
        RECT 628.950 252.450 631.050 253.050 ;
        RECT 604.950 251.550 631.050 252.450 ;
        RECT 604.950 250.650 607.050 251.550 ;
        RECT 610.950 250.950 613.050 251.550 ;
        RECT 628.950 250.950 631.050 251.550 ;
        RECT 583.500 237.600 585.300 248.100 ;
        RECT 592.950 247.950 597.000 248.550 ;
        RECT 592.950 247.800 595.050 247.950 ;
        RECT 586.200 245.100 588.000 246.900 ;
        RECT 586.500 237.000 588.300 243.600 ;
        RECT 602.100 237.600 603.900 249.600 ;
        RECT 605.100 248.700 612.900 249.600 ;
        RECT 605.100 237.600 606.900 248.700 ;
        RECT 608.100 237.000 609.900 247.800 ;
        RECT 611.100 237.600 612.900 248.700 ;
        RECT 632.100 243.600 633.300 256.950 ;
        RECT 656.100 243.600 657.300 256.950 ;
        RECT 677.700 243.600 678.900 256.950 ;
        RECT 680.100 255.150 681.900 256.950 ;
        RECT 695.700 243.600 696.900 256.950 ;
        RECT 698.100 255.150 699.900 256.950 ;
        RECT 700.950 249.450 703.050 250.050 ;
        RECT 709.950 249.450 712.050 253.050 ;
        RECT 700.950 249.000 712.050 249.450 ;
        RECT 700.950 248.550 711.450 249.000 ;
        RECT 700.950 247.950 703.050 248.550 ;
        RECT 713.700 243.600 714.900 256.950 ;
        RECT 716.100 255.150 717.900 256.950 ;
        RECT 731.700 249.600 732.600 256.950 ;
        RECT 735.000 255.150 736.800 256.950 ;
        RECT 629.100 237.000 630.900 243.600 ;
        RECT 632.100 237.600 633.900 243.600 ;
        RECT 635.100 237.000 636.900 243.600 ;
        RECT 653.100 237.000 654.900 243.600 ;
        RECT 656.100 237.600 657.900 243.600 ;
        RECT 659.100 237.000 660.900 243.600 ;
        RECT 677.100 237.600 678.900 243.600 ;
        RECT 680.100 237.000 681.900 243.600 ;
        RECT 695.100 237.600 696.900 243.600 ;
        RECT 698.100 237.000 699.900 243.600 ;
        RECT 713.100 237.600 714.900 243.600 ;
        RECT 716.100 237.000 717.900 243.600 ;
        RECT 731.100 237.600 732.900 249.600 ;
        RECT 734.100 237.000 735.900 249.000 ;
        RECT 738.000 243.600 738.900 263.700 ;
        RECT 739.950 259.050 741.750 260.850 ;
        RECT 755.700 259.050 756.900 269.400 ;
        RECT 773.100 267.300 774.900 272.400 ;
        RECT 776.100 268.200 777.900 273.000 ;
        RECT 779.100 267.300 780.900 272.400 ;
        RECT 773.100 265.950 780.900 267.300 ;
        RECT 782.100 266.400 783.900 272.400 ;
        RECT 800.100 269.400 801.900 273.000 ;
        RECT 803.100 269.400 804.900 272.400 ;
        RECT 818.100 269.400 819.900 273.000 ;
        RECT 821.100 269.400 822.900 272.400 ;
        RECT 839.700 269.400 841.500 273.000 ;
        RECT 782.100 264.300 783.300 266.400 ;
        RECT 779.700 263.400 783.300 264.300 ;
        RECT 776.100 259.050 777.900 260.850 ;
        RECT 779.700 259.050 780.900 263.400 ;
        RECT 782.100 259.050 783.900 260.850 ;
        RECT 803.100 259.050 804.300 269.400 ;
        RECT 821.100 259.050 822.300 269.400 ;
        RECT 842.700 267.600 844.500 272.400 ;
        RECT 839.400 266.400 844.500 267.600 ;
        RECT 847.200 266.400 849.000 273.000 ;
        RECT 839.400 259.050 840.300 266.400 ;
        RECT 863.100 263.400 864.900 273.000 ;
        RECT 869.700 264.000 871.500 272.400 ;
        RECT 869.700 262.800 873.000 264.000 ;
        RECT 887.100 263.400 888.900 273.000 ;
        RECT 893.700 264.000 895.500 272.400 ;
        RECT 912.000 266.400 913.800 273.000 ;
        RECT 916.500 267.600 918.300 272.400 ;
        RECT 919.500 269.400 921.300 273.000 ;
        RECT 916.500 266.400 921.600 267.600 ;
        RECT 935.100 266.400 936.900 272.400 ;
        RECT 893.700 262.800 897.000 264.000 ;
        RECT 841.950 259.050 843.750 260.850 ;
        RECT 848.100 259.050 849.900 260.850 ;
        RECT 863.100 259.050 864.900 260.850 ;
        RECT 869.100 259.050 870.900 260.850 ;
        RECT 872.100 259.050 873.000 262.800 ;
        RECT 887.100 259.050 888.900 260.850 ;
        RECT 893.100 259.050 894.900 260.850 ;
        RECT 896.100 259.050 897.000 262.800 ;
        RECT 911.100 259.050 912.900 260.850 ;
        RECT 917.250 259.050 919.050 260.850 ;
        RECT 920.700 259.050 921.600 266.400 ;
        RECT 935.700 264.300 936.900 266.400 ;
        RECT 938.100 267.300 939.900 272.400 ;
        RECT 941.100 268.200 942.900 273.000 ;
        RECT 944.100 267.300 945.900 272.400 ;
        RECT 938.100 265.950 945.900 267.300 ;
        RECT 962.100 266.400 963.900 272.400 ;
        RECT 962.700 264.300 963.900 266.400 ;
        RECT 965.100 267.300 966.900 272.400 ;
        RECT 968.100 268.200 969.900 273.000 ;
        RECT 971.100 267.300 972.900 272.400 ;
        RECT 965.100 265.950 972.900 267.300 ;
        RECT 987.000 266.400 988.800 273.000 ;
        RECT 991.500 267.600 993.300 272.400 ;
        RECT 994.500 269.400 996.300 273.000 ;
        RECT 991.500 266.400 996.600 267.600 ;
        RECT 973.950 264.450 976.050 265.050 ;
        RECT 991.950 264.450 994.050 265.050 ;
        RECT 935.700 263.400 939.300 264.300 ;
        RECT 962.700 263.400 966.300 264.300 ;
        RECT 935.100 259.050 936.900 260.850 ;
        RECT 938.100 259.050 939.300 263.400 ;
        RECT 946.950 261.450 949.050 262.050 ;
        RECT 958.950 261.450 961.050 262.050 ;
        RECT 941.100 259.050 942.900 260.850 ;
        RECT 946.950 260.550 961.050 261.450 ;
        RECT 946.950 259.950 949.050 260.550 ;
        RECT 958.950 259.950 961.050 260.550 ;
        RECT 962.100 259.050 963.900 260.850 ;
        RECT 965.100 259.050 966.300 263.400 ;
        RECT 973.950 263.550 994.050 264.450 ;
        RECT 973.950 262.950 976.050 263.550 ;
        RECT 991.950 262.950 994.050 263.550 ;
        RECT 968.100 259.050 969.900 260.850 ;
        RECT 986.100 259.050 987.900 260.850 ;
        RECT 992.250 259.050 994.050 260.850 ;
        RECT 995.700 259.050 996.600 266.400 ;
        RECT 997.950 261.450 1000.050 262.050 ;
        RECT 1009.950 261.450 1012.050 262.050 ;
        RECT 997.950 260.550 1012.050 261.450 ;
        RECT 997.950 259.950 1000.050 260.550 ;
        RECT 1009.950 259.950 1012.050 260.550 ;
        RECT 739.800 256.950 741.900 259.050 ;
        RECT 754.950 256.950 757.050 259.050 ;
        RECT 757.950 256.950 760.050 259.050 ;
        RECT 772.950 256.950 775.050 259.050 ;
        RECT 775.950 256.950 778.050 259.050 ;
        RECT 778.950 256.950 781.050 259.050 ;
        RECT 781.950 256.950 784.050 259.050 ;
        RECT 799.950 256.950 802.050 259.050 ;
        RECT 802.950 256.950 805.050 259.050 ;
        RECT 817.950 256.950 820.050 259.050 ;
        RECT 820.950 256.950 823.050 259.050 ;
        RECT 838.950 256.950 841.050 259.050 ;
        RECT 841.950 256.950 844.050 259.050 ;
        RECT 844.950 256.950 847.050 259.050 ;
        RECT 847.950 256.950 850.050 259.050 ;
        RECT 862.950 256.950 865.050 259.050 ;
        RECT 865.950 256.950 868.050 259.050 ;
        RECT 868.950 256.950 871.050 259.050 ;
        RECT 871.950 256.950 874.050 259.050 ;
        RECT 886.950 256.950 889.050 259.050 ;
        RECT 889.950 256.950 892.050 259.050 ;
        RECT 892.950 256.950 895.050 259.050 ;
        RECT 895.950 256.950 898.050 259.050 ;
        RECT 910.950 256.950 913.050 259.050 ;
        RECT 913.950 256.950 916.050 259.050 ;
        RECT 916.950 256.950 919.050 259.050 ;
        RECT 919.950 256.950 922.050 259.050 ;
        RECT 934.950 256.950 937.050 259.050 ;
        RECT 937.950 256.950 940.050 259.050 ;
        RECT 940.950 256.950 943.050 259.050 ;
        RECT 943.950 256.950 946.050 259.050 ;
        RECT 961.950 256.950 964.050 259.050 ;
        RECT 964.950 256.950 967.050 259.050 ;
        RECT 967.950 256.950 970.050 259.050 ;
        RECT 970.950 256.950 973.050 259.050 ;
        RECT 985.950 256.950 988.050 259.050 ;
        RECT 988.950 256.950 991.050 259.050 ;
        RECT 991.950 256.950 994.050 259.050 ;
        RECT 994.950 256.950 997.050 259.050 ;
        RECT 755.700 243.600 756.900 256.950 ;
        RECT 758.100 255.150 759.900 256.950 ;
        RECT 773.100 255.150 774.900 256.950 ;
        RECT 779.700 249.600 780.900 256.950 ;
        RECT 800.100 255.150 801.900 256.950 ;
        RECT 737.100 237.600 738.900 243.600 ;
        RECT 740.100 237.000 741.900 243.600 ;
        RECT 755.100 237.600 756.900 243.600 ;
        RECT 758.100 237.000 759.900 243.600 ;
        RECT 773.400 237.000 775.200 249.600 ;
        RECT 778.500 248.100 780.900 249.600 ;
        RECT 778.500 237.600 780.300 248.100 ;
        RECT 781.200 245.100 783.000 246.900 ;
        RECT 803.100 243.600 804.300 256.950 ;
        RECT 818.100 255.150 819.900 256.950 ;
        RECT 821.100 243.600 822.300 256.950 ;
        RECT 839.400 249.600 840.300 256.950 ;
        RECT 844.950 255.150 846.750 256.950 ;
        RECT 866.100 255.150 867.900 256.950 ;
        RECT 847.950 252.450 850.050 253.050 ;
        RECT 868.950 252.450 871.050 253.050 ;
        RECT 847.950 251.550 871.050 252.450 ;
        RECT 847.950 250.950 850.050 251.550 ;
        RECT 868.950 250.950 871.050 251.550 ;
        RECT 781.500 237.000 783.300 243.600 ;
        RECT 800.100 237.000 801.900 243.600 ;
        RECT 803.100 237.600 804.900 243.600 ;
        RECT 818.100 237.000 819.900 243.600 ;
        RECT 821.100 237.600 822.900 243.600 ;
        RECT 839.100 237.600 840.900 249.600 ;
        RECT 842.100 248.700 849.900 249.600 ;
        RECT 842.100 237.600 843.900 248.700 ;
        RECT 845.100 237.000 846.900 247.800 ;
        RECT 848.100 237.600 849.900 248.700 ;
        RECT 872.100 244.800 873.000 256.950 ;
        RECT 890.100 255.150 891.900 256.950 ;
        RECT 896.100 244.800 897.000 256.950 ;
        RECT 914.250 255.150 916.050 256.950 ;
        RECT 920.700 249.600 921.600 256.950 ;
        RECT 938.100 249.600 939.300 256.950 ;
        RECT 944.100 255.150 945.900 256.950 ;
        RECT 965.100 249.600 966.300 256.950 ;
        RECT 971.100 255.150 972.900 256.950 ;
        RECT 989.250 255.150 991.050 256.950 ;
        RECT 995.700 249.600 996.600 256.950 ;
        RECT 866.400 243.900 873.000 244.800 ;
        RECT 866.400 243.600 867.900 243.900 ;
        RECT 863.100 237.000 864.900 243.600 ;
        RECT 866.100 237.600 867.900 243.600 ;
        RECT 872.100 243.600 873.000 243.900 ;
        RECT 890.400 243.900 897.000 244.800 ;
        RECT 890.400 243.600 891.900 243.900 ;
        RECT 869.100 237.000 870.900 243.000 ;
        RECT 872.100 237.600 873.900 243.600 ;
        RECT 887.100 237.000 888.900 243.600 ;
        RECT 890.100 237.600 891.900 243.600 ;
        RECT 896.100 243.600 897.000 243.900 ;
        RECT 911.100 248.700 918.900 249.600 ;
        RECT 893.100 237.000 894.900 243.000 ;
        RECT 896.100 237.600 897.900 243.600 ;
        RECT 911.100 237.600 912.900 248.700 ;
        RECT 914.100 237.000 915.900 247.800 ;
        RECT 917.100 237.600 918.900 248.700 ;
        RECT 920.100 237.600 921.900 249.600 ;
        RECT 938.100 248.100 940.500 249.600 ;
        RECT 936.000 245.100 937.800 246.900 ;
        RECT 935.700 237.000 937.500 243.600 ;
        RECT 938.700 237.600 940.500 248.100 ;
        RECT 943.800 237.000 945.600 249.600 ;
        RECT 965.100 248.100 967.500 249.600 ;
        RECT 963.000 245.100 964.800 246.900 ;
        RECT 962.700 237.000 964.500 243.600 ;
        RECT 965.700 237.600 967.500 248.100 ;
        RECT 970.800 237.000 972.600 249.600 ;
        RECT 986.100 248.700 993.900 249.600 ;
        RECT 986.100 237.600 987.900 248.700 ;
        RECT 989.100 237.000 990.900 247.800 ;
        RECT 992.100 237.600 993.900 248.700 ;
        RECT 995.100 237.600 996.900 249.600 ;
        RECT 14.100 227.400 15.900 233.400 ;
        RECT 14.100 220.500 15.300 227.400 ;
        RECT 17.100 223.200 18.900 234.000 ;
        RECT 20.100 221.400 21.900 233.400 ;
        RECT 38.100 227.400 39.900 234.000 ;
        RECT 41.100 227.400 42.900 233.400 ;
        RECT 56.100 227.400 57.900 234.000 ;
        RECT 59.100 227.400 60.900 233.400 ;
        RECT 62.100 228.000 63.900 234.000 ;
        RECT 14.100 219.600 19.800 220.500 ;
        RECT 18.000 218.700 19.800 219.600 ;
        RECT 14.400 214.050 16.200 215.850 ;
        RECT 14.400 211.950 16.500 214.050 ;
        RECT 18.000 207.300 18.900 218.700 ;
        RECT 20.700 214.050 21.900 221.400 ;
        RECT 38.100 214.050 39.900 215.850 ;
        RECT 41.100 214.050 42.300 227.400 ;
        RECT 59.400 227.100 60.900 227.400 ;
        RECT 65.100 227.400 66.900 233.400 ;
        RECT 83.700 227.400 85.500 234.000 ;
        RECT 65.100 227.100 66.000 227.400 ;
        RECT 59.400 226.200 66.000 227.100 ;
        RECT 59.100 214.050 60.900 215.850 ;
        RECT 65.100 214.050 66.000 226.200 ;
        RECT 84.000 224.100 85.800 225.900 ;
        RECT 86.700 222.900 88.500 233.400 ;
        RECT 86.100 221.400 88.500 222.900 ;
        RECT 91.800 221.400 93.600 234.000 ;
        RECT 107.100 222.300 108.900 233.400 ;
        RECT 110.100 223.200 111.900 234.000 ;
        RECT 113.100 222.300 114.900 233.400 ;
        RECT 107.100 221.400 114.900 222.300 ;
        RECT 116.100 221.400 117.900 233.400 ;
        RECT 131.100 221.400 132.900 233.400 ;
        RECT 134.100 222.300 135.900 233.400 ;
        RECT 137.100 223.200 138.900 234.000 ;
        RECT 140.100 222.300 141.900 233.400 ;
        RECT 155.100 227.400 156.900 234.000 ;
        RECT 158.100 227.400 159.900 233.400 ;
        RECT 176.100 227.400 177.900 234.000 ;
        RECT 179.100 227.400 180.900 233.400 ;
        RECT 182.100 227.400 183.900 234.000 ;
        RECT 200.700 227.400 202.500 234.000 ;
        RECT 134.100 221.400 141.900 222.300 ;
        RECT 86.100 214.050 87.300 221.400 ;
        RECT 92.100 214.050 93.900 215.850 ;
        RECT 110.250 214.050 112.050 215.850 ;
        RECT 116.700 214.050 117.600 221.400 ;
        RECT 131.400 214.050 132.300 221.400 ;
        RECT 136.950 214.050 138.750 215.850 ;
        RECT 155.100 214.050 156.900 215.850 ;
        RECT 158.100 214.050 159.300 227.400 ;
        RECT 179.100 214.050 180.300 227.400 ;
        RECT 201.000 224.100 202.800 225.900 ;
        RECT 203.700 222.900 205.500 233.400 ;
        RECT 203.100 221.400 205.500 222.900 ;
        RECT 208.800 221.400 210.600 234.000 ;
        RECT 224.100 227.400 225.900 234.000 ;
        RECT 227.100 227.400 228.900 233.400 ;
        RECT 230.100 227.400 231.900 234.000 ;
        RECT 245.100 227.400 246.900 234.000 ;
        RECT 248.100 227.400 249.900 233.400 ;
        RECT 251.100 228.000 252.900 234.000 ;
        RECT 203.100 214.050 204.300 221.400 ;
        RECT 209.100 214.050 210.900 215.850 ;
        RECT 227.700 214.050 228.900 227.400 ;
        RECT 248.400 227.100 249.900 227.400 ;
        RECT 254.100 227.400 255.900 233.400 ;
        RECT 254.100 227.100 255.000 227.400 ;
        RECT 248.400 226.200 255.000 227.100 ;
        RECT 248.100 214.050 249.900 215.850 ;
        RECT 254.100 214.050 255.000 226.200 ;
        RECT 272.100 221.400 273.900 233.400 ;
        RECT 275.100 222.300 276.900 233.400 ;
        RECT 278.100 223.200 279.900 234.000 ;
        RECT 281.100 222.300 282.900 233.400 ;
        RECT 296.700 227.400 298.500 234.000 ;
        RECT 297.000 224.100 298.800 225.900 ;
        RECT 299.700 222.900 301.500 233.400 ;
        RECT 275.100 221.400 282.900 222.300 ;
        RECT 299.100 221.400 301.500 222.900 ;
        RECT 304.800 221.400 306.600 234.000 ;
        RECT 309.150 223.200 310.950 233.400 ;
        RECT 308.550 221.400 310.950 223.200 ;
        RECT 312.150 221.400 313.950 234.000 ;
        RECT 317.550 224.400 319.350 233.400 ;
        RECT 322.350 227.400 324.150 234.000 ;
        RECT 325.350 226.500 327.150 233.400 ;
        RECT 328.350 227.400 330.150 234.000 ;
        RECT 332.850 227.400 334.650 233.400 ;
        RECT 321.450 225.450 328.050 226.500 ;
        RECT 321.450 224.700 323.250 225.450 ;
        RECT 326.250 224.700 328.050 225.450 ;
        RECT 332.550 225.300 334.650 227.400 ;
        RECT 317.250 223.500 319.350 224.400 ;
        RECT 329.850 223.800 331.650 224.400 ;
        RECT 317.250 222.300 325.050 223.500 ;
        RECT 323.250 221.700 325.050 222.300 ;
        RECT 325.950 222.900 331.650 223.800 ;
        RECT 272.400 214.050 273.300 221.400 ;
        RECT 277.950 214.050 279.750 215.850 ;
        RECT 299.100 214.050 300.300 221.400 ;
        RECT 308.550 220.500 309.450 221.400 ;
        RECT 325.950 220.800 326.850 222.900 ;
        RECT 329.850 222.600 331.650 222.900 ;
        RECT 332.550 222.600 335.550 224.400 ;
        RECT 332.550 221.700 333.750 222.600 ;
        RECT 318.450 220.500 326.850 220.800 ;
        RECT 308.550 219.900 326.850 220.500 ;
        RECT 328.950 220.800 333.750 221.700 ;
        RECT 337.650 221.400 339.450 234.000 ;
        RECT 340.650 221.400 342.450 233.400 ;
        RECT 359.100 227.400 360.900 234.000 ;
        RECT 362.100 227.400 363.900 233.400 ;
        RECT 308.550 219.300 320.250 219.900 ;
        RECT 305.100 214.050 306.900 215.850 ;
        RECT 19.800 211.950 21.900 214.050 ;
        RECT 37.950 211.950 40.050 214.050 ;
        RECT 40.950 211.950 43.050 214.050 ;
        RECT 55.950 211.950 58.050 214.050 ;
        RECT 58.950 211.950 61.050 214.050 ;
        RECT 61.950 211.950 64.050 214.050 ;
        RECT 64.950 211.950 67.050 214.050 ;
        RECT 82.950 211.950 85.050 214.050 ;
        RECT 85.950 211.950 88.050 214.050 ;
        RECT 88.950 211.950 91.050 214.050 ;
        RECT 91.950 211.950 94.050 214.050 ;
        RECT 106.950 211.950 109.050 214.050 ;
        RECT 109.950 211.950 112.050 214.050 ;
        RECT 112.950 211.950 115.050 214.050 ;
        RECT 115.950 211.950 118.050 214.050 ;
        RECT 130.950 211.950 133.050 214.050 ;
        RECT 133.950 211.950 136.050 214.050 ;
        RECT 136.950 211.950 139.050 214.050 ;
        RECT 139.950 211.950 142.050 214.050 ;
        RECT 154.950 211.950 157.050 214.050 ;
        RECT 157.950 211.950 160.050 214.050 ;
        RECT 175.950 211.950 178.050 214.050 ;
        RECT 178.950 211.950 181.050 214.050 ;
        RECT 181.950 211.950 184.050 214.050 ;
        RECT 199.950 211.950 202.050 214.050 ;
        RECT 202.950 211.950 205.050 214.050 ;
        RECT 205.950 211.950 208.050 214.050 ;
        RECT 208.950 211.950 211.050 214.050 ;
        RECT 223.950 211.950 226.050 214.050 ;
        RECT 226.950 211.950 229.050 214.050 ;
        RECT 229.950 211.950 232.050 214.050 ;
        RECT 244.950 211.950 247.050 214.050 ;
        RECT 247.950 211.950 250.050 214.050 ;
        RECT 250.950 211.950 253.050 214.050 ;
        RECT 253.950 211.950 256.050 214.050 ;
        RECT 271.950 211.950 274.050 214.050 ;
        RECT 274.950 211.950 277.050 214.050 ;
        RECT 277.950 211.950 280.050 214.050 ;
        RECT 280.950 211.950 283.050 214.050 ;
        RECT 295.950 211.950 298.050 214.050 ;
        RECT 298.950 211.950 301.050 214.050 ;
        RECT 301.950 211.950 304.050 214.050 ;
        RECT 304.950 211.950 307.050 214.050 ;
        RECT 18.000 206.400 19.800 207.300 ;
        RECT 14.100 205.500 19.800 206.400 ;
        RECT 14.100 201.600 15.300 205.500 ;
        RECT 20.700 204.600 21.900 211.950 ;
        RECT 14.100 198.600 15.900 201.600 ;
        RECT 17.100 198.000 18.900 204.600 ;
        RECT 20.100 198.600 21.900 204.600 ;
        RECT 41.100 201.600 42.300 211.950 ;
        RECT 56.100 210.150 57.900 211.950 ;
        RECT 62.100 210.150 63.900 211.950 ;
        RECT 65.100 208.200 66.000 211.950 ;
        RECT 83.100 210.150 84.900 211.950 ;
        RECT 38.100 198.000 39.900 201.600 ;
        RECT 41.100 198.600 42.900 201.600 ;
        RECT 56.100 198.000 57.900 207.600 ;
        RECT 62.700 207.000 66.000 208.200 ;
        RECT 86.100 207.600 87.300 211.950 ;
        RECT 89.100 210.150 90.900 211.950 ;
        RECT 107.100 210.150 108.900 211.950 ;
        RECT 113.250 210.150 115.050 211.950 ;
        RECT 62.700 198.600 64.500 207.000 ;
        RECT 83.700 206.700 87.300 207.600 ;
        RECT 83.700 204.600 84.900 206.700 ;
        RECT 83.100 198.600 84.900 204.600 ;
        RECT 86.100 203.700 93.900 205.050 ;
        RECT 116.700 204.600 117.600 211.950 ;
        RECT 86.100 198.600 87.900 203.700 ;
        RECT 89.100 198.000 90.900 202.800 ;
        RECT 92.100 198.600 93.900 203.700 ;
        RECT 108.000 198.000 109.800 204.600 ;
        RECT 112.500 203.400 117.600 204.600 ;
        RECT 131.400 204.600 132.300 211.950 ;
        RECT 133.950 210.150 135.750 211.950 ;
        RECT 140.100 210.150 141.900 211.950 ;
        RECT 131.400 203.400 136.500 204.600 ;
        RECT 112.500 198.600 114.300 203.400 ;
        RECT 115.500 198.000 117.300 201.600 ;
        RECT 131.700 198.000 133.500 201.600 ;
        RECT 134.700 198.600 136.500 203.400 ;
        RECT 139.200 198.000 141.000 204.600 ;
        RECT 158.100 201.600 159.300 211.950 ;
        RECT 176.250 210.150 178.050 211.950 ;
        RECT 179.100 206.700 180.300 211.950 ;
        RECT 182.100 210.150 183.900 211.950 ;
        RECT 200.100 210.150 201.900 211.950 ;
        RECT 203.100 207.600 204.300 211.950 ;
        RECT 206.100 210.150 207.900 211.950 ;
        RECT 224.100 210.150 225.900 211.950 ;
        RECT 200.700 206.700 204.300 207.600 ;
        RECT 227.700 206.700 228.900 211.950 ;
        RECT 229.950 210.150 231.750 211.950 ;
        RECT 245.100 210.150 246.900 211.950 ;
        RECT 251.100 210.150 252.900 211.950 ;
        RECT 254.100 208.200 255.000 211.950 ;
        RECT 179.100 205.800 183.300 206.700 ;
        RECT 155.100 198.000 156.900 201.600 ;
        RECT 158.100 198.600 159.900 201.600 ;
        RECT 176.400 198.000 178.200 204.600 ;
        RECT 181.500 198.600 183.300 205.800 ;
        RECT 200.700 204.600 201.900 206.700 ;
        RECT 224.700 205.800 228.900 206.700 ;
        RECT 200.100 198.600 201.900 204.600 ;
        RECT 203.100 203.700 210.900 205.050 ;
        RECT 203.100 198.600 204.900 203.700 ;
        RECT 206.100 198.000 207.900 202.800 ;
        RECT 209.100 198.600 210.900 203.700 ;
        RECT 224.700 198.600 226.500 205.800 ;
        RECT 229.800 198.000 231.600 204.600 ;
        RECT 245.100 198.000 246.900 207.600 ;
        RECT 251.700 207.000 255.000 208.200 ;
        RECT 251.700 198.600 253.500 207.000 ;
        RECT 272.400 204.600 273.300 211.950 ;
        RECT 274.950 210.150 276.750 211.950 ;
        RECT 281.100 210.150 282.900 211.950 ;
        RECT 296.100 210.150 297.900 211.950 ;
        RECT 299.100 207.600 300.300 211.950 ;
        RECT 302.100 210.150 303.900 211.950 ;
        RECT 296.700 206.700 300.300 207.600 ;
        RECT 296.700 204.600 297.900 206.700 ;
        RECT 272.400 203.400 277.500 204.600 ;
        RECT 272.700 198.000 274.500 201.600 ;
        RECT 275.700 198.600 277.500 203.400 ;
        RECT 280.200 198.000 282.000 204.600 ;
        RECT 296.100 198.600 297.900 204.600 ;
        RECT 299.100 203.700 306.900 205.050 ;
        RECT 299.100 198.600 300.900 203.700 ;
        RECT 302.100 198.000 303.900 202.800 ;
        RECT 305.100 198.600 306.900 203.700 ;
        RECT 308.550 204.600 309.450 219.300 ;
        RECT 318.450 219.000 320.250 219.300 ;
        RECT 310.950 211.950 313.050 214.050 ;
        RECT 320.100 212.400 322.200 214.050 ;
        RECT 310.950 209.400 312.750 211.950 ;
        RECT 314.100 211.200 322.200 212.400 ;
        RECT 314.100 210.600 315.900 211.200 ;
        RECT 317.100 209.400 318.900 210.000 ;
        RECT 310.950 208.200 318.900 209.400 ;
        RECT 328.950 208.200 329.850 220.800 ;
        RECT 332.550 218.100 334.650 218.700 ;
        RECT 338.550 218.100 340.350 218.550 ;
        RECT 332.550 216.900 340.350 218.100 ;
        RECT 332.550 216.600 334.650 216.900 ;
        RECT 338.550 216.750 340.350 216.900 ;
        RECT 341.250 214.050 342.450 221.400 ;
        RECT 359.100 214.050 360.900 215.850 ;
        RECT 362.100 214.050 363.300 227.400 ;
        RECT 380.100 221.400 381.900 233.400 ;
        RECT 383.100 223.200 384.900 234.000 ;
        RECT 386.100 227.400 387.900 233.400 ;
        RECT 380.100 214.050 381.300 221.400 ;
        RECT 386.700 220.500 387.900 227.400 ;
        RECT 390.150 223.200 391.950 233.400 ;
        RECT 382.200 219.600 387.900 220.500 ;
        RECT 389.550 221.400 391.950 223.200 ;
        RECT 393.150 221.400 394.950 234.000 ;
        RECT 398.550 224.400 400.350 233.400 ;
        RECT 403.350 227.400 405.150 234.000 ;
        RECT 406.350 226.500 408.150 233.400 ;
        RECT 409.350 227.400 411.150 234.000 ;
        RECT 413.850 227.400 415.650 233.400 ;
        RECT 402.450 225.450 409.050 226.500 ;
        RECT 402.450 224.700 404.250 225.450 ;
        RECT 407.250 224.700 409.050 225.450 ;
        RECT 413.550 225.300 415.650 227.400 ;
        RECT 398.250 223.500 400.350 224.400 ;
        RECT 410.850 223.800 412.650 224.400 ;
        RECT 398.250 222.300 406.050 223.500 ;
        RECT 404.250 221.700 406.050 222.300 ;
        RECT 406.950 222.900 412.650 223.800 ;
        RECT 389.550 220.500 390.450 221.400 ;
        RECT 406.950 220.800 407.850 222.900 ;
        RECT 410.850 222.600 412.650 222.900 ;
        RECT 413.550 222.600 416.550 224.400 ;
        RECT 413.550 221.700 414.750 222.600 ;
        RECT 399.450 220.500 407.850 220.800 ;
        RECT 389.550 219.900 407.850 220.500 ;
        RECT 409.950 220.800 414.750 221.700 ;
        RECT 418.650 221.400 420.450 234.000 ;
        RECT 421.650 221.400 423.450 233.400 ;
        RECT 440.100 227.400 441.900 234.000 ;
        RECT 443.100 227.400 444.900 233.400 ;
        RECT 446.100 227.400 447.900 234.000 ;
        RECT 382.200 218.700 384.000 219.600 ;
        RECT 337.950 213.750 342.450 214.050 ;
        RECT 336.150 211.950 342.450 213.750 ;
        RECT 358.950 211.950 361.050 214.050 ;
        RECT 361.950 211.950 364.050 214.050 ;
        RECT 380.100 211.950 382.200 214.050 ;
        RECT 317.850 207.000 329.850 208.200 ;
        RECT 317.850 205.200 318.900 207.000 ;
        RECT 328.050 206.400 329.850 207.000 ;
        RECT 308.550 202.800 310.950 204.600 ;
        RECT 309.150 198.600 310.950 202.800 ;
        RECT 312.150 198.000 313.950 204.600 ;
        RECT 314.850 202.200 316.950 203.700 ;
        RECT 317.850 203.400 319.650 205.200 ;
        RECT 341.250 204.600 342.450 211.950 ;
        RECT 320.850 203.550 322.650 204.300 ;
        RECT 320.850 202.500 325.800 203.550 ;
        RECT 314.850 201.600 318.750 202.200 ;
        RECT 324.750 201.600 325.800 202.500 ;
        RECT 332.250 201.600 334.650 203.700 ;
        RECT 315.150 200.700 318.750 201.600 ;
        RECT 316.950 198.600 318.750 200.700 ;
        RECT 321.450 198.000 323.250 201.600 ;
        RECT 324.750 198.600 326.550 201.600 ;
        RECT 327.750 198.000 329.550 201.600 ;
        RECT 332.250 198.600 334.050 201.600 ;
        RECT 337.350 198.000 339.150 204.600 ;
        RECT 340.650 198.600 342.450 204.600 ;
        RECT 362.100 201.600 363.300 211.950 ;
        RECT 380.100 204.600 381.300 211.950 ;
        RECT 383.100 207.300 384.000 218.700 ;
        RECT 389.550 219.300 401.250 219.900 ;
        RECT 385.800 214.050 387.600 215.850 ;
        RECT 385.500 211.950 387.600 214.050 ;
        RECT 382.200 206.400 384.000 207.300 ;
        RECT 382.200 205.500 387.900 206.400 ;
        RECT 359.100 198.000 360.900 201.600 ;
        RECT 362.100 198.600 363.900 201.600 ;
        RECT 380.100 198.600 381.900 204.600 ;
        RECT 383.100 198.000 384.900 204.600 ;
        RECT 386.700 201.600 387.900 205.500 ;
        RECT 389.550 204.600 390.450 219.300 ;
        RECT 399.450 219.000 401.250 219.300 ;
        RECT 391.950 211.950 394.050 214.050 ;
        RECT 401.100 212.400 403.200 214.050 ;
        RECT 391.950 209.400 393.750 211.950 ;
        RECT 395.100 211.200 403.200 212.400 ;
        RECT 395.100 210.600 396.900 211.200 ;
        RECT 398.100 209.400 399.900 210.000 ;
        RECT 391.950 208.200 399.900 209.400 ;
        RECT 409.950 208.200 410.850 220.800 ;
        RECT 413.550 218.100 415.650 218.700 ;
        RECT 419.550 218.100 421.350 218.550 ;
        RECT 413.550 216.900 421.350 218.100 ;
        RECT 413.550 216.600 415.650 216.900 ;
        RECT 419.550 216.750 421.350 216.900 ;
        RECT 422.250 214.050 423.450 221.400 ;
        RECT 443.700 214.050 444.900 227.400 ;
        RECT 449.550 221.400 451.350 233.400 ;
        RECT 452.550 221.400 454.350 234.000 ;
        RECT 457.350 227.400 459.150 233.400 ;
        RECT 461.850 227.400 463.650 234.000 ;
        RECT 457.350 225.300 459.450 227.400 ;
        RECT 464.850 226.500 466.650 233.400 ;
        RECT 467.850 227.400 469.650 234.000 ;
        RECT 463.950 225.450 470.550 226.500 ;
        RECT 463.950 224.700 465.750 225.450 ;
        RECT 468.750 224.700 470.550 225.450 ;
        RECT 472.650 224.400 474.450 233.400 ;
        RECT 456.450 222.600 459.450 224.400 ;
        RECT 460.350 223.800 462.150 224.400 ;
        RECT 460.350 222.900 466.050 223.800 ;
        RECT 472.650 223.500 474.750 224.400 ;
        RECT 460.350 222.600 462.150 222.900 ;
        RECT 458.250 221.700 459.450 222.600 ;
        RECT 449.550 214.050 450.750 221.400 ;
        RECT 458.250 220.800 463.050 221.700 ;
        RECT 451.650 218.100 453.450 218.550 ;
        RECT 457.350 218.100 459.450 218.700 ;
        RECT 451.650 216.900 459.450 218.100 ;
        RECT 451.650 216.750 453.450 216.900 ;
        RECT 457.350 216.600 459.450 216.900 ;
        RECT 418.950 213.750 423.450 214.050 ;
        RECT 417.150 211.950 423.450 213.750 ;
        RECT 439.950 211.950 442.050 214.050 ;
        RECT 442.950 211.950 445.050 214.050 ;
        RECT 445.950 211.950 448.050 214.050 ;
        RECT 449.550 213.750 454.050 214.050 ;
        RECT 449.550 211.950 455.850 213.750 ;
        RECT 398.850 207.000 410.850 208.200 ;
        RECT 398.850 205.200 399.900 207.000 ;
        RECT 409.050 206.400 410.850 207.000 ;
        RECT 389.550 202.800 391.950 204.600 ;
        RECT 386.100 198.600 387.900 201.600 ;
        RECT 390.150 198.600 391.950 202.800 ;
        RECT 393.150 198.000 394.950 204.600 ;
        RECT 395.850 202.200 397.950 203.700 ;
        RECT 398.850 203.400 400.650 205.200 ;
        RECT 422.250 204.600 423.450 211.950 ;
        RECT 440.100 210.150 441.900 211.950 ;
        RECT 443.700 206.700 444.900 211.950 ;
        RECT 445.950 210.150 447.750 211.950 ;
        RECT 401.850 203.550 403.650 204.300 ;
        RECT 401.850 202.500 406.800 203.550 ;
        RECT 395.850 201.600 399.750 202.200 ;
        RECT 405.750 201.600 406.800 202.500 ;
        RECT 413.250 201.600 415.650 203.700 ;
        RECT 396.150 200.700 399.750 201.600 ;
        RECT 397.950 198.600 399.750 200.700 ;
        RECT 402.450 198.000 404.250 201.600 ;
        RECT 405.750 198.600 407.550 201.600 ;
        RECT 408.750 198.000 410.550 201.600 ;
        RECT 413.250 198.600 415.050 201.600 ;
        RECT 418.350 198.000 420.150 204.600 ;
        RECT 421.650 198.600 423.450 204.600 ;
        RECT 440.700 205.800 444.900 206.700 ;
        RECT 440.700 198.600 442.500 205.800 ;
        RECT 449.550 204.600 450.750 211.950 ;
        RECT 462.150 208.200 463.050 220.800 ;
        RECT 465.150 220.800 466.050 222.900 ;
        RECT 466.950 222.300 474.750 223.500 ;
        RECT 466.950 221.700 468.750 222.300 ;
        RECT 478.050 221.400 479.850 234.000 ;
        RECT 481.050 223.200 482.850 233.400 ;
        RECT 497.100 227.400 498.900 234.000 ;
        RECT 500.100 227.400 501.900 233.400 ;
        RECT 503.100 227.400 504.900 234.000 ;
        RECT 518.100 227.400 519.900 233.400 ;
        RECT 521.100 227.400 522.900 234.000 ;
        RECT 481.050 221.400 483.450 223.200 ;
        RECT 465.150 220.500 473.550 220.800 ;
        RECT 482.550 220.500 483.450 221.400 ;
        RECT 465.150 219.900 483.450 220.500 ;
        RECT 471.750 219.300 483.450 219.900 ;
        RECT 471.750 219.000 473.550 219.300 ;
        RECT 469.800 212.400 471.900 214.050 ;
        RECT 469.800 211.200 477.900 212.400 ;
        RECT 478.950 211.950 481.050 214.050 ;
        RECT 476.100 210.600 477.900 211.200 ;
        RECT 473.100 209.400 474.900 210.000 ;
        RECT 479.250 209.400 481.050 211.950 ;
        RECT 473.100 208.200 481.050 209.400 ;
        RECT 462.150 207.000 474.150 208.200 ;
        RECT 462.150 206.400 463.950 207.000 ;
        RECT 473.100 205.200 474.150 207.000 ;
        RECT 445.800 198.000 447.600 204.600 ;
        RECT 449.550 198.600 451.350 204.600 ;
        RECT 452.850 198.000 454.650 204.600 ;
        RECT 457.350 201.600 459.750 203.700 ;
        RECT 469.350 203.550 471.150 204.300 ;
        RECT 466.200 202.500 471.150 203.550 ;
        RECT 472.350 203.400 474.150 205.200 ;
        RECT 482.550 204.600 483.450 219.300 ;
        RECT 487.950 219.450 490.050 220.050 ;
        RECT 496.950 219.450 499.050 219.900 ;
        RECT 487.950 218.550 499.050 219.450 ;
        RECT 487.950 217.950 490.050 218.550 ;
        RECT 496.950 217.800 499.050 218.550 ;
        RECT 500.100 214.050 501.300 227.400 ;
        RECT 518.700 214.050 519.900 227.400 ;
        RECT 539.400 221.400 541.200 234.000 ;
        RECT 544.500 222.900 546.300 233.400 ;
        RECT 547.500 227.400 549.300 234.000 ;
        RECT 547.200 224.100 549.000 225.900 ;
        RECT 544.500 221.400 546.900 222.900 ;
        RECT 566.100 222.300 567.900 233.400 ;
        RECT 569.100 223.200 570.900 234.000 ;
        RECT 572.100 222.300 573.900 233.400 ;
        RECT 566.100 221.400 573.900 222.300 ;
        RECT 575.100 221.400 576.900 233.400 ;
        RECT 590.100 227.400 591.900 234.000 ;
        RECT 593.100 227.400 594.900 233.400 ;
        RECT 596.100 227.400 597.900 234.000 ;
        RECT 611.100 227.400 612.900 234.000 ;
        RECT 614.100 227.400 615.900 233.400 ;
        RECT 617.100 227.400 618.900 234.000 ;
        RECT 526.950 219.450 529.050 220.050 ;
        RECT 541.950 219.450 544.050 220.200 ;
        RECT 526.950 218.550 544.050 219.450 ;
        RECT 526.950 217.950 529.050 218.550 ;
        RECT 541.950 218.100 544.050 218.550 ;
        RECT 523.950 216.450 526.050 217.050 ;
        RECT 529.950 216.450 532.050 217.050 ;
        RECT 521.100 214.050 522.900 215.850 ;
        RECT 523.950 215.550 532.050 216.450 ;
        RECT 523.950 214.950 526.050 215.550 ;
        RECT 529.950 214.950 532.050 215.550 ;
        RECT 539.100 214.050 540.900 215.850 ;
        RECT 545.700 214.050 546.900 221.400 ;
        RECT 547.950 219.450 550.050 220.050 ;
        RECT 571.950 219.450 574.050 220.050 ;
        RECT 547.950 218.550 574.050 219.450 ;
        RECT 547.950 217.950 550.050 218.550 ;
        RECT 571.950 217.950 574.050 218.550 ;
        RECT 569.250 214.050 571.050 215.850 ;
        RECT 575.700 214.050 576.600 221.400 ;
        RECT 593.100 214.050 594.300 227.400 ;
        RECT 595.950 225.450 598.050 226.050 ;
        RECT 610.950 225.450 613.050 226.050 ;
        RECT 595.950 224.550 613.050 225.450 ;
        RECT 595.950 223.950 598.050 224.550 ;
        RECT 610.950 223.950 613.050 224.550 ;
        RECT 614.700 214.050 615.900 227.400 ;
        RECT 632.400 221.400 634.200 234.000 ;
        RECT 637.500 222.900 639.300 233.400 ;
        RECT 640.500 227.400 642.300 234.000 ;
        RECT 659.100 227.400 660.900 233.400 ;
        RECT 662.100 228.000 663.900 234.000 ;
        RECT 660.000 227.100 660.900 227.400 ;
        RECT 665.100 227.400 666.900 233.400 ;
        RECT 668.100 227.400 669.900 234.000 ;
        RECT 665.100 227.100 666.600 227.400 ;
        RECT 660.000 226.200 666.600 227.100 ;
        RECT 640.200 224.100 642.000 225.900 ;
        RECT 637.500 221.400 639.900 222.900 ;
        RECT 632.100 214.050 633.900 215.850 ;
        RECT 638.700 214.050 639.900 221.400 ;
        RECT 660.000 214.050 660.900 226.200 ;
        RECT 686.400 221.400 688.200 234.000 ;
        RECT 691.500 222.900 693.300 233.400 ;
        RECT 694.500 227.400 696.300 234.000 ;
        RECT 694.200 224.100 696.000 225.900 ;
        RECT 697.950 225.450 700.050 229.050 ;
        RECT 713.100 227.400 714.900 233.400 ;
        RECT 716.100 227.400 717.900 234.000 ;
        RECT 731.100 227.400 732.900 234.000 ;
        RECT 734.100 227.400 735.900 233.400 ;
        RECT 737.100 227.400 738.900 234.000 ;
        RECT 706.950 225.450 709.050 226.050 ;
        RECT 697.950 225.000 709.050 225.450 ;
        RECT 698.550 224.550 709.050 225.000 ;
        RECT 706.950 223.950 709.050 224.550 ;
        RECT 691.500 221.400 693.900 222.900 ;
        RECT 665.100 214.050 666.900 215.850 ;
        RECT 686.100 214.050 687.900 215.850 ;
        RECT 692.700 214.050 693.900 221.400 ;
        RECT 694.950 219.450 697.050 220.050 ;
        RECT 706.950 219.450 709.050 220.050 ;
        RECT 694.950 218.550 709.050 219.450 ;
        RECT 694.950 217.950 697.050 218.550 ;
        RECT 706.950 217.950 709.050 218.550 ;
        RECT 713.700 214.050 714.900 227.400 ;
        RECT 716.100 214.050 717.900 215.850 ;
        RECT 734.700 214.050 735.900 227.400 ;
        RECT 752.100 221.400 753.900 233.400 ;
        RECT 755.100 222.000 756.900 234.000 ;
        RECT 758.100 227.400 759.900 233.400 ;
        RECT 761.100 227.400 762.900 234.000 ;
        RECT 779.100 227.400 780.900 233.400 ;
        RECT 782.100 227.400 783.900 234.000 ;
        RECT 797.700 227.400 799.500 234.000 ;
        RECT 752.700 214.050 753.600 221.400 ;
        RECT 756.000 214.050 757.800 215.850 ;
        RECT 496.950 211.950 499.050 214.050 ;
        RECT 499.950 211.950 502.050 214.050 ;
        RECT 502.950 211.950 505.050 214.050 ;
        RECT 517.950 211.950 520.050 214.050 ;
        RECT 520.950 211.950 523.050 214.050 ;
        RECT 538.950 211.950 541.050 214.050 ;
        RECT 541.950 211.950 544.050 214.050 ;
        RECT 544.950 211.950 547.050 214.050 ;
        RECT 547.950 211.950 550.050 214.050 ;
        RECT 565.950 211.950 568.050 214.050 ;
        RECT 568.950 211.950 571.050 214.050 ;
        RECT 571.950 211.950 574.050 214.050 ;
        RECT 574.950 211.950 577.050 214.050 ;
        RECT 589.950 211.950 592.050 214.050 ;
        RECT 592.950 211.950 595.050 214.050 ;
        RECT 595.950 211.950 598.050 214.050 ;
        RECT 610.950 211.950 613.050 214.050 ;
        RECT 613.950 211.950 616.050 214.050 ;
        RECT 616.950 211.950 619.050 214.050 ;
        RECT 631.950 211.950 634.050 214.050 ;
        RECT 634.950 211.950 637.050 214.050 ;
        RECT 637.950 211.950 640.050 214.050 ;
        RECT 640.950 211.950 643.050 214.050 ;
        RECT 658.950 211.950 661.050 214.050 ;
        RECT 661.950 211.950 664.050 214.050 ;
        RECT 664.950 211.950 667.050 214.050 ;
        RECT 667.950 211.950 670.050 214.050 ;
        RECT 685.950 211.950 688.050 214.050 ;
        RECT 688.950 211.950 691.050 214.050 ;
        RECT 691.950 211.950 694.050 214.050 ;
        RECT 694.950 211.950 697.050 214.050 ;
        RECT 712.950 211.950 715.050 214.050 ;
        RECT 715.950 211.950 718.050 214.050 ;
        RECT 730.950 211.950 733.050 214.050 ;
        RECT 733.950 211.950 736.050 214.050 ;
        RECT 736.950 211.950 739.050 214.050 ;
        RECT 752.100 211.950 754.200 214.050 ;
        RECT 755.400 211.950 757.500 214.050 ;
        RECT 497.250 210.150 499.050 211.950 ;
        RECT 500.100 206.700 501.300 211.950 ;
        RECT 503.100 210.150 504.900 211.950 ;
        RECT 500.100 205.800 504.300 206.700 ;
        RECT 466.200 201.600 467.250 202.500 ;
        RECT 475.050 202.200 477.150 203.700 ;
        RECT 473.250 201.600 477.150 202.200 ;
        RECT 457.950 198.600 459.750 201.600 ;
        RECT 462.450 198.000 464.250 201.600 ;
        RECT 465.450 198.600 467.250 201.600 ;
        RECT 468.750 198.000 470.550 201.600 ;
        RECT 473.250 200.700 476.850 201.600 ;
        RECT 473.250 198.600 475.050 200.700 ;
        RECT 478.050 198.000 479.850 204.600 ;
        RECT 481.050 202.800 483.450 204.600 ;
        RECT 481.050 198.600 482.850 202.800 ;
        RECT 497.400 198.000 499.200 204.600 ;
        RECT 502.500 198.600 504.300 205.800 ;
        RECT 518.700 201.600 519.900 211.950 ;
        RECT 542.100 210.150 543.900 211.950 ;
        RECT 520.950 207.450 523.050 208.050 ;
        RECT 529.950 207.450 532.050 208.050 ;
        RECT 520.950 206.550 532.050 207.450 ;
        RECT 545.700 207.600 546.900 211.950 ;
        RECT 548.100 210.150 549.900 211.950 ;
        RECT 566.100 210.150 567.900 211.950 ;
        RECT 572.250 210.150 574.050 211.950 ;
        RECT 545.700 206.700 549.300 207.600 ;
        RECT 520.950 205.950 523.050 206.550 ;
        RECT 529.950 205.950 532.050 206.550 ;
        RECT 539.100 203.700 546.900 205.050 ;
        RECT 518.100 198.600 519.900 201.600 ;
        RECT 521.100 198.000 522.900 201.600 ;
        RECT 539.100 198.600 540.900 203.700 ;
        RECT 542.100 198.000 543.900 202.800 ;
        RECT 545.100 198.600 546.900 203.700 ;
        RECT 548.100 204.600 549.300 206.700 ;
        RECT 575.700 204.600 576.600 211.950 ;
        RECT 590.250 210.150 592.050 211.950 ;
        RECT 593.100 206.700 594.300 211.950 ;
        RECT 596.100 210.150 597.900 211.950 ;
        RECT 611.100 210.150 612.900 211.950 ;
        RECT 614.700 206.700 615.900 211.950 ;
        RECT 616.950 210.150 618.750 211.950 ;
        RECT 635.100 210.150 636.900 211.950 ;
        RECT 638.700 207.600 639.900 211.950 ;
        RECT 641.100 210.150 642.900 211.950 ;
        RECT 660.000 208.200 660.900 211.950 ;
        RECT 662.100 210.150 663.900 211.950 ;
        RECT 668.100 210.150 669.900 211.950 ;
        RECT 673.950 210.450 676.050 211.050 ;
        RECT 682.950 210.450 685.050 211.050 ;
        RECT 673.950 209.550 685.050 210.450 ;
        RECT 689.100 210.150 690.900 211.950 ;
        RECT 673.950 208.950 676.050 209.550 ;
        RECT 682.950 208.950 685.050 209.550 ;
        RECT 638.700 206.700 642.300 207.600 ;
        RECT 660.000 207.000 663.300 208.200 ;
        RECT 692.700 207.600 693.900 211.950 ;
        RECT 695.100 210.150 696.900 211.950 ;
        RECT 593.100 205.800 597.300 206.700 ;
        RECT 548.100 198.600 549.900 204.600 ;
        RECT 567.000 198.000 568.800 204.600 ;
        RECT 571.500 203.400 576.600 204.600 ;
        RECT 571.500 198.600 573.300 203.400 ;
        RECT 574.500 198.000 576.300 201.600 ;
        RECT 590.400 198.000 592.200 204.600 ;
        RECT 595.500 198.600 597.300 205.800 ;
        RECT 611.700 205.800 615.900 206.700 ;
        RECT 611.700 198.600 613.500 205.800 ;
        RECT 616.800 198.000 618.600 204.600 ;
        RECT 632.100 203.700 639.900 205.050 ;
        RECT 632.100 198.600 633.900 203.700 ;
        RECT 635.100 198.000 636.900 202.800 ;
        RECT 638.100 198.600 639.900 203.700 ;
        RECT 641.100 204.600 642.300 206.700 ;
        RECT 641.100 198.600 642.900 204.600 ;
        RECT 661.500 198.600 663.300 207.000 ;
        RECT 668.100 198.000 669.900 207.600 ;
        RECT 692.700 206.700 696.300 207.600 ;
        RECT 686.100 203.700 693.900 205.050 ;
        RECT 686.100 198.600 687.900 203.700 ;
        RECT 689.100 198.000 690.900 202.800 ;
        RECT 692.100 198.600 693.900 203.700 ;
        RECT 695.100 204.600 696.300 206.700 ;
        RECT 695.100 198.600 696.900 204.600 ;
        RECT 713.700 201.600 714.900 211.950 ;
        RECT 731.100 210.150 732.900 211.950 ;
        RECT 734.700 206.700 735.900 211.950 ;
        RECT 736.950 210.150 738.750 211.950 ;
        RECT 731.700 205.800 735.900 206.700 ;
        RECT 713.100 198.600 714.900 201.600 ;
        RECT 716.100 198.000 717.900 201.600 ;
        RECT 731.700 198.600 733.500 205.800 ;
        RECT 752.700 204.600 753.600 211.950 ;
        RECT 759.000 207.300 759.900 227.400 ;
        RECT 779.700 214.050 780.900 227.400 ;
        RECT 798.000 224.100 799.800 225.900 ;
        RECT 800.700 222.900 802.500 233.400 ;
        RECT 800.100 221.400 802.500 222.900 ;
        RECT 805.800 221.400 807.600 234.000 ;
        RECT 824.400 221.400 826.200 234.000 ;
        RECT 829.500 222.900 831.300 233.400 ;
        RECT 832.500 227.400 834.300 234.000 ;
        RECT 848.100 227.400 849.900 234.000 ;
        RECT 851.100 227.400 852.900 233.400 ;
        RECT 866.100 227.400 867.900 233.400 ;
        RECT 869.100 228.000 870.900 234.000 ;
        RECT 832.200 224.100 834.000 225.900 ;
        RECT 829.500 221.400 831.900 222.900 ;
        RECT 782.100 214.050 783.900 215.850 ;
        RECT 800.100 214.050 801.300 221.400 ;
        RECT 802.950 219.450 805.050 220.050 ;
        RECT 826.950 219.450 829.050 220.050 ;
        RECT 802.950 218.550 829.050 219.450 ;
        RECT 802.950 217.950 805.050 218.550 ;
        RECT 826.950 217.950 829.050 218.550 ;
        RECT 806.100 214.050 807.900 215.850 ;
        RECT 824.100 214.050 825.900 215.850 ;
        RECT 830.700 214.050 831.900 221.400 ;
        RECT 848.100 214.050 849.900 215.850 ;
        RECT 851.100 214.050 852.300 227.400 ;
        RECT 867.000 227.100 867.900 227.400 ;
        RECT 872.100 227.400 873.900 233.400 ;
        RECT 875.100 227.400 876.900 234.000 ;
        RECT 872.100 227.100 873.600 227.400 ;
        RECT 867.000 226.200 873.600 227.100 ;
        RECT 867.000 214.050 867.900 226.200 ;
        RECT 893.100 221.400 894.900 233.400 ;
        RECT 896.100 222.300 897.900 233.400 ;
        RECT 899.100 223.200 900.900 234.000 ;
        RECT 902.100 222.300 903.900 233.400 ;
        RECT 920.100 227.400 921.900 233.400 ;
        RECT 923.100 228.000 924.900 234.000 ;
        RECT 896.100 221.400 903.900 222.300 ;
        RECT 921.000 227.100 921.900 227.400 ;
        RECT 926.100 227.400 927.900 233.400 ;
        RECT 929.100 227.400 930.900 234.000 ;
        RECT 947.100 227.400 948.900 233.400 ;
        RECT 950.100 228.000 951.900 234.000 ;
        RECT 926.100 227.100 927.600 227.400 ;
        RECT 921.000 226.200 927.600 227.100 ;
        RECT 948.000 227.100 948.900 227.400 ;
        RECT 953.100 227.400 954.900 233.400 ;
        RECT 956.100 227.400 957.900 234.000 ;
        RECT 971.100 227.400 972.900 233.400 ;
        RECT 974.100 228.000 975.900 234.000 ;
        RECT 953.100 227.100 954.600 227.400 ;
        RECT 948.000 226.200 954.600 227.100 ;
        RECT 972.000 227.100 972.900 227.400 ;
        RECT 977.100 227.400 978.900 233.400 ;
        RECT 980.100 227.400 981.900 234.000 ;
        RECT 977.100 227.100 978.600 227.400 ;
        RECT 972.000 226.200 978.600 227.100 ;
        RECT 872.100 214.050 873.900 215.850 ;
        RECT 893.400 214.050 894.300 221.400 ;
        RECT 898.950 214.050 900.750 215.850 ;
        RECT 921.000 214.050 921.900 226.200 ;
        RECT 926.100 214.050 927.900 215.850 ;
        RECT 948.000 214.050 948.900 226.200 ;
        RECT 949.950 219.450 952.050 219.900 ;
        RECT 961.800 219.450 963.900 220.050 ;
        RECT 949.950 218.550 963.900 219.450 ;
        RECT 949.950 217.800 952.050 218.550 ;
        RECT 961.800 217.950 963.900 218.550 ;
        RECT 964.950 217.950 967.050 220.050 ;
        RECT 953.100 214.050 954.900 215.850 ;
        RECT 760.800 211.950 762.900 214.050 ;
        RECT 778.950 211.950 781.050 214.050 ;
        RECT 781.950 211.950 784.050 214.050 ;
        RECT 796.950 211.950 799.050 214.050 ;
        RECT 799.950 211.950 802.050 214.050 ;
        RECT 802.950 211.950 805.050 214.050 ;
        RECT 805.950 211.950 808.050 214.050 ;
        RECT 823.950 211.950 826.050 214.050 ;
        RECT 826.950 211.950 829.050 214.050 ;
        RECT 829.950 211.950 832.050 214.050 ;
        RECT 832.950 211.950 835.050 214.050 ;
        RECT 847.950 211.950 850.050 214.050 ;
        RECT 850.950 211.950 853.050 214.050 ;
        RECT 865.950 211.950 868.050 214.050 ;
        RECT 868.950 211.950 871.050 214.050 ;
        RECT 871.950 211.950 874.050 214.050 ;
        RECT 874.950 211.950 877.050 214.050 ;
        RECT 892.950 211.950 895.050 214.050 ;
        RECT 895.950 211.950 898.050 214.050 ;
        RECT 898.950 211.950 901.050 214.050 ;
        RECT 901.950 211.950 904.050 214.050 ;
        RECT 919.950 211.950 922.050 214.050 ;
        RECT 922.950 211.950 925.050 214.050 ;
        RECT 925.950 211.950 928.050 214.050 ;
        RECT 928.950 211.950 931.050 214.050 ;
        RECT 946.950 211.950 949.050 214.050 ;
        RECT 949.950 211.950 952.050 214.050 ;
        RECT 952.950 211.950 955.050 214.050 ;
        RECT 955.950 211.950 958.050 214.050 ;
        RECT 760.950 210.150 762.750 211.950 ;
        RECT 754.500 206.400 762.900 207.300 ;
        RECT 754.500 205.500 756.300 206.400 ;
        RECT 736.800 198.000 738.600 204.600 ;
        RECT 752.700 202.800 755.400 204.600 ;
        RECT 753.600 198.600 755.400 202.800 ;
        RECT 756.600 198.000 758.400 204.600 ;
        RECT 761.100 198.600 762.900 206.400 ;
        RECT 779.700 201.600 780.900 211.950 ;
        RECT 797.100 210.150 798.900 211.950 ;
        RECT 800.100 207.600 801.300 211.950 ;
        RECT 803.100 210.150 804.900 211.950 ;
        RECT 827.100 210.150 828.900 211.950 ;
        RECT 797.700 206.700 801.300 207.600 ;
        RECT 830.700 207.600 831.900 211.950 ;
        RECT 833.100 210.150 834.900 211.950 ;
        RECT 830.700 206.700 834.300 207.600 ;
        RECT 797.700 204.600 798.900 206.700 ;
        RECT 779.100 198.600 780.900 201.600 ;
        RECT 782.100 198.000 783.900 201.600 ;
        RECT 797.100 198.600 798.900 204.600 ;
        RECT 800.100 203.700 807.900 205.050 ;
        RECT 800.100 198.600 801.900 203.700 ;
        RECT 803.100 198.000 804.900 202.800 ;
        RECT 806.100 198.600 807.900 203.700 ;
        RECT 824.100 203.700 831.900 205.050 ;
        RECT 811.950 201.450 814.050 202.050 ;
        RECT 817.950 201.450 820.050 201.900 ;
        RECT 811.950 200.550 820.050 201.450 ;
        RECT 811.950 199.950 814.050 200.550 ;
        RECT 817.950 199.800 820.050 200.550 ;
        RECT 824.100 198.600 825.900 203.700 ;
        RECT 827.100 198.000 828.900 202.800 ;
        RECT 830.100 198.600 831.900 203.700 ;
        RECT 833.100 204.600 834.300 206.700 ;
        RECT 838.950 207.450 841.050 208.050 ;
        RECT 847.950 207.450 850.050 208.050 ;
        RECT 838.950 206.550 850.050 207.450 ;
        RECT 838.950 205.950 841.050 206.550 ;
        RECT 847.950 205.950 850.050 206.550 ;
        RECT 833.100 198.600 834.900 204.600 ;
        RECT 851.100 201.600 852.300 211.950 ;
        RECT 867.000 208.200 867.900 211.950 ;
        RECT 869.100 210.150 870.900 211.950 ;
        RECT 875.100 210.150 876.900 211.950 ;
        RECT 867.000 207.000 870.300 208.200 ;
        RECT 848.100 198.000 849.900 201.600 ;
        RECT 851.100 198.600 852.900 201.600 ;
        RECT 856.950 201.450 859.050 202.050 ;
        RECT 862.950 201.450 865.050 202.050 ;
        RECT 856.950 200.550 865.050 201.450 ;
        RECT 856.950 199.950 859.050 200.550 ;
        RECT 862.950 199.950 865.050 200.550 ;
        RECT 868.500 198.600 870.300 207.000 ;
        RECT 875.100 198.000 876.900 207.600 ;
        RECT 893.400 204.600 894.300 211.950 ;
        RECT 895.950 210.150 897.750 211.950 ;
        RECT 902.100 210.150 903.900 211.950 ;
        RECT 921.000 208.200 921.900 211.950 ;
        RECT 923.100 210.150 924.900 211.950 ;
        RECT 929.100 210.150 930.900 211.950 ;
        RECT 948.000 208.200 948.900 211.950 ;
        RECT 950.100 210.150 951.900 211.950 ;
        RECT 956.100 210.150 957.900 211.950 ;
        RECT 965.550 211.050 966.450 217.950 ;
        RECT 972.000 214.050 972.900 226.200 ;
        RECT 998.100 221.400 999.900 233.400 ;
        RECT 1001.100 222.300 1002.900 233.400 ;
        RECT 1004.100 223.200 1005.900 234.000 ;
        RECT 1007.100 222.300 1008.900 233.400 ;
        RECT 1001.100 221.400 1008.900 222.300 ;
        RECT 977.100 214.050 978.900 215.850 ;
        RECT 998.400 214.050 999.300 221.400 ;
        RECT 1009.950 216.450 1014.000 217.050 ;
        RECT 1003.950 214.050 1005.750 215.850 ;
        RECT 1009.950 214.950 1014.450 216.450 ;
        RECT 970.950 211.950 973.050 214.050 ;
        RECT 973.950 211.950 976.050 214.050 ;
        RECT 976.950 211.950 979.050 214.050 ;
        RECT 979.950 211.950 982.050 214.050 ;
        RECT 997.950 211.950 1000.050 214.050 ;
        RECT 1000.950 211.950 1003.050 214.050 ;
        RECT 1003.950 211.950 1006.050 214.050 ;
        RECT 1006.950 211.950 1009.050 214.050 ;
        RECT 965.550 209.550 970.050 211.050 ;
        RECT 966.000 208.950 970.050 209.550 ;
        RECT 972.000 208.200 972.900 211.950 ;
        RECT 974.100 210.150 975.900 211.950 ;
        RECT 980.100 210.150 981.900 211.950 ;
        RECT 982.950 210.450 985.050 211.050 ;
        RECT 991.950 210.450 994.050 211.050 ;
        RECT 982.950 209.550 994.050 210.450 ;
        RECT 982.950 208.950 985.050 209.550 ;
        RECT 991.950 208.950 994.050 209.550 ;
        RECT 921.000 207.000 924.300 208.200 ;
        RECT 893.400 203.400 898.500 204.600 ;
        RECT 893.700 198.000 895.500 201.600 ;
        RECT 896.700 198.600 898.500 203.400 ;
        RECT 901.200 198.000 903.000 204.600 ;
        RECT 922.500 198.600 924.300 207.000 ;
        RECT 929.100 198.000 930.900 207.600 ;
        RECT 948.000 207.000 951.300 208.200 ;
        RECT 949.500 198.600 951.300 207.000 ;
        RECT 956.100 198.000 957.900 207.600 ;
        RECT 972.000 207.000 975.300 208.200 ;
        RECT 973.500 198.600 975.300 207.000 ;
        RECT 980.100 198.000 981.900 207.600 ;
        RECT 998.400 204.600 999.300 211.950 ;
        RECT 1000.950 210.150 1002.750 211.950 ;
        RECT 1007.100 210.150 1008.900 211.950 ;
        RECT 1013.550 211.050 1014.450 214.950 ;
        RECT 1009.950 209.550 1014.450 211.050 ;
        RECT 1009.950 208.950 1014.000 209.550 ;
        RECT 998.400 203.400 1003.500 204.600 ;
        RECT 998.700 198.000 1000.500 201.600 ;
        RECT 1001.700 198.600 1003.500 203.400 ;
        RECT 1006.200 198.000 1008.000 204.600 ;
        RECT 14.700 187.200 16.500 194.400 ;
        RECT 19.800 188.400 21.600 195.000 ;
        RECT 38.700 187.200 40.500 194.400 ;
        RECT 43.800 188.400 45.600 195.000 ;
        RECT 59.700 191.400 61.500 195.000 ;
        RECT 62.700 189.600 64.500 194.400 ;
        RECT 59.400 188.400 64.500 189.600 ;
        RECT 67.200 188.400 69.000 195.000 ;
        RECT 14.700 186.300 18.900 187.200 ;
        RECT 38.700 186.300 42.900 187.200 ;
        RECT 14.100 181.050 15.900 182.850 ;
        RECT 17.700 181.050 18.900 186.300 ;
        RECT 19.950 181.050 21.750 182.850 ;
        RECT 38.100 181.050 39.900 182.850 ;
        RECT 41.700 181.050 42.900 186.300 ;
        RECT 49.950 183.450 52.050 184.050 ;
        RECT 55.950 183.450 58.050 184.050 ;
        RECT 43.950 181.050 45.750 182.850 ;
        RECT 49.950 182.550 58.050 183.450 ;
        RECT 49.950 181.950 52.050 182.550 ;
        RECT 55.950 181.950 58.050 182.550 ;
        RECT 59.400 181.050 60.300 188.400 ;
        RECT 83.100 185.400 84.900 195.000 ;
        RECT 89.700 186.000 91.500 194.400 ;
        RECT 107.100 191.400 108.900 195.000 ;
        RECT 110.100 191.400 111.900 194.400 ;
        RECT 113.100 191.400 114.900 195.000 ;
        RECT 89.700 184.800 93.000 186.000 ;
        RECT 61.950 181.050 63.750 182.850 ;
        RECT 68.100 181.050 69.900 182.850 ;
        RECT 83.100 181.050 84.900 182.850 ;
        RECT 89.100 181.050 90.900 182.850 ;
        RECT 92.100 181.050 93.000 184.800 ;
        RECT 110.700 181.050 111.600 191.400 ;
        RECT 128.100 189.300 129.900 194.400 ;
        RECT 131.100 190.200 132.900 195.000 ;
        RECT 134.100 189.300 135.900 194.400 ;
        RECT 128.100 187.950 135.900 189.300 ;
        RECT 137.100 188.400 138.900 194.400 ;
        RECT 137.100 186.300 138.300 188.400 ;
        RECT 152.700 187.200 154.500 194.400 ;
        RECT 157.800 188.400 159.600 195.000 ;
        RECT 173.100 191.400 174.900 195.000 ;
        RECT 176.100 191.400 177.900 194.400 ;
        RECT 152.700 186.300 156.900 187.200 ;
        RECT 134.700 185.400 138.300 186.300 ;
        RECT 131.100 181.050 132.900 182.850 ;
        RECT 134.700 181.050 135.900 185.400 ;
        RECT 137.100 181.050 138.900 182.850 ;
        RECT 152.100 181.050 153.900 182.850 ;
        RECT 155.700 181.050 156.900 186.300 ;
        RECT 160.950 183.450 163.050 184.050 ;
        RECT 166.950 183.450 169.050 184.050 ;
        RECT 157.950 181.050 159.750 182.850 ;
        RECT 160.950 182.550 169.050 183.450 ;
        RECT 160.950 181.950 163.050 182.550 ;
        RECT 166.950 181.950 169.050 182.550 ;
        RECT 176.100 181.050 177.300 191.400 ;
        RECT 194.100 185.400 195.900 195.000 ;
        RECT 200.700 186.000 202.500 194.400 ;
        RECT 218.100 188.400 219.900 194.400 ;
        RECT 218.700 186.300 219.900 188.400 ;
        RECT 221.100 189.300 222.900 194.400 ;
        RECT 224.100 190.200 225.900 195.000 ;
        RECT 227.100 189.300 228.900 194.400 ;
        RECT 245.100 191.400 246.900 194.400 ;
        RECT 248.100 191.400 249.900 195.000 ;
        RECT 221.100 187.950 228.900 189.300 ;
        RECT 200.700 184.800 204.000 186.000 ;
        RECT 218.700 185.400 222.300 186.300 ;
        RECT 194.100 181.050 195.900 182.850 ;
        RECT 200.100 181.050 201.900 182.850 ;
        RECT 203.100 181.050 204.000 184.800 ;
        RECT 205.950 183.450 208.050 184.050 ;
        RECT 211.950 183.450 214.050 184.050 ;
        RECT 205.950 182.550 214.050 183.450 ;
        RECT 205.950 181.950 208.050 182.550 ;
        RECT 211.950 181.950 214.050 182.550 ;
        RECT 218.100 181.050 219.900 182.850 ;
        RECT 221.100 181.050 222.300 185.400 ;
        RECT 224.100 181.050 225.900 182.850 ;
        RECT 245.700 181.050 246.900 191.400 ;
        RECT 263.700 187.200 265.500 194.400 ;
        RECT 268.800 188.400 270.600 195.000 ;
        RECT 287.400 188.400 289.200 195.000 ;
        RECT 292.500 187.200 294.300 194.400 ;
        RECT 308.100 189.300 309.900 194.400 ;
        RECT 311.100 190.200 312.900 195.000 ;
        RECT 314.100 189.300 315.900 194.400 ;
        RECT 308.100 187.950 315.900 189.300 ;
        RECT 317.100 188.400 318.900 194.400 ;
        RECT 332.400 188.400 334.200 195.000 ;
        RECT 263.700 186.300 267.900 187.200 ;
        RECT 263.100 181.050 264.900 182.850 ;
        RECT 266.700 181.050 267.900 186.300 ;
        RECT 290.100 186.300 294.300 187.200 ;
        RECT 317.100 186.300 318.300 188.400 ;
        RECT 337.500 187.200 339.300 194.400 ;
        RECT 353.100 188.400 354.900 194.400 ;
        RECT 268.950 181.050 270.750 182.850 ;
        RECT 287.250 181.050 289.050 182.850 ;
        RECT 290.100 181.050 291.300 186.300 ;
        RECT 314.700 185.400 318.300 186.300 ;
        RECT 335.100 186.300 339.300 187.200 ;
        RECT 353.700 186.300 354.900 188.400 ;
        RECT 356.100 189.300 357.900 194.400 ;
        RECT 359.100 190.200 360.900 195.000 ;
        RECT 362.100 189.300 363.900 194.400 ;
        RECT 356.100 187.950 363.900 189.300 ;
        RECT 380.400 188.400 382.200 195.000 ;
        RECT 385.500 187.200 387.300 194.400 ;
        RECT 401.100 188.400 402.900 194.400 ;
        RECT 383.100 186.300 387.300 187.200 ;
        RECT 401.700 186.300 402.900 188.400 ;
        RECT 404.100 189.300 405.900 194.400 ;
        RECT 407.100 190.200 408.900 195.000 ;
        RECT 410.100 189.300 411.900 194.400 ;
        RECT 404.100 187.950 411.900 189.300 ;
        RECT 428.700 187.200 430.500 194.400 ;
        RECT 433.800 188.400 435.600 195.000 ;
        RECT 449.700 187.200 451.500 194.400 ;
        RECT 454.800 188.400 456.600 195.000 ;
        RECT 473.100 188.400 474.900 194.400 ;
        RECT 428.700 186.300 432.900 187.200 ;
        RECT 449.700 186.300 453.900 187.200 ;
        RECT 293.100 181.050 294.900 182.850 ;
        RECT 311.100 181.050 312.900 182.850 ;
        RECT 314.700 181.050 315.900 185.400 ;
        RECT 317.100 181.050 318.900 182.850 ;
        RECT 332.250 181.050 334.050 182.850 ;
        RECT 335.100 181.050 336.300 186.300 ;
        RECT 353.700 185.400 357.300 186.300 ;
        RECT 338.100 181.050 339.900 182.850 ;
        RECT 353.100 181.050 354.900 182.850 ;
        RECT 356.100 181.050 357.300 185.400 ;
        RECT 359.100 181.050 360.900 182.850 ;
        RECT 380.250 181.050 382.050 182.850 ;
        RECT 383.100 181.050 384.300 186.300 ;
        RECT 401.700 185.400 405.300 186.300 ;
        RECT 386.100 181.050 387.900 182.850 ;
        RECT 401.100 181.050 402.900 182.850 ;
        RECT 404.100 181.050 405.300 185.400 ;
        RECT 407.100 181.050 408.900 182.850 ;
        RECT 428.100 181.050 429.900 182.850 ;
        RECT 431.700 181.050 432.900 186.300 ;
        RECT 433.950 181.050 435.750 182.850 ;
        RECT 449.100 181.050 450.900 182.850 ;
        RECT 452.700 181.050 453.900 186.300 ;
        RECT 473.700 186.300 474.900 188.400 ;
        RECT 476.100 189.300 477.900 194.400 ;
        RECT 479.100 190.200 480.900 195.000 ;
        RECT 482.100 189.300 483.900 194.400 ;
        RECT 497.100 191.400 498.900 195.000 ;
        RECT 500.100 191.400 501.900 194.400 ;
        RECT 476.100 187.950 483.900 189.300 ;
        RECT 473.700 185.400 477.300 186.300 ;
        RECT 454.950 181.050 456.750 182.850 ;
        RECT 473.100 181.050 474.900 182.850 ;
        RECT 476.100 181.050 477.300 185.400 ;
        RECT 479.100 181.050 480.900 182.850 ;
        RECT 500.100 181.050 501.300 191.400 ;
        RECT 515.100 188.400 516.900 194.400 ;
        RECT 515.700 186.300 516.900 188.400 ;
        RECT 518.100 189.300 519.900 194.400 ;
        RECT 521.100 190.200 522.900 195.000 ;
        RECT 524.100 189.300 525.900 194.400 ;
        RECT 539.100 191.400 540.900 195.000 ;
        RECT 542.100 191.400 543.900 194.400 ;
        RECT 518.100 187.950 525.900 189.300 ;
        RECT 515.700 185.400 519.300 186.300 ;
        RECT 515.100 181.050 516.900 182.850 ;
        RECT 518.100 181.050 519.300 185.400 ;
        RECT 521.100 181.050 522.900 182.850 ;
        RECT 542.100 181.050 543.300 191.400 ;
        RECT 557.100 189.300 558.900 194.400 ;
        RECT 560.100 190.200 561.900 195.000 ;
        RECT 563.100 189.300 564.900 194.400 ;
        RECT 557.100 187.950 564.900 189.300 ;
        RECT 566.100 188.400 567.900 194.400 ;
        RECT 566.100 186.300 567.300 188.400 ;
        RECT 563.700 185.400 567.300 186.300 ;
        RECT 583.500 186.000 585.300 194.400 ;
        RECT 560.100 181.050 561.900 182.850 ;
        RECT 563.700 181.050 564.900 185.400 ;
        RECT 582.000 184.800 585.300 186.000 ;
        RECT 590.100 185.400 591.900 195.000 ;
        RECT 608.100 189.300 609.900 194.400 ;
        RECT 611.100 190.200 612.900 195.000 ;
        RECT 614.100 189.300 615.900 194.400 ;
        RECT 608.100 187.950 615.900 189.300 ;
        RECT 617.100 188.400 618.900 194.400 ;
        RECT 635.100 189.000 636.900 194.400 ;
        RECT 638.100 189.900 639.900 195.000 ;
        RECT 641.100 193.500 648.900 194.400 ;
        RECT 641.100 189.000 642.900 193.500 ;
        RECT 617.100 186.300 618.300 188.400 ;
        RECT 635.100 188.100 642.900 189.000 ;
        RECT 644.100 188.400 645.900 192.600 ;
        RECT 647.100 188.400 648.900 193.500 ;
        RECT 644.400 186.900 645.300 188.400 ;
        RECT 614.700 185.400 618.300 186.300 ;
        RECT 640.950 185.700 645.300 186.900 ;
        RECT 662.100 186.600 663.900 194.400 ;
        RECT 666.600 188.400 668.400 195.000 ;
        RECT 669.600 190.200 671.400 194.400 ;
        RECT 686.100 191.400 687.900 195.000 ;
        RECT 689.100 191.400 690.900 194.400 ;
        RECT 669.600 188.400 672.300 190.200 ;
        RECT 668.700 186.600 670.500 187.500 ;
        RECT 662.100 185.700 670.500 186.600 ;
        RECT 566.100 181.050 567.900 182.850 ;
        RECT 582.000 181.050 582.900 184.800 ;
        RECT 604.950 183.450 607.050 184.050 ;
        RECT 584.100 181.050 585.900 182.850 ;
        RECT 590.100 181.050 591.900 182.850 ;
        RECT 596.550 182.550 607.050 183.450 ;
        RECT 13.950 178.950 16.050 181.050 ;
        RECT 16.950 178.950 19.050 181.050 ;
        RECT 19.950 178.950 22.050 181.050 ;
        RECT 37.950 178.950 40.050 181.050 ;
        RECT 40.950 178.950 43.050 181.050 ;
        RECT 43.950 178.950 46.050 181.050 ;
        RECT 58.950 178.950 61.050 181.050 ;
        RECT 61.950 178.950 64.050 181.050 ;
        RECT 64.950 178.950 67.050 181.050 ;
        RECT 67.950 178.950 70.050 181.050 ;
        RECT 82.950 178.950 85.050 181.050 ;
        RECT 85.950 178.950 88.050 181.050 ;
        RECT 88.950 178.950 91.050 181.050 ;
        RECT 91.950 178.950 94.050 181.050 ;
        RECT 106.950 178.950 109.050 181.050 ;
        RECT 109.950 178.950 112.050 181.050 ;
        RECT 112.950 178.950 115.050 181.050 ;
        RECT 127.950 178.950 130.050 181.050 ;
        RECT 130.950 178.950 133.050 181.050 ;
        RECT 133.950 178.950 136.050 181.050 ;
        RECT 136.950 178.950 139.050 181.050 ;
        RECT 151.950 178.950 154.050 181.050 ;
        RECT 154.950 178.950 157.050 181.050 ;
        RECT 157.950 178.950 160.050 181.050 ;
        RECT 172.950 178.950 175.050 181.050 ;
        RECT 175.950 178.950 178.050 181.050 ;
        RECT 193.950 178.950 196.050 181.050 ;
        RECT 196.950 178.950 199.050 181.050 ;
        RECT 199.950 178.950 202.050 181.050 ;
        RECT 202.950 178.950 205.050 181.050 ;
        RECT 217.950 178.950 220.050 181.050 ;
        RECT 220.950 178.950 223.050 181.050 ;
        RECT 223.950 178.950 226.050 181.050 ;
        RECT 226.950 178.950 229.050 181.050 ;
        RECT 244.950 178.950 247.050 181.050 ;
        RECT 247.950 178.950 250.050 181.050 ;
        RECT 262.950 178.950 265.050 181.050 ;
        RECT 265.950 178.950 268.050 181.050 ;
        RECT 268.950 178.950 271.050 181.050 ;
        RECT 286.950 178.950 289.050 181.050 ;
        RECT 289.950 178.950 292.050 181.050 ;
        RECT 292.950 178.950 295.050 181.050 ;
        RECT 307.950 178.950 310.050 181.050 ;
        RECT 310.950 178.950 313.050 181.050 ;
        RECT 313.950 178.950 316.050 181.050 ;
        RECT 316.950 178.950 319.050 181.050 ;
        RECT 331.950 178.950 334.050 181.050 ;
        RECT 334.950 178.950 337.050 181.050 ;
        RECT 337.950 178.950 340.050 181.050 ;
        RECT 352.950 178.950 355.050 181.050 ;
        RECT 355.950 178.950 358.050 181.050 ;
        RECT 358.950 178.950 361.050 181.050 ;
        RECT 361.950 178.950 364.050 181.050 ;
        RECT 379.950 178.950 382.050 181.050 ;
        RECT 382.950 178.950 385.050 181.050 ;
        RECT 385.950 178.950 388.050 181.050 ;
        RECT 400.950 178.950 403.050 181.050 ;
        RECT 403.950 178.950 406.050 181.050 ;
        RECT 406.950 178.950 409.050 181.050 ;
        RECT 409.950 178.950 412.050 181.050 ;
        RECT 427.950 178.950 430.050 181.050 ;
        RECT 430.950 178.950 433.050 181.050 ;
        RECT 433.950 178.950 436.050 181.050 ;
        RECT 448.950 178.950 451.050 181.050 ;
        RECT 451.950 178.950 454.050 181.050 ;
        RECT 454.950 178.950 457.050 181.050 ;
        RECT 472.950 178.950 475.050 181.050 ;
        RECT 475.950 178.950 478.050 181.050 ;
        RECT 478.950 178.950 481.050 181.050 ;
        RECT 481.950 178.950 484.050 181.050 ;
        RECT 496.950 178.950 499.050 181.050 ;
        RECT 499.950 178.950 502.050 181.050 ;
        RECT 514.950 178.950 517.050 181.050 ;
        RECT 517.950 178.950 520.050 181.050 ;
        RECT 520.950 178.950 523.050 181.050 ;
        RECT 523.950 178.950 526.050 181.050 ;
        RECT 538.950 178.950 541.050 181.050 ;
        RECT 541.950 178.950 544.050 181.050 ;
        RECT 556.950 178.950 559.050 181.050 ;
        RECT 559.950 178.950 562.050 181.050 ;
        RECT 562.950 178.950 565.050 181.050 ;
        RECT 565.950 178.950 568.050 181.050 ;
        RECT 580.950 178.950 583.050 181.050 ;
        RECT 583.950 178.950 586.050 181.050 ;
        RECT 586.950 178.950 589.050 181.050 ;
        RECT 589.950 178.950 592.050 181.050 ;
        RECT 17.700 165.600 18.900 178.950 ;
        RECT 41.700 165.600 42.900 178.950 ;
        RECT 59.400 171.600 60.300 178.950 ;
        RECT 64.950 177.150 66.750 178.950 ;
        RECT 86.100 177.150 87.900 178.950 ;
        RECT 76.950 174.450 79.050 175.050 ;
        RECT 88.950 174.450 91.050 175.050 ;
        RECT 76.950 173.550 91.050 174.450 ;
        RECT 76.950 172.950 79.050 173.550 ;
        RECT 88.950 172.950 91.050 173.550 ;
        RECT 14.100 159.000 15.900 165.600 ;
        RECT 17.100 159.600 18.900 165.600 ;
        RECT 20.100 159.000 21.900 165.600 ;
        RECT 38.100 159.000 39.900 165.600 ;
        RECT 41.100 159.600 42.900 165.600 ;
        RECT 44.100 159.000 45.900 165.600 ;
        RECT 59.100 159.600 60.900 171.600 ;
        RECT 62.100 170.700 69.900 171.600 ;
        RECT 62.100 159.600 63.900 170.700 ;
        RECT 65.100 159.000 66.900 169.800 ;
        RECT 68.100 159.600 69.900 170.700 ;
        RECT 92.100 166.800 93.000 178.950 ;
        RECT 107.100 177.150 108.900 178.950 ;
        RECT 110.700 171.600 111.600 178.950 ;
        RECT 112.950 177.150 114.750 178.950 ;
        RECT 128.100 177.150 129.900 178.950 ;
        RECT 134.700 171.600 135.900 178.950 ;
        RECT 86.400 165.900 93.000 166.800 ;
        RECT 86.400 165.600 87.900 165.900 ;
        RECT 83.100 159.000 84.900 165.600 ;
        RECT 86.100 159.600 87.900 165.600 ;
        RECT 92.100 165.600 93.000 165.900 ;
        RECT 108.000 170.400 111.600 171.600 ;
        RECT 89.100 159.000 90.900 165.000 ;
        RECT 92.100 159.600 93.900 165.600 ;
        RECT 108.000 159.600 109.800 170.400 ;
        RECT 113.100 159.000 114.900 171.600 ;
        RECT 128.400 159.000 130.200 171.600 ;
        RECT 133.500 170.100 135.900 171.600 ;
        RECT 133.500 159.600 135.300 170.100 ;
        RECT 136.200 167.100 138.000 168.900 ;
        RECT 155.700 165.600 156.900 178.950 ;
        RECT 173.100 177.150 174.900 178.950 ;
        RECT 176.100 165.600 177.300 178.950 ;
        RECT 197.100 177.150 198.900 178.950 ;
        RECT 203.100 166.800 204.000 178.950 ;
        RECT 221.100 171.600 222.300 178.950 ;
        RECT 227.100 177.150 228.900 178.950 ;
        RECT 221.100 170.100 223.500 171.600 ;
        RECT 219.000 167.100 220.800 168.900 ;
        RECT 197.400 165.900 204.000 166.800 ;
        RECT 197.400 165.600 198.900 165.900 ;
        RECT 136.500 159.000 138.300 165.600 ;
        RECT 152.100 159.000 153.900 165.600 ;
        RECT 155.100 159.600 156.900 165.600 ;
        RECT 158.100 159.000 159.900 165.600 ;
        RECT 173.100 159.000 174.900 165.600 ;
        RECT 176.100 159.600 177.900 165.600 ;
        RECT 194.100 159.000 195.900 165.600 ;
        RECT 197.100 159.600 198.900 165.600 ;
        RECT 203.100 165.600 204.000 165.900 ;
        RECT 200.100 159.000 201.900 165.000 ;
        RECT 203.100 159.600 204.900 165.600 ;
        RECT 218.700 159.000 220.500 165.600 ;
        RECT 221.700 159.600 223.500 170.100 ;
        RECT 226.800 159.000 228.600 171.600 ;
        RECT 245.700 165.600 246.900 178.950 ;
        RECT 248.100 177.150 249.900 178.950 ;
        RECT 266.700 165.600 267.900 178.950 ;
        RECT 290.100 165.600 291.300 178.950 ;
        RECT 308.100 177.150 309.900 178.950 ;
        RECT 298.950 174.450 301.050 175.050 ;
        RECT 310.950 174.450 313.050 174.750 ;
        RECT 298.950 173.550 313.050 174.450 ;
        RECT 298.950 172.950 301.050 173.550 ;
        RECT 310.950 172.650 313.050 173.550 ;
        RECT 314.700 171.600 315.900 178.950 ;
        RECT 322.950 177.450 325.050 178.050 ;
        RECT 328.950 177.450 331.050 178.050 ;
        RECT 322.950 176.550 331.050 177.450 ;
        RECT 322.950 175.950 325.050 176.550 ;
        RECT 328.950 175.950 331.050 176.550 ;
        RECT 245.100 159.600 246.900 165.600 ;
        RECT 248.100 159.000 249.900 165.600 ;
        RECT 263.100 159.000 264.900 165.600 ;
        RECT 266.100 159.600 267.900 165.600 ;
        RECT 269.100 159.000 270.900 165.600 ;
        RECT 287.100 159.000 288.900 165.600 ;
        RECT 290.100 159.600 291.900 165.600 ;
        RECT 293.100 159.000 294.900 165.600 ;
        RECT 308.400 159.000 310.200 171.600 ;
        RECT 313.500 170.100 315.900 171.600 ;
        RECT 313.500 159.600 315.300 170.100 ;
        RECT 316.200 167.100 318.000 168.900 ;
        RECT 335.100 165.600 336.300 178.950 ;
        RECT 343.950 174.450 346.050 175.050 ;
        RECT 352.950 174.450 355.050 175.050 ;
        RECT 343.950 173.550 355.050 174.450 ;
        RECT 343.950 172.950 346.050 173.550 ;
        RECT 352.950 172.950 355.050 173.550 ;
        RECT 356.100 171.600 357.300 178.950 ;
        RECT 362.100 177.150 363.900 178.950 ;
        RECT 356.100 170.100 358.500 171.600 ;
        RECT 354.000 167.100 355.800 168.900 ;
        RECT 316.500 159.000 318.300 165.600 ;
        RECT 332.100 159.000 333.900 165.600 ;
        RECT 335.100 159.600 336.900 165.600 ;
        RECT 338.100 159.000 339.900 165.600 ;
        RECT 353.700 159.000 355.500 165.600 ;
        RECT 356.700 159.600 358.500 170.100 ;
        RECT 361.800 159.000 363.600 171.600 ;
        RECT 383.100 165.600 384.300 178.950 ;
        RECT 391.950 174.450 394.050 175.050 ;
        RECT 400.950 174.450 403.050 175.050 ;
        RECT 391.950 173.550 403.050 174.450 ;
        RECT 391.950 172.950 394.050 173.550 ;
        RECT 400.950 172.950 403.050 173.550 ;
        RECT 404.100 171.600 405.300 178.950 ;
        RECT 410.100 177.150 411.900 178.950 ;
        RECT 404.100 170.100 406.500 171.600 ;
        RECT 402.000 167.100 403.800 168.900 ;
        RECT 380.100 159.000 381.900 165.600 ;
        RECT 383.100 159.600 384.900 165.600 ;
        RECT 386.100 159.000 387.900 165.600 ;
        RECT 401.700 159.000 403.500 165.600 ;
        RECT 404.700 159.600 406.500 170.100 ;
        RECT 409.800 159.000 411.600 171.600 ;
        RECT 431.700 165.600 432.900 178.950 ;
        RECT 452.700 165.600 453.900 178.950 ;
        RECT 476.100 171.600 477.300 178.950 ;
        RECT 482.100 177.150 483.900 178.950 ;
        RECT 497.100 177.150 498.900 178.950 ;
        RECT 476.100 170.100 478.500 171.600 ;
        RECT 474.000 167.100 475.800 168.900 ;
        RECT 428.100 159.000 429.900 165.600 ;
        RECT 431.100 159.600 432.900 165.600 ;
        RECT 434.100 159.000 435.900 165.600 ;
        RECT 449.100 159.000 450.900 165.600 ;
        RECT 452.100 159.600 453.900 165.600 ;
        RECT 455.100 159.000 456.900 165.600 ;
        RECT 473.700 159.000 475.500 165.600 ;
        RECT 476.700 159.600 478.500 170.100 ;
        RECT 481.800 159.000 483.600 171.600 ;
        RECT 500.100 165.600 501.300 178.950 ;
        RECT 518.100 171.600 519.300 178.950 ;
        RECT 524.100 177.150 525.900 178.950 ;
        RECT 539.100 177.150 540.900 178.950 ;
        RECT 520.950 174.450 523.050 175.050 ;
        RECT 532.950 174.450 535.050 175.050 ;
        RECT 520.950 173.550 535.050 174.450 ;
        RECT 520.950 172.950 523.050 173.550 ;
        RECT 532.950 172.950 535.050 173.550 ;
        RECT 518.100 170.100 520.500 171.600 ;
        RECT 516.000 167.100 517.800 168.900 ;
        RECT 497.100 159.000 498.900 165.600 ;
        RECT 500.100 159.600 501.900 165.600 ;
        RECT 515.700 159.000 517.500 165.600 ;
        RECT 518.700 159.600 520.500 170.100 ;
        RECT 523.800 159.000 525.600 171.600 ;
        RECT 542.100 165.600 543.300 178.950 ;
        RECT 557.100 177.150 558.900 178.950 ;
        RECT 563.700 171.600 564.900 178.950 ;
        RECT 539.100 159.000 540.900 165.600 ;
        RECT 542.100 159.600 543.900 165.600 ;
        RECT 557.400 159.000 559.200 171.600 ;
        RECT 562.500 170.100 564.900 171.600 ;
        RECT 562.500 159.600 564.300 170.100 ;
        RECT 565.200 167.100 567.000 168.900 ;
        RECT 582.000 166.800 582.900 178.950 ;
        RECT 587.100 177.150 588.900 178.950 ;
        RECT 596.550 177.450 597.450 182.550 ;
        RECT 604.950 181.950 607.050 182.550 ;
        RECT 611.100 181.050 612.900 182.850 ;
        RECT 614.700 181.050 615.900 185.400 ;
        RECT 619.950 183.450 624.000 184.050 ;
        RECT 617.100 181.050 618.900 182.850 ;
        RECT 619.950 181.950 624.450 183.450 ;
        RECT 607.950 178.950 610.050 181.050 ;
        RECT 610.950 178.950 613.050 181.050 ;
        RECT 613.950 178.950 616.050 181.050 ;
        RECT 616.950 178.950 619.050 181.050 ;
        RECT 593.550 176.550 597.450 177.450 ;
        RECT 608.100 177.150 609.900 178.950 ;
        RECT 583.950 174.450 586.050 175.050 ;
        RECT 593.550 174.450 594.450 176.550 ;
        RECT 583.950 173.550 594.450 174.450 ;
        RECT 583.950 172.950 586.050 173.550 ;
        RECT 614.700 171.600 615.900 178.950 ;
        RECT 623.550 178.050 624.450 181.950 ;
        RECT 638.250 181.050 640.050 182.850 ;
        RECT 634.950 178.950 637.050 181.050 ;
        RECT 637.950 178.950 640.050 181.050 ;
        RECT 640.950 181.050 642.000 185.700 ;
        RECT 643.950 181.050 645.750 182.850 ;
        RECT 662.250 181.050 664.050 182.850 ;
        RECT 640.950 178.950 643.050 181.050 ;
        RECT 643.950 178.950 646.050 181.050 ;
        RECT 646.950 178.950 649.050 181.050 ;
        RECT 654.000 180.450 658.050 181.050 ;
        RECT 653.550 178.950 658.050 180.450 ;
        RECT 662.100 178.950 664.200 181.050 ;
        RECT 619.950 176.550 624.450 178.050 ;
        RECT 635.100 177.150 636.900 178.950 ;
        RECT 619.950 175.950 624.000 176.550 ;
        RECT 640.950 171.600 642.000 178.950 ;
        RECT 646.950 177.150 648.750 178.950 ;
        RECT 653.550 178.050 654.450 178.950 ;
        RECT 649.950 176.550 654.450 178.050 ;
        RECT 649.950 175.950 654.000 176.550 ;
        RECT 643.950 174.450 646.050 175.050 ;
        RECT 655.950 174.450 658.050 175.050 ;
        RECT 643.950 173.550 658.050 174.450 ;
        RECT 643.950 172.950 646.050 173.550 ;
        RECT 655.950 172.950 658.050 173.550 ;
        RECT 592.950 168.450 595.050 169.050 ;
        RECT 601.950 168.450 604.050 169.050 ;
        RECT 592.950 167.550 604.050 168.450 ;
        RECT 592.950 166.950 595.050 167.550 ;
        RECT 601.950 166.950 604.050 167.550 ;
        RECT 582.000 165.900 588.600 166.800 ;
        RECT 582.000 165.600 582.900 165.900 ;
        RECT 565.500 159.000 567.300 165.600 ;
        RECT 581.100 159.600 582.900 165.600 ;
        RECT 587.100 165.600 588.600 165.900 ;
        RECT 584.100 159.000 585.900 165.000 ;
        RECT 587.100 159.600 588.900 165.600 ;
        RECT 590.100 159.000 591.900 165.600 ;
        RECT 608.400 159.000 610.200 171.600 ;
        RECT 613.500 170.100 615.900 171.600 ;
        RECT 613.500 159.600 615.300 170.100 ;
        RECT 616.200 167.100 618.000 168.900 ;
        RECT 616.500 159.000 618.300 165.600 ;
        RECT 635.100 159.000 636.900 171.600 ;
        RECT 639.600 159.600 642.900 171.600 ;
        RECT 645.600 159.000 647.400 171.600 ;
        RECT 665.100 165.600 666.000 185.700 ;
        RECT 671.400 181.050 672.300 188.400 ;
        RECT 689.100 181.050 690.300 191.400 ;
        RECT 704.100 189.300 705.900 194.400 ;
        RECT 707.100 190.200 708.900 195.000 ;
        RECT 710.100 189.300 711.900 194.400 ;
        RECT 704.100 187.950 711.900 189.300 ;
        RECT 713.100 188.400 714.900 194.400 ;
        RECT 713.100 186.300 714.300 188.400 ;
        RECT 710.700 185.400 714.300 186.300 ;
        RECT 728.100 185.400 729.900 195.000 ;
        RECT 734.700 186.000 736.500 194.400 ;
        RECT 752.100 193.500 759.900 194.400 ;
        RECT 752.100 188.400 753.900 193.500 ;
        RECT 755.100 188.400 756.900 192.600 ;
        RECT 758.100 189.000 759.900 193.500 ;
        RECT 761.100 189.900 762.900 195.000 ;
        RECT 764.100 189.000 765.900 194.400 ;
        RECT 780.600 190.200 782.400 194.400 ;
        RECT 755.700 186.900 756.600 188.400 ;
        RECT 758.100 188.100 765.900 189.000 ;
        RECT 779.700 188.400 782.400 190.200 ;
        RECT 783.600 188.400 785.400 195.000 ;
        RECT 707.100 181.050 708.900 182.850 ;
        RECT 710.700 181.050 711.900 185.400 ;
        RECT 734.700 184.800 738.000 186.000 ;
        RECT 755.700 185.700 760.050 186.900 ;
        RECT 713.100 181.050 714.900 182.850 ;
        RECT 728.100 181.050 729.900 182.850 ;
        RECT 734.100 181.050 735.900 182.850 ;
        RECT 737.100 181.050 738.000 184.800 ;
        RECT 755.250 181.050 757.050 182.850 ;
        RECT 759.000 181.050 760.050 185.700 ;
        RECT 667.500 178.950 669.600 181.050 ;
        RECT 670.800 178.950 672.900 181.050 ;
        RECT 685.950 178.950 688.050 181.050 ;
        RECT 688.950 178.950 691.050 181.050 ;
        RECT 703.950 178.950 706.050 181.050 ;
        RECT 706.950 178.950 709.050 181.050 ;
        RECT 709.950 178.950 712.050 181.050 ;
        RECT 712.950 178.950 715.050 181.050 ;
        RECT 727.950 178.950 730.050 181.050 ;
        RECT 730.950 178.950 733.050 181.050 ;
        RECT 733.950 178.950 736.050 181.050 ;
        RECT 736.950 178.950 739.050 181.050 ;
        RECT 751.950 178.950 754.050 181.050 ;
        RECT 754.950 178.950 757.050 181.050 ;
        RECT 757.950 178.950 760.050 181.050 ;
        RECT 760.950 181.050 762.750 182.850 ;
        RECT 779.700 181.050 780.600 188.400 ;
        RECT 781.500 186.600 783.300 187.500 ;
        RECT 788.100 186.600 789.900 194.400 ;
        RECT 803.400 188.400 805.200 195.000 ;
        RECT 808.500 187.200 810.300 194.400 ;
        RECT 825.000 188.400 826.800 195.000 ;
        RECT 829.500 189.600 831.300 194.400 ;
        RECT 832.500 191.400 834.300 195.000 ;
        RECT 829.500 188.400 834.600 189.600 ;
        RECT 781.500 185.700 789.900 186.600 ;
        RECT 806.100 186.300 810.300 187.200 ;
        RECT 760.950 178.950 763.050 181.050 ;
        RECT 763.950 178.950 766.050 181.050 ;
        RECT 779.100 178.950 781.200 181.050 ;
        RECT 782.400 178.950 784.500 181.050 ;
        RECT 667.200 177.150 669.000 178.950 ;
        RECT 671.400 171.600 672.300 178.950 ;
        RECT 686.100 177.150 687.900 178.950 ;
        RECT 662.100 159.000 663.900 165.600 ;
        RECT 665.100 159.600 666.900 165.600 ;
        RECT 668.100 159.000 669.900 171.000 ;
        RECT 671.100 159.600 672.900 171.600 ;
        RECT 689.100 165.600 690.300 178.950 ;
        RECT 704.100 177.150 705.900 178.950 ;
        RECT 710.700 171.600 711.900 178.950 ;
        RECT 731.100 177.150 732.900 178.950 ;
        RECT 712.950 174.450 715.050 175.050 ;
        RECT 730.950 174.450 733.050 175.050 ;
        RECT 712.950 173.550 733.050 174.450 ;
        RECT 712.950 172.950 715.050 173.550 ;
        RECT 730.950 172.950 733.050 173.550 ;
        RECT 686.100 159.000 687.900 165.600 ;
        RECT 689.100 159.600 690.900 165.600 ;
        RECT 704.400 159.000 706.200 171.600 ;
        RECT 709.500 170.100 711.900 171.600 ;
        RECT 709.500 159.600 711.300 170.100 ;
        RECT 712.200 167.100 714.000 168.900 ;
        RECT 737.100 166.800 738.000 178.950 ;
        RECT 752.250 177.150 754.050 178.950 ;
        RECT 759.000 171.600 760.050 178.950 ;
        RECT 764.100 177.150 765.900 178.950 ;
        RECT 779.700 171.600 780.600 178.950 ;
        RECT 783.000 177.150 784.800 178.950 ;
        RECT 731.400 165.900 738.000 166.800 ;
        RECT 731.400 165.600 732.900 165.900 ;
        RECT 712.500 159.000 714.300 165.600 ;
        RECT 728.100 159.000 729.900 165.600 ;
        RECT 731.100 159.600 732.900 165.600 ;
        RECT 737.100 165.600 738.000 165.900 ;
        RECT 734.100 159.000 735.900 165.000 ;
        RECT 737.100 159.600 738.900 165.600 ;
        RECT 753.600 159.000 755.400 171.600 ;
        RECT 758.100 159.600 761.400 171.600 ;
        RECT 764.100 159.000 765.900 171.600 ;
        RECT 779.100 159.600 780.900 171.600 ;
        RECT 782.100 159.000 783.900 171.000 ;
        RECT 786.000 165.600 786.900 185.700 ;
        RECT 787.950 181.050 789.750 182.850 ;
        RECT 803.250 181.050 805.050 182.850 ;
        RECT 806.100 181.050 807.300 186.300 ;
        RECT 809.100 181.050 810.900 182.850 ;
        RECT 824.100 181.050 825.900 182.850 ;
        RECT 830.250 181.050 832.050 182.850 ;
        RECT 833.700 181.050 834.600 188.400 ;
        RECT 848.100 185.400 849.900 195.000 ;
        RECT 854.700 186.000 856.500 194.400 ;
        RECT 872.100 188.400 873.900 194.400 ;
        RECT 872.700 186.300 873.900 188.400 ;
        RECT 875.100 189.300 876.900 194.400 ;
        RECT 878.100 190.200 879.900 195.000 ;
        RECT 881.100 189.300 882.900 194.400 ;
        RECT 875.100 187.950 882.900 189.300 ;
        RECT 896.400 188.400 898.200 195.000 ;
        RECT 901.500 187.200 903.300 194.400 ;
        RECT 899.100 186.300 903.300 187.200 ;
        RECT 854.700 184.800 858.000 186.000 ;
        RECT 872.700 185.400 876.300 186.300 ;
        RECT 848.100 181.050 849.900 182.850 ;
        RECT 854.100 181.050 855.900 182.850 ;
        RECT 857.100 181.050 858.000 184.800 ;
        RECT 859.950 183.450 864.000 184.050 ;
        RECT 859.950 181.950 864.450 183.450 ;
        RECT 787.800 178.950 789.900 181.050 ;
        RECT 802.950 178.950 805.050 181.050 ;
        RECT 805.950 178.950 808.050 181.050 ;
        RECT 808.950 178.950 811.050 181.050 ;
        RECT 823.950 178.950 826.050 181.050 ;
        RECT 826.950 178.950 829.050 181.050 ;
        RECT 829.950 178.950 832.050 181.050 ;
        RECT 832.950 178.950 835.050 181.050 ;
        RECT 847.950 178.950 850.050 181.050 ;
        RECT 850.950 178.950 853.050 181.050 ;
        RECT 853.950 178.950 856.050 181.050 ;
        RECT 856.950 178.950 859.050 181.050 ;
        RECT 806.100 165.600 807.300 178.950 ;
        RECT 827.250 177.150 829.050 178.950 ;
        RECT 833.700 171.600 834.600 178.950 ;
        RECT 851.100 177.150 852.900 178.950 ;
        RECT 824.100 170.700 831.900 171.600 ;
        RECT 785.100 159.600 786.900 165.600 ;
        RECT 788.100 159.000 789.900 165.600 ;
        RECT 803.100 159.000 804.900 165.600 ;
        RECT 806.100 159.600 807.900 165.600 ;
        RECT 809.100 159.000 810.900 165.600 ;
        RECT 824.100 159.600 825.900 170.700 ;
        RECT 827.100 159.000 828.900 169.800 ;
        RECT 830.100 159.600 831.900 170.700 ;
        RECT 833.100 159.600 834.900 171.600 ;
        RECT 857.100 166.800 858.000 178.950 ;
        RECT 863.550 178.050 864.450 181.950 ;
        RECT 872.100 181.050 873.900 182.850 ;
        RECT 875.100 181.050 876.300 185.400 ;
        RECT 892.950 183.450 895.050 184.050 ;
        RECT 878.100 181.050 879.900 182.850 ;
        RECT 887.550 182.550 895.050 183.450 ;
        RECT 871.950 178.950 874.050 181.050 ;
        RECT 874.950 178.950 877.050 181.050 ;
        RECT 877.950 178.950 880.050 181.050 ;
        RECT 880.950 178.950 883.050 181.050 ;
        RECT 859.950 176.550 864.450 178.050 ;
        RECT 859.950 175.950 864.000 176.550 ;
        RECT 875.100 171.600 876.300 178.950 ;
        RECT 881.100 177.150 882.900 178.950 ;
        RECT 887.550 177.450 888.450 182.550 ;
        RECT 892.950 181.950 895.050 182.550 ;
        RECT 896.250 181.050 898.050 182.850 ;
        RECT 899.100 181.050 900.300 186.300 ;
        RECT 919.500 186.000 921.300 194.400 ;
        RECT 918.000 184.800 921.300 186.000 ;
        RECT 926.100 185.400 927.900 195.000 ;
        RECT 941.700 191.400 943.500 195.000 ;
        RECT 944.700 189.600 946.500 194.400 ;
        RECT 941.400 188.400 946.500 189.600 ;
        RECT 949.200 188.400 951.000 195.000 ;
        RECT 902.100 181.050 903.900 182.850 ;
        RECT 918.000 181.050 918.900 184.800 ;
        RECT 928.950 183.450 931.050 184.050 ;
        RECT 937.950 183.450 940.050 183.900 ;
        RECT 920.100 181.050 921.900 182.850 ;
        RECT 926.100 181.050 927.900 182.850 ;
        RECT 928.950 182.550 940.050 183.450 ;
        RECT 928.950 181.950 931.050 182.550 ;
        RECT 937.950 181.800 940.050 182.550 ;
        RECT 941.400 181.050 942.300 188.400 ;
        RECT 967.500 186.000 969.300 194.400 ;
        RECT 966.000 184.800 969.300 186.000 ;
        RECT 974.100 185.400 975.900 195.000 ;
        RECT 989.100 191.400 990.900 195.000 ;
        RECT 992.100 191.400 993.900 194.400 ;
        RECT 943.950 181.050 945.750 182.850 ;
        RECT 950.100 181.050 951.900 182.850 ;
        RECT 966.000 181.050 966.900 184.800 ;
        RECT 968.100 181.050 969.900 182.850 ;
        RECT 974.100 181.050 975.900 182.850 ;
        RECT 992.100 181.050 993.300 191.400 ;
        RECT 895.950 178.950 898.050 181.050 ;
        RECT 898.950 178.950 901.050 181.050 ;
        RECT 901.950 178.950 904.050 181.050 ;
        RECT 916.950 178.950 919.050 181.050 ;
        RECT 919.950 178.950 922.050 181.050 ;
        RECT 922.950 178.950 925.050 181.050 ;
        RECT 925.950 178.950 928.050 181.050 ;
        RECT 940.950 178.950 943.050 181.050 ;
        RECT 943.950 178.950 946.050 181.050 ;
        RECT 946.950 178.950 949.050 181.050 ;
        RECT 949.950 178.950 952.050 181.050 ;
        RECT 964.950 178.950 967.050 181.050 ;
        RECT 967.950 178.950 970.050 181.050 ;
        RECT 970.950 178.950 973.050 181.050 ;
        RECT 973.950 178.950 976.050 181.050 ;
        RECT 988.950 178.950 991.050 181.050 ;
        RECT 991.950 178.950 994.050 181.050 ;
        RECT 884.550 176.550 888.450 177.450 ;
        RECT 877.950 174.450 880.050 175.050 ;
        RECT 884.550 174.450 885.450 176.550 ;
        RECT 877.950 173.550 885.450 174.450 ;
        RECT 877.950 172.950 880.050 173.550 ;
        RECT 875.100 170.100 877.500 171.600 ;
        RECT 873.000 167.100 874.800 168.900 ;
        RECT 851.400 165.900 858.000 166.800 ;
        RECT 851.400 165.600 852.900 165.900 ;
        RECT 848.100 159.000 849.900 165.600 ;
        RECT 851.100 159.600 852.900 165.600 ;
        RECT 857.100 165.600 858.000 165.900 ;
        RECT 854.100 159.000 855.900 165.000 ;
        RECT 857.100 159.600 858.900 165.600 ;
        RECT 872.700 159.000 874.500 165.600 ;
        RECT 875.700 159.600 877.500 170.100 ;
        RECT 880.800 159.000 882.600 171.600 ;
        RECT 899.100 165.600 900.300 178.950 ;
        RECT 918.000 166.800 918.900 178.950 ;
        RECT 923.100 177.150 924.900 178.950 ;
        RECT 941.400 171.600 942.300 178.950 ;
        RECT 946.950 177.150 948.750 178.950 ;
        RECT 918.000 165.900 924.600 166.800 ;
        RECT 918.000 165.600 918.900 165.900 ;
        RECT 896.100 159.000 897.900 165.600 ;
        RECT 899.100 159.600 900.900 165.600 ;
        RECT 902.100 159.000 903.900 165.600 ;
        RECT 917.100 159.600 918.900 165.600 ;
        RECT 923.100 165.600 924.600 165.900 ;
        RECT 920.100 159.000 921.900 165.000 ;
        RECT 923.100 159.600 924.900 165.600 ;
        RECT 926.100 159.000 927.900 165.600 ;
        RECT 941.100 159.600 942.900 171.600 ;
        RECT 944.100 170.700 951.900 171.600 ;
        RECT 944.100 159.600 945.900 170.700 ;
        RECT 947.100 159.000 948.900 169.800 ;
        RECT 950.100 159.600 951.900 170.700 ;
        RECT 966.000 166.800 966.900 178.950 ;
        RECT 971.100 177.150 972.900 178.950 ;
        RECT 989.100 177.150 990.900 178.950 ;
        RECT 966.000 165.900 972.600 166.800 ;
        RECT 966.000 165.600 966.900 165.900 ;
        RECT 965.100 159.600 966.900 165.600 ;
        RECT 971.100 165.600 972.600 165.900 ;
        RECT 992.100 165.600 993.300 178.950 ;
        RECT 968.100 159.000 969.900 165.000 ;
        RECT 971.100 159.600 972.900 165.600 ;
        RECT 974.100 159.000 975.900 165.600 ;
        RECT 989.100 159.000 990.900 165.600 ;
        RECT 992.100 159.600 993.900 165.600 ;
        RECT 17.100 143.400 18.900 155.400 ;
        RECT 20.100 144.300 21.900 155.400 ;
        RECT 23.100 145.200 24.900 156.000 ;
        RECT 26.100 144.300 27.900 155.400 ;
        RECT 41.100 149.400 42.900 155.400 ;
        RECT 44.100 149.400 45.900 156.000 ;
        RECT 59.100 149.400 60.900 155.400 ;
        RECT 62.100 150.000 63.900 156.000 ;
        RECT 20.100 143.400 27.900 144.300 ;
        RECT 17.400 136.050 18.300 143.400 ;
        RECT 22.950 136.050 24.750 137.850 ;
        RECT 41.700 136.050 42.900 149.400 ;
        RECT 60.000 149.100 60.900 149.400 ;
        RECT 65.100 149.400 66.900 155.400 ;
        RECT 68.100 149.400 69.900 156.000 ;
        RECT 65.100 149.100 66.600 149.400 ;
        RECT 60.000 148.200 66.600 149.100 ;
        RECT 44.100 136.050 45.900 137.850 ;
        RECT 60.000 136.050 60.900 148.200 ;
        RECT 83.400 143.400 85.200 156.000 ;
        RECT 88.500 144.900 90.300 155.400 ;
        RECT 91.500 149.400 93.300 156.000 ;
        RECT 107.100 149.400 108.900 156.000 ;
        RECT 110.100 149.400 111.900 155.400 ;
        RECT 128.100 149.400 129.900 156.000 ;
        RECT 131.100 149.400 132.900 155.400 ;
        RECT 146.700 149.400 148.500 156.000 ;
        RECT 91.200 146.100 93.000 147.900 ;
        RECT 88.500 143.400 90.900 144.900 ;
        RECT 65.100 136.050 66.900 137.850 ;
        RECT 83.100 136.050 84.900 137.850 ;
        RECT 89.700 136.050 90.900 143.400 ;
        RECT 107.100 136.050 108.900 137.850 ;
        RECT 110.100 136.050 111.300 149.400 ;
        RECT 128.100 136.050 129.900 137.850 ;
        RECT 131.100 136.050 132.300 149.400 ;
        RECT 147.000 146.100 148.800 147.900 ;
        RECT 149.700 144.900 151.500 155.400 ;
        RECT 149.100 143.400 151.500 144.900 ;
        RECT 154.800 143.400 156.600 156.000 ;
        RECT 170.400 143.400 172.200 156.000 ;
        RECT 175.500 144.900 177.300 155.400 ;
        RECT 178.500 149.400 180.300 156.000 ;
        RECT 178.200 146.100 180.000 147.900 ;
        RECT 175.500 143.400 177.900 144.900 ;
        RECT 194.100 144.300 195.900 155.400 ;
        RECT 197.100 145.200 198.900 156.000 ;
        RECT 200.100 144.300 201.900 155.400 ;
        RECT 194.100 143.400 201.900 144.300 ;
        RECT 203.100 143.400 204.900 155.400 ;
        RECT 221.100 149.400 222.900 156.000 ;
        RECT 224.100 149.400 225.900 155.400 ;
        RECT 227.100 150.000 228.900 156.000 ;
        RECT 224.400 149.100 225.900 149.400 ;
        RECT 230.100 149.400 231.900 155.400 ;
        RECT 245.100 149.400 246.900 155.400 ;
        RECT 248.100 150.000 249.900 156.000 ;
        RECT 230.100 149.100 231.000 149.400 ;
        RECT 224.400 148.200 231.000 149.100 ;
        RECT 149.100 136.050 150.300 143.400 ;
        RECT 151.950 141.450 154.050 142.050 ;
        RECT 160.950 141.450 163.050 142.050 ;
        RECT 151.950 140.550 163.050 141.450 ;
        RECT 151.950 139.950 154.050 140.550 ;
        RECT 160.950 139.950 163.050 140.550 ;
        RECT 155.100 136.050 156.900 137.850 ;
        RECT 170.100 136.050 171.900 137.850 ;
        RECT 176.700 136.050 177.900 143.400 ;
        RECT 184.950 141.450 187.050 142.050 ;
        RECT 193.950 141.450 196.050 142.050 ;
        RECT 184.950 140.550 196.050 141.450 ;
        RECT 184.950 139.950 187.050 140.550 ;
        RECT 193.950 139.950 196.050 140.550 ;
        RECT 197.250 136.050 199.050 137.850 ;
        RECT 203.700 136.050 204.600 143.400 ;
        RECT 214.950 141.450 217.050 142.050 ;
        RECT 220.950 141.450 223.050 142.200 ;
        RECT 214.950 140.550 223.050 141.450 ;
        RECT 214.950 139.950 217.050 140.550 ;
        RECT 220.950 140.100 223.050 140.550 ;
        RECT 224.100 136.050 225.900 137.850 ;
        RECT 230.100 136.050 231.000 148.200 ;
        RECT 246.000 149.100 246.900 149.400 ;
        RECT 251.100 149.400 252.900 155.400 ;
        RECT 254.100 149.400 255.900 156.000 ;
        RECT 272.700 149.400 274.500 156.000 ;
        RECT 251.100 149.100 252.600 149.400 ;
        RECT 246.000 148.200 252.600 149.100 ;
        RECT 246.000 136.050 246.900 148.200 ;
        RECT 273.000 146.100 274.800 147.900 ;
        RECT 250.950 144.450 253.050 145.050 ;
        RECT 271.950 144.450 274.050 145.050 ;
        RECT 275.700 144.900 277.500 155.400 ;
        RECT 250.950 143.550 274.050 144.450 ;
        RECT 250.950 142.950 253.050 143.550 ;
        RECT 271.950 142.950 274.050 143.550 ;
        RECT 275.100 143.400 277.500 144.900 ;
        RECT 280.800 143.400 282.600 156.000 ;
        RECT 296.100 149.400 297.900 155.400 ;
        RECT 299.100 149.400 300.900 156.000 ;
        RECT 314.100 149.400 315.900 156.000 ;
        RECT 317.100 149.400 318.900 155.400 ;
        RECT 320.100 149.400 321.900 156.000 ;
        RECT 338.100 149.400 339.900 155.400 ;
        RECT 341.100 149.400 342.900 156.000 ;
        RECT 359.100 149.400 360.900 156.000 ;
        RECT 362.100 149.400 363.900 155.400 ;
        RECT 365.100 149.400 366.900 156.000 ;
        RECT 383.100 154.500 390.900 155.400 ;
        RECT 251.100 136.050 252.900 137.850 ;
        RECT 275.100 136.050 276.300 143.400 ;
        RECT 281.100 136.050 282.900 137.850 ;
        RECT 296.700 136.050 297.900 149.400 ;
        RECT 299.100 136.050 300.900 137.850 ;
        RECT 317.100 136.050 318.300 149.400 ;
        RECT 338.700 136.050 339.900 149.400 ;
        RECT 341.100 136.050 342.900 137.850 ;
        RECT 362.100 136.050 363.300 149.400 ;
        RECT 383.100 143.400 384.900 154.500 ;
        RECT 386.100 142.500 387.900 153.600 ;
        RECT 389.100 144.600 390.900 154.500 ;
        RECT 392.100 145.500 393.900 156.000 ;
        RECT 395.100 144.600 396.900 155.400 ;
        RECT 413.100 149.400 414.900 156.000 ;
        RECT 416.100 149.400 417.900 155.400 ;
        RECT 419.100 150.000 420.900 156.000 ;
        RECT 416.400 149.100 417.900 149.400 ;
        RECT 422.100 149.400 423.900 155.400 ;
        RECT 422.100 149.100 423.000 149.400 ;
        RECT 416.400 148.200 423.000 149.100 ;
        RECT 389.100 143.700 396.900 144.600 ;
        RECT 386.100 141.600 390.900 142.500 ;
        RECT 386.100 136.050 387.900 137.850 ;
        RECT 390.000 136.050 390.900 141.600 ;
        RECT 391.950 136.050 393.750 137.850 ;
        RECT 416.100 136.050 417.900 137.850 ;
        RECT 422.100 136.050 423.000 148.200 ;
        RECT 437.100 144.300 438.900 155.400 ;
        RECT 440.100 145.200 441.900 156.000 ;
        RECT 443.100 144.300 444.900 155.400 ;
        RECT 437.100 143.400 444.900 144.300 ;
        RECT 446.100 143.400 447.900 155.400 ;
        RECT 461.400 143.400 463.200 156.000 ;
        RECT 466.500 144.900 468.300 155.400 ;
        RECT 469.500 149.400 471.300 156.000 ;
        RECT 485.100 149.400 486.900 156.000 ;
        RECT 488.100 149.400 489.900 155.400 ;
        RECT 491.100 149.400 492.900 156.000 ;
        RECT 469.200 146.100 471.000 147.900 ;
        RECT 466.500 143.400 468.900 144.900 ;
        RECT 440.250 136.050 442.050 137.850 ;
        RECT 446.700 136.050 447.600 143.400 ;
        RECT 461.100 136.050 462.900 137.850 ;
        RECT 467.700 136.050 468.900 143.400 ;
        RECT 488.100 136.050 489.300 149.400 ;
        RECT 495.150 145.200 496.950 155.400 ;
        RECT 494.550 143.400 496.950 145.200 ;
        RECT 498.150 143.400 499.950 156.000 ;
        RECT 503.550 146.400 505.350 155.400 ;
        RECT 508.350 149.400 510.150 156.000 ;
        RECT 511.350 148.500 513.150 155.400 ;
        RECT 514.350 149.400 516.150 156.000 ;
        RECT 518.850 149.400 520.650 155.400 ;
        RECT 507.450 147.450 514.050 148.500 ;
        RECT 507.450 146.700 509.250 147.450 ;
        RECT 512.250 146.700 514.050 147.450 ;
        RECT 518.550 147.300 520.650 149.400 ;
        RECT 503.250 145.500 505.350 146.400 ;
        RECT 515.850 145.800 517.650 146.400 ;
        RECT 503.250 144.300 511.050 145.500 ;
        RECT 509.250 143.700 511.050 144.300 ;
        RECT 511.950 144.900 517.650 145.800 ;
        RECT 494.550 142.500 495.450 143.400 ;
        RECT 511.950 142.800 512.850 144.900 ;
        RECT 515.850 144.600 517.650 144.900 ;
        RECT 518.550 144.600 521.550 146.400 ;
        RECT 518.550 143.700 519.750 144.600 ;
        RECT 504.450 142.500 512.850 142.800 ;
        RECT 494.550 141.900 512.850 142.500 ;
        RECT 514.950 142.800 519.750 143.700 ;
        RECT 523.650 143.400 525.450 156.000 ;
        RECT 526.650 143.400 528.450 155.400 ;
        RECT 542.100 149.400 543.900 156.000 ;
        RECT 545.100 149.400 546.900 155.400 ;
        RECT 548.100 149.400 549.900 156.000 ;
        RECT 566.100 149.400 567.900 156.000 ;
        RECT 569.100 149.400 570.900 155.400 ;
        RECT 572.100 150.000 573.900 156.000 ;
        RECT 494.550 141.300 506.250 141.900 ;
        RECT 16.950 133.950 19.050 136.050 ;
        RECT 19.950 133.950 22.050 136.050 ;
        RECT 22.950 133.950 25.050 136.050 ;
        RECT 25.950 133.950 28.050 136.050 ;
        RECT 40.950 133.950 43.050 136.050 ;
        RECT 43.950 133.950 46.050 136.050 ;
        RECT 58.950 133.950 61.050 136.050 ;
        RECT 61.950 133.950 64.050 136.050 ;
        RECT 64.950 133.950 67.050 136.050 ;
        RECT 67.950 133.950 70.050 136.050 ;
        RECT 82.950 133.950 85.050 136.050 ;
        RECT 85.950 133.950 88.050 136.050 ;
        RECT 88.950 133.950 91.050 136.050 ;
        RECT 91.950 133.950 94.050 136.050 ;
        RECT 106.950 133.950 109.050 136.050 ;
        RECT 109.950 133.950 112.050 136.050 ;
        RECT 127.950 133.950 130.050 136.050 ;
        RECT 130.950 133.950 133.050 136.050 ;
        RECT 145.950 133.950 148.050 136.050 ;
        RECT 148.950 133.950 151.050 136.050 ;
        RECT 151.950 133.950 154.050 136.050 ;
        RECT 154.950 133.950 157.050 136.050 ;
        RECT 169.950 133.950 172.050 136.050 ;
        RECT 172.950 133.950 175.050 136.050 ;
        RECT 175.950 133.950 178.050 136.050 ;
        RECT 178.950 133.950 181.050 136.050 ;
        RECT 193.950 133.950 196.050 136.050 ;
        RECT 196.950 133.950 199.050 136.050 ;
        RECT 199.950 133.950 202.050 136.050 ;
        RECT 202.950 133.950 205.050 136.050 ;
        RECT 220.950 133.950 223.050 136.050 ;
        RECT 223.950 133.950 226.050 136.050 ;
        RECT 226.950 133.950 229.050 136.050 ;
        RECT 229.950 133.950 232.050 136.050 ;
        RECT 244.950 133.950 247.050 136.050 ;
        RECT 247.950 133.950 250.050 136.050 ;
        RECT 250.950 133.950 253.050 136.050 ;
        RECT 253.950 133.950 256.050 136.050 ;
        RECT 271.950 133.950 274.050 136.050 ;
        RECT 274.950 133.950 277.050 136.050 ;
        RECT 277.950 133.950 280.050 136.050 ;
        RECT 280.950 133.950 283.050 136.050 ;
        RECT 295.950 133.950 298.050 136.050 ;
        RECT 298.950 133.950 301.050 136.050 ;
        RECT 313.950 133.950 316.050 136.050 ;
        RECT 316.950 133.950 319.050 136.050 ;
        RECT 319.950 133.950 322.050 136.050 ;
        RECT 337.950 133.950 340.050 136.050 ;
        RECT 340.950 133.950 343.050 136.050 ;
        RECT 358.950 133.950 361.050 136.050 ;
        RECT 361.950 133.950 364.050 136.050 ;
        RECT 364.950 133.950 367.050 136.050 ;
        RECT 382.950 133.950 385.050 136.050 ;
        RECT 385.950 133.950 388.050 136.050 ;
        RECT 388.950 133.950 391.050 136.050 ;
        RECT 391.950 133.950 394.050 136.050 ;
        RECT 394.950 133.950 397.050 136.050 ;
        RECT 412.950 133.950 415.050 136.050 ;
        RECT 415.950 133.950 418.050 136.050 ;
        RECT 418.950 133.950 421.050 136.050 ;
        RECT 421.950 133.950 424.050 136.050 ;
        RECT 436.950 133.950 439.050 136.050 ;
        RECT 439.950 133.950 442.050 136.050 ;
        RECT 442.950 133.950 445.050 136.050 ;
        RECT 445.950 133.950 448.050 136.050 ;
        RECT 460.950 133.950 463.050 136.050 ;
        RECT 463.950 133.950 466.050 136.050 ;
        RECT 466.950 133.950 469.050 136.050 ;
        RECT 469.950 133.950 472.050 136.050 ;
        RECT 484.950 133.950 487.050 136.050 ;
        RECT 487.950 133.950 490.050 136.050 ;
        RECT 490.950 133.950 493.050 136.050 ;
        RECT 17.400 126.600 18.300 133.950 ;
        RECT 19.950 132.150 21.750 133.950 ;
        RECT 26.100 132.150 27.900 133.950 ;
        RECT 17.400 125.400 22.500 126.600 ;
        RECT 17.700 120.000 19.500 123.600 ;
        RECT 20.700 120.600 22.500 125.400 ;
        RECT 25.200 120.000 27.000 126.600 ;
        RECT 41.700 123.600 42.900 133.950 ;
        RECT 60.000 130.200 60.900 133.950 ;
        RECT 62.100 132.150 63.900 133.950 ;
        RECT 68.100 132.150 69.900 133.950 ;
        RECT 86.100 132.150 87.900 133.950 ;
        RECT 60.000 129.000 63.300 130.200 ;
        RECT 89.700 129.600 90.900 133.950 ;
        RECT 92.100 132.150 93.900 133.950 ;
        RECT 41.100 120.600 42.900 123.600 ;
        RECT 44.100 120.000 45.900 123.600 ;
        RECT 61.500 120.600 63.300 129.000 ;
        RECT 68.100 120.000 69.900 129.600 ;
        RECT 89.700 128.700 93.300 129.600 ;
        RECT 83.100 125.700 90.900 127.050 ;
        RECT 83.100 120.600 84.900 125.700 ;
        RECT 86.100 120.000 87.900 124.800 ;
        RECT 89.100 120.600 90.900 125.700 ;
        RECT 92.100 126.600 93.300 128.700 ;
        RECT 92.100 120.600 93.900 126.600 ;
        RECT 110.100 123.600 111.300 133.950 ;
        RECT 131.100 123.600 132.300 133.950 ;
        RECT 146.100 132.150 147.900 133.950 ;
        RECT 149.100 129.600 150.300 133.950 ;
        RECT 152.100 132.150 153.900 133.950 ;
        RECT 173.100 132.150 174.900 133.950 ;
        RECT 146.700 128.700 150.300 129.600 ;
        RECT 176.700 129.600 177.900 133.950 ;
        RECT 179.100 132.150 180.900 133.950 ;
        RECT 194.100 132.150 195.900 133.950 ;
        RECT 200.250 132.150 202.050 133.950 ;
        RECT 176.700 128.700 180.300 129.600 ;
        RECT 146.700 126.600 147.900 128.700 ;
        RECT 107.100 120.000 108.900 123.600 ;
        RECT 110.100 120.600 111.900 123.600 ;
        RECT 128.100 120.000 129.900 123.600 ;
        RECT 131.100 120.600 132.900 123.600 ;
        RECT 146.100 120.600 147.900 126.600 ;
        RECT 149.100 125.700 156.900 127.050 ;
        RECT 149.100 120.600 150.900 125.700 ;
        RECT 152.100 120.000 153.900 124.800 ;
        RECT 155.100 120.600 156.900 125.700 ;
        RECT 170.100 125.700 177.900 127.050 ;
        RECT 170.100 120.600 171.900 125.700 ;
        RECT 173.100 120.000 174.900 124.800 ;
        RECT 176.100 120.600 177.900 125.700 ;
        RECT 179.100 126.600 180.300 128.700 ;
        RECT 203.700 126.600 204.600 133.950 ;
        RECT 221.100 132.150 222.900 133.950 ;
        RECT 227.100 132.150 228.900 133.950 ;
        RECT 230.100 130.200 231.000 133.950 ;
        RECT 179.100 120.600 180.900 126.600 ;
        RECT 195.000 120.000 196.800 126.600 ;
        RECT 199.500 125.400 204.600 126.600 ;
        RECT 199.500 120.600 201.300 125.400 ;
        RECT 202.500 120.000 204.300 123.600 ;
        RECT 221.100 120.000 222.900 129.600 ;
        RECT 227.700 129.000 231.000 130.200 ;
        RECT 246.000 130.200 246.900 133.950 ;
        RECT 248.100 132.150 249.900 133.950 ;
        RECT 254.100 132.150 255.900 133.950 ;
        RECT 272.100 132.150 273.900 133.950 ;
        RECT 246.000 129.000 249.300 130.200 ;
        RECT 275.100 129.600 276.300 133.950 ;
        RECT 278.100 132.150 279.900 133.950 ;
        RECT 227.700 120.600 229.500 129.000 ;
        RECT 247.500 120.600 249.300 129.000 ;
        RECT 254.100 120.000 255.900 129.600 ;
        RECT 272.700 128.700 276.300 129.600 ;
        RECT 272.700 126.600 273.900 128.700 ;
        RECT 272.100 120.600 273.900 126.600 ;
        RECT 275.100 125.700 282.900 127.050 ;
        RECT 275.100 120.600 276.900 125.700 ;
        RECT 278.100 120.000 279.900 124.800 ;
        RECT 281.100 120.600 282.900 125.700 ;
        RECT 296.700 123.600 297.900 133.950 ;
        RECT 314.250 132.150 316.050 133.950 ;
        RECT 317.100 128.700 318.300 133.950 ;
        RECT 320.100 132.150 321.900 133.950 ;
        RECT 317.100 127.800 321.300 128.700 ;
        RECT 296.100 120.600 297.900 123.600 ;
        RECT 299.100 120.000 300.900 123.600 ;
        RECT 314.400 120.000 316.200 126.600 ;
        RECT 319.500 120.600 321.300 127.800 ;
        RECT 338.700 123.600 339.900 133.950 ;
        RECT 359.250 132.150 361.050 133.950 ;
        RECT 362.100 128.700 363.300 133.950 ;
        RECT 365.100 132.150 366.900 133.950 ;
        RECT 383.100 132.150 384.900 133.950 ;
        RECT 362.100 127.800 366.300 128.700 ;
        RECT 338.100 120.600 339.900 123.600 ;
        RECT 341.100 120.000 342.900 123.600 ;
        RECT 359.400 120.000 361.200 126.600 ;
        RECT 364.500 120.600 366.300 127.800 ;
        RECT 389.700 126.600 390.900 133.950 ;
        RECT 394.950 132.150 396.750 133.950 ;
        RECT 413.100 132.150 414.900 133.950 ;
        RECT 419.100 132.150 420.900 133.950 ;
        RECT 422.100 130.200 423.000 133.950 ;
        RECT 437.100 132.150 438.900 133.950 ;
        RECT 443.250 132.150 445.050 133.950 ;
        RECT 385.500 120.000 387.300 126.600 ;
        RECT 390.000 120.600 391.800 126.600 ;
        RECT 394.500 120.000 396.300 126.600 ;
        RECT 413.100 120.000 414.900 129.600 ;
        RECT 419.700 129.000 423.000 130.200 ;
        RECT 427.950 129.450 430.050 130.050 ;
        RECT 442.950 129.450 445.050 130.050 ;
        RECT 419.700 120.600 421.500 129.000 ;
        RECT 427.950 128.550 445.050 129.450 ;
        RECT 427.950 127.950 430.050 128.550 ;
        RECT 442.950 127.950 445.050 128.550 ;
        RECT 446.700 126.600 447.600 133.950 ;
        RECT 464.100 132.150 465.900 133.950 ;
        RECT 467.700 129.600 468.900 133.950 ;
        RECT 470.100 132.150 471.900 133.950 ;
        RECT 485.250 132.150 487.050 133.950 ;
        RECT 467.700 128.700 471.300 129.600 ;
        RECT 438.000 120.000 439.800 126.600 ;
        RECT 442.500 125.400 447.600 126.600 ;
        RECT 461.100 125.700 468.900 127.050 ;
        RECT 442.500 120.600 444.300 125.400 ;
        RECT 445.500 120.000 447.300 123.600 ;
        RECT 461.100 120.600 462.900 125.700 ;
        RECT 464.100 120.000 465.900 124.800 ;
        RECT 467.100 120.600 468.900 125.700 ;
        RECT 470.100 126.600 471.300 128.700 ;
        RECT 488.100 128.700 489.300 133.950 ;
        RECT 491.100 132.150 492.900 133.950 ;
        RECT 488.100 127.800 492.300 128.700 ;
        RECT 470.100 120.600 471.900 126.600 ;
        RECT 485.400 120.000 487.200 126.600 ;
        RECT 490.500 120.600 492.300 127.800 ;
        RECT 494.550 126.600 495.450 141.300 ;
        RECT 504.450 141.000 506.250 141.300 ;
        RECT 496.950 133.950 499.050 136.050 ;
        RECT 506.100 134.400 508.200 136.050 ;
        RECT 496.950 131.400 498.750 133.950 ;
        RECT 500.100 133.200 508.200 134.400 ;
        RECT 500.100 132.600 501.900 133.200 ;
        RECT 503.100 131.400 504.900 132.000 ;
        RECT 496.950 130.200 504.900 131.400 ;
        RECT 514.950 130.200 515.850 142.800 ;
        RECT 518.550 140.100 520.650 140.700 ;
        RECT 524.550 140.100 526.350 140.550 ;
        RECT 518.550 138.900 526.350 140.100 ;
        RECT 518.550 138.600 520.650 138.900 ;
        RECT 524.550 138.750 526.350 138.900 ;
        RECT 527.250 136.050 528.450 143.400 ;
        RECT 545.700 136.050 546.900 149.400 ;
        RECT 569.400 149.100 570.900 149.400 ;
        RECT 575.100 149.400 576.900 155.400 ;
        RECT 575.100 149.100 576.000 149.400 ;
        RECT 569.400 148.200 576.000 149.100 ;
        RECT 569.100 136.050 570.900 137.850 ;
        RECT 575.100 136.050 576.000 148.200 ;
        RECT 590.100 144.300 591.900 155.400 ;
        RECT 593.100 145.200 594.900 156.000 ;
        RECT 596.100 144.300 597.900 155.400 ;
        RECT 590.100 143.400 597.900 144.300 ;
        RECT 599.100 143.400 600.900 155.400 ;
        RECT 614.700 149.400 616.500 156.000 ;
        RECT 615.000 146.100 616.800 147.900 ;
        RECT 617.700 144.900 619.500 155.400 ;
        RECT 617.100 143.400 619.500 144.900 ;
        RECT 622.800 143.400 624.600 156.000 ;
        RECT 638.400 143.400 640.200 156.000 ;
        RECT 643.500 144.900 645.300 155.400 ;
        RECT 646.500 149.400 648.300 156.000 ;
        RECT 662.100 149.400 663.900 156.000 ;
        RECT 665.100 149.400 666.900 155.400 ;
        RECT 646.200 146.100 648.000 147.900 ;
        RECT 643.500 143.400 645.900 144.900 ;
        RECT 593.250 136.050 595.050 137.850 ;
        RECT 599.700 136.050 600.600 143.400 ;
        RECT 617.100 136.050 618.300 143.400 ;
        RECT 619.950 141.450 622.050 142.050 ;
        RECT 640.950 141.450 643.050 142.050 ;
        RECT 619.950 140.550 643.050 141.450 ;
        RECT 619.950 139.950 622.050 140.550 ;
        RECT 640.950 139.950 643.050 140.550 ;
        RECT 623.100 136.050 624.900 137.850 ;
        RECT 638.100 136.050 639.900 137.850 ;
        RECT 644.700 136.050 645.900 143.400 ;
        RECT 523.950 135.750 528.450 136.050 ;
        RECT 522.150 133.950 528.450 135.750 ;
        RECT 541.950 133.950 544.050 136.050 ;
        RECT 544.950 133.950 547.050 136.050 ;
        RECT 547.950 133.950 550.050 136.050 ;
        RECT 565.950 133.950 568.050 136.050 ;
        RECT 568.950 133.950 571.050 136.050 ;
        RECT 571.950 133.950 574.050 136.050 ;
        RECT 574.950 133.950 577.050 136.050 ;
        RECT 589.950 133.950 592.050 136.050 ;
        RECT 592.950 133.950 595.050 136.050 ;
        RECT 595.950 133.950 598.050 136.050 ;
        RECT 598.950 133.950 601.050 136.050 ;
        RECT 613.950 133.950 616.050 136.050 ;
        RECT 616.950 133.950 619.050 136.050 ;
        RECT 619.950 133.950 622.050 136.050 ;
        RECT 622.950 133.950 625.050 136.050 ;
        RECT 637.950 133.950 640.050 136.050 ;
        RECT 640.950 133.950 643.050 136.050 ;
        RECT 643.950 133.950 646.050 136.050 ;
        RECT 646.950 133.950 649.050 136.050 ;
        RECT 662.100 133.950 664.200 136.050 ;
        RECT 503.850 129.000 515.850 130.200 ;
        RECT 503.850 127.200 504.900 129.000 ;
        RECT 514.050 128.400 515.850 129.000 ;
        RECT 494.550 124.800 496.950 126.600 ;
        RECT 495.150 120.600 496.950 124.800 ;
        RECT 498.150 120.000 499.950 126.600 ;
        RECT 500.850 124.200 502.950 125.700 ;
        RECT 503.850 125.400 505.650 127.200 ;
        RECT 527.250 126.600 528.450 133.950 ;
        RECT 542.100 132.150 543.900 133.950 ;
        RECT 545.700 128.700 546.900 133.950 ;
        RECT 547.950 132.150 549.750 133.950 ;
        RECT 566.100 132.150 567.900 133.950 ;
        RECT 572.100 132.150 573.900 133.950 ;
        RECT 575.100 130.200 576.000 133.950 ;
        RECT 590.100 132.150 591.900 133.950 ;
        RECT 596.250 132.150 598.050 133.950 ;
        RECT 506.850 125.550 508.650 126.300 ;
        RECT 506.850 124.500 511.800 125.550 ;
        RECT 500.850 123.600 504.750 124.200 ;
        RECT 510.750 123.600 511.800 124.500 ;
        RECT 518.250 123.600 520.650 125.700 ;
        RECT 501.150 122.700 504.750 123.600 ;
        RECT 502.950 120.600 504.750 122.700 ;
        RECT 507.450 120.000 509.250 123.600 ;
        RECT 510.750 120.600 512.550 123.600 ;
        RECT 513.750 120.000 515.550 123.600 ;
        RECT 518.250 120.600 520.050 123.600 ;
        RECT 523.350 120.000 525.150 126.600 ;
        RECT 526.650 120.600 528.450 126.600 ;
        RECT 542.700 127.800 546.900 128.700 ;
        RECT 542.700 120.600 544.500 127.800 ;
        RECT 547.800 120.000 549.600 126.600 ;
        RECT 566.100 120.000 567.900 129.600 ;
        RECT 572.700 129.000 576.000 130.200 ;
        RECT 572.700 120.600 574.500 129.000 ;
        RECT 599.700 126.600 600.600 133.950 ;
        RECT 614.100 132.150 615.900 133.950 ;
        RECT 617.100 129.600 618.300 133.950 ;
        RECT 620.100 132.150 621.900 133.950 ;
        RECT 641.100 132.150 642.900 133.950 ;
        RECT 614.700 128.700 618.300 129.600 ;
        RECT 644.700 129.600 645.900 133.950 ;
        RECT 647.100 132.150 648.900 133.950 ;
        RECT 662.250 132.150 664.050 133.950 ;
        RECT 644.700 128.700 648.300 129.600 ;
        RECT 665.100 129.300 666.000 149.400 ;
        RECT 668.100 144.000 669.900 156.000 ;
        RECT 671.100 143.400 672.900 155.400 ;
        RECT 689.100 149.400 690.900 156.000 ;
        RECT 692.100 149.400 693.900 155.400 ;
        RECT 695.100 149.400 696.900 156.000 ;
        RECT 713.100 149.400 714.900 156.000 ;
        RECT 716.100 149.400 717.900 155.400 ;
        RECT 719.100 150.000 720.900 156.000 ;
        RECT 667.200 136.050 669.000 137.850 ;
        RECT 671.400 136.050 672.300 143.400 ;
        RECT 692.100 136.050 693.300 149.400 ;
        RECT 716.400 149.100 717.900 149.400 ;
        RECT 722.100 149.400 723.900 155.400 ;
        RECT 740.100 149.400 741.900 155.400 ;
        RECT 743.100 149.400 744.900 156.000 ;
        RECT 758.100 149.400 759.900 156.000 ;
        RECT 761.100 149.400 762.900 155.400 ;
        RECT 764.100 149.400 765.900 156.000 ;
        RECT 722.100 149.100 723.000 149.400 ;
        RECT 716.400 148.200 723.000 149.100 ;
        RECT 716.100 136.050 717.900 137.850 ;
        RECT 722.100 136.050 723.000 148.200 ;
        RECT 740.700 136.050 741.900 149.400 ;
        RECT 742.950 141.450 745.050 142.050 ;
        RECT 748.950 141.450 751.050 142.050 ;
        RECT 742.950 140.550 751.050 141.450 ;
        RECT 742.950 139.950 745.050 140.550 ;
        RECT 748.950 139.950 751.050 140.550 ;
        RECT 743.100 136.050 744.900 137.850 ;
        RECT 761.100 136.050 762.300 149.400 ;
        RECT 782.100 143.400 783.900 155.400 ;
        RECT 785.100 144.000 786.900 156.000 ;
        RECT 788.100 149.400 789.900 155.400 ;
        RECT 791.100 149.400 792.900 156.000 ;
        RECT 809.100 149.400 810.900 156.000 ;
        RECT 812.100 149.400 813.900 155.400 ;
        RECT 815.100 149.400 816.900 156.000 ;
        RECT 833.100 149.400 834.900 155.400 ;
        RECT 836.100 149.400 837.900 156.000 ;
        RECT 782.700 136.050 783.600 143.400 ;
        RECT 786.000 136.050 787.800 137.850 ;
        RECT 667.500 133.950 669.600 136.050 ;
        RECT 670.800 133.950 672.900 136.050 ;
        RECT 688.950 133.950 691.050 136.050 ;
        RECT 691.950 133.950 694.050 136.050 ;
        RECT 694.950 133.950 697.050 136.050 ;
        RECT 712.950 133.950 715.050 136.050 ;
        RECT 715.950 133.950 718.050 136.050 ;
        RECT 718.950 133.950 721.050 136.050 ;
        RECT 721.950 133.950 724.050 136.050 ;
        RECT 739.950 133.950 742.050 136.050 ;
        RECT 742.950 133.950 745.050 136.050 ;
        RECT 757.950 133.950 760.050 136.050 ;
        RECT 760.950 133.950 763.050 136.050 ;
        RECT 763.950 133.950 766.050 136.050 ;
        RECT 782.100 133.950 784.200 136.050 ;
        RECT 785.400 133.950 787.500 136.050 ;
        RECT 614.700 126.600 615.900 128.700 ;
        RECT 591.000 120.000 592.800 126.600 ;
        RECT 595.500 125.400 600.600 126.600 ;
        RECT 595.500 120.600 597.300 125.400 ;
        RECT 598.500 120.000 600.300 123.600 ;
        RECT 614.100 120.600 615.900 126.600 ;
        RECT 617.100 125.700 624.900 127.050 ;
        RECT 617.100 120.600 618.900 125.700 ;
        RECT 620.100 120.000 621.900 124.800 ;
        RECT 623.100 120.600 624.900 125.700 ;
        RECT 638.100 125.700 645.900 127.050 ;
        RECT 638.100 120.600 639.900 125.700 ;
        RECT 641.100 120.000 642.900 124.800 ;
        RECT 644.100 120.600 645.900 125.700 ;
        RECT 647.100 126.600 648.300 128.700 ;
        RECT 662.100 128.400 670.500 129.300 ;
        RECT 647.100 120.600 648.900 126.600 ;
        RECT 662.100 120.600 663.900 128.400 ;
        RECT 668.700 127.500 670.500 128.400 ;
        RECT 671.400 126.600 672.300 133.950 ;
        RECT 689.250 132.150 691.050 133.950 ;
        RECT 692.100 128.700 693.300 133.950 ;
        RECT 695.100 132.150 696.900 133.950 ;
        RECT 713.100 132.150 714.900 133.950 ;
        RECT 719.100 132.150 720.900 133.950 ;
        RECT 722.100 130.200 723.000 133.950 ;
        RECT 692.100 127.800 696.300 128.700 ;
        RECT 666.600 120.000 668.400 126.600 ;
        RECT 669.600 124.800 672.300 126.600 ;
        RECT 669.600 120.600 671.400 124.800 ;
        RECT 689.400 120.000 691.200 126.600 ;
        RECT 694.500 120.600 696.300 127.800 ;
        RECT 713.100 120.000 714.900 129.600 ;
        RECT 719.700 129.000 723.000 130.200 ;
        RECT 719.700 120.600 721.500 129.000 ;
        RECT 740.700 123.600 741.900 133.950 ;
        RECT 758.250 132.150 760.050 133.950 ;
        RECT 761.100 128.700 762.300 133.950 ;
        RECT 764.100 132.150 765.900 133.950 ;
        RECT 761.100 127.800 765.300 128.700 ;
        RECT 740.100 120.600 741.900 123.600 ;
        RECT 743.100 120.000 744.900 123.600 ;
        RECT 758.400 120.000 760.200 126.600 ;
        RECT 763.500 120.600 765.300 127.800 ;
        RECT 782.700 126.600 783.600 133.950 ;
        RECT 789.000 129.300 789.900 149.400 ;
        RECT 812.700 136.050 813.900 149.400 ;
        RECT 833.700 136.050 834.900 149.400 ;
        RECT 851.400 143.400 853.200 156.000 ;
        RECT 856.500 144.900 858.300 155.400 ;
        RECT 859.500 149.400 861.300 156.000 ;
        RECT 859.200 146.100 861.000 147.900 ;
        RECT 856.500 143.400 858.900 144.900 ;
        RECT 878.100 143.400 879.900 155.400 ;
        RECT 881.100 144.300 882.900 155.400 ;
        RECT 884.100 145.200 885.900 156.000 ;
        RECT 887.100 144.300 888.900 155.400 ;
        RECT 905.100 149.400 906.900 156.000 ;
        RECT 908.100 149.400 909.900 155.400 ;
        RECT 911.100 150.000 912.900 156.000 ;
        RECT 908.400 149.100 909.900 149.400 ;
        RECT 914.100 149.400 915.900 155.400 ;
        RECT 914.100 149.100 915.000 149.400 ;
        RECT 908.400 148.200 915.000 149.100 ;
        RECT 881.100 143.400 888.900 144.300 ;
        RECT 836.100 136.050 837.900 137.850 ;
        RECT 851.100 136.050 852.900 137.850 ;
        RECT 857.700 136.050 858.900 143.400 ;
        RECT 878.400 136.050 879.300 143.400 ;
        RECT 886.950 141.450 889.050 142.050 ;
        RECT 910.950 141.450 913.050 142.050 ;
        RECT 886.950 140.550 913.050 141.450 ;
        RECT 886.950 139.950 889.050 140.550 ;
        RECT 910.950 139.950 913.050 140.550 ;
        RECT 883.950 136.050 885.750 137.850 ;
        RECT 908.100 136.050 909.900 137.850 ;
        RECT 914.100 136.050 915.000 148.200 ;
        RECT 929.100 144.300 930.900 155.400 ;
        RECT 932.100 145.200 933.900 156.000 ;
        RECT 935.100 144.300 936.900 155.400 ;
        RECT 929.100 143.400 936.900 144.300 ;
        RECT 938.100 143.400 939.900 155.400 ;
        RECT 953.100 144.600 954.900 155.400 ;
        RECT 956.100 145.500 958.200 156.000 ;
        RECT 953.100 143.400 958.200 144.600 ;
        RECT 960.600 144.300 962.400 155.400 ;
        RECT 965.100 145.500 966.900 156.000 ;
        RECT 968.100 144.300 969.900 155.400 ;
        RECT 932.250 136.050 934.050 137.850 ;
        RECT 938.700 136.050 939.600 143.400 ;
        RECT 956.100 142.500 958.200 143.400 ;
        RECT 959.100 143.400 962.400 144.300 ;
        RECT 959.100 139.050 960.300 143.400 ;
        RECT 965.100 143.100 969.900 144.300 ;
        RECT 986.100 144.600 987.900 155.400 ;
        RECT 989.100 145.500 990.900 156.000 ;
        RECT 986.100 143.400 990.900 144.600 ;
        RECT 965.100 142.200 967.200 143.100 ;
        RECT 988.800 142.500 990.900 143.400 ;
        RECT 993.600 143.400 995.400 155.400 ;
        RECT 998.100 145.500 999.900 156.000 ;
        RECT 1001.100 144.300 1002.900 155.400 ;
        RECT 998.400 143.400 1002.900 144.300 ;
        RECT 961.800 141.300 967.200 142.200 ;
        RECT 993.600 142.050 994.800 143.400 ;
        RECT 961.800 139.500 963.600 141.300 ;
        RECT 993.300 141.000 994.800 142.050 ;
        RECT 998.400 141.300 1000.500 143.400 ;
        RECT 993.300 139.050 994.200 141.000 ;
        RECT 958.800 138.300 960.900 139.050 ;
        RECT 953.400 136.050 955.200 137.850 ;
        RECT 958.800 136.950 961.800 138.300 ;
        RECT 790.800 133.950 792.900 136.050 ;
        RECT 808.950 133.950 811.050 136.050 ;
        RECT 811.950 133.950 814.050 136.050 ;
        RECT 814.950 133.950 817.050 136.050 ;
        RECT 832.950 133.950 835.050 136.050 ;
        RECT 835.950 133.950 838.050 136.050 ;
        RECT 850.950 133.950 853.050 136.050 ;
        RECT 853.950 133.950 856.050 136.050 ;
        RECT 856.950 133.950 859.050 136.050 ;
        RECT 859.950 133.950 862.050 136.050 ;
        RECT 877.950 133.950 880.050 136.050 ;
        RECT 880.950 133.950 883.050 136.050 ;
        RECT 883.950 133.950 886.050 136.050 ;
        RECT 886.950 133.950 889.050 136.050 ;
        RECT 904.950 133.950 907.050 136.050 ;
        RECT 907.950 133.950 910.050 136.050 ;
        RECT 910.950 133.950 913.050 136.050 ;
        RECT 913.950 133.950 916.050 136.050 ;
        RECT 928.950 133.950 931.050 136.050 ;
        RECT 931.950 133.950 934.050 136.050 ;
        RECT 934.950 133.950 937.050 136.050 ;
        RECT 937.950 133.950 940.050 136.050 ;
        RECT 953.100 133.950 955.200 136.050 ;
        RECT 958.200 134.100 960.000 135.900 ;
        RECT 790.950 132.150 792.750 133.950 ;
        RECT 809.100 132.150 810.900 133.950 ;
        RECT 784.500 128.400 792.900 129.300 ;
        RECT 812.700 128.700 813.900 133.950 ;
        RECT 814.950 132.150 816.750 133.950 ;
        RECT 784.500 127.500 786.300 128.400 ;
        RECT 782.700 124.800 785.400 126.600 ;
        RECT 783.600 120.600 785.400 124.800 ;
        RECT 786.600 120.000 788.400 126.600 ;
        RECT 791.100 120.600 792.900 128.400 ;
        RECT 809.700 127.800 813.900 128.700 ;
        RECT 809.700 120.600 811.500 127.800 ;
        RECT 814.800 120.000 816.600 126.600 ;
        RECT 833.700 123.600 834.900 133.950 ;
        RECT 854.100 132.150 855.900 133.950 ;
        RECT 857.700 129.600 858.900 133.950 ;
        RECT 860.100 132.150 861.900 133.950 ;
        RECT 857.700 128.700 861.300 129.600 ;
        RECT 851.100 125.700 858.900 127.050 ;
        RECT 833.100 120.600 834.900 123.600 ;
        RECT 836.100 120.000 837.900 123.600 ;
        RECT 851.100 120.600 852.900 125.700 ;
        RECT 854.100 120.000 855.900 124.800 ;
        RECT 857.100 120.600 858.900 125.700 ;
        RECT 860.100 126.600 861.300 128.700 ;
        RECT 878.400 126.600 879.300 133.950 ;
        RECT 880.950 132.150 882.750 133.950 ;
        RECT 887.100 132.150 888.900 133.950 ;
        RECT 905.100 132.150 906.900 133.950 ;
        RECT 911.100 132.150 912.900 133.950 ;
        RECT 914.100 130.200 915.000 133.950 ;
        RECT 929.100 132.150 930.900 133.950 ;
        RECT 935.250 132.150 937.050 133.950 ;
        RECT 860.100 120.600 861.900 126.600 ;
        RECT 878.400 125.400 883.500 126.600 ;
        RECT 878.700 120.000 880.500 123.600 ;
        RECT 881.700 120.600 883.500 125.400 ;
        RECT 886.200 120.000 888.000 126.600 ;
        RECT 905.100 120.000 906.900 129.600 ;
        RECT 911.700 129.000 915.000 130.200 ;
        RECT 922.950 129.450 925.050 130.050 ;
        RECT 934.950 129.450 937.050 130.050 ;
        RECT 911.700 120.600 913.500 129.000 ;
        RECT 922.950 128.550 937.050 129.450 ;
        RECT 922.950 127.950 925.050 128.550 ;
        RECT 934.950 127.950 937.050 128.550 ;
        RECT 938.700 126.600 939.600 133.950 ;
        RECT 957.900 132.000 960.000 134.100 ;
        RECT 960.900 130.200 961.800 136.950 ;
        RECT 963.300 136.200 965.100 138.000 ;
        RECT 963.000 134.100 965.100 136.200 ;
        RECT 986.400 136.050 988.200 137.850 ;
        RECT 992.100 136.950 994.200 139.050 ;
        RECT 995.100 139.500 997.200 139.800 ;
        RECT 995.100 137.700 999.000 139.500 ;
        RECT 967.800 133.800 969.900 136.050 ;
        RECT 986.100 133.950 988.200 136.050 ;
        RECT 992.700 136.800 994.200 136.950 ;
        RECT 992.700 135.900 995.100 136.800 ;
        RECT 967.800 133.200 969.600 133.800 ;
        RECT 963.000 132.000 969.600 133.200 ;
        RECT 990.900 133.200 992.700 135.000 ;
        RECT 963.000 131.100 965.100 132.000 ;
        RECT 990.900 131.100 993.000 133.200 ;
        RECT 955.500 127.500 957.600 129.900 ;
        RECT 958.800 128.100 961.800 130.200 ;
        RECT 962.700 129.300 964.500 131.100 ;
        RECT 993.900 130.200 995.100 135.900 ;
        RECT 996.000 136.050 997.800 136.500 ;
        RECT 996.000 134.700 1002.900 136.050 ;
        RECT 1000.800 133.950 1002.900 134.700 ;
        RECT 930.000 120.000 931.800 126.600 ;
        RECT 934.500 125.400 939.600 126.600 ;
        RECT 953.100 126.600 957.600 127.500 ;
        RECT 934.500 120.600 936.300 125.400 ;
        RECT 937.500 120.000 939.300 123.600 ;
        RECT 953.100 120.600 954.900 126.600 ;
        RECT 960.900 126.000 961.800 128.100 ;
        RECT 965.400 129.000 967.500 129.600 ;
        RECT 965.400 127.500 969.900 129.000 ;
        RECT 988.800 127.500 990.900 128.700 ;
        RECT 992.100 128.100 995.100 130.200 ;
        RECT 996.000 131.400 997.800 133.200 ;
        RECT 1000.800 132.150 1002.600 133.950 ;
        RECT 996.000 129.300 998.100 131.400 ;
        RECT 996.000 128.400 1002.300 129.300 ;
        RECT 968.400 126.600 969.900 127.500 ;
        RECT 956.400 120.000 958.200 125.700 ;
        RECT 960.900 120.600 962.700 126.000 ;
        RECT 965.100 120.000 966.900 125.700 ;
        RECT 968.100 120.600 969.900 126.600 ;
        RECT 986.100 126.600 990.900 127.500 ;
        RECT 993.900 126.600 995.100 128.100 ;
        RECT 1001.100 126.600 1002.300 128.400 ;
        RECT 986.100 120.600 987.900 126.600 ;
        RECT 989.100 120.000 990.900 125.700 ;
        RECT 993.600 120.600 995.400 126.600 ;
        RECT 998.100 120.000 999.900 125.700 ;
        RECT 1001.100 120.600 1002.900 126.600 ;
        RECT 17.100 113.400 18.900 117.000 ;
        RECT 20.100 113.400 21.900 116.400 ;
        RECT 20.100 103.050 21.300 113.400 ;
        RECT 36.000 110.400 37.800 117.000 ;
        RECT 40.500 111.600 42.300 116.400 ;
        RECT 43.500 113.400 45.300 117.000 ;
        RECT 40.500 110.400 45.600 111.600 ;
        RECT 35.100 103.050 36.900 104.850 ;
        RECT 41.250 103.050 43.050 104.850 ;
        RECT 44.700 103.050 45.600 110.400 ;
        RECT 59.100 107.400 60.900 117.000 ;
        RECT 65.700 108.000 67.500 116.400 ;
        RECT 85.500 108.000 87.300 116.400 ;
        RECT 65.700 106.800 69.000 108.000 ;
        RECT 59.100 103.050 60.900 104.850 ;
        RECT 65.100 103.050 66.900 104.850 ;
        RECT 68.100 103.050 69.000 106.800 ;
        RECT 84.000 106.800 87.300 108.000 ;
        RECT 92.100 107.400 93.900 117.000 ;
        RECT 108.000 110.400 109.800 117.000 ;
        RECT 112.500 111.600 114.300 116.400 ;
        RECT 115.500 113.400 117.300 117.000 ;
        RECT 112.500 110.400 117.600 111.600 ;
        RECT 84.000 103.050 84.900 106.800 ;
        RECT 86.100 103.050 87.900 104.850 ;
        RECT 92.100 103.050 93.900 104.850 ;
        RECT 107.100 103.050 108.900 104.850 ;
        RECT 113.250 103.050 115.050 104.850 ;
        RECT 116.700 103.050 117.600 110.400 ;
        RECT 134.100 111.300 135.900 116.400 ;
        RECT 137.100 112.200 138.900 117.000 ;
        RECT 140.100 111.300 141.900 116.400 ;
        RECT 134.100 109.950 141.900 111.300 ;
        RECT 143.100 110.400 144.900 116.400 ;
        RECT 161.100 113.400 162.900 117.000 ;
        RECT 164.100 113.400 165.900 116.400 ;
        RECT 143.100 108.300 144.300 110.400 ;
        RECT 140.700 107.400 144.300 108.300 ;
        RECT 137.100 103.050 138.900 104.850 ;
        RECT 140.700 103.050 141.900 107.400 ;
        RECT 143.100 103.050 144.900 104.850 ;
        RECT 164.100 103.050 165.300 113.400 ;
        RECT 179.100 111.300 180.900 116.400 ;
        RECT 182.100 112.200 183.900 117.000 ;
        RECT 185.100 111.300 186.900 116.400 ;
        RECT 179.100 109.950 186.900 111.300 ;
        RECT 188.100 110.400 189.900 116.400 ;
        RECT 207.000 110.400 208.800 117.000 ;
        RECT 211.500 111.600 213.300 116.400 ;
        RECT 214.500 113.400 216.300 117.000 ;
        RECT 211.500 110.400 216.600 111.600 ;
        RECT 230.400 110.400 232.200 117.000 ;
        RECT 188.100 108.300 189.300 110.400 ;
        RECT 185.700 107.400 189.300 108.300 ;
        RECT 205.950 108.450 208.050 109.050 ;
        RECT 211.950 108.450 214.050 109.050 ;
        RECT 205.950 107.550 214.050 108.450 ;
        RECT 182.100 103.050 183.900 104.850 ;
        RECT 185.700 103.050 186.900 107.400 ;
        RECT 205.950 106.950 208.050 107.550 ;
        RECT 211.950 106.950 214.050 107.550 ;
        RECT 188.100 103.050 189.900 104.850 ;
        RECT 206.100 103.050 207.900 104.850 ;
        RECT 212.250 103.050 214.050 104.850 ;
        RECT 215.700 103.050 216.600 110.400 ;
        RECT 235.500 109.200 237.300 116.400 ;
        RECT 256.500 110.400 258.300 117.000 ;
        RECT 261.000 110.400 262.800 116.400 ;
        RECT 265.500 110.400 267.300 117.000 ;
        RECT 281.100 113.400 282.900 117.000 ;
        RECT 284.100 113.400 285.900 116.400 ;
        RECT 287.100 113.400 288.900 117.000 ;
        RECT 233.100 108.300 237.300 109.200 ;
        RECT 230.250 103.050 232.050 104.850 ;
        RECT 233.100 103.050 234.300 108.300 ;
        RECT 236.100 103.050 237.900 104.850 ;
        RECT 254.100 103.050 255.900 104.850 ;
        RECT 260.700 103.050 261.900 110.400 ;
        RECT 265.950 103.050 267.750 104.850 ;
        RECT 284.400 103.050 285.300 113.400 ;
        RECT 302.100 111.300 303.900 116.400 ;
        RECT 305.100 112.200 306.900 117.000 ;
        RECT 308.100 111.300 309.900 116.400 ;
        RECT 302.100 109.950 309.900 111.300 ;
        RECT 311.100 110.400 312.900 116.400 ;
        RECT 328.800 113.400 330.900 117.000 ;
        RECT 332.100 113.400 333.900 116.400 ;
        RECT 335.100 113.400 336.900 117.000 ;
        RECT 338.100 113.400 340.800 116.400 ;
        RECT 362.100 113.400 363.900 117.000 ;
        RECT 365.100 113.400 366.900 116.400 ;
        RECT 368.100 113.400 369.900 117.000 ;
        RECT 383.100 113.400 384.900 117.000 ;
        RECT 386.100 113.400 387.900 116.400 ;
        RECT 389.100 113.400 390.900 117.000 ;
        RECT 404.100 113.400 405.900 117.000 ;
        RECT 407.100 113.400 408.900 116.400 ;
        RECT 422.100 113.400 423.900 117.000 ;
        RECT 425.100 113.400 426.900 116.400 ;
        RECT 332.700 112.500 333.600 113.400 ;
        RECT 339.900 112.500 340.800 113.400 ;
        RECT 332.700 111.600 345.300 112.500 ;
        RECT 311.100 108.300 312.300 110.400 ;
        RECT 308.700 107.400 312.300 108.300 ;
        RECT 316.950 108.450 319.050 109.050 ;
        RECT 337.950 108.450 340.050 109.050 ;
        RECT 316.950 107.550 340.050 108.450 ;
        RECT 305.100 103.050 306.900 104.850 ;
        RECT 308.700 103.050 309.900 107.400 ;
        RECT 316.950 106.950 319.050 107.550 ;
        RECT 337.950 106.950 340.050 107.550 ;
        RECT 311.100 103.050 312.900 104.850 ;
        RECT 334.950 103.050 336.750 104.850 ;
        RECT 344.100 103.050 345.300 111.600 ;
        RECT 365.400 103.050 366.300 113.400 ;
        RECT 367.950 108.450 370.050 109.050 ;
        RECT 376.950 108.450 379.050 109.050 ;
        RECT 367.950 107.550 379.050 108.450 ;
        RECT 367.950 106.950 370.050 107.550 ;
        RECT 376.950 106.950 379.050 107.550 ;
        RECT 386.400 103.050 387.300 113.400 ;
        RECT 407.100 103.050 408.300 113.400 ;
        RECT 425.100 103.050 426.300 113.400 ;
        RECT 440.400 110.400 442.200 117.000 ;
        RECT 445.500 109.200 447.300 116.400 ;
        RECT 464.100 110.400 465.900 116.400 ;
        RECT 467.100 111.300 468.900 117.000 ;
        RECT 471.600 110.400 473.400 116.400 ;
        RECT 476.100 111.300 477.900 117.000 ;
        RECT 479.100 110.400 480.900 116.400 ;
        RECT 494.100 113.400 495.900 117.000 ;
        RECT 497.100 113.400 498.900 116.400 ;
        RECT 512.100 113.400 513.900 117.000 ;
        RECT 515.100 113.400 516.900 116.400 ;
        RECT 518.100 113.400 519.900 117.000 ;
        RECT 464.100 109.500 468.900 110.400 ;
        RECT 443.100 108.300 447.300 109.200 ;
        RECT 466.800 108.300 468.900 109.500 ;
        RECT 471.900 108.900 473.100 110.400 ;
        RECT 440.250 103.050 442.050 104.850 ;
        RECT 443.100 103.050 444.300 108.300 ;
        RECT 470.100 106.800 473.100 108.900 ;
        RECT 479.100 108.600 480.300 110.400 ;
        RECT 446.100 103.050 447.900 104.850 ;
        RECT 468.900 103.800 471.000 105.900 ;
        RECT 16.950 100.950 19.050 103.050 ;
        RECT 19.950 100.950 22.050 103.050 ;
        RECT 34.950 100.950 37.050 103.050 ;
        RECT 37.950 100.950 40.050 103.050 ;
        RECT 40.950 100.950 43.050 103.050 ;
        RECT 43.950 100.950 46.050 103.050 ;
        RECT 58.950 100.950 61.050 103.050 ;
        RECT 61.950 100.950 64.050 103.050 ;
        RECT 64.950 100.950 67.050 103.050 ;
        RECT 67.950 100.950 70.050 103.050 ;
        RECT 82.950 100.950 85.050 103.050 ;
        RECT 85.950 100.950 88.050 103.050 ;
        RECT 88.950 100.950 91.050 103.050 ;
        RECT 91.950 100.950 94.050 103.050 ;
        RECT 106.950 100.950 109.050 103.050 ;
        RECT 109.950 100.950 112.050 103.050 ;
        RECT 112.950 100.950 115.050 103.050 ;
        RECT 115.950 100.950 118.050 103.050 ;
        RECT 133.950 100.950 136.050 103.050 ;
        RECT 136.950 100.950 139.050 103.050 ;
        RECT 139.950 100.950 142.050 103.050 ;
        RECT 142.950 100.950 145.050 103.050 ;
        RECT 160.950 100.950 163.050 103.050 ;
        RECT 163.950 100.950 166.050 103.050 ;
        RECT 178.950 100.950 181.050 103.050 ;
        RECT 181.950 100.950 184.050 103.050 ;
        RECT 184.950 100.950 187.050 103.050 ;
        RECT 187.950 100.950 190.050 103.050 ;
        RECT 205.950 100.950 208.050 103.050 ;
        RECT 208.950 100.950 211.050 103.050 ;
        RECT 211.950 100.950 214.050 103.050 ;
        RECT 214.950 100.950 217.050 103.050 ;
        RECT 229.950 100.950 232.050 103.050 ;
        RECT 232.950 100.950 235.050 103.050 ;
        RECT 235.950 100.950 238.050 103.050 ;
        RECT 253.950 100.950 256.050 103.050 ;
        RECT 256.950 100.950 259.050 103.050 ;
        RECT 259.950 100.950 262.050 103.050 ;
        RECT 262.950 100.950 265.050 103.050 ;
        RECT 265.950 100.950 268.050 103.050 ;
        RECT 280.950 100.950 283.050 103.050 ;
        RECT 283.950 100.950 286.050 103.050 ;
        RECT 286.950 100.950 289.050 103.050 ;
        RECT 301.950 100.950 304.050 103.050 ;
        RECT 304.950 100.950 307.050 103.050 ;
        RECT 307.950 100.950 310.050 103.050 ;
        RECT 310.950 100.950 313.050 103.050 ;
        RECT 328.800 100.950 330.900 103.050 ;
        RECT 334.950 100.950 337.050 103.050 ;
        RECT 337.950 100.950 340.050 103.050 ;
        RECT 343.500 100.950 345.600 103.050 ;
        RECT 361.950 100.950 364.050 103.050 ;
        RECT 364.950 100.950 367.050 103.050 ;
        RECT 367.950 100.950 370.050 103.050 ;
        RECT 382.950 100.950 385.050 103.050 ;
        RECT 385.950 100.950 388.050 103.050 ;
        RECT 388.950 100.950 391.050 103.050 ;
        RECT 403.950 100.950 406.050 103.050 ;
        RECT 406.950 100.950 409.050 103.050 ;
        RECT 421.950 100.950 424.050 103.050 ;
        RECT 424.950 100.950 427.050 103.050 ;
        RECT 439.950 100.950 442.050 103.050 ;
        RECT 442.950 100.950 445.050 103.050 ;
        RECT 445.950 100.950 448.050 103.050 ;
        RECT 464.100 100.950 466.200 103.050 ;
        RECT 468.900 102.000 470.700 103.800 ;
        RECT 471.900 101.100 473.100 106.800 ;
        RECT 474.000 107.700 480.300 108.600 ;
        RECT 474.000 105.600 476.100 107.700 ;
        RECT 474.000 103.800 475.800 105.600 ;
        RECT 478.800 103.050 480.600 104.850 ;
        RECT 497.100 103.050 498.300 113.400 ;
        RECT 515.700 103.050 516.600 113.400 ;
        RECT 533.100 111.300 534.900 116.400 ;
        RECT 536.100 112.200 537.900 117.000 ;
        RECT 539.100 111.300 540.900 116.400 ;
        RECT 533.100 109.950 540.900 111.300 ;
        RECT 542.100 110.400 543.900 116.400 ;
        RECT 557.100 113.400 558.900 117.000 ;
        RECT 560.100 113.400 561.900 116.400 ;
        RECT 542.100 108.300 543.300 110.400 ;
        RECT 539.700 107.400 543.300 108.300 ;
        RECT 536.100 103.050 537.900 104.850 ;
        RECT 539.700 103.050 540.900 107.400 ;
        RECT 542.100 103.050 543.900 104.850 ;
        RECT 560.100 103.050 561.300 113.400 ;
        RECT 571.950 109.950 574.050 112.050 ;
        RECT 579.000 110.400 580.800 117.000 ;
        RECT 583.500 111.600 585.300 116.400 ;
        RECT 586.500 113.400 588.300 117.000 ;
        RECT 583.500 110.400 588.600 111.600 ;
        RECT 572.550 106.050 573.450 109.950 ;
        RECT 574.950 108.450 577.050 109.050 ;
        RECT 580.950 108.450 583.050 109.050 ;
        RECT 574.950 107.550 583.050 108.450 ;
        RECT 574.950 106.950 577.050 107.550 ;
        RECT 580.950 106.950 583.050 107.550 ;
        RECT 571.950 103.950 574.050 106.050 ;
        RECT 578.100 103.050 579.900 104.850 ;
        RECT 584.250 103.050 586.050 104.850 ;
        RECT 587.700 103.050 588.600 110.400 ;
        RECT 602.100 107.400 603.900 117.000 ;
        RECT 608.700 108.000 610.500 116.400 ;
        RECT 608.700 106.800 612.000 108.000 ;
        RECT 626.100 107.400 627.900 117.000 ;
        RECT 632.700 108.000 634.500 116.400 ;
        RECT 654.000 110.400 655.800 117.000 ;
        RECT 658.500 111.600 660.300 116.400 ;
        RECT 661.500 113.400 663.300 117.000 ;
        RECT 658.500 110.400 663.600 111.600 ;
        RECT 643.950 108.450 646.050 109.050 ;
        RECT 655.950 108.450 658.050 109.050 ;
        RECT 632.700 106.800 636.000 108.000 ;
        RECT 643.950 107.550 658.050 108.450 ;
        RECT 643.950 106.950 646.050 107.550 ;
        RECT 655.950 106.950 658.050 107.550 ;
        RECT 602.100 103.050 603.900 104.850 ;
        RECT 608.100 103.050 609.900 104.850 ;
        RECT 611.100 103.050 612.000 106.800 ;
        RECT 613.950 105.450 616.050 106.050 ;
        RECT 613.950 104.550 621.450 105.450 ;
        RECT 613.950 103.950 616.050 104.550 ;
        RECT 478.800 102.300 480.900 103.050 ;
        RECT 17.100 99.150 18.900 100.950 ;
        RECT 20.100 87.600 21.300 100.950 ;
        RECT 38.250 99.150 40.050 100.950 ;
        RECT 44.700 93.600 45.600 100.950 ;
        RECT 62.100 99.150 63.900 100.950 ;
        RECT 35.100 92.700 42.900 93.600 ;
        RECT 17.100 81.000 18.900 87.600 ;
        RECT 20.100 81.600 21.900 87.600 ;
        RECT 35.100 81.600 36.900 92.700 ;
        RECT 38.100 81.000 39.900 91.800 ;
        RECT 41.100 81.600 42.900 92.700 ;
        RECT 44.100 81.600 45.900 93.600 ;
        RECT 68.100 88.800 69.000 100.950 ;
        RECT 62.400 87.900 69.000 88.800 ;
        RECT 62.400 87.600 63.900 87.900 ;
        RECT 59.100 81.000 60.900 87.600 ;
        RECT 62.100 81.600 63.900 87.600 ;
        RECT 68.100 87.600 69.000 87.900 ;
        RECT 84.000 88.800 84.900 100.950 ;
        RECT 89.100 99.150 90.900 100.950 ;
        RECT 110.250 99.150 112.050 100.950 ;
        RECT 91.950 96.450 94.050 97.050 ;
        RECT 112.950 96.450 115.050 97.050 ;
        RECT 91.950 95.550 115.050 96.450 ;
        RECT 91.950 94.950 94.050 95.550 ;
        RECT 112.950 94.950 115.050 95.550 ;
        RECT 85.950 93.450 88.050 94.050 ;
        RECT 103.950 93.450 106.050 94.050 ;
        RECT 116.700 93.600 117.600 100.950 ;
        RECT 134.100 99.150 135.900 100.950 ;
        RECT 140.700 93.600 141.900 100.950 ;
        RECT 161.100 99.150 162.900 100.950 ;
        RECT 85.950 92.550 106.050 93.450 ;
        RECT 85.950 91.950 88.050 92.550 ;
        RECT 103.950 91.950 106.050 92.550 ;
        RECT 107.100 92.700 114.900 93.600 ;
        RECT 84.000 87.900 90.600 88.800 ;
        RECT 84.000 87.600 84.900 87.900 ;
        RECT 65.100 81.000 66.900 87.000 ;
        RECT 68.100 81.600 69.900 87.600 ;
        RECT 83.100 81.600 84.900 87.600 ;
        RECT 89.100 87.600 90.600 87.900 ;
        RECT 86.100 81.000 87.900 87.000 ;
        RECT 89.100 81.600 90.900 87.600 ;
        RECT 92.100 81.000 93.900 87.600 ;
        RECT 107.100 81.600 108.900 92.700 ;
        RECT 110.100 81.000 111.900 91.800 ;
        RECT 113.100 81.600 114.900 92.700 ;
        RECT 116.100 81.600 117.900 93.600 ;
        RECT 134.400 81.000 136.200 93.600 ;
        RECT 139.500 92.100 141.900 93.600 ;
        RECT 139.500 81.600 141.300 92.100 ;
        RECT 142.200 89.100 144.000 90.900 ;
        RECT 164.100 87.600 165.300 100.950 ;
        RECT 179.100 99.150 180.900 100.950 ;
        RECT 185.700 93.600 186.900 100.950 ;
        RECT 209.250 99.150 211.050 100.950 ;
        RECT 215.700 93.600 216.600 100.950 ;
        RECT 142.500 81.000 144.300 87.600 ;
        RECT 161.100 81.000 162.900 87.600 ;
        RECT 164.100 81.600 165.900 87.600 ;
        RECT 179.400 81.000 181.200 93.600 ;
        RECT 184.500 92.100 186.900 93.600 ;
        RECT 206.100 92.700 213.900 93.600 ;
        RECT 184.500 81.600 186.300 92.100 ;
        RECT 187.200 89.100 189.000 90.900 ;
        RECT 187.500 81.000 189.300 87.600 ;
        RECT 206.100 81.600 207.900 92.700 ;
        RECT 209.100 81.000 210.900 91.800 ;
        RECT 212.100 81.600 213.900 92.700 ;
        RECT 215.100 81.600 216.900 93.600 ;
        RECT 233.100 87.600 234.300 100.950 ;
        RECT 257.100 99.150 258.900 100.950 ;
        RECT 261.000 95.400 261.900 100.950 ;
        RECT 262.950 99.150 264.750 100.950 ;
        RECT 281.250 99.150 283.050 100.950 ;
        RECT 257.100 94.500 261.900 95.400 ;
        RECT 230.100 81.000 231.900 87.600 ;
        RECT 233.100 81.600 234.900 87.600 ;
        RECT 236.100 81.000 237.900 87.600 ;
        RECT 254.100 82.500 255.900 93.600 ;
        RECT 257.100 83.400 258.900 94.500 ;
        RECT 284.400 93.600 285.300 100.950 ;
        RECT 287.100 99.150 288.900 100.950 ;
        RECT 302.100 99.150 303.900 100.950 ;
        RECT 292.950 96.450 295.050 97.050 ;
        RECT 301.950 96.450 304.050 96.750 ;
        RECT 292.950 95.550 304.050 96.450 ;
        RECT 292.950 94.950 295.050 95.550 ;
        RECT 301.950 94.650 304.050 95.550 ;
        RECT 308.700 93.600 309.900 100.950 ;
        RECT 329.100 99.150 330.900 100.950 ;
        RECT 338.250 99.150 340.050 100.950 ;
        RECT 260.100 92.400 267.900 93.300 ;
        RECT 260.100 82.500 261.900 92.400 ;
        RECT 254.100 81.600 261.900 82.500 ;
        RECT 263.100 81.000 264.900 91.500 ;
        RECT 266.100 81.600 267.900 92.400 ;
        RECT 281.100 81.000 282.900 93.600 ;
        RECT 284.400 92.400 288.000 93.600 ;
        RECT 286.200 81.600 288.000 92.400 ;
        RECT 302.400 81.000 304.200 93.600 ;
        RECT 307.500 92.100 309.900 93.600 ;
        RECT 307.500 81.600 309.300 92.100 ;
        RECT 326.100 91.500 333.900 92.400 ;
        RECT 310.200 89.100 312.000 90.900 ;
        RECT 310.500 81.000 312.300 87.600 ;
        RECT 326.100 81.600 327.900 91.500 ;
        RECT 329.100 81.000 330.900 90.600 ;
        RECT 332.100 82.500 333.900 91.500 ;
        RECT 335.100 91.200 342.900 92.100 ;
        RECT 335.100 83.400 336.900 91.200 ;
        RECT 338.100 82.500 339.900 90.300 ;
        RECT 332.100 81.600 339.900 82.500 ;
        RECT 341.100 82.500 342.900 91.200 ;
        RECT 344.100 91.200 345.300 100.950 ;
        RECT 362.250 99.150 364.050 100.950 ;
        RECT 365.400 93.600 366.300 100.950 ;
        RECT 368.100 99.150 369.900 100.950 ;
        RECT 383.250 99.150 385.050 100.950 ;
        RECT 386.400 93.600 387.300 100.950 ;
        RECT 389.100 99.150 390.900 100.950 ;
        RECT 404.100 99.150 405.900 100.950 ;
        RECT 344.100 83.400 345.900 91.200 ;
        RECT 347.100 82.500 348.900 91.800 ;
        RECT 341.100 81.600 348.900 82.500 ;
        RECT 362.100 81.000 363.900 93.600 ;
        RECT 365.400 92.400 369.000 93.600 ;
        RECT 367.200 81.600 369.000 92.400 ;
        RECT 383.100 81.000 384.900 93.600 ;
        RECT 386.400 92.400 390.000 93.600 ;
        RECT 388.200 81.600 390.000 92.400 ;
        RECT 407.100 87.600 408.300 100.950 ;
        RECT 422.100 99.150 423.900 100.950 ;
        RECT 425.100 87.600 426.300 100.950 ;
        RECT 443.100 87.600 444.300 100.950 ;
        RECT 464.400 99.150 466.200 100.950 ;
        RECT 470.700 100.200 473.100 101.100 ;
        RECT 474.000 100.950 480.900 102.300 ;
        RECT 493.950 100.950 496.050 103.050 ;
        RECT 496.950 100.950 499.050 103.050 ;
        RECT 511.950 100.950 514.050 103.050 ;
        RECT 514.950 100.950 517.050 103.050 ;
        RECT 517.950 100.950 520.050 103.050 ;
        RECT 532.950 100.950 535.050 103.050 ;
        RECT 535.950 100.950 538.050 103.050 ;
        RECT 538.950 100.950 541.050 103.050 ;
        RECT 541.950 100.950 544.050 103.050 ;
        RECT 556.950 100.950 559.050 103.050 ;
        RECT 559.950 100.950 562.050 103.050 ;
        RECT 577.950 100.950 580.050 103.050 ;
        RECT 580.950 100.950 583.050 103.050 ;
        RECT 583.950 100.950 586.050 103.050 ;
        RECT 586.950 100.950 589.050 103.050 ;
        RECT 601.950 100.950 604.050 103.050 ;
        RECT 604.950 100.950 607.050 103.050 ;
        RECT 607.950 100.950 610.050 103.050 ;
        RECT 610.950 100.950 613.050 103.050 ;
        RECT 474.000 100.500 475.800 100.950 ;
        RECT 470.700 100.050 472.200 100.200 ;
        RECT 470.100 97.950 472.200 100.050 ;
        RECT 471.300 96.000 472.200 97.950 ;
        RECT 473.100 97.500 477.000 99.300 ;
        RECT 494.100 99.150 495.900 100.950 ;
        RECT 473.100 97.200 475.200 97.500 ;
        RECT 471.300 94.950 472.800 96.000 ;
        RECT 466.800 93.600 468.900 94.500 ;
        RECT 464.100 92.400 468.900 93.600 ;
        RECT 471.600 93.600 472.800 94.950 ;
        RECT 476.400 93.600 478.500 95.700 ;
        RECT 404.100 81.000 405.900 87.600 ;
        RECT 407.100 81.600 408.900 87.600 ;
        RECT 422.100 81.000 423.900 87.600 ;
        RECT 425.100 81.600 426.900 87.600 ;
        RECT 440.100 81.000 441.900 87.600 ;
        RECT 443.100 81.600 444.900 87.600 ;
        RECT 446.100 81.000 447.900 87.600 ;
        RECT 464.100 81.600 465.900 92.400 ;
        RECT 467.100 81.000 468.900 91.500 ;
        RECT 471.600 81.600 473.400 93.600 ;
        RECT 476.400 92.700 480.900 93.600 ;
        RECT 476.100 81.000 477.900 91.500 ;
        RECT 479.100 81.600 480.900 92.700 ;
        RECT 497.100 87.600 498.300 100.950 ;
        RECT 512.100 99.150 513.900 100.950 ;
        RECT 515.700 93.600 516.600 100.950 ;
        RECT 517.950 99.150 519.750 100.950 ;
        RECT 533.100 99.150 534.900 100.950 ;
        RECT 539.700 93.600 540.900 100.950 ;
        RECT 557.100 99.150 558.900 100.950 ;
        RECT 513.000 92.400 516.600 93.600 ;
        RECT 494.100 81.000 495.900 87.600 ;
        RECT 497.100 81.600 498.900 87.600 ;
        RECT 513.000 81.600 514.800 92.400 ;
        RECT 518.100 81.000 519.900 93.600 ;
        RECT 533.400 81.000 535.200 93.600 ;
        RECT 538.500 92.100 540.900 93.600 ;
        RECT 538.500 81.600 540.300 92.100 ;
        RECT 541.200 89.100 543.000 90.900 ;
        RECT 560.100 87.600 561.300 100.950 ;
        RECT 581.250 99.150 583.050 100.950 ;
        RECT 565.950 96.450 568.050 97.050 ;
        RECT 577.950 96.450 580.050 97.050 ;
        RECT 565.950 95.550 580.050 96.450 ;
        RECT 565.950 94.950 568.050 95.550 ;
        RECT 577.950 94.950 580.050 95.550 ;
        RECT 587.700 93.600 588.600 100.950 ;
        RECT 605.100 99.150 606.900 100.950 ;
        RECT 589.950 96.450 592.050 97.050 ;
        RECT 607.950 96.450 610.050 97.050 ;
        RECT 589.950 95.550 610.050 96.450 ;
        RECT 589.950 94.950 592.050 95.550 ;
        RECT 607.950 94.950 610.050 95.550 ;
        RECT 578.100 92.700 585.900 93.600 ;
        RECT 541.500 81.000 543.300 87.600 ;
        RECT 557.100 81.000 558.900 87.600 ;
        RECT 560.100 81.600 561.900 87.600 ;
        RECT 578.100 81.600 579.900 92.700 ;
        RECT 581.100 81.000 582.900 91.800 ;
        RECT 584.100 81.600 585.900 92.700 ;
        RECT 587.100 81.600 588.900 93.600 ;
        RECT 611.100 88.800 612.000 100.950 ;
        RECT 620.550 100.050 621.450 104.550 ;
        RECT 626.100 103.050 627.900 104.850 ;
        RECT 632.100 103.050 633.900 104.850 ;
        RECT 635.100 103.050 636.000 106.800 ;
        RECT 653.100 103.050 654.900 104.850 ;
        RECT 659.250 103.050 661.050 104.850 ;
        RECT 662.700 103.050 663.600 110.400 ;
        RECT 682.500 108.000 684.300 116.400 ;
        RECT 681.000 106.800 684.300 108.000 ;
        RECT 689.100 107.400 690.900 117.000 ;
        RECT 704.100 111.300 705.900 116.400 ;
        RECT 707.100 112.200 708.900 117.000 ;
        RECT 710.100 111.300 711.900 116.400 ;
        RECT 704.100 109.950 711.900 111.300 ;
        RECT 713.100 110.400 714.900 116.400 ;
        RECT 728.100 110.400 729.900 116.400 ;
        RECT 713.100 108.300 714.300 110.400 ;
        RECT 710.700 107.400 714.300 108.300 ;
        RECT 728.700 108.300 729.900 110.400 ;
        RECT 731.100 111.300 732.900 116.400 ;
        RECT 734.100 112.200 735.900 117.000 ;
        RECT 737.100 111.300 738.900 116.400 ;
        RECT 755.100 113.400 756.900 117.000 ;
        RECT 758.100 113.400 759.900 116.400 ;
        RECT 731.100 109.950 738.900 111.300 ;
        RECT 728.700 107.400 732.300 108.300 ;
        RECT 681.000 103.050 681.900 106.800 ;
        RECT 683.100 103.050 684.900 104.850 ;
        RECT 689.100 103.050 690.900 104.850 ;
        RECT 707.100 103.050 708.900 104.850 ;
        RECT 710.700 103.050 711.900 107.400 ;
        RECT 713.100 103.050 714.900 104.850 ;
        RECT 728.100 103.050 729.900 104.850 ;
        RECT 731.100 103.050 732.300 107.400 ;
        RECT 734.100 103.050 735.900 104.850 ;
        RECT 758.100 103.050 759.300 113.400 ;
        RECT 774.000 110.400 775.800 117.000 ;
        RECT 778.500 111.600 780.300 116.400 ;
        RECT 781.500 113.400 783.300 117.000 ;
        RECT 797.700 113.400 799.500 117.000 ;
        RECT 800.700 111.600 802.500 116.400 ;
        RECT 778.500 110.400 783.600 111.600 ;
        RECT 766.950 108.450 769.050 109.050 ;
        RECT 778.950 108.450 781.050 109.050 ;
        RECT 766.950 107.550 781.050 108.450 ;
        RECT 766.950 106.950 769.050 107.550 ;
        RECT 778.950 106.950 781.050 107.550 ;
        RECT 773.100 103.050 774.900 104.850 ;
        RECT 779.250 103.050 781.050 104.850 ;
        RECT 782.700 103.050 783.600 110.400 ;
        RECT 797.400 110.400 802.500 111.600 ;
        RECT 805.200 110.400 807.000 117.000 ;
        RECT 797.400 103.050 798.300 110.400 ;
        RECT 821.100 107.400 822.900 117.000 ;
        RECT 827.700 108.000 829.500 116.400 ;
        RECT 845.100 110.400 846.900 116.400 ;
        RECT 845.700 108.300 846.900 110.400 ;
        RECT 848.100 111.300 849.900 116.400 ;
        RECT 851.100 112.200 852.900 117.000 ;
        RECT 854.100 111.300 855.900 116.400 ;
        RECT 848.100 109.950 855.900 111.300 ;
        RECT 869.100 111.300 870.900 116.400 ;
        RECT 872.100 112.200 873.900 117.000 ;
        RECT 875.100 111.300 876.900 116.400 ;
        RECT 869.100 109.950 876.900 111.300 ;
        RECT 878.100 110.400 879.900 116.400 ;
        RECT 878.100 108.300 879.300 110.400 ;
        RECT 827.700 106.800 831.000 108.000 ;
        RECT 845.700 107.400 849.300 108.300 ;
        RECT 799.950 103.050 801.750 104.850 ;
        RECT 806.100 103.050 807.900 104.850 ;
        RECT 821.100 103.050 822.900 104.850 ;
        RECT 827.100 103.050 828.900 104.850 ;
        RECT 830.100 103.050 831.000 106.800 ;
        RECT 845.100 103.050 846.900 104.850 ;
        RECT 848.100 103.050 849.300 107.400 ;
        RECT 875.700 107.400 879.300 108.300 ;
        RECT 895.500 108.000 897.300 116.400 ;
        RECT 851.100 103.050 852.900 104.850 ;
        RECT 872.100 103.050 873.900 104.850 ;
        RECT 875.700 103.050 876.900 107.400 ;
        RECT 894.000 106.800 897.300 108.000 ;
        RECT 902.100 107.400 903.900 117.000 ;
        RECT 917.100 107.400 918.900 117.000 ;
        RECT 923.700 108.000 925.500 116.400 ;
        RECT 941.100 111.300 942.900 116.400 ;
        RECT 944.100 112.200 945.900 117.000 ;
        RECT 947.100 111.300 948.900 116.400 ;
        RECT 941.100 109.950 948.900 111.300 ;
        RECT 950.100 110.400 951.900 116.400 ;
        RECT 965.100 113.400 966.900 117.000 ;
        RECT 968.100 113.400 969.900 116.400 ;
        RECT 986.700 113.400 988.500 117.000 ;
        RECT 950.100 108.300 951.300 110.400 ;
        RECT 923.700 106.800 927.000 108.000 ;
        RECT 878.100 103.050 879.900 104.850 ;
        RECT 894.000 103.050 894.900 106.800 ;
        RECT 896.100 103.050 897.900 104.850 ;
        RECT 902.100 103.050 903.900 104.850 ;
        RECT 917.100 103.050 918.900 104.850 ;
        RECT 923.100 103.050 924.900 104.850 ;
        RECT 926.100 103.050 927.000 106.800 ;
        RECT 947.700 107.400 951.300 108.300 ;
        RECT 944.100 103.050 945.900 104.850 ;
        RECT 947.700 103.050 948.900 107.400 ;
        RECT 950.100 103.050 951.900 104.850 ;
        RECT 968.100 103.050 969.300 113.400 ;
        RECT 989.700 111.600 991.500 116.400 ;
        RECT 986.400 110.400 991.500 111.600 ;
        RECT 994.200 110.400 996.000 117.000 ;
        RECT 986.400 103.050 987.300 110.400 ;
        RECT 988.950 103.050 990.750 104.850 ;
        RECT 995.100 103.050 996.900 104.850 ;
        RECT 625.950 100.950 628.050 103.050 ;
        RECT 628.950 100.950 631.050 103.050 ;
        RECT 631.950 100.950 634.050 103.050 ;
        RECT 634.950 100.950 637.050 103.050 ;
        RECT 652.950 100.950 655.050 103.050 ;
        RECT 655.950 100.950 658.050 103.050 ;
        RECT 658.950 100.950 661.050 103.050 ;
        RECT 661.950 100.950 664.050 103.050 ;
        RECT 679.950 100.950 682.050 103.050 ;
        RECT 682.950 100.950 685.050 103.050 ;
        RECT 685.950 100.950 688.050 103.050 ;
        RECT 688.950 100.950 691.050 103.050 ;
        RECT 703.950 100.950 706.050 103.050 ;
        RECT 706.950 100.950 709.050 103.050 ;
        RECT 709.950 100.950 712.050 103.050 ;
        RECT 712.950 100.950 715.050 103.050 ;
        RECT 727.950 100.950 730.050 103.050 ;
        RECT 730.950 100.950 733.050 103.050 ;
        RECT 733.950 100.950 736.050 103.050 ;
        RECT 736.950 100.950 739.050 103.050 ;
        RECT 754.950 100.950 757.050 103.050 ;
        RECT 757.950 100.950 760.050 103.050 ;
        RECT 772.950 100.950 775.050 103.050 ;
        RECT 775.950 100.950 778.050 103.050 ;
        RECT 778.950 100.950 781.050 103.050 ;
        RECT 781.950 100.950 784.050 103.050 ;
        RECT 796.950 100.950 799.050 103.050 ;
        RECT 799.950 100.950 802.050 103.050 ;
        RECT 802.950 100.950 805.050 103.050 ;
        RECT 805.950 100.950 808.050 103.050 ;
        RECT 820.950 100.950 823.050 103.050 ;
        RECT 823.950 100.950 826.050 103.050 ;
        RECT 826.950 100.950 829.050 103.050 ;
        RECT 829.950 100.950 832.050 103.050 ;
        RECT 844.950 100.950 847.050 103.050 ;
        RECT 847.950 100.950 850.050 103.050 ;
        RECT 850.950 100.950 853.050 103.050 ;
        RECT 853.950 100.950 856.050 103.050 ;
        RECT 868.950 100.950 871.050 103.050 ;
        RECT 871.950 100.950 874.050 103.050 ;
        RECT 874.950 100.950 877.050 103.050 ;
        RECT 877.950 100.950 880.050 103.050 ;
        RECT 892.950 100.950 895.050 103.050 ;
        RECT 895.950 100.950 898.050 103.050 ;
        RECT 898.950 100.950 901.050 103.050 ;
        RECT 901.950 100.950 904.050 103.050 ;
        RECT 916.950 100.950 919.050 103.050 ;
        RECT 919.950 100.950 922.050 103.050 ;
        RECT 922.950 100.950 925.050 103.050 ;
        RECT 925.950 100.950 928.050 103.050 ;
        RECT 940.950 100.950 943.050 103.050 ;
        RECT 943.950 100.950 946.050 103.050 ;
        RECT 946.950 100.950 949.050 103.050 ;
        RECT 949.950 100.950 952.050 103.050 ;
        RECT 964.950 100.950 967.050 103.050 ;
        RECT 967.950 100.950 970.050 103.050 ;
        RECT 985.950 100.950 988.050 103.050 ;
        RECT 988.950 100.950 991.050 103.050 ;
        RECT 991.950 100.950 994.050 103.050 ;
        RECT 994.950 100.950 997.050 103.050 ;
        RECT 620.550 98.550 625.050 100.050 ;
        RECT 629.100 99.150 630.900 100.950 ;
        RECT 621.000 97.950 625.050 98.550 ;
        RECT 635.100 88.800 636.000 100.950 ;
        RECT 656.250 99.150 658.050 100.950 ;
        RECT 637.950 96.450 640.050 97.050 ;
        RECT 655.950 96.450 658.050 97.050 ;
        RECT 637.950 95.550 658.050 96.450 ;
        RECT 637.950 94.950 640.050 95.550 ;
        RECT 655.950 94.950 658.050 95.550 ;
        RECT 637.950 90.450 640.050 90.900 ;
        RECT 646.950 90.450 649.050 94.050 ;
        RECT 662.700 93.600 663.600 100.950 ;
        RECT 637.950 90.000 649.050 90.450 ;
        RECT 653.100 92.700 660.900 93.600 ;
        RECT 637.950 89.550 648.450 90.000 ;
        RECT 637.950 88.800 640.050 89.550 ;
        RECT 605.400 87.900 612.000 88.800 ;
        RECT 605.400 87.600 606.900 87.900 ;
        RECT 602.100 81.000 603.900 87.600 ;
        RECT 605.100 81.600 606.900 87.600 ;
        RECT 611.100 87.600 612.000 87.900 ;
        RECT 629.400 87.900 636.000 88.800 ;
        RECT 629.400 87.600 630.900 87.900 ;
        RECT 608.100 81.000 609.900 87.000 ;
        RECT 611.100 81.600 612.900 87.600 ;
        RECT 626.100 81.000 627.900 87.600 ;
        RECT 629.100 81.600 630.900 87.600 ;
        RECT 635.100 87.600 636.000 87.900 ;
        RECT 632.100 81.000 633.900 87.000 ;
        RECT 635.100 81.600 636.900 87.600 ;
        RECT 653.100 81.600 654.900 92.700 ;
        RECT 656.100 81.000 657.900 91.800 ;
        RECT 659.100 81.600 660.900 92.700 ;
        RECT 662.100 81.600 663.900 93.600 ;
        RECT 681.000 88.800 681.900 100.950 ;
        RECT 686.100 99.150 687.900 100.950 ;
        RECT 704.100 99.150 705.900 100.950 ;
        RECT 685.950 96.450 688.050 97.050 ;
        RECT 706.950 96.450 709.050 96.750 ;
        RECT 685.950 95.550 709.050 96.450 ;
        RECT 685.950 94.950 688.050 95.550 ;
        RECT 706.950 94.650 709.050 95.550 ;
        RECT 710.700 93.600 711.900 100.950 ;
        RECT 681.000 87.900 687.600 88.800 ;
        RECT 681.000 87.600 681.900 87.900 ;
        RECT 680.100 81.600 681.900 87.600 ;
        RECT 686.100 87.600 687.600 87.900 ;
        RECT 683.100 81.000 684.900 87.000 ;
        RECT 686.100 81.600 687.900 87.600 ;
        RECT 689.100 81.000 690.900 87.600 ;
        RECT 704.400 81.000 706.200 93.600 ;
        RECT 709.500 92.100 711.900 93.600 ;
        RECT 731.100 93.600 732.300 100.950 ;
        RECT 737.100 99.150 738.900 100.950 ;
        RECT 755.100 99.150 756.900 100.950 ;
        RECT 731.100 92.100 733.500 93.600 ;
        RECT 709.500 81.600 711.300 92.100 ;
        RECT 712.200 89.100 714.000 90.900 ;
        RECT 729.000 89.100 730.800 90.900 ;
        RECT 712.500 81.000 714.300 87.600 ;
        RECT 728.700 81.000 730.500 87.600 ;
        RECT 731.700 81.600 733.500 92.100 ;
        RECT 736.800 81.000 738.600 93.600 ;
        RECT 758.100 87.600 759.300 100.950 ;
        RECT 776.250 99.150 778.050 100.950 ;
        RECT 760.950 96.450 763.050 97.050 ;
        RECT 778.950 96.450 781.050 97.050 ;
        RECT 760.950 95.550 781.050 96.450 ;
        RECT 760.950 94.950 763.050 95.550 ;
        RECT 778.950 94.950 781.050 95.550 ;
        RECT 782.700 93.600 783.600 100.950 ;
        RECT 797.400 93.600 798.300 100.950 ;
        RECT 802.950 99.150 804.750 100.950 ;
        RECT 824.100 99.150 825.900 100.950 ;
        RECT 805.950 96.450 808.050 97.050 ;
        RECT 826.950 96.450 829.050 97.050 ;
        RECT 805.950 95.550 829.050 96.450 ;
        RECT 805.950 94.950 808.050 95.550 ;
        RECT 826.950 94.950 829.050 95.550 ;
        RECT 773.100 92.700 780.900 93.600 ;
        RECT 755.100 81.000 756.900 87.600 ;
        RECT 758.100 81.600 759.900 87.600 ;
        RECT 773.100 81.600 774.900 92.700 ;
        RECT 776.100 81.000 777.900 91.800 ;
        RECT 779.100 81.600 780.900 92.700 ;
        RECT 782.100 81.600 783.900 93.600 ;
        RECT 797.100 81.600 798.900 93.600 ;
        RECT 800.100 92.700 807.900 93.600 ;
        RECT 800.100 81.600 801.900 92.700 ;
        RECT 803.100 81.000 804.900 91.800 ;
        RECT 806.100 81.600 807.900 92.700 ;
        RECT 808.950 93.450 811.050 94.050 ;
        RECT 823.950 93.450 826.050 93.900 ;
        RECT 808.950 92.550 826.050 93.450 ;
        RECT 808.950 91.950 811.050 92.550 ;
        RECT 823.950 91.800 826.050 92.550 ;
        RECT 830.100 88.800 831.000 100.950 ;
        RECT 848.100 93.600 849.300 100.950 ;
        RECT 854.100 99.150 855.900 100.950 ;
        RECT 869.100 99.150 870.900 100.950 ;
        RECT 875.700 93.600 876.900 100.950 ;
        RECT 848.100 92.100 850.500 93.600 ;
        RECT 846.000 89.100 847.800 90.900 ;
        RECT 824.400 87.900 831.000 88.800 ;
        RECT 824.400 87.600 825.900 87.900 ;
        RECT 821.100 81.000 822.900 87.600 ;
        RECT 824.100 81.600 825.900 87.600 ;
        RECT 830.100 87.600 831.000 87.900 ;
        RECT 827.100 81.000 828.900 87.000 ;
        RECT 830.100 81.600 831.900 87.600 ;
        RECT 845.700 81.000 847.500 87.600 ;
        RECT 848.700 81.600 850.500 92.100 ;
        RECT 853.800 81.000 855.600 93.600 ;
        RECT 869.400 81.000 871.200 93.600 ;
        RECT 874.500 92.100 876.900 93.600 ;
        RECT 874.500 81.600 876.300 92.100 ;
        RECT 877.200 89.100 879.000 90.900 ;
        RECT 894.000 88.800 894.900 100.950 ;
        RECT 899.100 99.150 900.900 100.950 ;
        RECT 920.100 99.150 921.900 100.950 ;
        RECT 907.950 96.450 910.050 97.050 ;
        RECT 922.950 96.450 925.050 97.050 ;
        RECT 907.950 95.550 925.050 96.450 ;
        RECT 907.950 94.950 910.050 95.550 ;
        RECT 922.950 94.950 925.050 95.550 ;
        RECT 926.100 88.800 927.000 100.950 ;
        RECT 941.100 99.150 942.900 100.950 ;
        RECT 947.700 93.600 948.900 100.950 ;
        RECT 965.100 99.150 966.900 100.950 ;
        RECT 894.000 87.900 900.600 88.800 ;
        RECT 894.000 87.600 894.900 87.900 ;
        RECT 877.500 81.000 879.300 87.600 ;
        RECT 893.100 81.600 894.900 87.600 ;
        RECT 899.100 87.600 900.600 87.900 ;
        RECT 920.400 87.900 927.000 88.800 ;
        RECT 920.400 87.600 921.900 87.900 ;
        RECT 896.100 81.000 897.900 87.000 ;
        RECT 899.100 81.600 900.900 87.600 ;
        RECT 902.100 81.000 903.900 87.600 ;
        RECT 917.100 81.000 918.900 87.600 ;
        RECT 920.100 81.600 921.900 87.600 ;
        RECT 926.100 87.600 927.000 87.900 ;
        RECT 923.100 81.000 924.900 87.000 ;
        RECT 926.100 81.600 927.900 87.600 ;
        RECT 941.400 81.000 943.200 93.600 ;
        RECT 946.500 92.100 948.900 93.600 ;
        RECT 946.500 81.600 948.300 92.100 ;
        RECT 949.200 89.100 951.000 90.900 ;
        RECT 968.100 87.600 969.300 100.950 ;
        RECT 986.400 93.600 987.300 100.950 ;
        RECT 991.950 99.150 993.750 100.950 ;
        RECT 994.950 96.450 997.050 97.050 ;
        RECT 1000.950 96.450 1003.050 97.050 ;
        RECT 994.950 95.550 1003.050 96.450 ;
        RECT 994.950 94.950 997.050 95.550 ;
        RECT 1000.950 94.950 1003.050 95.550 ;
        RECT 949.500 81.000 951.300 87.600 ;
        RECT 965.100 81.000 966.900 87.600 ;
        RECT 968.100 81.600 969.900 87.600 ;
        RECT 986.100 81.600 987.900 93.600 ;
        RECT 989.100 92.700 996.900 93.600 ;
        RECT 989.100 81.600 990.900 92.700 ;
        RECT 992.100 81.000 993.900 91.800 ;
        RECT 995.100 81.600 996.900 92.700 ;
        RECT 17.400 65.400 19.200 78.000 ;
        RECT 22.500 66.900 24.300 77.400 ;
        RECT 25.500 71.400 27.300 78.000 ;
        RECT 41.100 71.400 42.900 78.000 ;
        RECT 44.100 71.400 45.900 77.400 ;
        RECT 25.200 68.100 27.000 69.900 ;
        RECT 22.500 65.400 24.900 66.900 ;
        RECT 17.100 58.050 18.900 59.850 ;
        RECT 23.700 58.050 24.900 65.400 ;
        RECT 41.100 58.050 42.900 59.850 ;
        RECT 44.100 58.050 45.300 71.400 ;
        RECT 59.400 65.400 61.200 78.000 ;
        RECT 64.500 66.900 66.300 77.400 ;
        RECT 67.500 71.400 69.300 78.000 ;
        RECT 86.100 71.400 87.900 78.000 ;
        RECT 89.100 71.400 90.900 77.400 ;
        RECT 107.100 71.400 108.900 78.000 ;
        RECT 110.100 71.400 111.900 77.400 ;
        RECT 113.100 72.000 114.900 78.000 ;
        RECT 67.200 68.100 69.000 69.900 ;
        RECT 64.500 65.400 66.900 66.900 ;
        RECT 46.950 63.450 49.050 64.050 ;
        RECT 61.950 63.450 64.050 64.050 ;
        RECT 46.950 62.550 64.050 63.450 ;
        RECT 46.950 61.950 49.050 62.550 ;
        RECT 61.950 61.950 64.050 62.550 ;
        RECT 59.100 58.050 60.900 59.850 ;
        RECT 65.700 58.050 66.900 65.400 ;
        RECT 86.100 58.050 87.900 59.850 ;
        RECT 89.100 58.050 90.300 71.400 ;
        RECT 110.400 71.100 111.900 71.400 ;
        RECT 116.100 71.400 117.900 77.400 ;
        RECT 131.700 71.400 133.500 78.000 ;
        RECT 116.100 71.100 117.000 71.400 ;
        RECT 110.400 70.200 117.000 71.100 ;
        RECT 110.100 58.050 111.900 59.850 ;
        RECT 116.100 58.050 117.000 70.200 ;
        RECT 132.000 68.100 133.800 69.900 ;
        RECT 134.700 66.900 136.500 77.400 ;
        RECT 134.100 65.400 136.500 66.900 ;
        RECT 139.800 65.400 141.600 78.000 ;
        RECT 158.100 71.400 159.900 77.400 ;
        RECT 161.100 71.400 162.900 78.000 ;
        RECT 179.100 71.400 180.900 78.000 ;
        RECT 182.100 71.400 183.900 77.400 ;
        RECT 185.100 72.000 186.900 78.000 ;
        RECT 134.100 58.050 135.300 65.400 ;
        RECT 140.100 58.050 141.900 59.850 ;
        RECT 158.700 58.050 159.900 71.400 ;
        RECT 182.400 71.100 183.900 71.400 ;
        RECT 188.100 71.400 189.900 77.400 ;
        RECT 203.100 71.400 204.900 78.000 ;
        RECT 206.100 71.400 207.900 77.400 ;
        RECT 209.100 72.000 210.900 78.000 ;
        RECT 188.100 71.100 189.000 71.400 ;
        RECT 182.400 70.200 189.000 71.100 ;
        RECT 206.400 71.100 207.900 71.400 ;
        RECT 212.100 71.400 213.900 77.400 ;
        RECT 212.100 71.100 213.000 71.400 ;
        RECT 206.400 70.200 213.000 71.100 ;
        RECT 161.100 58.050 162.900 59.850 ;
        RECT 182.100 58.050 183.900 59.850 ;
        RECT 188.100 58.050 189.000 70.200 ;
        RECT 206.100 58.050 207.900 59.850 ;
        RECT 212.100 58.050 213.000 70.200 ;
        RECT 227.100 66.600 228.900 77.400 ;
        RECT 230.100 67.500 231.900 78.000 ;
        RECT 233.100 76.500 240.900 77.400 ;
        RECT 233.100 66.600 234.900 76.500 ;
        RECT 227.100 65.700 234.900 66.600 ;
        RECT 236.100 64.500 237.900 75.600 ;
        RECT 239.100 65.400 240.900 76.500 ;
        RECT 254.100 71.400 255.900 78.000 ;
        RECT 257.100 71.400 258.900 77.400 ;
        RECT 260.100 72.000 261.900 78.000 ;
        RECT 257.400 71.100 258.900 71.400 ;
        RECT 263.100 71.400 264.900 77.400 ;
        RECT 281.100 71.400 282.900 78.000 ;
        RECT 284.100 71.400 285.900 77.400 ;
        RECT 287.100 72.000 288.900 78.000 ;
        RECT 263.100 71.100 264.000 71.400 ;
        RECT 257.400 70.200 264.000 71.100 ;
        RECT 284.400 71.100 285.900 71.400 ;
        RECT 290.100 71.400 291.900 77.400 ;
        RECT 305.100 71.400 306.900 78.000 ;
        RECT 308.100 71.400 309.900 77.400 ;
        RECT 311.100 72.000 312.900 78.000 ;
        RECT 290.100 71.100 291.000 71.400 ;
        RECT 284.400 70.200 291.000 71.100 ;
        RECT 308.400 71.100 309.900 71.400 ;
        RECT 314.100 71.400 315.900 77.400 ;
        RECT 314.100 71.100 315.000 71.400 ;
        RECT 308.400 70.200 315.000 71.100 ;
        RECT 233.100 63.600 237.900 64.500 ;
        RECT 230.250 58.050 232.050 59.850 ;
        RECT 233.100 58.050 234.000 63.600 ;
        RECT 236.100 58.050 237.900 59.850 ;
        RECT 257.100 58.050 258.900 59.850 ;
        RECT 263.100 58.050 264.000 70.200 ;
        RECT 284.100 58.050 285.900 59.850 ;
        RECT 290.100 58.050 291.000 70.200 ;
        RECT 308.100 58.050 309.900 59.850 ;
        RECT 314.100 58.050 315.000 70.200 ;
        RECT 332.100 66.300 333.900 77.400 ;
        RECT 335.100 67.200 336.900 78.000 ;
        RECT 338.100 66.300 339.900 77.400 ;
        RECT 332.100 65.400 339.900 66.300 ;
        RECT 341.100 65.400 342.900 77.400 ;
        RECT 359.100 71.400 360.900 78.000 ;
        RECT 362.100 71.400 363.900 77.400 ;
        RECT 365.100 72.000 366.900 78.000 ;
        RECT 362.400 71.100 363.900 71.400 ;
        RECT 368.100 71.400 369.900 77.400 ;
        RECT 368.100 71.100 369.000 71.400 ;
        RECT 362.400 70.200 369.000 71.100 ;
        RECT 335.250 58.050 337.050 59.850 ;
        RECT 341.700 58.050 342.600 65.400 ;
        RECT 362.100 58.050 363.900 59.850 ;
        RECT 368.100 58.050 369.000 70.200 ;
        RECT 386.100 66.300 387.900 77.400 ;
        RECT 389.100 67.200 390.900 78.000 ;
        RECT 392.100 66.300 393.900 77.400 ;
        RECT 386.100 65.400 393.900 66.300 ;
        RECT 395.100 65.400 396.900 77.400 ;
        RECT 410.400 65.400 412.200 78.000 ;
        RECT 415.500 66.900 417.300 77.400 ;
        RECT 418.500 71.400 420.300 78.000 ;
        RECT 418.200 68.100 420.000 69.900 ;
        RECT 415.500 65.400 417.900 66.900 ;
        RECT 434.400 65.400 436.200 78.000 ;
        RECT 439.500 66.900 441.300 77.400 ;
        RECT 442.500 71.400 444.300 78.000 ;
        RECT 458.100 71.400 459.900 77.400 ;
        RECT 461.100 72.000 462.900 78.000 ;
        RECT 459.000 71.100 459.900 71.400 ;
        RECT 464.100 71.400 465.900 77.400 ;
        RECT 467.100 71.400 468.900 78.000 ;
        RECT 485.100 71.400 486.900 78.000 ;
        RECT 488.100 71.400 489.900 77.400 ;
        RECT 491.100 71.400 492.900 78.000 ;
        RECT 509.100 71.400 510.900 78.000 ;
        RECT 512.100 71.400 513.900 77.400 ;
        RECT 464.100 71.100 465.600 71.400 ;
        RECT 459.000 70.200 465.600 71.100 ;
        RECT 442.200 68.100 444.000 69.900 ;
        RECT 439.500 65.400 441.900 66.900 ;
        RECT 389.250 58.050 391.050 59.850 ;
        RECT 395.700 58.050 396.600 65.400 ;
        RECT 410.100 58.050 411.900 59.850 ;
        RECT 416.700 58.050 417.900 65.400 ;
        RECT 430.950 60.450 433.050 61.050 ;
        RECT 425.550 59.550 433.050 60.450 ;
        RECT 16.950 55.950 19.050 58.050 ;
        RECT 19.950 55.950 22.050 58.050 ;
        RECT 22.950 55.950 25.050 58.050 ;
        RECT 25.950 55.950 28.050 58.050 ;
        RECT 40.950 55.950 43.050 58.050 ;
        RECT 43.950 55.950 46.050 58.050 ;
        RECT 58.950 55.950 61.050 58.050 ;
        RECT 61.950 55.950 64.050 58.050 ;
        RECT 64.950 55.950 67.050 58.050 ;
        RECT 67.950 55.950 70.050 58.050 ;
        RECT 85.950 55.950 88.050 58.050 ;
        RECT 88.950 55.950 91.050 58.050 ;
        RECT 106.950 55.950 109.050 58.050 ;
        RECT 109.950 55.950 112.050 58.050 ;
        RECT 112.950 55.950 115.050 58.050 ;
        RECT 115.950 55.950 118.050 58.050 ;
        RECT 130.950 55.950 133.050 58.050 ;
        RECT 133.950 55.950 136.050 58.050 ;
        RECT 136.950 55.950 139.050 58.050 ;
        RECT 139.950 55.950 142.050 58.050 ;
        RECT 157.950 55.950 160.050 58.050 ;
        RECT 160.950 55.950 163.050 58.050 ;
        RECT 178.950 55.950 181.050 58.050 ;
        RECT 181.950 55.950 184.050 58.050 ;
        RECT 184.950 55.950 187.050 58.050 ;
        RECT 187.950 55.950 190.050 58.050 ;
        RECT 202.950 55.950 205.050 58.050 ;
        RECT 205.950 55.950 208.050 58.050 ;
        RECT 208.950 55.950 211.050 58.050 ;
        RECT 211.950 55.950 214.050 58.050 ;
        RECT 226.950 55.950 229.050 58.050 ;
        RECT 229.950 55.950 232.050 58.050 ;
        RECT 232.950 55.950 235.050 58.050 ;
        RECT 235.950 55.950 238.050 58.050 ;
        RECT 238.950 55.950 241.050 58.050 ;
        RECT 253.950 55.950 256.050 58.050 ;
        RECT 256.950 55.950 259.050 58.050 ;
        RECT 259.950 55.950 262.050 58.050 ;
        RECT 262.950 55.950 265.050 58.050 ;
        RECT 280.950 55.950 283.050 58.050 ;
        RECT 283.950 55.950 286.050 58.050 ;
        RECT 286.950 55.950 289.050 58.050 ;
        RECT 289.950 55.950 292.050 58.050 ;
        RECT 304.950 55.950 307.050 58.050 ;
        RECT 307.950 55.950 310.050 58.050 ;
        RECT 310.950 55.950 313.050 58.050 ;
        RECT 313.950 55.950 316.050 58.050 ;
        RECT 331.950 55.950 334.050 58.050 ;
        RECT 334.950 55.950 337.050 58.050 ;
        RECT 337.950 55.950 340.050 58.050 ;
        RECT 340.950 55.950 343.050 58.050 ;
        RECT 358.950 55.950 361.050 58.050 ;
        RECT 361.950 55.950 364.050 58.050 ;
        RECT 364.950 55.950 367.050 58.050 ;
        RECT 367.950 55.950 370.050 58.050 ;
        RECT 385.950 55.950 388.050 58.050 ;
        RECT 388.950 55.950 391.050 58.050 ;
        RECT 391.950 55.950 394.050 58.050 ;
        RECT 394.950 55.950 397.050 58.050 ;
        RECT 409.950 55.950 412.050 58.050 ;
        RECT 412.950 55.950 415.050 58.050 ;
        RECT 415.950 55.950 418.050 58.050 ;
        RECT 418.950 55.950 421.050 58.050 ;
        RECT 20.100 54.150 21.900 55.950 ;
        RECT 23.700 51.600 24.900 55.950 ;
        RECT 26.100 54.150 27.900 55.950 ;
        RECT 23.700 50.700 27.300 51.600 ;
        RECT 17.100 47.700 24.900 49.050 ;
        RECT 17.100 42.600 18.900 47.700 ;
        RECT 20.100 42.000 21.900 46.800 ;
        RECT 23.100 42.600 24.900 47.700 ;
        RECT 26.100 48.600 27.300 50.700 ;
        RECT 26.100 42.600 27.900 48.600 ;
        RECT 44.100 45.600 45.300 55.950 ;
        RECT 62.100 54.150 63.900 55.950 ;
        RECT 65.700 51.600 66.900 55.950 ;
        RECT 68.100 54.150 69.900 55.950 ;
        RECT 65.700 50.700 69.300 51.600 ;
        RECT 59.100 47.700 66.900 49.050 ;
        RECT 41.100 42.000 42.900 45.600 ;
        RECT 44.100 42.600 45.900 45.600 ;
        RECT 59.100 42.600 60.900 47.700 ;
        RECT 62.100 42.000 63.900 46.800 ;
        RECT 65.100 42.600 66.900 47.700 ;
        RECT 68.100 48.600 69.300 50.700 ;
        RECT 68.100 42.600 69.900 48.600 ;
        RECT 89.100 45.600 90.300 55.950 ;
        RECT 107.100 54.150 108.900 55.950 ;
        RECT 113.100 54.150 114.900 55.950 ;
        RECT 116.100 52.200 117.000 55.950 ;
        RECT 131.100 54.150 132.900 55.950 ;
        RECT 86.100 42.000 87.900 45.600 ;
        RECT 89.100 42.600 90.900 45.600 ;
        RECT 107.100 42.000 108.900 51.600 ;
        RECT 113.700 51.000 117.000 52.200 ;
        RECT 134.100 51.600 135.300 55.950 ;
        RECT 137.100 54.150 138.900 55.950 ;
        RECT 113.700 42.600 115.500 51.000 ;
        RECT 131.700 50.700 135.300 51.600 ;
        RECT 131.700 48.600 132.900 50.700 ;
        RECT 131.100 42.600 132.900 48.600 ;
        RECT 134.100 47.700 141.900 49.050 ;
        RECT 134.100 42.600 135.900 47.700 ;
        RECT 137.100 42.000 138.900 46.800 ;
        RECT 140.100 42.600 141.900 47.700 ;
        RECT 158.700 45.600 159.900 55.950 ;
        RECT 179.100 54.150 180.900 55.950 ;
        RECT 185.100 54.150 186.900 55.950 ;
        RECT 188.100 52.200 189.000 55.950 ;
        RECT 203.100 54.150 204.900 55.950 ;
        RECT 209.100 54.150 210.900 55.950 ;
        RECT 212.100 52.200 213.000 55.950 ;
        RECT 227.250 54.150 229.050 55.950 ;
        RECT 158.100 42.600 159.900 45.600 ;
        RECT 161.100 42.000 162.900 45.600 ;
        RECT 179.100 42.000 180.900 51.600 ;
        RECT 185.700 51.000 189.000 52.200 ;
        RECT 185.700 42.600 187.500 51.000 ;
        RECT 203.100 42.000 204.900 51.600 ;
        RECT 209.700 51.000 213.000 52.200 ;
        RECT 209.700 42.600 211.500 51.000 ;
        RECT 233.100 48.600 234.300 55.950 ;
        RECT 239.100 54.150 240.900 55.950 ;
        RECT 254.100 54.150 255.900 55.950 ;
        RECT 260.100 54.150 261.900 55.950 ;
        RECT 263.100 52.200 264.000 55.950 ;
        RECT 281.100 54.150 282.900 55.950 ;
        RECT 287.100 54.150 288.900 55.950 ;
        RECT 290.100 52.200 291.000 55.950 ;
        RECT 305.100 54.150 306.900 55.950 ;
        RECT 311.100 54.150 312.900 55.950 ;
        RECT 314.100 52.200 315.000 55.950 ;
        RECT 332.100 54.150 333.900 55.950 ;
        RECT 338.250 54.150 340.050 55.950 ;
        RECT 227.700 42.000 229.500 48.600 ;
        RECT 232.200 42.600 234.000 48.600 ;
        RECT 236.700 42.000 238.500 48.600 ;
        RECT 254.100 42.000 255.900 51.600 ;
        RECT 260.700 51.000 264.000 52.200 ;
        RECT 260.700 42.600 262.500 51.000 ;
        RECT 281.100 42.000 282.900 51.600 ;
        RECT 287.700 51.000 291.000 52.200 ;
        RECT 287.700 42.600 289.500 51.000 ;
        RECT 305.100 42.000 306.900 51.600 ;
        RECT 311.700 51.000 315.000 52.200 ;
        RECT 311.700 42.600 313.500 51.000 ;
        RECT 341.700 48.600 342.600 55.950 ;
        RECT 359.100 54.150 360.900 55.950 ;
        RECT 365.100 54.150 366.900 55.950 ;
        RECT 368.100 52.200 369.000 55.950 ;
        RECT 386.100 54.150 387.900 55.950 ;
        RECT 392.250 54.150 394.050 55.950 ;
        RECT 333.000 42.000 334.800 48.600 ;
        RECT 337.500 47.400 342.600 48.600 ;
        RECT 337.500 42.600 339.300 47.400 ;
        RECT 340.500 42.000 342.300 45.600 ;
        RECT 359.100 42.000 360.900 51.600 ;
        RECT 365.700 51.000 369.000 52.200 ;
        RECT 365.700 42.600 367.500 51.000 ;
        RECT 395.700 48.600 396.600 55.950 ;
        RECT 413.100 54.150 414.900 55.950 ;
        RECT 416.700 51.600 417.900 55.950 ;
        RECT 419.100 54.150 420.900 55.950 ;
        RECT 425.550 55.050 426.450 59.550 ;
        RECT 430.950 58.950 433.050 59.550 ;
        RECT 434.100 58.050 435.900 59.850 ;
        RECT 440.700 58.050 441.900 65.400 ;
        RECT 459.000 58.050 459.900 70.200 ;
        RECT 464.100 58.050 465.900 59.850 ;
        RECT 488.100 58.050 489.300 71.400 ;
        RECT 433.950 55.950 436.050 58.050 ;
        RECT 436.950 55.950 439.050 58.050 ;
        RECT 439.950 55.950 442.050 58.050 ;
        RECT 442.950 55.950 445.050 58.050 ;
        RECT 457.950 55.950 460.050 58.050 ;
        RECT 460.950 55.950 463.050 58.050 ;
        RECT 463.950 55.950 466.050 58.050 ;
        RECT 466.950 55.950 469.050 58.050 ;
        RECT 484.950 55.950 487.050 58.050 ;
        RECT 487.950 55.950 490.050 58.050 ;
        RECT 490.950 55.950 493.050 58.050 ;
        RECT 509.100 55.950 511.200 58.050 ;
        RECT 421.950 53.550 426.450 55.050 ;
        RECT 437.100 54.150 438.900 55.950 ;
        RECT 421.950 52.950 426.000 53.550 ;
        RECT 440.700 51.600 441.900 55.950 ;
        RECT 443.100 54.150 444.900 55.950 ;
        RECT 459.000 52.200 459.900 55.950 ;
        RECT 461.100 54.150 462.900 55.950 ;
        RECT 467.100 54.150 468.900 55.950 ;
        RECT 485.250 54.150 487.050 55.950 ;
        RECT 416.700 50.700 420.300 51.600 ;
        RECT 440.700 50.700 444.300 51.600 ;
        RECT 459.000 51.000 462.300 52.200 ;
        RECT 387.000 42.000 388.800 48.600 ;
        RECT 391.500 47.400 396.600 48.600 ;
        RECT 410.100 47.700 417.900 49.050 ;
        RECT 391.500 42.600 393.300 47.400 ;
        RECT 394.500 42.000 396.300 45.600 ;
        RECT 410.100 42.600 411.900 47.700 ;
        RECT 413.100 42.000 414.900 46.800 ;
        RECT 416.100 42.600 417.900 47.700 ;
        RECT 419.100 48.600 420.300 50.700 ;
        RECT 419.100 42.600 420.900 48.600 ;
        RECT 434.100 47.700 441.900 49.050 ;
        RECT 434.100 42.600 435.900 47.700 ;
        RECT 437.100 42.000 438.900 46.800 ;
        RECT 440.100 42.600 441.900 47.700 ;
        RECT 443.100 48.600 444.300 50.700 ;
        RECT 443.100 42.600 444.900 48.600 ;
        RECT 460.500 42.600 462.300 51.000 ;
        RECT 467.100 42.000 468.900 51.600 ;
        RECT 488.100 50.700 489.300 55.950 ;
        RECT 491.100 54.150 492.900 55.950 ;
        RECT 509.250 54.150 511.050 55.950 ;
        RECT 512.100 51.300 513.000 71.400 ;
        RECT 515.100 66.000 516.900 78.000 ;
        RECT 518.100 65.400 519.900 77.400 ;
        RECT 533.100 66.600 534.900 77.400 ;
        RECT 536.100 67.500 537.900 78.000 ;
        RECT 539.100 76.500 546.900 77.400 ;
        RECT 539.100 66.600 540.900 76.500 ;
        RECT 533.100 65.700 540.900 66.600 ;
        RECT 514.200 58.050 516.000 59.850 ;
        RECT 518.400 58.050 519.300 65.400 ;
        RECT 542.100 64.500 543.900 75.600 ;
        RECT 545.100 65.400 546.900 76.500 ;
        RECT 560.100 65.400 561.900 77.400 ;
        RECT 563.100 66.000 564.900 78.000 ;
        RECT 566.100 71.400 567.900 77.400 ;
        RECT 569.100 71.400 570.900 78.000 ;
        RECT 587.100 71.400 588.900 78.000 ;
        RECT 590.100 71.400 591.900 77.400 ;
        RECT 593.100 71.400 594.900 78.000 ;
        RECT 608.100 71.400 609.900 78.000 ;
        RECT 611.100 71.400 612.900 77.400 ;
        RECT 614.100 72.000 615.900 78.000 ;
        RECT 539.100 63.600 543.900 64.500 ;
        RECT 536.250 58.050 538.050 59.850 ;
        RECT 539.100 58.050 540.000 63.600 ;
        RECT 542.100 58.050 543.900 59.850 ;
        RECT 560.700 58.050 561.600 65.400 ;
        RECT 564.000 58.050 565.800 59.850 ;
        RECT 514.500 55.950 516.600 58.050 ;
        RECT 517.800 55.950 519.900 58.050 ;
        RECT 532.950 55.950 535.050 58.050 ;
        RECT 535.950 55.950 538.050 58.050 ;
        RECT 538.950 55.950 541.050 58.050 ;
        RECT 541.950 55.950 544.050 58.050 ;
        RECT 544.950 55.950 547.050 58.050 ;
        RECT 560.100 55.950 562.200 58.050 ;
        RECT 563.400 55.950 565.500 58.050 ;
        RECT 488.100 49.800 492.300 50.700 ;
        RECT 485.400 42.000 487.200 48.600 ;
        RECT 490.500 42.600 492.300 49.800 ;
        RECT 509.100 50.400 517.500 51.300 ;
        RECT 509.100 42.600 510.900 50.400 ;
        RECT 515.700 49.500 517.500 50.400 ;
        RECT 518.400 48.600 519.300 55.950 ;
        RECT 533.250 54.150 535.050 55.950 ;
        RECT 539.100 48.600 540.300 55.950 ;
        RECT 545.100 54.150 546.900 55.950 ;
        RECT 541.950 51.450 544.050 51.750 ;
        RECT 556.950 51.450 559.050 52.050 ;
        RECT 541.950 50.550 559.050 51.450 ;
        RECT 541.950 49.650 544.050 50.550 ;
        RECT 556.950 49.950 559.050 50.550 ;
        RECT 560.700 48.600 561.600 55.950 ;
        RECT 567.000 51.300 567.900 71.400 ;
        RECT 590.700 58.050 591.900 71.400 ;
        RECT 611.400 71.100 612.900 71.400 ;
        RECT 617.100 71.400 618.900 77.400 ;
        RECT 617.100 71.100 618.000 71.400 ;
        RECT 611.400 70.200 618.000 71.100 ;
        RECT 611.100 58.050 612.900 59.850 ;
        RECT 617.100 58.050 618.000 70.200 ;
        RECT 632.100 65.400 633.900 77.400 ;
        RECT 635.100 66.300 636.900 77.400 ;
        RECT 638.100 67.200 639.900 78.000 ;
        RECT 641.100 66.300 642.900 77.400 ;
        RECT 656.100 71.400 657.900 78.000 ;
        RECT 659.100 71.400 660.900 77.400 ;
        RECT 662.100 72.000 663.900 78.000 ;
        RECT 659.400 71.100 660.900 71.400 ;
        RECT 665.100 71.400 666.900 77.400 ;
        RECT 680.100 71.400 681.900 78.000 ;
        RECT 683.100 71.400 684.900 77.400 ;
        RECT 686.100 72.000 687.900 78.000 ;
        RECT 665.100 71.100 666.000 71.400 ;
        RECT 659.400 70.200 666.000 71.100 ;
        RECT 683.400 71.100 684.900 71.400 ;
        RECT 689.100 71.400 690.900 77.400 ;
        RECT 704.100 71.400 705.900 77.400 ;
        RECT 707.100 72.000 708.900 78.000 ;
        RECT 689.100 71.100 690.000 71.400 ;
        RECT 683.400 70.200 690.000 71.100 ;
        RECT 635.100 65.400 642.900 66.300 ;
        RECT 649.950 66.450 652.050 67.050 ;
        RECT 658.950 66.450 661.050 67.050 ;
        RECT 649.950 65.550 661.050 66.450 ;
        RECT 632.400 58.050 633.300 65.400 ;
        RECT 649.950 64.950 652.050 65.550 ;
        RECT 658.950 64.950 661.050 65.550 ;
        RECT 640.950 63.450 643.050 64.050 ;
        RECT 661.950 63.450 664.050 63.900 ;
        RECT 640.950 62.550 664.050 63.450 ;
        RECT 640.950 61.950 643.050 62.550 ;
        RECT 661.950 61.800 664.050 62.550 ;
        RECT 637.950 58.050 639.750 59.850 ;
        RECT 659.100 58.050 660.900 59.850 ;
        RECT 665.100 58.050 666.000 70.200 ;
        RECT 670.950 63.450 673.050 64.050 ;
        RECT 685.950 63.450 688.050 64.050 ;
        RECT 670.950 62.550 688.050 63.450 ;
        RECT 670.950 61.950 673.050 62.550 ;
        RECT 685.950 61.950 688.050 62.550 ;
        RECT 683.100 58.050 684.900 59.850 ;
        RECT 689.100 58.050 690.000 70.200 ;
        RECT 705.000 71.100 705.900 71.400 ;
        RECT 710.100 71.400 711.900 77.400 ;
        RECT 713.100 71.400 714.900 78.000 ;
        RECT 710.100 71.100 711.600 71.400 ;
        RECT 705.000 70.200 711.600 71.100 ;
        RECT 705.000 58.050 705.900 70.200 ;
        RECT 728.100 66.300 729.900 77.400 ;
        RECT 731.100 67.500 732.900 78.000 ;
        RECT 728.100 65.400 732.600 66.300 ;
        RECT 735.600 65.400 737.400 77.400 ;
        RECT 740.100 67.500 741.900 78.000 ;
        RECT 743.100 66.600 744.900 77.400 ;
        RECT 758.100 71.400 759.900 77.400 ;
        RECT 761.100 71.400 762.900 78.000 ;
        RECT 776.100 71.400 777.900 78.000 ;
        RECT 779.100 71.400 780.900 77.400 ;
        RECT 782.100 71.400 783.900 78.000 ;
        RECT 800.700 71.400 802.500 78.000 ;
        RECT 730.500 63.300 732.600 65.400 ;
        RECT 736.200 64.050 737.400 65.400 ;
        RECT 740.100 65.400 744.900 66.600 ;
        RECT 740.100 64.500 742.200 65.400 ;
        RECT 736.200 63.000 737.700 64.050 ;
        RECT 733.800 61.500 735.900 61.800 ;
        RECT 710.100 58.050 711.900 59.850 ;
        RECT 732.000 59.700 735.900 61.500 ;
        RECT 736.800 61.050 737.700 63.000 ;
        RECT 736.800 58.950 738.900 61.050 ;
        RECT 745.950 60.450 748.050 61.050 ;
        RECT 754.950 60.450 757.050 61.050 ;
        RECT 736.800 58.800 738.300 58.950 ;
        RECT 733.200 58.050 735.000 58.500 ;
        RECT 568.800 55.950 570.900 58.050 ;
        RECT 586.950 55.950 589.050 58.050 ;
        RECT 589.950 55.950 592.050 58.050 ;
        RECT 592.950 55.950 595.050 58.050 ;
        RECT 607.950 55.950 610.050 58.050 ;
        RECT 610.950 55.950 613.050 58.050 ;
        RECT 613.950 55.950 616.050 58.050 ;
        RECT 616.950 55.950 619.050 58.050 ;
        RECT 631.950 55.950 634.050 58.050 ;
        RECT 634.950 55.950 637.050 58.050 ;
        RECT 637.950 55.950 640.050 58.050 ;
        RECT 640.950 55.950 643.050 58.050 ;
        RECT 655.950 55.950 658.050 58.050 ;
        RECT 658.950 55.950 661.050 58.050 ;
        RECT 661.950 55.950 664.050 58.050 ;
        RECT 664.950 55.950 667.050 58.050 ;
        RECT 679.950 55.950 682.050 58.050 ;
        RECT 682.950 55.950 685.050 58.050 ;
        RECT 685.950 55.950 688.050 58.050 ;
        RECT 688.950 55.950 691.050 58.050 ;
        RECT 703.950 55.950 706.050 58.050 ;
        RECT 706.950 55.950 709.050 58.050 ;
        RECT 709.950 55.950 712.050 58.050 ;
        RECT 712.950 55.950 715.050 58.050 ;
        RECT 728.100 56.700 735.000 58.050 ;
        RECT 735.900 57.900 738.300 58.800 ;
        RECT 742.800 58.050 744.600 59.850 ;
        RECT 745.950 59.550 757.050 60.450 ;
        RECT 745.950 58.950 748.050 59.550 ;
        RECT 754.950 58.950 757.050 59.550 ;
        RECT 758.700 58.050 759.900 71.400 ;
        RECT 761.100 58.050 762.900 59.850 ;
        RECT 779.700 58.050 780.900 71.400 ;
        RECT 801.000 68.100 802.800 69.900 ;
        RECT 803.700 66.900 805.500 77.400 ;
        RECT 803.100 65.400 805.500 66.900 ;
        RECT 808.800 65.400 810.600 78.000 ;
        RECT 824.100 71.400 825.900 78.000 ;
        RECT 827.100 71.400 828.900 77.400 ;
        RECT 803.100 58.050 804.300 65.400 ;
        RECT 805.950 63.450 808.050 64.050 ;
        RECT 805.950 62.550 816.450 63.450 ;
        RECT 805.950 61.950 808.050 62.550 ;
        RECT 809.100 58.050 810.900 59.850 ;
        RECT 728.100 55.950 730.200 56.700 ;
        RECT 568.950 54.150 570.750 55.950 ;
        RECT 587.100 54.150 588.900 55.950 ;
        RECT 562.500 50.400 570.900 51.300 ;
        RECT 590.700 50.700 591.900 55.950 ;
        RECT 592.950 54.150 594.750 55.950 ;
        RECT 608.100 54.150 609.900 55.950 ;
        RECT 614.100 54.150 615.900 55.950 ;
        RECT 617.100 52.200 618.000 55.950 ;
        RECT 562.500 49.500 564.300 50.400 ;
        RECT 513.600 42.000 515.400 48.600 ;
        RECT 516.600 46.800 519.300 48.600 ;
        RECT 516.600 42.600 518.400 46.800 ;
        RECT 533.700 42.000 535.500 48.600 ;
        RECT 538.200 42.600 540.000 48.600 ;
        RECT 542.700 42.000 544.500 48.600 ;
        RECT 560.700 46.800 563.400 48.600 ;
        RECT 561.600 42.600 563.400 46.800 ;
        RECT 564.600 42.000 566.400 48.600 ;
        RECT 569.100 42.600 570.900 50.400 ;
        RECT 587.700 49.800 591.900 50.700 ;
        RECT 587.700 42.600 589.500 49.800 ;
        RECT 592.800 42.000 594.600 48.600 ;
        RECT 608.100 42.000 609.900 51.600 ;
        RECT 614.700 51.000 618.000 52.200 ;
        RECT 614.700 42.600 616.500 51.000 ;
        RECT 632.400 48.600 633.300 55.950 ;
        RECT 634.950 54.150 636.750 55.950 ;
        RECT 641.100 54.150 642.900 55.950 ;
        RECT 656.100 54.150 657.900 55.950 ;
        RECT 662.100 54.150 663.900 55.950 ;
        RECT 665.100 52.200 666.000 55.950 ;
        RECT 680.100 54.150 681.900 55.950 ;
        RECT 686.100 54.150 687.900 55.950 ;
        RECT 689.100 52.200 690.000 55.950 ;
        RECT 637.950 51.450 640.050 52.050 ;
        RECT 646.950 51.450 649.050 52.050 ;
        RECT 652.950 51.450 655.050 52.050 ;
        RECT 637.950 50.550 655.050 51.450 ;
        RECT 637.950 49.950 640.050 50.550 ;
        RECT 646.950 49.950 649.050 50.550 ;
        RECT 652.950 49.950 655.050 50.550 ;
        RECT 632.400 47.400 637.500 48.600 ;
        RECT 632.700 42.000 634.500 45.600 ;
        RECT 635.700 42.600 637.500 47.400 ;
        RECT 640.200 42.000 642.000 48.600 ;
        RECT 656.100 42.000 657.900 51.600 ;
        RECT 662.700 51.000 666.000 52.200 ;
        RECT 662.700 42.600 664.500 51.000 ;
        RECT 680.100 42.000 681.900 51.600 ;
        RECT 686.700 51.000 690.000 52.200 ;
        RECT 705.000 52.200 705.900 55.950 ;
        RECT 707.100 54.150 708.900 55.950 ;
        RECT 713.100 54.150 714.900 55.950 ;
        RECT 728.400 54.150 730.200 55.950 ;
        RECT 733.200 53.400 735.000 55.200 ;
        RECT 705.000 51.000 708.300 52.200 ;
        RECT 686.700 42.600 688.500 51.000 ;
        RECT 706.500 42.600 708.300 51.000 ;
        RECT 713.100 42.000 714.900 51.600 ;
        RECT 732.900 51.300 735.000 53.400 ;
        RECT 728.700 50.400 735.000 51.300 ;
        RECT 735.900 52.200 737.100 57.900 ;
        RECT 738.300 55.200 740.100 57.000 ;
        RECT 742.800 55.950 744.900 58.050 ;
        RECT 757.950 55.950 760.050 58.050 ;
        RECT 760.950 55.950 763.050 58.050 ;
        RECT 775.950 55.950 778.050 58.050 ;
        RECT 778.950 55.950 781.050 58.050 ;
        RECT 781.950 55.950 784.050 58.050 ;
        RECT 799.950 55.950 802.050 58.050 ;
        RECT 802.950 55.950 805.050 58.050 ;
        RECT 805.950 55.950 808.050 58.050 ;
        RECT 808.950 55.950 811.050 58.050 ;
        RECT 738.000 53.100 740.100 55.200 ;
        RECT 728.700 48.600 729.900 50.400 ;
        RECT 735.900 50.100 738.900 52.200 ;
        RECT 735.900 48.600 737.100 50.100 ;
        RECT 740.100 49.500 742.200 50.700 ;
        RECT 740.100 48.600 744.900 49.500 ;
        RECT 728.100 42.600 729.900 48.600 ;
        RECT 731.100 42.000 732.900 47.700 ;
        RECT 735.600 42.600 737.400 48.600 ;
        RECT 740.100 42.000 741.900 47.700 ;
        RECT 743.100 42.600 744.900 48.600 ;
        RECT 758.700 45.600 759.900 55.950 ;
        RECT 776.100 54.150 777.900 55.950 ;
        RECT 779.700 50.700 780.900 55.950 ;
        RECT 781.950 54.150 783.750 55.950 ;
        RECT 800.100 54.150 801.900 55.950 ;
        RECT 803.100 51.600 804.300 55.950 ;
        RECT 806.100 54.150 807.900 55.950 ;
        RECT 815.550 55.050 816.450 62.550 ;
        RECT 824.100 58.050 825.900 59.850 ;
        RECT 827.100 58.050 828.300 71.400 ;
        RECT 842.100 65.400 843.900 77.400 ;
        RECT 845.100 66.300 846.900 77.400 ;
        RECT 848.100 67.200 849.900 78.000 ;
        RECT 851.100 66.300 852.900 77.400 ;
        RECT 845.100 65.400 852.900 66.300 ;
        RECT 869.100 65.400 870.900 77.400 ;
        RECT 872.100 66.300 873.900 77.400 ;
        RECT 875.100 67.200 876.900 78.000 ;
        RECT 878.100 66.300 879.900 77.400 ;
        RECT 893.100 71.400 894.900 77.400 ;
        RECT 896.100 72.000 897.900 78.000 ;
        RECT 872.100 65.400 879.900 66.300 ;
        RECT 894.000 71.100 894.900 71.400 ;
        RECT 899.100 71.400 900.900 77.400 ;
        RECT 902.100 71.400 903.900 78.000 ;
        RECT 899.100 71.100 900.600 71.400 ;
        RECT 894.000 70.200 900.600 71.100 ;
        RECT 842.400 58.050 843.300 65.400 ;
        RECT 847.950 58.050 849.750 59.850 ;
        RECT 869.400 58.050 870.300 65.400 ;
        RECT 874.950 58.050 876.750 59.850 ;
        RECT 894.000 58.050 894.900 70.200 ;
        RECT 917.100 65.400 918.900 77.400 ;
        RECT 920.100 66.300 921.900 77.400 ;
        RECT 923.100 67.200 924.900 78.000 ;
        RECT 926.100 66.300 927.900 77.400 ;
        RECT 941.100 71.400 942.900 78.000 ;
        RECT 944.100 71.400 945.900 77.400 ;
        RECT 947.100 72.000 948.900 78.000 ;
        RECT 944.400 71.100 945.900 71.400 ;
        RECT 950.100 71.400 951.900 77.400 ;
        RECT 965.700 71.400 967.500 78.000 ;
        RECT 950.100 71.100 951.000 71.400 ;
        RECT 944.400 70.200 951.000 71.100 ;
        RECT 920.100 65.400 927.900 66.300 ;
        RECT 899.100 58.050 900.900 59.850 ;
        RECT 917.400 58.050 918.300 65.400 ;
        RECT 922.950 58.050 924.750 59.850 ;
        RECT 944.100 58.050 945.900 59.850 ;
        RECT 950.100 58.050 951.000 70.200 ;
        RECT 966.000 68.100 967.800 69.900 ;
        RECT 968.700 66.900 970.500 77.400 ;
        RECT 968.100 65.400 970.500 66.900 ;
        RECT 973.800 65.400 975.600 78.000 ;
        RECT 989.100 65.400 990.900 77.400 ;
        RECT 992.100 66.300 993.900 77.400 ;
        RECT 995.100 67.200 996.900 78.000 ;
        RECT 998.100 66.300 999.900 77.400 ;
        RECT 992.100 65.400 999.900 66.300 ;
        RECT 968.100 58.050 969.300 65.400 ;
        RECT 970.950 63.450 973.050 64.050 ;
        RECT 970.950 62.550 978.450 63.450 ;
        RECT 970.950 61.950 973.050 62.550 ;
        RECT 977.550 60.450 978.450 62.550 ;
        RECT 974.100 58.050 975.900 59.850 ;
        RECT 977.550 59.550 981.450 60.450 ;
        RECT 823.950 55.950 826.050 58.050 ;
        RECT 826.950 55.950 829.050 58.050 ;
        RECT 841.950 55.950 844.050 58.050 ;
        RECT 844.950 55.950 847.050 58.050 ;
        RECT 847.950 55.950 850.050 58.050 ;
        RECT 850.950 55.950 853.050 58.050 ;
        RECT 868.950 55.950 871.050 58.050 ;
        RECT 871.950 55.950 874.050 58.050 ;
        RECT 874.950 55.950 877.050 58.050 ;
        RECT 877.950 55.950 880.050 58.050 ;
        RECT 892.950 55.950 895.050 58.050 ;
        RECT 895.950 55.950 898.050 58.050 ;
        RECT 898.950 55.950 901.050 58.050 ;
        RECT 901.950 55.950 904.050 58.050 ;
        RECT 916.950 55.950 919.050 58.050 ;
        RECT 919.950 55.950 922.050 58.050 ;
        RECT 922.950 55.950 925.050 58.050 ;
        RECT 925.950 55.950 928.050 58.050 ;
        RECT 940.950 55.950 943.050 58.050 ;
        RECT 943.950 55.950 946.050 58.050 ;
        RECT 946.950 55.950 949.050 58.050 ;
        RECT 949.950 55.950 952.050 58.050 ;
        RECT 964.950 55.950 967.050 58.050 ;
        RECT 967.950 55.950 970.050 58.050 ;
        RECT 970.950 55.950 973.050 58.050 ;
        RECT 973.950 55.950 976.050 58.050 ;
        RECT 811.950 53.550 816.450 55.050 ;
        RECT 811.950 52.950 816.000 53.550 ;
        RECT 776.700 49.800 780.900 50.700 ;
        RECT 800.700 50.700 804.300 51.600 ;
        RECT 758.100 42.600 759.900 45.600 ;
        RECT 761.100 42.000 762.900 45.600 ;
        RECT 776.700 42.600 778.500 49.800 ;
        RECT 800.700 48.600 801.900 50.700 ;
        RECT 781.800 42.000 783.600 48.600 ;
        RECT 800.100 42.600 801.900 48.600 ;
        RECT 803.100 47.700 810.900 49.050 ;
        RECT 803.100 42.600 804.900 47.700 ;
        RECT 806.100 42.000 807.900 46.800 ;
        RECT 809.100 42.600 810.900 47.700 ;
        RECT 827.100 45.600 828.300 55.950 ;
        RECT 842.400 48.600 843.300 55.950 ;
        RECT 844.950 54.150 846.750 55.950 ;
        RECT 851.100 54.150 852.900 55.950 ;
        RECT 844.950 51.450 847.050 52.050 ;
        RECT 856.950 51.450 859.050 52.050 ;
        RECT 844.950 50.550 859.050 51.450 ;
        RECT 844.950 49.950 847.050 50.550 ;
        RECT 856.950 49.950 859.050 50.550 ;
        RECT 869.400 48.600 870.300 55.950 ;
        RECT 871.950 54.150 873.750 55.950 ;
        RECT 878.100 54.150 879.900 55.950 ;
        RECT 894.000 52.200 894.900 55.950 ;
        RECT 896.100 54.150 897.900 55.950 ;
        RECT 902.100 54.150 903.900 55.950 ;
        RECT 894.000 51.000 897.300 52.200 ;
        RECT 842.400 47.400 847.500 48.600 ;
        RECT 824.100 42.000 825.900 45.600 ;
        RECT 827.100 42.600 828.900 45.600 ;
        RECT 842.700 42.000 844.500 45.600 ;
        RECT 845.700 42.600 847.500 47.400 ;
        RECT 850.200 42.000 852.000 48.600 ;
        RECT 869.400 47.400 874.500 48.600 ;
        RECT 869.700 42.000 871.500 45.600 ;
        RECT 872.700 42.600 874.500 47.400 ;
        RECT 877.200 42.000 879.000 48.600 ;
        RECT 895.500 42.600 897.300 51.000 ;
        RECT 902.100 42.000 903.900 51.600 ;
        RECT 917.400 48.600 918.300 55.950 ;
        RECT 919.950 54.150 921.750 55.950 ;
        RECT 926.100 54.150 927.900 55.950 ;
        RECT 941.100 54.150 942.900 55.950 ;
        RECT 947.100 54.150 948.900 55.950 ;
        RECT 950.100 52.200 951.000 55.950 ;
        RECT 965.100 54.150 966.900 55.950 ;
        RECT 917.400 47.400 922.500 48.600 ;
        RECT 917.700 42.000 919.500 45.600 ;
        RECT 920.700 42.600 922.500 47.400 ;
        RECT 925.200 42.000 927.000 48.600 ;
        RECT 941.100 42.000 942.900 51.600 ;
        RECT 947.700 51.000 951.000 52.200 ;
        RECT 968.100 51.600 969.300 55.950 ;
        RECT 971.100 54.150 972.900 55.950 ;
        RECT 980.550 54.450 981.450 59.550 ;
        RECT 989.400 58.050 990.300 65.400 ;
        RECT 994.950 58.050 996.750 59.850 ;
        RECT 988.950 55.950 991.050 58.050 ;
        RECT 991.950 55.950 994.050 58.050 ;
        RECT 994.950 55.950 997.050 58.050 ;
        RECT 997.950 55.950 1000.050 58.050 ;
        RECT 985.950 54.450 988.050 55.050 ;
        RECT 980.550 53.550 988.050 54.450 ;
        RECT 985.950 52.950 988.050 53.550 ;
        RECT 947.700 42.600 949.500 51.000 ;
        RECT 965.700 50.700 969.300 51.600 ;
        RECT 965.700 48.600 966.900 50.700 ;
        RECT 965.100 42.600 966.900 48.600 ;
        RECT 968.100 47.700 975.900 49.050 ;
        RECT 968.100 42.600 969.900 47.700 ;
        RECT 971.100 42.000 972.900 46.800 ;
        RECT 974.100 42.600 975.900 47.700 ;
        RECT 989.400 48.600 990.300 55.950 ;
        RECT 991.950 54.150 993.750 55.950 ;
        RECT 998.100 54.150 999.900 55.950 ;
        RECT 989.400 47.400 994.500 48.600 ;
        RECT 989.700 42.000 991.500 45.600 ;
        RECT 992.700 42.600 994.500 47.400 ;
        RECT 997.200 42.000 999.000 48.600 ;
        RECT 14.100 35.400 15.900 38.400 ;
        RECT 17.100 35.400 18.900 39.000 ;
        RECT 32.100 35.400 33.900 39.000 ;
        RECT 35.100 35.400 36.900 38.400 ;
        RECT 14.700 25.050 15.900 35.400 ;
        RECT 35.100 25.050 36.300 35.400 ;
        RECT 53.100 32.400 54.900 38.400 ;
        RECT 53.700 30.300 54.900 32.400 ;
        RECT 56.100 33.300 57.900 38.400 ;
        RECT 59.100 34.200 60.900 39.000 ;
        RECT 62.100 33.300 63.900 38.400 ;
        RECT 56.100 31.950 63.900 33.300 ;
        RECT 80.100 33.300 81.900 38.400 ;
        RECT 83.100 34.200 84.900 39.000 ;
        RECT 86.100 33.300 87.900 38.400 ;
        RECT 80.100 31.950 87.900 33.300 ;
        RECT 89.100 32.400 90.900 38.400 ;
        RECT 94.950 36.450 97.050 37.050 ;
        RECT 94.950 36.000 102.450 36.450 ;
        RECT 94.950 35.550 103.050 36.000 ;
        RECT 94.950 34.950 97.050 35.550 ;
        RECT 89.100 30.300 90.300 32.400 ;
        RECT 100.950 31.950 103.050 35.550 ;
        RECT 53.700 29.400 57.300 30.300 ;
        RECT 53.100 25.050 54.900 26.850 ;
        RECT 56.100 25.050 57.300 29.400 ;
        RECT 86.700 29.400 90.300 30.300 ;
        RECT 104.100 29.400 105.900 39.000 ;
        RECT 110.700 30.000 112.500 38.400 ;
        RECT 59.100 25.050 60.900 26.850 ;
        RECT 83.100 25.050 84.900 26.850 ;
        RECT 86.700 25.050 87.900 29.400 ;
        RECT 110.700 28.800 114.000 30.000 ;
        RECT 128.100 29.400 129.900 39.000 ;
        RECT 134.700 30.000 136.500 38.400 ;
        RECT 153.000 32.400 154.800 39.000 ;
        RECT 157.500 33.600 159.300 38.400 ;
        RECT 160.500 35.400 162.300 39.000 ;
        RECT 176.100 35.400 177.900 39.000 ;
        RECT 179.100 35.400 180.900 38.400 ;
        RECT 157.500 32.400 162.600 33.600 ;
        RECT 134.700 28.800 138.000 30.000 ;
        RECT 89.100 25.050 90.900 26.850 ;
        RECT 104.100 25.050 105.900 26.850 ;
        RECT 110.100 25.050 111.900 26.850 ;
        RECT 113.100 25.050 114.000 28.800 ;
        RECT 128.100 25.050 129.900 26.850 ;
        RECT 134.100 25.050 135.900 26.850 ;
        RECT 137.100 25.050 138.000 28.800 ;
        RECT 152.100 25.050 153.900 26.850 ;
        RECT 158.250 25.050 160.050 26.850 ;
        RECT 161.700 25.050 162.600 32.400 ;
        RECT 179.100 25.050 180.300 35.400 ;
        RECT 195.000 32.400 196.800 39.000 ;
        RECT 199.500 33.600 201.300 38.400 ;
        RECT 202.500 35.400 204.300 39.000 ;
        RECT 199.500 32.400 204.600 33.600 ;
        RECT 194.100 25.050 195.900 26.850 ;
        RECT 200.250 25.050 202.050 26.850 ;
        RECT 203.700 25.050 204.600 32.400 ;
        RECT 218.100 29.400 219.900 39.000 ;
        RECT 224.700 30.000 226.500 38.400 ;
        RECT 245.100 33.300 246.900 38.400 ;
        RECT 248.100 34.200 249.900 39.000 ;
        RECT 251.100 33.300 252.900 38.400 ;
        RECT 245.100 31.950 252.900 33.300 ;
        RECT 254.100 32.400 255.900 38.400 ;
        RECT 254.100 30.300 255.300 32.400 ;
        RECT 224.700 28.800 228.000 30.000 ;
        RECT 218.100 25.050 219.900 26.850 ;
        RECT 224.100 25.050 225.900 26.850 ;
        RECT 227.100 25.050 228.000 28.800 ;
        RECT 251.700 29.400 255.300 30.300 ;
        RECT 271.500 30.000 273.300 38.400 ;
        RECT 248.100 25.050 249.900 26.850 ;
        RECT 251.700 25.050 252.900 29.400 ;
        RECT 270.000 28.800 273.300 30.000 ;
        RECT 278.100 29.400 279.900 39.000 ;
        RECT 293.100 32.400 294.900 38.400 ;
        RECT 293.700 30.300 294.900 32.400 ;
        RECT 296.100 33.300 297.900 38.400 ;
        RECT 299.100 34.200 300.900 39.000 ;
        RECT 302.100 33.300 303.900 38.400 ;
        RECT 296.100 31.950 303.900 33.300 ;
        RECT 317.100 33.300 318.900 38.400 ;
        RECT 320.100 34.200 321.900 39.000 ;
        RECT 323.100 33.300 324.900 38.400 ;
        RECT 317.100 31.950 324.900 33.300 ;
        RECT 326.100 32.400 327.900 38.400 ;
        RECT 345.000 32.400 346.800 39.000 ;
        RECT 349.500 33.600 351.300 38.400 ;
        RECT 352.500 35.400 354.300 39.000 ;
        RECT 368.100 35.400 369.900 38.400 ;
        RECT 349.500 32.400 354.600 33.600 ;
        RECT 326.100 30.300 327.300 32.400 ;
        RECT 293.700 29.400 297.300 30.300 ;
        RECT 254.100 25.050 255.900 26.850 ;
        RECT 270.000 25.050 270.900 28.800 ;
        RECT 272.100 25.050 273.900 26.850 ;
        RECT 278.100 25.050 279.900 26.850 ;
        RECT 293.100 25.050 294.900 26.850 ;
        RECT 296.100 25.050 297.300 29.400 ;
        RECT 323.700 29.400 327.300 30.300 ;
        RECT 299.100 25.050 300.900 26.850 ;
        RECT 320.100 25.050 321.900 26.850 ;
        RECT 323.700 25.050 324.900 29.400 ;
        RECT 326.100 25.050 327.900 26.850 ;
        RECT 344.100 25.050 345.900 26.850 ;
        RECT 350.250 25.050 352.050 26.850 ;
        RECT 353.700 25.050 354.600 32.400 ;
        RECT 368.100 31.500 369.300 35.400 ;
        RECT 371.100 32.400 372.900 39.000 ;
        RECT 374.100 32.400 375.900 38.400 ;
        RECT 368.100 30.600 373.800 31.500 ;
        RECT 372.000 29.700 373.800 30.600 ;
        RECT 13.950 22.950 16.050 25.050 ;
        RECT 16.950 22.950 19.050 25.050 ;
        RECT 31.950 22.950 34.050 25.050 ;
        RECT 34.950 22.950 37.050 25.050 ;
        RECT 52.950 22.950 55.050 25.050 ;
        RECT 55.950 22.950 58.050 25.050 ;
        RECT 58.950 22.950 61.050 25.050 ;
        RECT 61.950 22.950 64.050 25.050 ;
        RECT 79.950 22.950 82.050 25.050 ;
        RECT 82.950 22.950 85.050 25.050 ;
        RECT 85.950 22.950 88.050 25.050 ;
        RECT 88.950 22.950 91.050 25.050 ;
        RECT 103.950 22.950 106.050 25.050 ;
        RECT 106.950 22.950 109.050 25.050 ;
        RECT 109.950 22.950 112.050 25.050 ;
        RECT 112.950 22.950 115.050 25.050 ;
        RECT 127.950 22.950 130.050 25.050 ;
        RECT 130.950 22.950 133.050 25.050 ;
        RECT 133.950 22.950 136.050 25.050 ;
        RECT 136.950 22.950 139.050 25.050 ;
        RECT 151.950 22.950 154.050 25.050 ;
        RECT 154.950 22.950 157.050 25.050 ;
        RECT 157.950 22.950 160.050 25.050 ;
        RECT 160.950 22.950 163.050 25.050 ;
        RECT 175.950 22.950 178.050 25.050 ;
        RECT 178.950 22.950 181.050 25.050 ;
        RECT 193.950 22.950 196.050 25.050 ;
        RECT 196.950 22.950 199.050 25.050 ;
        RECT 199.950 22.950 202.050 25.050 ;
        RECT 202.950 22.950 205.050 25.050 ;
        RECT 208.950 24.450 213.000 25.050 ;
        RECT 208.950 22.950 213.450 24.450 ;
        RECT 217.950 22.950 220.050 25.050 ;
        RECT 220.950 22.950 223.050 25.050 ;
        RECT 223.950 22.950 226.050 25.050 ;
        RECT 226.950 22.950 229.050 25.050 ;
        RECT 244.950 22.950 247.050 25.050 ;
        RECT 247.950 22.950 250.050 25.050 ;
        RECT 250.950 22.950 253.050 25.050 ;
        RECT 253.950 22.950 256.050 25.050 ;
        RECT 268.950 22.950 271.050 25.050 ;
        RECT 271.950 22.950 274.050 25.050 ;
        RECT 274.950 22.950 277.050 25.050 ;
        RECT 277.950 22.950 280.050 25.050 ;
        RECT 292.950 22.950 295.050 25.050 ;
        RECT 295.950 22.950 298.050 25.050 ;
        RECT 298.950 22.950 301.050 25.050 ;
        RECT 301.950 22.950 304.050 25.050 ;
        RECT 316.950 22.950 319.050 25.050 ;
        RECT 319.950 22.950 322.050 25.050 ;
        RECT 322.950 22.950 325.050 25.050 ;
        RECT 325.950 22.950 328.050 25.050 ;
        RECT 343.950 22.950 346.050 25.050 ;
        RECT 346.950 22.950 349.050 25.050 ;
        RECT 349.950 22.950 352.050 25.050 ;
        RECT 352.950 22.950 355.050 25.050 ;
        RECT 368.400 22.950 370.500 25.050 ;
        RECT 14.700 9.600 15.900 22.950 ;
        RECT 17.100 21.150 18.900 22.950 ;
        RECT 32.100 21.150 33.900 22.950 ;
        RECT 35.100 9.600 36.300 22.950 ;
        RECT 56.100 15.600 57.300 22.950 ;
        RECT 62.100 21.150 63.900 22.950 ;
        RECT 80.100 21.150 81.900 22.950 ;
        RECT 58.950 18.450 61.050 19.050 ;
        RECT 82.950 18.450 85.050 19.050 ;
        RECT 58.950 17.550 85.050 18.450 ;
        RECT 58.950 16.950 61.050 17.550 ;
        RECT 82.950 16.950 85.050 17.550 ;
        RECT 86.700 15.600 87.900 22.950 ;
        RECT 107.100 21.150 108.900 22.950 ;
        RECT 56.100 14.100 58.500 15.600 ;
        RECT 54.000 11.100 55.800 12.900 ;
        RECT 14.100 3.600 15.900 9.600 ;
        RECT 17.100 3.000 18.900 9.600 ;
        RECT 32.100 3.000 33.900 9.600 ;
        RECT 35.100 3.600 36.900 9.600 ;
        RECT 53.700 3.000 55.500 9.600 ;
        RECT 56.700 3.600 58.500 14.100 ;
        RECT 61.800 3.000 63.600 15.600 ;
        RECT 80.400 3.000 82.200 15.600 ;
        RECT 85.500 14.100 87.900 15.600 ;
        RECT 91.950 15.450 94.050 16.050 ;
        RECT 106.950 15.450 109.050 16.050 ;
        RECT 91.950 14.550 109.050 15.450 ;
        RECT 85.500 3.600 87.300 14.100 ;
        RECT 91.950 13.950 94.050 14.550 ;
        RECT 106.950 13.950 109.050 14.550 ;
        RECT 88.200 11.100 90.000 12.900 ;
        RECT 113.100 10.800 114.000 22.950 ;
        RECT 131.100 21.150 132.900 22.950 ;
        RECT 137.100 10.800 138.000 22.950 ;
        RECT 155.250 21.150 157.050 22.950 ;
        RECT 161.700 15.600 162.600 22.950 ;
        RECT 176.100 21.150 177.900 22.950 ;
        RECT 107.400 9.900 114.000 10.800 ;
        RECT 107.400 9.600 108.900 9.900 ;
        RECT 88.500 3.000 90.300 9.600 ;
        RECT 104.100 3.000 105.900 9.600 ;
        RECT 107.100 3.600 108.900 9.600 ;
        RECT 113.100 9.600 114.000 9.900 ;
        RECT 131.400 9.900 138.000 10.800 ;
        RECT 131.400 9.600 132.900 9.900 ;
        RECT 110.100 3.000 111.900 9.000 ;
        RECT 113.100 3.600 114.900 9.600 ;
        RECT 128.100 3.000 129.900 9.600 ;
        RECT 131.100 3.600 132.900 9.600 ;
        RECT 137.100 9.600 138.000 9.900 ;
        RECT 152.100 14.700 159.900 15.600 ;
        RECT 134.100 3.000 135.900 9.000 ;
        RECT 137.100 3.600 138.900 9.600 ;
        RECT 152.100 3.600 153.900 14.700 ;
        RECT 155.100 3.000 156.900 13.800 ;
        RECT 158.100 3.600 159.900 14.700 ;
        RECT 161.100 3.600 162.900 15.600 ;
        RECT 179.100 9.600 180.300 22.950 ;
        RECT 197.250 21.150 199.050 22.950 ;
        RECT 203.700 15.600 204.600 22.950 ;
        RECT 212.550 22.050 213.450 22.950 ;
        RECT 212.550 20.550 217.050 22.050 ;
        RECT 221.100 21.150 222.900 22.950 ;
        RECT 213.000 19.950 217.050 20.550 ;
        RECT 208.950 18.450 211.050 19.050 ;
        RECT 223.950 18.450 226.050 19.050 ;
        RECT 208.950 17.550 226.050 18.450 ;
        RECT 208.950 16.950 211.050 17.550 ;
        RECT 223.950 16.950 226.050 17.550 ;
        RECT 194.100 14.700 201.900 15.600 ;
        RECT 176.100 3.000 177.900 9.600 ;
        RECT 179.100 3.600 180.900 9.600 ;
        RECT 194.100 3.600 195.900 14.700 ;
        RECT 197.100 3.000 198.900 13.800 ;
        RECT 200.100 3.600 201.900 14.700 ;
        RECT 203.100 3.600 204.900 15.600 ;
        RECT 227.100 10.800 228.000 22.950 ;
        RECT 245.100 21.150 246.900 22.950 ;
        RECT 251.700 15.600 252.900 22.950 ;
        RECT 256.950 21.450 259.050 22.050 ;
        RECT 262.950 21.450 265.050 22.050 ;
        RECT 256.950 20.550 265.050 21.450 ;
        RECT 256.950 19.950 259.050 20.550 ;
        RECT 262.950 19.950 265.050 20.550 ;
        RECT 221.400 9.900 228.000 10.800 ;
        RECT 221.400 9.600 222.900 9.900 ;
        RECT 218.100 3.000 219.900 9.600 ;
        RECT 221.100 3.600 222.900 9.600 ;
        RECT 227.100 9.600 228.000 9.900 ;
        RECT 224.100 3.000 225.900 9.000 ;
        RECT 227.100 3.600 228.900 9.600 ;
        RECT 245.400 3.000 247.200 15.600 ;
        RECT 250.500 14.100 252.900 15.600 ;
        RECT 250.500 3.600 252.300 14.100 ;
        RECT 253.200 11.100 255.000 12.900 ;
        RECT 270.000 10.800 270.900 22.950 ;
        RECT 275.100 21.150 276.900 22.950 ;
        RECT 296.100 15.600 297.300 22.950 ;
        RECT 302.100 21.150 303.900 22.950 ;
        RECT 317.100 21.150 318.900 22.950 ;
        RECT 323.700 15.600 324.900 22.950 ;
        RECT 347.250 21.150 349.050 22.950 ;
        RECT 353.700 15.600 354.600 22.950 ;
        RECT 368.400 21.150 370.200 22.950 ;
        RECT 372.000 18.300 372.900 29.700 ;
        RECT 374.700 25.050 375.900 32.400 ;
        RECT 373.800 22.950 375.900 25.050 ;
        RECT 372.000 17.400 373.800 18.300 ;
        RECT 368.100 16.500 373.800 17.400 ;
        RECT 296.100 14.100 298.500 15.600 ;
        RECT 294.000 11.100 295.800 12.900 ;
        RECT 270.000 9.900 276.600 10.800 ;
        RECT 270.000 9.600 270.900 9.900 ;
        RECT 253.500 3.000 255.300 9.600 ;
        RECT 269.100 3.600 270.900 9.600 ;
        RECT 275.100 9.600 276.600 9.900 ;
        RECT 272.100 3.000 273.900 9.000 ;
        RECT 275.100 3.600 276.900 9.600 ;
        RECT 278.100 3.000 279.900 9.600 ;
        RECT 293.700 3.000 295.500 9.600 ;
        RECT 296.700 3.600 298.500 14.100 ;
        RECT 301.800 3.000 303.600 15.600 ;
        RECT 317.400 3.000 319.200 15.600 ;
        RECT 322.500 14.100 324.900 15.600 ;
        RECT 344.100 14.700 351.900 15.600 ;
        RECT 322.500 3.600 324.300 14.100 ;
        RECT 325.200 11.100 327.000 12.900 ;
        RECT 325.500 3.000 327.300 9.600 ;
        RECT 344.100 3.600 345.900 14.700 ;
        RECT 347.100 3.000 348.900 13.800 ;
        RECT 350.100 3.600 351.900 14.700 ;
        RECT 353.100 3.600 354.900 15.600 ;
        RECT 368.100 9.600 369.300 16.500 ;
        RECT 374.700 15.600 375.900 22.950 ;
        RECT 368.100 3.600 369.900 9.600 ;
        RECT 371.100 3.000 372.900 13.800 ;
        RECT 374.100 3.600 375.900 15.600 ;
        RECT 389.100 32.400 390.900 38.400 ;
        RECT 392.100 32.400 393.900 39.000 ;
        RECT 395.100 35.400 396.900 38.400 ;
        RECT 389.100 25.050 390.300 32.400 ;
        RECT 395.700 31.500 396.900 35.400 ;
        RECT 391.200 30.600 396.900 31.500 ;
        RECT 413.100 32.400 414.900 38.400 ;
        RECT 416.100 32.400 417.900 39.000 ;
        RECT 419.100 35.400 420.900 38.400 ;
        RECT 434.100 35.400 435.900 38.400 ;
        RECT 437.100 35.400 438.900 39.000 ;
        RECT 391.200 29.700 393.000 30.600 ;
        RECT 389.100 22.950 391.200 25.050 ;
        RECT 389.100 15.600 390.300 22.950 ;
        RECT 392.100 18.300 393.000 29.700 ;
        RECT 413.100 25.050 414.300 32.400 ;
        RECT 419.700 31.500 420.900 35.400 ;
        RECT 415.200 30.600 420.900 31.500 ;
        RECT 415.200 29.700 417.000 30.600 ;
        RECT 394.500 22.950 396.600 25.050 ;
        RECT 394.800 21.150 396.600 22.950 ;
        RECT 413.100 22.950 415.200 25.050 ;
        RECT 391.200 17.400 393.000 18.300 ;
        RECT 391.200 16.500 396.900 17.400 ;
        RECT 389.100 3.600 390.900 15.600 ;
        RECT 392.100 3.000 393.900 13.800 ;
        RECT 395.700 9.600 396.900 16.500 ;
        RECT 395.100 3.600 396.900 9.600 ;
        RECT 413.100 15.600 414.300 22.950 ;
        RECT 416.100 18.300 417.000 29.700 ;
        RECT 434.700 25.050 435.900 35.400 ;
        RECT 455.100 32.400 456.900 38.400 ;
        RECT 455.700 30.300 456.900 32.400 ;
        RECT 458.100 33.300 459.900 38.400 ;
        RECT 461.100 34.200 462.900 39.000 ;
        RECT 464.100 33.300 465.900 38.400 ;
        RECT 458.100 31.950 465.900 33.300 ;
        RECT 455.700 29.400 459.300 30.300 ;
        RECT 481.500 30.000 483.300 38.400 ;
        RECT 455.100 25.050 456.900 26.850 ;
        RECT 458.100 25.050 459.300 29.400 ;
        RECT 480.000 28.800 483.300 30.000 ;
        RECT 488.100 29.400 489.900 39.000 ;
        RECT 503.700 35.400 505.500 39.000 ;
        RECT 506.700 33.600 508.500 38.400 ;
        RECT 503.400 32.400 508.500 33.600 ;
        RECT 511.200 32.400 513.000 39.000 ;
        RECT 461.100 25.050 462.900 26.850 ;
        RECT 480.000 25.050 480.900 28.800 ;
        RECT 482.100 25.050 483.900 26.850 ;
        RECT 488.100 25.050 489.900 26.850 ;
        RECT 503.400 25.050 504.300 32.400 ;
        RECT 530.100 29.400 531.900 39.000 ;
        RECT 536.700 30.000 538.500 38.400 ;
        RECT 554.100 32.400 555.900 38.400 ;
        RECT 554.700 30.300 555.900 32.400 ;
        RECT 557.100 33.300 558.900 38.400 ;
        RECT 560.100 34.200 561.900 39.000 ;
        RECT 563.100 33.300 564.900 38.400 ;
        RECT 557.100 31.950 564.900 33.300 ;
        RECT 581.100 33.300 582.900 38.400 ;
        RECT 584.100 34.200 585.900 39.000 ;
        RECT 587.100 33.300 588.900 38.400 ;
        RECT 581.100 31.950 588.900 33.300 ;
        RECT 590.100 32.400 591.900 38.400 ;
        RECT 590.100 30.300 591.300 32.400 ;
        RECT 536.700 28.800 540.000 30.000 ;
        RECT 554.700 29.400 558.300 30.300 ;
        RECT 505.950 25.050 507.750 26.850 ;
        RECT 512.100 25.050 513.900 26.850 ;
        RECT 530.100 25.050 531.900 26.850 ;
        RECT 536.100 25.050 537.900 26.850 ;
        RECT 539.100 25.050 540.000 28.800 ;
        RECT 554.100 25.050 555.900 26.850 ;
        RECT 557.100 25.050 558.300 29.400 ;
        RECT 587.700 29.400 591.300 30.300 ;
        RECT 607.500 30.000 609.300 38.400 ;
        RECT 560.100 25.050 561.900 26.850 ;
        RECT 584.100 25.050 585.900 26.850 ;
        RECT 587.700 25.050 588.900 29.400 ;
        RECT 606.000 28.800 609.300 30.000 ;
        RECT 614.100 29.400 615.900 39.000 ;
        RECT 629.700 35.400 631.500 39.000 ;
        RECT 632.700 33.600 634.500 38.400 ;
        RECT 629.400 32.400 634.500 33.600 ;
        RECT 637.200 32.400 639.000 39.000 ;
        RECT 653.100 35.400 654.900 39.000 ;
        RECT 656.100 35.400 657.900 38.400 ;
        RECT 590.100 25.050 591.900 26.850 ;
        RECT 606.000 25.050 606.900 28.800 ;
        RECT 608.100 25.050 609.900 26.850 ;
        RECT 614.100 25.050 615.900 26.850 ;
        RECT 629.400 25.050 630.300 32.400 ;
        RECT 631.950 25.050 633.750 26.850 ;
        RECT 638.100 25.050 639.900 26.850 ;
        RECT 656.100 25.050 657.300 35.400 ;
        RECT 672.000 32.400 673.800 39.000 ;
        RECT 676.500 33.600 678.300 38.400 ;
        RECT 679.500 35.400 681.300 39.000 ;
        RECT 676.500 32.400 681.600 33.600 ;
        RECT 699.000 32.400 700.800 39.000 ;
        RECT 703.500 33.600 705.300 38.400 ;
        RECT 706.500 35.400 708.300 39.000 ;
        RECT 722.100 35.400 723.900 38.400 ;
        RECT 725.100 35.400 726.900 39.000 ;
        RECT 703.500 32.400 708.600 33.600 ;
        RECT 667.950 27.450 670.050 31.050 ;
        RECT 665.550 27.000 670.050 27.450 ;
        RECT 665.550 26.550 669.450 27.000 ;
        RECT 418.500 22.950 420.600 25.050 ;
        RECT 433.950 22.950 436.050 25.050 ;
        RECT 436.950 22.950 439.050 25.050 ;
        RECT 454.950 22.950 457.050 25.050 ;
        RECT 457.950 22.950 460.050 25.050 ;
        RECT 460.950 22.950 463.050 25.050 ;
        RECT 463.950 22.950 466.050 25.050 ;
        RECT 478.950 22.950 481.050 25.050 ;
        RECT 481.950 22.950 484.050 25.050 ;
        RECT 484.950 22.950 487.050 25.050 ;
        RECT 487.950 22.950 490.050 25.050 ;
        RECT 502.950 22.950 505.050 25.050 ;
        RECT 505.950 22.950 508.050 25.050 ;
        RECT 508.950 22.950 511.050 25.050 ;
        RECT 511.950 22.950 514.050 25.050 ;
        RECT 529.950 22.950 532.050 25.050 ;
        RECT 532.950 22.950 535.050 25.050 ;
        RECT 535.950 22.950 538.050 25.050 ;
        RECT 538.950 22.950 541.050 25.050 ;
        RECT 553.950 22.950 556.050 25.050 ;
        RECT 556.950 22.950 559.050 25.050 ;
        RECT 559.950 22.950 562.050 25.050 ;
        RECT 562.950 22.950 565.050 25.050 ;
        RECT 580.950 22.950 583.050 25.050 ;
        RECT 583.950 22.950 586.050 25.050 ;
        RECT 586.950 22.950 589.050 25.050 ;
        RECT 589.950 22.950 592.050 25.050 ;
        RECT 604.950 22.950 607.050 25.050 ;
        RECT 607.950 22.950 610.050 25.050 ;
        RECT 610.950 22.950 613.050 25.050 ;
        RECT 613.950 22.950 616.050 25.050 ;
        RECT 628.950 22.950 631.050 25.050 ;
        RECT 631.950 22.950 634.050 25.050 ;
        RECT 634.950 22.950 637.050 25.050 ;
        RECT 637.950 22.950 640.050 25.050 ;
        RECT 652.950 22.950 655.050 25.050 ;
        RECT 655.950 22.950 658.050 25.050 ;
        RECT 418.800 21.150 420.600 22.950 ;
        RECT 415.200 17.400 417.000 18.300 ;
        RECT 415.200 16.500 420.900 17.400 ;
        RECT 413.100 3.600 414.900 15.600 ;
        RECT 416.100 3.000 417.900 13.800 ;
        RECT 419.700 9.600 420.900 16.500 ;
        RECT 434.700 9.600 435.900 22.950 ;
        RECT 437.100 21.150 438.900 22.950 ;
        RECT 458.100 15.600 459.300 22.950 ;
        RECT 464.100 21.150 465.900 22.950 ;
        RECT 458.100 14.100 460.500 15.600 ;
        RECT 456.000 11.100 457.800 12.900 ;
        RECT 419.100 3.600 420.900 9.600 ;
        RECT 434.100 3.600 435.900 9.600 ;
        RECT 437.100 3.000 438.900 9.600 ;
        RECT 455.700 3.000 457.500 9.600 ;
        RECT 458.700 3.600 460.500 14.100 ;
        RECT 463.800 3.000 465.600 15.600 ;
        RECT 480.000 10.800 480.900 22.950 ;
        RECT 485.100 21.150 486.900 22.950 ;
        RECT 490.950 21.450 493.050 22.050 ;
        RECT 496.950 21.450 499.050 22.050 ;
        RECT 490.950 20.550 499.050 21.450 ;
        RECT 490.950 19.950 493.050 20.550 ;
        RECT 496.950 19.950 499.050 20.550 ;
        RECT 503.400 15.600 504.300 22.950 ;
        RECT 508.950 21.150 510.750 22.950 ;
        RECT 533.100 21.150 534.900 22.950 ;
        RECT 480.000 9.900 486.600 10.800 ;
        RECT 480.000 9.600 480.900 9.900 ;
        RECT 479.100 3.600 480.900 9.600 ;
        RECT 485.100 9.600 486.600 9.900 ;
        RECT 482.100 3.000 483.900 9.000 ;
        RECT 485.100 3.600 486.900 9.600 ;
        RECT 488.100 3.000 489.900 9.600 ;
        RECT 503.100 3.600 504.900 15.600 ;
        RECT 506.100 14.700 513.900 15.600 ;
        RECT 506.100 3.600 507.900 14.700 ;
        RECT 509.100 3.000 510.900 13.800 ;
        RECT 512.100 3.600 513.900 14.700 ;
        RECT 539.100 10.800 540.000 22.950 ;
        RECT 557.100 15.600 558.300 22.950 ;
        RECT 563.100 21.150 564.900 22.950 ;
        RECT 581.100 21.150 582.900 22.950 ;
        RECT 587.700 15.600 588.900 22.950 ;
        RECT 557.100 14.100 559.500 15.600 ;
        RECT 555.000 11.100 556.800 12.900 ;
        RECT 533.400 9.900 540.000 10.800 ;
        RECT 533.400 9.600 534.900 9.900 ;
        RECT 530.100 3.000 531.900 9.600 ;
        RECT 533.100 3.600 534.900 9.600 ;
        RECT 539.100 9.600 540.000 9.900 ;
        RECT 536.100 3.000 537.900 9.000 ;
        RECT 539.100 3.600 540.900 9.600 ;
        RECT 554.700 3.000 556.500 9.600 ;
        RECT 557.700 3.600 559.500 14.100 ;
        RECT 562.800 3.000 564.600 15.600 ;
        RECT 581.400 3.000 583.200 15.600 ;
        RECT 586.500 14.100 588.900 15.600 ;
        RECT 586.500 3.600 588.300 14.100 ;
        RECT 589.200 11.100 591.000 12.900 ;
        RECT 606.000 10.800 606.900 22.950 ;
        RECT 611.100 21.150 612.900 22.950 ;
        RECT 629.400 15.600 630.300 22.950 ;
        RECT 634.950 21.150 636.750 22.950 ;
        RECT 653.100 21.150 654.900 22.950 ;
        RECT 637.950 18.450 640.050 19.050 ;
        RECT 643.950 18.450 646.050 19.050 ;
        RECT 637.950 17.550 646.050 18.450 ;
        RECT 637.950 16.950 640.050 17.550 ;
        RECT 643.950 16.950 646.050 17.550 ;
        RECT 606.000 9.900 612.600 10.800 ;
        RECT 606.000 9.600 606.900 9.900 ;
        RECT 589.500 3.000 591.300 9.600 ;
        RECT 605.100 3.600 606.900 9.600 ;
        RECT 611.100 9.600 612.600 9.900 ;
        RECT 608.100 3.000 609.900 9.000 ;
        RECT 611.100 3.600 612.900 9.600 ;
        RECT 614.100 3.000 615.900 9.600 ;
        RECT 629.100 3.600 630.900 15.600 ;
        RECT 632.100 14.700 639.900 15.600 ;
        RECT 632.100 3.600 633.900 14.700 ;
        RECT 635.100 3.000 636.900 13.800 ;
        RECT 638.100 3.600 639.900 14.700 ;
        RECT 656.100 9.600 657.300 22.950 ;
        RECT 658.950 21.450 661.050 22.050 ;
        RECT 665.550 21.450 666.450 26.550 ;
        RECT 671.100 25.050 672.900 26.850 ;
        RECT 677.250 25.050 679.050 26.850 ;
        RECT 680.700 25.050 681.600 32.400 ;
        RECT 698.100 25.050 699.900 26.850 ;
        RECT 704.250 25.050 706.050 26.850 ;
        RECT 707.700 25.050 708.600 32.400 ;
        RECT 722.700 25.050 723.900 35.400 ;
        RECT 743.100 33.300 744.900 38.400 ;
        RECT 746.100 34.200 747.900 39.000 ;
        RECT 749.100 33.300 750.900 38.400 ;
        RECT 743.100 31.950 750.900 33.300 ;
        RECT 752.100 32.400 753.900 38.400 ;
        RECT 770.100 35.400 771.900 39.000 ;
        RECT 773.100 35.400 774.900 38.400 ;
        RECT 752.100 30.300 753.300 32.400 ;
        RECT 749.700 29.400 753.300 30.300 ;
        RECT 746.100 25.050 747.900 26.850 ;
        RECT 749.700 25.050 750.900 29.400 ;
        RECT 752.100 25.050 753.900 26.850 ;
        RECT 773.100 25.050 774.300 35.400 ;
        RECT 791.100 29.400 792.900 39.000 ;
        RECT 797.700 30.000 799.500 38.400 ;
        RECT 815.700 35.400 817.500 39.000 ;
        RECT 818.700 33.600 820.500 38.400 ;
        RECT 815.400 32.400 820.500 33.600 ;
        RECT 823.200 32.400 825.000 39.000 ;
        RECT 797.700 28.800 801.000 30.000 ;
        RECT 791.100 25.050 792.900 26.850 ;
        RECT 797.100 25.050 798.900 26.850 ;
        RECT 800.100 25.050 801.000 28.800 ;
        RECT 815.400 25.050 816.300 32.400 ;
        RECT 841.500 30.000 843.300 38.400 ;
        RECT 840.000 28.800 843.300 30.000 ;
        RECT 848.100 29.400 849.900 39.000 ;
        RECT 863.100 35.400 864.900 39.000 ;
        RECT 866.100 35.400 867.900 38.400 ;
        RECT 817.950 25.050 819.750 26.850 ;
        RECT 824.100 25.050 825.900 26.850 ;
        RECT 840.000 25.050 840.900 28.800 ;
        RECT 842.100 25.050 843.900 26.850 ;
        RECT 848.100 25.050 849.900 26.850 ;
        RECT 866.100 25.050 867.300 35.400 ;
        RECT 884.100 32.400 885.900 38.400 ;
        RECT 884.700 30.300 885.900 32.400 ;
        RECT 887.100 33.300 888.900 38.400 ;
        RECT 890.100 34.200 891.900 39.000 ;
        RECT 893.100 33.300 894.900 38.400 ;
        RECT 887.100 31.950 894.900 33.300 ;
        RECT 908.100 32.400 909.900 38.400 ;
        RECT 908.700 30.300 909.900 32.400 ;
        RECT 911.100 33.300 912.900 38.400 ;
        RECT 914.100 34.200 915.900 39.000 ;
        RECT 917.100 33.300 918.900 38.400 ;
        RECT 911.100 31.950 918.900 33.300 ;
        RECT 884.700 29.400 888.300 30.300 ;
        RECT 908.700 29.400 912.300 30.300 ;
        RECT 934.500 30.000 936.300 38.400 ;
        RECT 884.100 25.050 885.900 26.850 ;
        RECT 887.100 25.050 888.300 29.400 ;
        RECT 890.100 25.050 891.900 26.850 ;
        RECT 908.100 25.050 909.900 26.850 ;
        RECT 911.100 25.050 912.300 29.400 ;
        RECT 933.000 28.800 936.300 30.000 ;
        RECT 941.100 29.400 942.900 39.000 ;
        RECT 961.500 30.000 963.300 38.400 ;
        RECT 960.000 28.800 963.300 30.000 ;
        RECT 968.100 29.400 969.900 39.000 ;
        RECT 986.700 35.400 988.500 39.000 ;
        RECT 989.700 33.600 991.500 38.400 ;
        RECT 986.400 32.400 991.500 33.600 ;
        RECT 994.200 32.400 996.000 39.000 ;
        RECT 914.100 25.050 915.900 26.850 ;
        RECT 933.000 25.050 933.900 28.800 ;
        RECT 935.100 25.050 936.900 26.850 ;
        RECT 941.100 25.050 942.900 26.850 ;
        RECT 960.000 25.050 960.900 28.800 ;
        RECT 962.100 25.050 963.900 26.850 ;
        RECT 968.100 25.050 969.900 26.850 ;
        RECT 986.400 25.050 987.300 32.400 ;
        RECT 988.950 25.050 990.750 26.850 ;
        RECT 995.100 25.050 996.900 26.850 ;
        RECT 670.950 22.950 673.050 25.050 ;
        RECT 673.950 22.950 676.050 25.050 ;
        RECT 676.950 22.950 679.050 25.050 ;
        RECT 679.950 22.950 682.050 25.050 ;
        RECT 697.950 22.950 700.050 25.050 ;
        RECT 700.950 22.950 703.050 25.050 ;
        RECT 703.950 22.950 706.050 25.050 ;
        RECT 706.950 22.950 709.050 25.050 ;
        RECT 721.950 22.950 724.050 25.050 ;
        RECT 724.950 22.950 727.050 25.050 ;
        RECT 742.950 22.950 745.050 25.050 ;
        RECT 745.950 22.950 748.050 25.050 ;
        RECT 748.950 22.950 751.050 25.050 ;
        RECT 751.950 22.950 754.050 25.050 ;
        RECT 769.950 22.950 772.050 25.050 ;
        RECT 772.950 22.950 775.050 25.050 ;
        RECT 790.950 22.950 793.050 25.050 ;
        RECT 793.950 22.950 796.050 25.050 ;
        RECT 796.950 22.950 799.050 25.050 ;
        RECT 799.950 22.950 802.050 25.050 ;
        RECT 814.950 22.950 817.050 25.050 ;
        RECT 817.950 22.950 820.050 25.050 ;
        RECT 820.950 22.950 823.050 25.050 ;
        RECT 823.950 22.950 826.050 25.050 ;
        RECT 838.950 22.950 841.050 25.050 ;
        RECT 841.950 22.950 844.050 25.050 ;
        RECT 844.950 22.950 847.050 25.050 ;
        RECT 847.950 22.950 850.050 25.050 ;
        RECT 862.950 22.950 865.050 25.050 ;
        RECT 865.950 22.950 868.050 25.050 ;
        RECT 883.950 22.950 886.050 25.050 ;
        RECT 886.950 22.950 889.050 25.050 ;
        RECT 889.950 22.950 892.050 25.050 ;
        RECT 892.950 22.950 895.050 25.050 ;
        RECT 907.950 22.950 910.050 25.050 ;
        RECT 910.950 22.950 913.050 25.050 ;
        RECT 913.950 22.950 916.050 25.050 ;
        RECT 916.950 22.950 919.050 25.050 ;
        RECT 931.950 22.950 934.050 25.050 ;
        RECT 934.950 22.950 937.050 25.050 ;
        RECT 937.950 22.950 940.050 25.050 ;
        RECT 940.950 22.950 943.050 25.050 ;
        RECT 958.950 22.950 961.050 25.050 ;
        RECT 961.950 22.950 964.050 25.050 ;
        RECT 964.950 22.950 967.050 25.050 ;
        RECT 967.950 22.950 970.050 25.050 ;
        RECT 985.950 22.950 988.050 25.050 ;
        RECT 988.950 22.950 991.050 25.050 ;
        RECT 991.950 22.950 994.050 25.050 ;
        RECT 994.950 22.950 997.050 25.050 ;
        RECT 658.950 20.550 666.450 21.450 ;
        RECT 674.250 21.150 676.050 22.950 ;
        RECT 658.950 19.950 661.050 20.550 ;
        RECT 664.950 18.450 667.050 19.050 ;
        RECT 676.950 18.450 679.050 19.050 ;
        RECT 664.950 17.550 679.050 18.450 ;
        RECT 664.950 16.950 667.050 17.550 ;
        RECT 676.950 16.950 679.050 17.550 ;
        RECT 680.700 15.600 681.600 22.950 ;
        RECT 701.250 21.150 703.050 22.950 ;
        RECT 707.700 15.600 708.600 22.950 ;
        RECT 671.100 14.700 678.900 15.600 ;
        RECT 653.100 3.000 654.900 9.600 ;
        RECT 656.100 3.600 657.900 9.600 ;
        RECT 671.100 3.600 672.900 14.700 ;
        RECT 674.100 3.000 675.900 13.800 ;
        RECT 677.100 3.600 678.900 14.700 ;
        RECT 680.100 3.600 681.900 15.600 ;
        RECT 698.100 14.700 705.900 15.600 ;
        RECT 698.100 3.600 699.900 14.700 ;
        RECT 701.100 3.000 702.900 13.800 ;
        RECT 704.100 3.600 705.900 14.700 ;
        RECT 707.100 3.600 708.900 15.600 ;
        RECT 722.700 9.600 723.900 22.950 ;
        RECT 725.100 21.150 726.900 22.950 ;
        RECT 743.100 21.150 744.900 22.950 ;
        RECT 749.700 15.600 750.900 22.950 ;
        RECT 770.100 21.150 771.900 22.950 ;
        RECT 722.100 3.600 723.900 9.600 ;
        RECT 725.100 3.000 726.900 9.600 ;
        RECT 743.400 3.000 745.200 15.600 ;
        RECT 748.500 14.100 750.900 15.600 ;
        RECT 748.500 3.600 750.300 14.100 ;
        RECT 751.200 11.100 753.000 12.900 ;
        RECT 773.100 9.600 774.300 22.950 ;
        RECT 794.100 21.150 795.900 22.950 ;
        RECT 800.100 10.800 801.000 22.950 ;
        RECT 815.400 15.600 816.300 22.950 ;
        RECT 820.950 21.150 822.750 22.950 ;
        RECT 794.400 9.900 801.000 10.800 ;
        RECT 794.400 9.600 795.900 9.900 ;
        RECT 751.500 3.000 753.300 9.600 ;
        RECT 770.100 3.000 771.900 9.600 ;
        RECT 773.100 3.600 774.900 9.600 ;
        RECT 791.100 3.000 792.900 9.600 ;
        RECT 794.100 3.600 795.900 9.600 ;
        RECT 800.100 9.600 801.000 9.900 ;
        RECT 797.100 3.000 798.900 9.000 ;
        RECT 800.100 3.600 801.900 9.600 ;
        RECT 815.100 3.600 816.900 15.600 ;
        RECT 818.100 14.700 825.900 15.600 ;
        RECT 818.100 3.600 819.900 14.700 ;
        RECT 821.100 3.000 822.900 13.800 ;
        RECT 824.100 3.600 825.900 14.700 ;
        RECT 840.000 10.800 840.900 22.950 ;
        RECT 845.100 21.150 846.900 22.950 ;
        RECT 863.100 21.150 864.900 22.950 ;
        RECT 840.000 9.900 846.600 10.800 ;
        RECT 840.000 9.600 840.900 9.900 ;
        RECT 839.100 3.600 840.900 9.600 ;
        RECT 845.100 9.600 846.600 9.900 ;
        RECT 866.100 9.600 867.300 22.950 ;
        RECT 887.100 15.600 888.300 22.950 ;
        RECT 893.100 21.150 894.900 22.950 ;
        RECT 898.950 18.450 901.050 18.900 ;
        RECT 907.950 18.450 910.050 19.050 ;
        RECT 898.950 17.550 910.050 18.450 ;
        RECT 898.950 16.800 901.050 17.550 ;
        RECT 907.950 16.950 910.050 17.550 ;
        RECT 911.100 15.600 912.300 22.950 ;
        RECT 917.100 21.150 918.900 22.950 ;
        RECT 887.100 14.100 889.500 15.600 ;
        RECT 885.000 11.100 886.800 12.900 ;
        RECT 842.100 3.000 843.900 9.000 ;
        RECT 845.100 3.600 846.900 9.600 ;
        RECT 848.100 3.000 849.900 9.600 ;
        RECT 863.100 3.000 864.900 9.600 ;
        RECT 866.100 3.600 867.900 9.600 ;
        RECT 884.700 3.000 886.500 9.600 ;
        RECT 887.700 3.600 889.500 14.100 ;
        RECT 892.800 3.000 894.600 15.600 ;
        RECT 911.100 14.100 913.500 15.600 ;
        RECT 909.000 11.100 910.800 12.900 ;
        RECT 908.700 3.000 910.500 9.600 ;
        RECT 911.700 3.600 913.500 14.100 ;
        RECT 916.800 3.000 918.600 15.600 ;
        RECT 933.000 10.800 933.900 22.950 ;
        RECT 938.100 21.150 939.900 22.950 ;
        RECT 943.950 21.450 946.050 22.050 ;
        RECT 949.950 21.450 952.050 22.050 ;
        RECT 943.950 20.550 952.050 21.450 ;
        RECT 943.950 19.950 946.050 20.550 ;
        RECT 949.950 19.950 952.050 20.550 ;
        RECT 960.000 10.800 960.900 22.950 ;
        RECT 965.100 21.150 966.900 22.950 ;
        RECT 986.400 15.600 987.300 22.950 ;
        RECT 991.950 21.150 993.750 22.950 ;
        RECT 933.000 9.900 939.600 10.800 ;
        RECT 933.000 9.600 933.900 9.900 ;
        RECT 932.100 3.600 933.900 9.600 ;
        RECT 938.100 9.600 939.600 9.900 ;
        RECT 960.000 9.900 966.600 10.800 ;
        RECT 960.000 9.600 960.900 9.900 ;
        RECT 935.100 3.000 936.900 9.000 ;
        RECT 938.100 3.600 939.900 9.600 ;
        RECT 941.100 3.000 942.900 9.600 ;
        RECT 959.100 3.600 960.900 9.600 ;
        RECT 965.100 9.600 966.600 9.900 ;
        RECT 962.100 3.000 963.900 9.000 ;
        RECT 965.100 3.600 966.900 9.600 ;
        RECT 968.100 3.000 969.900 9.600 ;
        RECT 986.100 3.600 987.900 15.600 ;
        RECT 989.100 14.700 996.900 15.600 ;
        RECT 989.100 3.600 990.900 14.700 ;
        RECT 992.100 3.000 993.900 13.800 ;
        RECT 995.100 3.600 996.900 14.700 ;
      LAYER via1 ;
        RECT 244.950 925.950 247.050 928.050 ;
        RECT 475.950 922.950 478.050 925.050 ;
        RECT 565.950 916.950 568.050 919.050 ;
        RECT 589.950 892.950 592.050 895.050 ;
        RECT 179.100 835.950 181.200 838.050 ;
        RECT 196.950 835.950 199.050 838.050 ;
        RECT 191.550 825.600 193.650 827.700 ;
        RECT 886.950 838.950 889.050 841.050 ;
        RECT 973.950 832.950 976.050 835.050 ;
        RECT 22.950 802.950 25.050 805.050 ;
        RECT 224.550 813.300 226.650 815.400 ;
        RECT 281.100 808.800 283.200 810.900 ;
        RECT 313.800 808.800 315.900 810.900 ;
        RECT 361.950 805.950 364.050 808.050 ;
        RECT 529.950 805.950 532.050 808.050 ;
        RECT 529.950 799.950 532.050 802.050 ;
        RECT 626.100 808.800 628.200 810.900 ;
        RECT 874.950 805.950 877.050 808.050 ;
        RECT 874.950 799.950 877.050 802.050 ;
        RECT 955.950 808.950 958.050 811.050 ;
        RECT 991.950 805.950 994.050 808.050 ;
        RECT 82.500 751.800 84.600 753.900 ;
        RECT 94.800 757.950 96.900 760.050 ;
        RECT 298.950 763.950 301.050 766.050 ;
        RECT 448.500 751.800 450.600 753.900 ;
        RECT 460.800 757.950 462.900 760.050 ;
        RECT 691.950 760.950 694.050 763.050 ;
        RECT 271.800 730.800 273.900 732.900 ;
        RECT 358.950 727.950 361.050 730.050 ;
        RECT 358.950 721.950 361.050 724.050 ;
        RECT 832.950 727.950 835.050 730.050 ;
        RECT 985.950 727.950 988.050 730.050 ;
        RECT 985.950 721.950 988.050 724.050 ;
        RECT 4.950 679.950 7.050 682.050 ;
        RECT 22.800 679.950 24.900 682.050 ;
        RECT 101.100 679.950 103.200 682.050 ;
        RECT 103.500 673.500 105.600 675.600 ;
        RECT 110.100 682.950 112.200 685.050 ;
        RECT 110.100 674.100 112.200 676.200 ;
        RECT 113.400 673.800 115.500 675.900 ;
        RECT 361.950 676.950 364.050 679.050 ;
        RECT 679.500 673.800 681.600 675.900 ;
        RECT 691.800 679.950 693.900 682.050 ;
        RECT 829.950 685.950 832.050 688.050 ;
        RECT 868.950 682.950 871.050 685.050 ;
        RECT 826.950 676.950 829.050 679.050 ;
        RECT 958.950 679.950 961.050 682.050 ;
        RECT 92.550 657.300 94.650 659.400 ;
        RECT 136.950 643.950 139.050 646.050 ;
        RECT 200.550 657.300 202.650 659.400 ;
        RECT 295.950 646.950 298.050 649.050 ;
        RECT 377.550 657.300 379.650 659.400 ;
        RECT 413.550 657.300 415.650 659.400 ;
        RECT 616.800 652.800 618.900 654.900 ;
        RECT 871.950 646.950 874.050 649.050 ;
        RECT 874.950 643.950 877.050 646.050 ;
        RECT 925.950 643.950 928.050 646.050 ;
        RECT 1000.950 649.950 1003.050 652.050 ;
        RECT 4.950 601.950 7.050 604.050 ;
        RECT 22.800 601.950 24.900 604.050 ;
        RECT 98.100 601.950 100.200 604.050 ;
        RECT 115.950 601.950 118.050 604.050 ;
        RECT 110.550 591.600 112.650 593.700 ;
        RECT 200.100 601.950 202.200 604.050 ;
        RECT 217.950 601.950 220.050 604.050 ;
        RECT 212.550 591.600 214.650 593.700 ;
        RECT 295.950 601.950 298.050 604.050 ;
        RECT 313.800 601.950 315.900 604.050 ;
        RECT 349.950 601.950 352.050 604.050 ;
        RECT 367.800 601.950 369.900 604.050 ;
        RECT 586.950 604.950 589.050 607.050 ;
        RECT 634.950 607.950 637.050 610.050 ;
        RECT 676.950 604.950 679.050 607.050 ;
        RECT 631.950 598.950 634.050 601.050 ;
        RECT 886.950 598.950 889.050 601.050 ;
        RECT 92.550 579.300 94.650 581.400 ;
        RECT 106.950 568.950 109.050 571.050 ;
        RECT 323.550 579.300 325.650 581.400 ;
        RECT 401.550 579.300 403.650 581.400 ;
        RECT 439.950 568.950 442.050 571.050 ;
        RECT 497.550 579.300 499.650 581.400 ;
        RECT 583.950 571.950 586.050 574.050 ;
        RECT 620.550 579.300 622.650 581.400 ;
        RECT 712.950 571.950 715.050 574.050 ;
        RECT 748.950 574.800 751.050 576.900 ;
        RECT 712.950 565.950 715.050 568.050 ;
        RECT 757.950 565.950 760.050 568.050 ;
        RECT 949.950 571.950 952.050 574.050 ;
        RECT 997.950 571.950 1000.050 574.050 ;
        RECT 160.950 526.950 163.050 529.050 ;
        RECT 64.950 523.950 67.050 526.050 ;
        RECT 191.100 523.950 193.200 526.050 ;
        RECT 208.950 523.950 211.050 526.050 ;
        RECT 203.550 513.600 205.650 515.700 ;
        RECT 418.950 526.950 421.050 529.050 ;
        RECT 436.950 523.950 439.050 526.050 ;
        RECT 418.950 520.950 421.050 523.050 ;
        RECT 454.800 523.950 456.900 526.050 ;
        RECT 535.950 523.950 538.050 526.050 ;
        RECT 553.800 523.950 555.900 526.050 ;
        RECT 883.950 526.950 886.050 529.050 ;
        RECT 934.950 526.950 937.050 529.050 ;
        RECT 86.550 501.300 88.650 503.400 ;
        RECT 122.550 501.300 124.650 503.400 ;
        RECT 266.550 501.300 268.650 503.400 ;
        RECT 302.550 501.300 304.650 503.400 ;
        RECT 362.550 501.300 364.650 503.400 ;
        RECT 559.950 490.950 562.050 493.050 ;
        RECT 874.950 499.950 877.050 502.050 ;
        RECT 907.950 493.950 910.050 496.050 ;
        RECT 955.950 493.950 958.050 496.050 ;
        RECT 982.950 493.950 985.050 496.050 ;
        RECT 982.950 487.950 985.050 490.050 ;
        RECT 191.100 445.950 193.200 448.050 ;
        RECT 208.950 445.950 211.050 448.050 ;
        RECT 203.550 435.600 205.650 437.700 ;
        RECT 227.100 445.950 229.200 448.050 ;
        RECT 244.950 445.950 247.050 448.050 ;
        RECT 523.950 445.950 526.050 448.050 ;
        RECT 239.550 435.600 241.650 437.700 ;
        RECT 541.800 445.950 543.900 448.050 ;
        RECT 559.950 445.950 562.050 448.050 ;
        RECT 577.800 445.950 579.900 448.050 ;
        RECT 961.950 442.950 964.050 445.050 ;
        RECT 26.550 423.300 28.650 425.400 ;
        RECT 62.550 423.300 64.650 425.400 ;
        RECT 122.550 423.300 124.650 425.400 ;
        RECT 332.550 423.300 334.650 425.400 ;
        RECT 368.550 423.300 370.650 425.400 ;
        RECT 571.950 412.950 574.050 415.050 ;
        RECT 559.950 409.950 562.050 412.050 ;
        RECT 919.950 415.950 922.050 418.050 ;
        RECT 943.950 415.950 946.050 418.050 ;
        RECT 919.950 409.950 922.050 412.050 ;
        RECT 943.950 409.950 946.050 412.050 ;
        RECT 80.100 367.950 82.200 370.050 ;
        RECT 97.950 367.950 100.050 370.050 ;
        RECT 92.550 357.600 94.650 359.700 ;
        RECT 200.100 367.950 202.200 370.050 ;
        RECT 217.950 367.950 220.050 370.050 ;
        RECT 212.550 357.600 214.650 359.700 ;
        RECT 302.100 367.950 304.200 370.050 ;
        RECT 319.950 367.950 322.050 370.050 ;
        RECT 358.950 370.950 361.050 373.050 ;
        RECT 463.950 367.950 466.050 370.050 ;
        RECT 358.950 364.950 361.050 367.050 ;
        RECT 314.550 357.600 316.650 359.700 ;
        RECT 481.800 367.950 483.900 370.050 ;
        RECT 509.100 367.950 511.200 370.050 ;
        RECT 526.950 367.950 529.050 370.050 ;
        RECT 871.950 376.950 874.050 379.050 ;
        RECT 889.950 370.950 892.050 373.050 ;
        RECT 592.500 367.950 594.600 370.050 ;
        RECT 521.550 357.600 523.650 359.700 ;
        RECT 913.950 370.950 916.050 373.050 ;
        RECT 988.950 370.950 991.050 373.050 ;
        RECT 913.950 364.950 916.050 367.050 ;
        RECT 988.950 364.950 991.050 367.050 ;
        RECT 119.550 345.300 121.650 347.400 ;
        RECT 362.550 345.300 364.650 347.400 ;
        RECT 599.550 345.300 601.650 347.400 ;
        RECT 874.950 346.950 877.050 349.050 ;
        RECT 898.950 337.950 901.050 340.050 ;
        RECT 772.950 331.950 775.050 334.050 ;
        RECT 919.950 331.950 922.050 334.050 ;
        RECT 35.100 289.950 37.200 292.050 ;
        RECT 52.950 289.950 55.050 292.050 ;
        RECT 47.550 279.600 49.650 281.700 ;
        RECT 284.100 289.950 286.200 292.050 ;
        RECT 301.950 289.950 304.050 292.050 ;
        RECT 355.950 289.950 358.050 292.050 ;
        RECT 296.550 279.600 298.650 281.700 ;
        RECT 373.800 289.950 375.900 292.050 ;
        RECT 401.100 289.950 403.200 292.050 ;
        RECT 475.950 292.950 478.050 295.050 ;
        RECT 418.950 289.950 421.050 292.050 ;
        RECT 413.550 279.600 415.650 281.700 ;
        RECT 511.950 289.950 514.050 292.050 ;
        RECT 529.800 289.950 531.900 292.050 ;
        RECT 568.950 289.950 571.050 292.050 ;
        RECT 586.800 289.950 588.900 292.050 ;
        RECT 74.550 267.300 76.650 269.400 ;
        RECT 329.550 267.300 331.650 269.400 ;
        RECT 421.950 259.950 424.050 262.050 ;
        RECT 421.950 253.950 424.050 256.050 ;
        RECT 482.550 267.300 484.650 269.400 ;
        RECT 550.950 253.950 553.050 256.050 ;
        RECT 709.950 250.950 712.050 253.050 ;
        RECT 320.100 211.950 322.200 214.050 ;
        RECT 337.950 211.950 340.050 214.050 ;
        RECT 332.550 201.600 334.650 203.700 ;
        RECT 401.100 211.950 403.200 214.050 ;
        RECT 418.950 211.950 421.050 214.050 ;
        RECT 451.950 211.950 454.050 214.050 ;
        RECT 413.550 201.600 415.650 203.700 ;
        RECT 469.800 211.950 471.900 214.050 ;
        RECT 697.950 226.950 700.050 229.050 ;
        RECT 967.950 208.950 970.050 211.050 ;
        RECT 655.950 178.950 658.050 181.050 ;
        RECT 506.100 133.950 508.200 136.050 ;
        RECT 523.950 133.950 526.050 136.050 ;
        RECT 518.550 123.600 520.650 125.700 ;
        RECT 955.500 127.800 957.600 129.900 ;
        RECT 967.800 133.950 969.900 136.050 ;
        RECT 622.950 97.950 625.050 100.050 ;
        RECT 646.950 91.950 649.050 94.050 ;
        RECT 733.800 59.700 735.900 61.800 ;
        RECT 736.800 50.100 738.900 52.200 ;
        RECT 214.950 19.950 217.050 22.050 ;
        RECT 667.950 28.950 670.050 31.050 ;
      LAYER metal2 ;
        RECT 79.950 973.950 82.050 976.050 ;
        RECT 190.950 973.950 193.050 976.050 ;
        RECT 349.950 973.950 352.050 976.050 ;
        RECT 553.950 973.950 556.050 976.050 ;
        RECT 595.950 973.950 598.050 976.050 ;
        RECT 835.950 973.950 838.050 976.050 ;
        RECT 919.950 973.950 922.050 976.050 ;
        RECT 25.950 967.950 28.050 970.050 ;
        RECT 16.950 962.100 19.050 964.200 ;
        RECT 17.400 961.350 18.600 962.100 ;
        RECT 14.100 958.950 16.200 961.050 ;
        RECT 17.400 958.950 19.500 961.050 ;
        RECT 22.800 958.950 24.900 961.050 ;
        RECT 14.400 957.450 15.600 958.650 ;
        RECT 11.400 956.400 15.600 957.450 ;
        RECT 23.400 956.400 24.600 958.650 ;
        RECT 11.400 955.050 12.450 956.400 ;
        RECT 10.950 952.950 13.050 955.050 ;
        RECT 11.400 904.050 12.450 952.950 ;
        RECT 23.400 949.050 24.450 956.400 ;
        RECT 22.950 946.950 25.050 949.050 ;
        RECT 19.950 917.100 22.050 919.200 ;
        RECT 26.400 918.600 27.450 967.950 ;
        RECT 31.950 962.100 34.050 964.200 ;
        RECT 40.950 962.100 43.050 964.200 ;
        RECT 32.400 919.200 33.450 962.100 ;
        RECT 41.400 961.350 42.600 962.100 ;
        RECT 55.950 961.950 58.050 964.050 ;
        RECT 64.950 962.100 67.050 964.200 ;
        RECT 80.400 964.050 81.450 973.950 ;
        RECT 85.950 967.950 88.050 970.050 ;
        RECT 37.950 958.950 40.050 961.050 ;
        RECT 40.950 958.950 43.050 961.050 ;
        RECT 43.950 958.950 46.050 961.050 ;
        RECT 38.400 956.400 39.600 958.650 ;
        RECT 44.400 957.000 45.600 958.650 ;
        RECT 56.400 957.900 57.450 961.950 ;
        RECT 65.400 961.350 66.600 962.100 ;
        RECT 79.950 961.950 82.050 964.050 ;
        RECT 86.400 963.600 87.450 967.950 ;
        RECT 86.400 961.350 87.600 963.600 ;
        RECT 91.950 962.100 94.050 964.200 ;
        RECT 109.950 962.100 112.050 964.200 ;
        RECT 92.400 961.350 93.600 962.100 ;
        RECT 110.400 961.350 111.600 962.100 ;
        RECT 118.950 961.950 121.050 964.050 ;
        RECT 128.400 963.450 129.600 963.600 ;
        RECT 122.400 962.400 129.600 963.450 ;
        RECT 61.950 958.950 64.050 961.050 ;
        RECT 64.950 958.950 67.050 961.050 ;
        RECT 67.950 958.950 70.050 961.050 ;
        RECT 82.950 958.950 85.050 961.050 ;
        RECT 85.950 958.950 88.050 961.050 ;
        RECT 88.950 958.950 91.050 961.050 ;
        RECT 91.950 958.950 94.050 961.050 ;
        RECT 109.950 958.950 112.050 961.050 ;
        RECT 112.950 958.950 115.050 961.050 ;
        RECT 62.400 957.900 63.600 958.650 ;
        RECT 68.400 957.900 69.600 958.650 ;
        RECT 83.400 957.900 84.600 958.650 ;
        RECT 20.400 916.350 21.600 917.100 ;
        RECT 26.400 916.350 27.600 918.600 ;
        RECT 31.950 917.100 34.050 919.200 ;
        RECT 38.400 919.050 39.450 956.400 ;
        RECT 43.950 952.950 46.050 957.000 ;
        RECT 55.950 955.800 58.050 957.900 ;
        RECT 61.950 955.800 64.050 957.900 ;
        RECT 67.950 955.800 70.050 957.900 ;
        RECT 82.950 955.800 85.050 957.900 ;
        RECT 89.400 956.400 90.600 958.650 ;
        RECT 113.400 957.900 114.600 958.650 ;
        RECT 68.400 949.050 69.450 955.800 ;
        RECT 67.950 946.950 70.050 949.050 ;
        RECT 89.400 934.050 90.450 956.400 ;
        RECT 112.950 955.800 115.050 957.900 ;
        RECT 82.950 931.950 85.050 934.050 ;
        RECT 88.950 931.950 91.050 934.050 ;
        RECT 43.950 922.950 46.050 925.050 ;
        RECT 16.950 913.950 19.050 916.050 ;
        RECT 19.950 913.950 22.050 916.050 ;
        RECT 22.950 913.950 25.050 916.050 ;
        RECT 25.950 913.950 28.050 916.050 ;
        RECT 17.400 911.400 18.600 913.650 ;
        RECT 23.400 912.900 24.600 913.650 ;
        RECT 17.400 904.050 18.450 911.400 ;
        RECT 22.950 910.800 25.050 912.900 ;
        RECT 10.950 901.950 13.050 904.050 ;
        RECT 16.950 901.950 19.050 904.050 ;
        RECT 22.950 884.100 25.050 886.200 ;
        RECT 23.400 883.350 24.600 884.100 ;
        RECT 17.100 880.950 19.200 883.050 ;
        RECT 22.500 880.950 24.600 883.050 ;
        RECT 25.800 880.950 27.900 883.050 ;
        RECT 17.400 878.400 18.600 880.650 ;
        RECT 26.400 879.900 27.600 880.650 ;
        RECT 17.400 874.050 18.450 878.400 ;
        RECT 25.950 877.800 28.050 879.900 ;
        RECT 32.400 876.450 33.450 917.100 ;
        RECT 37.950 916.950 40.050 919.050 ;
        RECT 44.400 918.600 45.450 922.950 ;
        RECT 44.400 916.350 45.600 918.600 ;
        RECT 49.950 917.100 52.050 919.200 ;
        RECT 67.950 918.000 70.050 922.050 ;
        RECT 74.400 918.450 75.600 918.600 ;
        RECT 50.400 916.350 51.600 917.100 ;
        RECT 68.400 916.350 69.600 918.000 ;
        RECT 74.400 917.400 81.450 918.450 ;
        RECT 74.400 916.350 75.600 917.400 ;
        RECT 80.400 916.050 81.450 917.400 ;
        RECT 43.950 913.950 46.050 916.050 ;
        RECT 46.950 913.950 49.050 916.050 ;
        RECT 49.950 913.950 52.050 916.050 ;
        RECT 52.950 913.950 55.050 916.050 ;
        RECT 67.950 913.950 70.050 916.050 ;
        RECT 70.950 913.950 73.050 916.050 ;
        RECT 73.950 913.950 76.050 916.050 ;
        RECT 79.950 913.950 82.050 916.050 ;
        RECT 47.400 912.900 48.600 913.650 ;
        RECT 46.950 910.800 49.050 912.900 ;
        RECT 53.400 912.000 54.600 913.650 ;
        RECT 71.400 912.900 72.600 913.650 ;
        RECT 52.950 907.950 55.050 912.000 ;
        RECT 70.950 910.800 73.050 912.900 ;
        RECT 52.950 901.950 55.050 904.050 ;
        RECT 34.950 884.100 37.050 886.200 ;
        RECT 43.950 884.100 46.050 886.200 ;
        RECT 35.400 879.450 36.450 884.100 ;
        RECT 44.400 883.350 45.600 884.100 ;
        RECT 40.950 880.950 43.050 883.050 ;
        RECT 43.950 880.950 46.050 883.050 ;
        RECT 46.950 880.950 49.050 883.050 ;
        RECT 41.400 879.450 42.600 880.650 ;
        RECT 47.400 879.900 48.600 880.650 ;
        RECT 35.400 878.400 42.600 879.450 ;
        RECT 32.400 875.400 36.450 876.450 ;
        RECT 16.950 871.950 19.050 874.050 ;
        RECT 19.800 844.500 21.900 846.600 ;
        RECT 17.100 835.950 19.200 838.050 ;
        RECT 20.100 837.300 21.300 844.500 ;
        RECT 23.400 841.350 24.600 843.600 ;
        RECT 29.400 843.300 31.500 845.400 ;
        RECT 35.400 844.050 36.450 875.400 ;
        RECT 23.100 838.950 25.200 841.050 ;
        RECT 26.100 839.700 28.200 841.800 ;
        RECT 26.100 837.300 27.000 839.700 ;
        RECT 20.100 836.100 27.000 837.300 ;
        RECT 17.400 834.900 18.600 835.650 ;
        RECT 7.950 832.800 10.050 834.900 ;
        RECT 16.950 832.800 19.050 834.900 ;
        RECT 8.400 802.050 9.450 832.800 ;
        RECT 20.100 830.700 21.000 836.100 ;
        RECT 21.900 834.300 24.000 835.200 ;
        RECT 29.700 834.300 30.600 843.300 ;
        RECT 34.950 841.950 37.050 844.050 ;
        RECT 32.400 840.450 33.600 840.600 ;
        RECT 32.400 839.400 36.450 840.450 ;
        RECT 32.400 838.350 33.600 839.400 ;
        RECT 31.800 835.950 33.900 838.050 ;
        RECT 21.900 833.100 30.600 834.300 ;
        RECT 19.800 828.600 21.900 830.700 ;
        RECT 23.100 830.100 25.200 832.200 ;
        RECT 27.000 831.300 29.100 833.100 ;
        RECT 31.950 829.950 34.050 832.050 ;
        RECT 23.400 829.050 24.600 829.800 ;
        RECT 22.950 826.950 25.050 829.050 ;
        RECT 28.350 813.300 30.450 815.400 ;
        RECT 16.950 806.100 19.050 808.200 ;
        RECT 22.950 806.100 25.050 808.200 ;
        RECT 17.400 805.350 18.600 806.100 ;
        RECT 23.400 805.350 24.600 806.100 ;
        RECT 13.950 802.950 16.050 805.050 ;
        RECT 16.950 802.950 19.050 805.050 ;
        RECT 22.950 802.950 25.050 805.050 ;
        RECT 7.950 799.950 10.050 802.050 ;
        RECT 14.400 801.900 15.600 802.650 ;
        RECT 13.950 801.450 16.050 801.900 ;
        RECT 11.400 800.400 16.050 801.450 ;
        RECT 29.250 800.400 30.450 813.300 ;
        RECT 32.400 808.050 33.450 829.950 ;
        RECT 35.400 826.050 36.450 839.400 ;
        RECT 34.950 823.950 37.050 826.050 ;
        RECT 38.400 822.450 39.450 878.400 ;
        RECT 46.950 877.800 49.050 879.900 ;
        RECT 47.400 856.050 48.450 877.800 ;
        RECT 53.400 859.050 54.450 901.950 ;
        RECT 80.400 898.050 81.450 913.950 ;
        RECT 83.400 913.050 84.450 931.950 ;
        RECT 88.950 925.950 91.050 928.050 ;
        RECT 89.400 918.600 90.450 925.950 ;
        RECT 109.950 922.950 112.050 925.050 ;
        RECT 97.950 919.950 100.050 922.050 ;
        RECT 89.400 916.350 90.600 918.600 ;
        RECT 88.950 913.950 91.050 916.050 ;
        RECT 91.950 913.950 94.050 916.050 ;
        RECT 82.950 910.950 85.050 913.050 ;
        RECT 92.400 912.900 93.600 913.650 ;
        RECT 91.950 910.800 94.050 912.900 ;
        RECT 79.950 895.950 82.050 898.050 ;
        RECT 85.950 895.950 88.050 898.050 ;
        RECT 64.950 889.950 67.050 892.050 ;
        RECT 76.950 889.950 79.050 892.050 ;
        RECT 55.950 883.950 58.050 886.050 ;
        RECT 65.400 885.600 66.450 889.950 ;
        RECT 56.400 879.900 57.450 883.950 ;
        RECT 65.400 883.350 66.600 885.600 ;
        RECT 61.950 880.950 64.050 883.050 ;
        RECT 64.950 880.950 67.050 883.050 ;
        RECT 67.950 880.950 70.050 883.050 ;
        RECT 62.400 879.900 63.600 880.650 ;
        RECT 55.950 877.800 58.050 879.900 ;
        RECT 61.950 877.800 64.050 879.900 ;
        RECT 68.400 878.400 69.600 880.650 ;
        RECT 77.400 879.900 78.450 889.950 ;
        RECT 86.400 885.600 87.450 895.950 ;
        RECT 98.400 895.050 99.450 919.950 ;
        RECT 110.400 918.600 111.450 922.950 ;
        RECT 119.400 921.450 120.450 961.950 ;
        RECT 122.400 928.050 123.450 962.400 ;
        RECT 128.400 961.350 129.600 962.400 ;
        RECT 133.950 962.100 136.050 964.200 ;
        RECT 134.400 961.350 135.600 962.100 ;
        RECT 142.950 961.950 145.050 964.050 ;
        RECT 154.950 962.100 157.050 964.200 ;
        RECT 172.950 962.100 175.050 964.200 ;
        RECT 191.400 963.600 192.450 973.950 ;
        RECT 208.950 967.950 211.050 970.050 ;
        RECT 220.950 967.950 223.050 970.050 ;
        RECT 226.950 967.950 229.050 970.050 ;
        RECT 259.950 967.950 262.050 970.050 ;
        RECT 127.950 958.950 130.050 961.050 ;
        RECT 130.950 958.950 133.050 961.050 ;
        RECT 133.950 958.950 136.050 961.050 ;
        RECT 136.950 958.950 139.050 961.050 ;
        RECT 131.400 957.900 132.600 958.650 ;
        RECT 130.950 955.800 133.050 957.900 ;
        RECT 137.400 957.000 138.600 958.650 ;
        RECT 136.950 952.950 139.050 957.000 ;
        RECT 121.950 925.950 124.050 928.050 ;
        RECT 139.950 925.950 142.050 928.050 ;
        RECT 127.950 922.950 130.050 925.050 ;
        RECT 116.400 920.400 120.450 921.450 ;
        RECT 116.400 919.200 117.450 920.400 ;
        RECT 110.400 916.350 111.600 918.600 ;
        RECT 115.950 917.100 118.050 919.200 ;
        RECT 116.400 916.350 117.600 917.100 ;
        RECT 109.950 913.950 112.050 916.050 ;
        RECT 112.950 913.950 115.050 916.050 ;
        RECT 115.950 913.950 118.050 916.050 ;
        RECT 118.950 913.950 121.050 916.050 ;
        RECT 113.400 912.900 114.600 913.650 ;
        RECT 112.950 910.800 115.050 912.900 ;
        RECT 119.400 911.400 120.600 913.650 ;
        RECT 128.400 912.900 129.450 922.950 ;
        RECT 133.950 917.100 136.050 919.200 ;
        RECT 140.400 918.600 141.450 925.950 ;
        RECT 143.400 925.050 144.450 961.950 ;
        RECT 155.400 961.350 156.600 962.100 ;
        RECT 173.400 961.350 174.600 962.100 ;
        RECT 191.400 961.350 192.600 963.600 ;
        RECT 199.950 961.950 202.050 964.050 ;
        RECT 209.400 963.600 210.450 967.950 ;
        RECT 151.950 958.950 154.050 961.050 ;
        RECT 154.950 958.950 157.050 961.050 ;
        RECT 169.950 958.950 172.050 961.050 ;
        RECT 172.950 958.950 175.050 961.050 ;
        RECT 175.950 958.950 178.050 961.050 ;
        RECT 190.950 958.950 193.050 961.050 ;
        RECT 193.950 958.950 196.050 961.050 ;
        RECT 152.400 957.000 153.600 958.650 ;
        RECT 151.950 952.950 154.050 957.000 ;
        RECT 157.950 955.950 160.050 958.050 ;
        RECT 170.400 956.400 171.600 958.650 ;
        RECT 176.400 957.000 177.600 958.650 ;
        RECT 194.400 957.900 195.600 958.650 ;
        RECT 158.400 931.050 159.450 955.950 ;
        RECT 170.400 952.050 171.450 956.400 ;
        RECT 175.950 952.950 178.050 957.000 ;
        RECT 193.950 955.800 196.050 957.900 ;
        RECT 200.400 955.050 201.450 961.950 ;
        RECT 209.400 961.350 210.600 963.600 ;
        RECT 214.950 962.100 217.050 964.200 ;
        RECT 221.400 964.050 222.450 967.950 ;
        RECT 215.400 961.350 216.600 962.100 ;
        RECT 220.950 961.950 223.050 964.050 ;
        RECT 208.950 958.950 211.050 961.050 ;
        RECT 211.950 958.950 214.050 961.050 ;
        RECT 214.950 958.950 217.050 961.050 ;
        RECT 217.950 958.950 220.050 961.050 ;
        RECT 212.400 957.900 213.600 958.650 ;
        RECT 218.400 957.900 219.600 958.650 ;
        RECT 227.400 957.900 228.450 967.950 ;
        RECT 229.950 961.950 232.050 964.050 ;
        RECT 235.950 962.100 238.050 964.200 ;
        RECT 241.950 962.100 244.050 964.200 ;
        RECT 250.950 962.100 253.050 964.200 ;
        RECT 260.400 963.600 261.450 967.950 ;
        RECT 211.950 955.800 214.050 957.900 ;
        RECT 217.950 955.800 220.050 957.900 ;
        RECT 226.950 955.800 229.050 957.900 ;
        RECT 230.400 955.050 231.450 961.950 ;
        RECT 236.400 961.350 237.600 962.100 ;
        RECT 242.400 961.350 243.600 962.100 ;
        RECT 235.950 958.950 238.050 961.050 ;
        RECT 238.950 958.950 241.050 961.050 ;
        RECT 241.950 958.950 244.050 961.050 ;
        RECT 244.950 958.950 247.050 961.050 ;
        RECT 239.400 956.400 240.600 958.650 ;
        RECT 245.400 957.900 246.600 958.650 ;
        RECT 199.950 952.950 202.050 955.050 ;
        RECT 229.950 952.950 232.050 955.050 ;
        RECT 169.950 949.950 172.050 952.050 ;
        RECT 239.400 943.050 240.450 956.400 ;
        RECT 244.950 955.800 247.050 957.900 ;
        RECT 251.400 952.050 252.450 962.100 ;
        RECT 260.400 961.350 261.600 963.600 ;
        RECT 265.950 962.100 268.050 964.200 ;
        RECT 274.950 962.100 277.050 964.200 ;
        RECT 286.950 962.100 289.050 964.200 ;
        RECT 292.950 962.100 295.050 964.200 ;
        RECT 266.400 961.350 267.600 962.100 ;
        RECT 259.950 958.950 262.050 961.050 ;
        RECT 262.950 958.950 265.050 961.050 ;
        RECT 265.950 958.950 268.050 961.050 ;
        RECT 268.950 958.950 271.050 961.050 ;
        RECT 253.950 955.800 256.050 957.900 ;
        RECT 263.400 956.400 264.600 958.650 ;
        RECT 269.400 957.900 270.600 958.650 ;
        RECT 250.950 949.950 253.050 952.050 ;
        RECT 238.950 940.950 241.050 943.050 ;
        RECT 220.950 934.950 223.050 937.050 ;
        RECT 157.950 928.950 160.050 931.050 ;
        RECT 184.950 928.950 187.050 931.050 ;
        RECT 193.950 928.950 196.050 931.050 ;
        RECT 142.950 922.950 145.050 925.050 ;
        RECT 134.400 916.350 135.600 917.100 ;
        RECT 140.400 916.350 141.600 918.600 ;
        RECT 151.950 917.100 154.050 919.200 ;
        RECT 158.400 918.600 159.450 928.950 ;
        RECT 178.950 925.950 181.050 928.050 ;
        RECT 133.950 913.950 136.050 916.050 ;
        RECT 136.950 913.950 139.050 916.050 ;
        RECT 139.950 913.950 142.050 916.050 ;
        RECT 142.950 913.950 145.050 916.050 ;
        RECT 137.400 912.900 138.600 913.650 ;
        RECT 119.400 910.050 120.450 911.400 ;
        RECT 127.950 910.800 130.050 912.900 ;
        RECT 136.950 910.800 139.050 912.900 ;
        RECT 143.400 912.450 144.600 913.650 ;
        RECT 143.400 911.400 147.450 912.450 ;
        RECT 119.400 908.400 124.050 910.050 ;
        RECT 120.000 907.950 124.050 908.400 ;
        RECT 139.950 907.950 145.050 910.050 ;
        RECT 97.950 892.950 100.050 895.050 ;
        RECT 124.950 892.950 127.050 895.050 ;
        RECT 86.400 883.350 87.600 885.600 ;
        RECT 91.950 884.100 94.050 886.200 ;
        RECT 92.400 883.350 93.600 884.100 ;
        RECT 82.950 880.950 85.050 883.050 ;
        RECT 85.950 880.950 88.050 883.050 ;
        RECT 88.950 880.950 91.050 883.050 ;
        RECT 91.950 880.950 94.050 883.050 ;
        RECT 83.400 879.900 84.600 880.650 ;
        RECT 68.400 874.050 69.450 878.400 ;
        RECT 76.950 877.800 79.050 879.900 ;
        RECT 82.950 877.800 85.050 879.900 ;
        RECT 89.400 878.400 90.600 880.650 ;
        RECT 89.400 874.050 90.450 878.400 ;
        RECT 67.950 871.950 70.050 874.050 ;
        RECT 88.950 871.950 91.050 874.050 ;
        RECT 52.950 856.950 55.050 859.050 ;
        RECT 40.950 853.950 43.050 856.050 ;
        RECT 46.950 853.950 49.050 856.050 ;
        RECT 41.400 835.050 42.450 853.950 ;
        RECT 68.400 850.050 69.450 871.950 ;
        RECT 61.950 847.950 64.050 850.050 ;
        RECT 67.950 847.950 70.050 850.050 ;
        RECT 91.950 847.950 94.050 850.050 ;
        RECT 46.950 839.100 49.050 841.200 ;
        RECT 53.400 840.450 54.600 840.600 ;
        RECT 53.400 839.400 60.450 840.450 ;
        RECT 47.400 838.350 48.600 839.100 ;
        RECT 53.400 838.350 54.600 839.400 ;
        RECT 46.950 835.950 49.050 838.050 ;
        RECT 49.950 835.950 52.050 838.050 ;
        RECT 52.950 835.950 55.050 838.050 ;
        RECT 40.950 832.950 43.050 835.050 ;
        RECT 50.400 834.900 51.600 835.650 ;
        RECT 49.950 832.800 52.050 834.900 ;
        RECT 59.400 826.050 60.450 839.400 ;
        RECT 62.400 834.900 63.450 847.950 ;
        RECT 67.950 840.000 70.050 844.050 ;
        RECT 68.400 838.350 69.600 840.000 ;
        RECT 73.950 839.100 76.050 841.200 ;
        RECT 82.950 839.100 85.050 841.200 ;
        RECT 92.400 840.600 93.450 847.950 ;
        RECT 98.400 844.050 99.450 892.950 ;
        RECT 106.950 889.950 109.050 892.050 ;
        RECT 107.400 885.600 108.450 889.950 ;
        RECT 118.950 886.950 121.050 889.050 ;
        RECT 107.400 883.350 108.600 885.600 ;
        RECT 106.950 880.950 109.050 883.050 ;
        RECT 109.950 880.950 112.050 883.050 ;
        RECT 110.400 879.900 111.600 880.650 ;
        RECT 119.400 880.050 120.450 886.950 ;
        RECT 125.400 885.600 126.450 892.950 ;
        RECT 125.400 883.350 126.600 885.600 ;
        RECT 130.950 885.000 133.050 889.050 ;
        RECT 131.400 883.350 132.600 885.000 ;
        RECT 124.950 880.950 127.050 883.050 ;
        RECT 127.950 880.950 130.050 883.050 ;
        RECT 130.950 880.950 133.050 883.050 ;
        RECT 133.950 880.950 136.050 883.050 ;
        RECT 109.950 877.800 112.050 879.900 ;
        RECT 118.950 877.950 121.050 880.050 ;
        RECT 128.400 879.900 129.600 880.650 ;
        RECT 127.950 877.800 130.050 879.900 ;
        RECT 134.400 879.000 135.600 880.650 ;
        RECT 124.950 874.950 127.050 877.050 ;
        RECT 133.950 874.950 136.050 879.000 ;
        RECT 142.950 874.950 145.050 877.050 ;
        RECT 115.950 871.950 118.050 874.050 ;
        RECT 97.950 841.950 100.050 844.050 ;
        RECT 98.400 840.600 99.450 841.950 ;
        RECT 116.400 841.200 117.450 871.950 ;
        RECT 74.400 838.350 75.600 839.100 ;
        RECT 67.950 835.950 70.050 838.050 ;
        RECT 70.950 835.950 73.050 838.050 ;
        RECT 73.950 835.950 76.050 838.050 ;
        RECT 76.950 835.950 79.050 838.050 ;
        RECT 71.400 834.900 72.600 835.650 ;
        RECT 61.950 832.800 64.050 834.900 ;
        RECT 70.950 832.800 73.050 834.900 ;
        RECT 77.400 833.400 78.600 835.650 ;
        RECT 77.400 832.050 78.450 833.400 ;
        RECT 76.950 829.950 79.050 832.050 ;
        RECT 58.950 823.950 61.050 826.050 ;
        RECT 35.400 821.400 39.450 822.450 ;
        RECT 31.950 805.950 34.050 808.050 ;
        RECT 7.950 763.950 10.050 766.050 ;
        RECT 8.400 706.050 9.450 763.950 ;
        RECT 11.400 763.050 12.450 800.400 ;
        RECT 13.950 799.800 16.050 800.400 ;
        RECT 28.350 798.300 30.450 800.400 ;
        RECT 31.950 799.800 34.050 801.900 ;
        RECT 29.250 791.700 30.450 798.300 ;
        RECT 28.350 789.600 30.450 791.700 ;
        RECT 16.950 769.950 19.050 772.050 ;
        RECT 17.400 766.050 18.450 769.950 ;
        RECT 10.950 760.950 13.050 763.050 ;
        RECT 16.950 762.000 19.050 766.050 ;
        RECT 17.400 760.350 18.600 762.000 ;
        RECT 22.950 761.100 25.050 763.200 ;
        RECT 28.950 761.100 31.050 763.200 ;
        RECT 23.400 760.350 24.600 761.100 ;
        RECT 13.950 757.950 16.050 760.050 ;
        RECT 16.950 757.950 19.050 760.050 ;
        RECT 19.950 757.950 22.050 760.050 ;
        RECT 22.950 757.950 25.050 760.050 ;
        RECT 14.400 756.900 15.600 757.650 ;
        RECT 20.400 756.900 21.600 757.650 ;
        RECT 13.950 754.800 16.050 756.900 ;
        RECT 19.950 754.800 22.050 756.900 ;
        RECT 16.950 751.950 19.050 754.050 ;
        RECT 17.400 729.600 18.450 751.950 ;
        RECT 25.950 748.950 28.050 751.050 ;
        RECT 17.400 727.350 18.600 729.600 ;
        RECT 13.950 724.950 16.050 727.050 ;
        RECT 16.950 724.950 19.050 727.050 ;
        RECT 19.950 724.950 22.050 727.050 ;
        RECT 20.400 722.400 21.600 724.650 ;
        RECT 20.400 706.050 21.450 722.400 ;
        RECT 7.950 703.950 10.050 706.050 ;
        RECT 19.950 703.950 22.050 706.050 ;
        RECT 26.400 697.050 27.450 748.950 ;
        RECT 29.400 715.050 30.450 761.100 ;
        RECT 32.400 757.050 33.450 799.800 ;
        RECT 35.400 790.050 36.450 821.400 ;
        RECT 46.050 813.300 48.150 815.400 ;
        RECT 40.800 802.950 42.900 805.050 ;
        RECT 41.400 801.900 42.600 802.650 ;
        RECT 40.950 799.800 43.050 801.900 ;
        RECT 46.650 794.700 47.850 813.300 ;
        RECT 74.400 807.450 75.600 807.600 ;
        RECT 77.400 807.450 78.450 829.950 ;
        RECT 79.950 822.450 82.050 823.050 ;
        RECT 83.400 822.450 84.450 839.100 ;
        RECT 92.400 838.350 93.600 840.600 ;
        RECT 98.400 838.350 99.600 840.600 ;
        RECT 109.950 838.950 112.050 841.050 ;
        RECT 115.950 839.100 118.050 841.200 ;
        RECT 91.950 835.950 94.050 838.050 ;
        RECT 94.950 835.950 97.050 838.050 ;
        RECT 97.950 835.950 100.050 838.050 ;
        RECT 100.950 835.950 103.050 838.050 ;
        RECT 95.400 833.400 96.600 835.650 ;
        RECT 101.400 833.400 102.600 835.650 ;
        RECT 95.400 823.050 96.450 833.400 ;
        RECT 79.950 821.400 84.450 822.450 ;
        RECT 79.950 820.950 82.050 821.400 ;
        RECT 94.950 820.950 97.050 823.050 ;
        RECT 74.400 806.400 78.450 807.450 ;
        RECT 74.400 805.350 75.600 806.400 ;
        RECT 49.950 802.950 52.050 805.050 ;
        RECT 70.950 802.950 73.050 805.050 ;
        RECT 73.950 802.950 76.050 805.050 ;
        RECT 43.650 793.500 47.850 794.700 ;
        RECT 50.400 800.400 51.600 802.650 ;
        RECT 71.400 800.400 72.600 802.650 ;
        RECT 43.650 792.600 45.750 793.500 ;
        RECT 34.950 787.950 37.050 790.050 ;
        RECT 43.950 787.950 46.050 790.050 ;
        RECT 34.950 778.950 37.050 781.050 ;
        RECT 31.950 754.950 34.050 757.050 ;
        RECT 35.400 754.050 36.450 778.950 ;
        RECT 44.400 762.600 45.450 787.950 ;
        RECT 50.400 787.050 51.450 800.400 ;
        RECT 71.400 799.050 72.450 800.400 ;
        RECT 71.400 797.400 76.050 799.050 ;
        RECT 72.000 796.950 76.050 797.400 ;
        RECT 80.400 795.450 81.450 820.950 ;
        RECT 101.400 811.050 102.450 833.400 ;
        RECT 91.950 807.000 94.050 811.050 ;
        RECT 100.950 808.950 103.050 811.050 ;
        RECT 98.400 807.450 99.600 807.600 ;
        RECT 92.400 805.350 93.600 807.000 ;
        RECT 98.400 806.400 105.450 807.450 ;
        RECT 98.400 805.350 99.600 806.400 ;
        RECT 88.950 802.950 91.050 805.050 ;
        RECT 91.950 802.950 94.050 805.050 ;
        RECT 94.950 802.950 97.050 805.050 ;
        RECT 97.950 802.950 100.050 805.050 ;
        RECT 89.400 801.900 90.600 802.650 ;
        RECT 88.950 799.800 91.050 801.900 ;
        RECT 95.400 801.000 96.600 802.650 ;
        RECT 94.950 796.950 97.050 801.000 ;
        RECT 104.400 796.050 105.450 806.400 ;
        RECT 110.400 801.900 111.450 838.950 ;
        RECT 116.400 838.350 117.600 839.100 ;
        RECT 115.950 835.950 118.050 838.050 ;
        RECT 118.950 835.950 121.050 838.050 ;
        RECT 119.400 834.450 120.600 835.650 ;
        RECT 125.400 834.450 126.450 874.950 ;
        RECT 136.950 839.100 139.050 841.200 ;
        RECT 143.400 840.600 144.450 874.950 ;
        RECT 137.400 838.350 138.600 839.100 ;
        RECT 143.400 838.350 144.600 840.600 ;
        RECT 146.400 840.450 147.450 911.400 ;
        RECT 152.400 910.050 153.450 917.100 ;
        RECT 158.400 916.350 159.600 918.600 ;
        RECT 163.950 917.100 166.050 919.200 ;
        RECT 179.400 918.600 180.450 925.950 ;
        RECT 185.400 918.600 186.450 928.950 ;
        RECT 164.400 916.350 165.600 917.100 ;
        RECT 179.400 916.350 180.600 918.600 ;
        RECT 185.400 916.350 186.600 918.600 ;
        RECT 157.950 913.950 160.050 916.050 ;
        RECT 160.950 913.950 163.050 916.050 ;
        RECT 163.950 913.950 166.050 916.050 ;
        RECT 178.950 913.950 181.050 916.050 ;
        RECT 181.950 913.950 184.050 916.050 ;
        RECT 184.950 913.950 187.050 916.050 ;
        RECT 187.950 913.950 190.050 916.050 ;
        RECT 161.400 911.400 162.600 913.650 ;
        RECT 182.400 912.000 183.600 913.650 ;
        RECT 151.950 907.950 154.050 910.050 ;
        RECT 161.400 907.050 162.450 911.400 ;
        RECT 181.950 907.950 184.050 912.000 ;
        RECT 188.400 911.400 189.600 913.650 ;
        RECT 160.950 904.950 163.050 907.050 ;
        RECT 157.950 889.950 160.050 892.050 ;
        RECT 184.950 889.950 187.050 892.050 ;
        RECT 158.400 885.600 159.450 889.950 ;
        RECT 158.400 883.350 159.600 885.600 ;
        RECT 163.950 884.100 166.050 886.200 ;
        RECT 172.950 884.100 175.050 886.200 ;
        RECT 178.950 884.100 181.050 886.200 ;
        RECT 185.400 885.600 186.450 889.950 ;
        RECT 152.100 880.950 154.200 883.050 ;
        RECT 157.500 880.950 159.600 883.050 ;
        RECT 160.800 880.950 162.900 883.050 ;
        RECT 152.400 879.900 153.600 880.650 ;
        RECT 151.950 877.800 154.050 879.900 ;
        RECT 161.400 878.400 162.600 880.650 ;
        RECT 164.400 880.050 165.450 884.100 ;
        RECT 161.400 871.050 162.450 878.400 ;
        RECT 163.950 877.950 166.050 880.050 ;
        RECT 173.400 871.050 174.450 884.100 ;
        RECT 179.400 883.350 180.600 884.100 ;
        RECT 185.400 883.350 186.600 885.600 ;
        RECT 188.400 885.450 189.450 911.400 ;
        RECT 194.400 907.050 195.450 928.950 ;
        RECT 205.950 922.950 208.050 925.050 ;
        RECT 206.400 918.600 207.450 922.950 ;
        RECT 206.400 916.350 207.600 918.600 ;
        RECT 211.950 917.100 214.050 919.200 ;
        RECT 217.950 917.100 220.050 919.200 ;
        RECT 212.400 916.350 213.600 917.100 ;
        RECT 202.950 913.950 205.050 916.050 ;
        RECT 205.950 913.950 208.050 916.050 ;
        RECT 208.950 913.950 211.050 916.050 ;
        RECT 211.950 913.950 214.050 916.050 ;
        RECT 203.400 911.400 204.600 913.650 ;
        RECT 209.400 912.900 210.600 913.650 ;
        RECT 193.950 904.950 196.050 907.050 ;
        RECT 203.400 901.050 204.450 911.400 ;
        RECT 208.950 910.800 211.050 912.900 ;
        RECT 202.950 898.950 205.050 901.050 ;
        RECT 218.400 892.050 219.450 917.100 ;
        RECT 221.400 913.050 222.450 934.950 ;
        RECT 254.400 934.050 255.450 955.800 ;
        RECT 263.400 955.050 264.450 956.400 ;
        RECT 268.950 955.800 271.050 957.900 ;
        RECT 262.950 952.950 265.050 955.050 ;
        RECT 259.950 940.950 262.050 943.050 ;
        RECT 253.950 931.950 256.050 934.050 ;
        RECT 235.950 928.950 238.050 931.050 ;
        RECT 250.950 928.950 253.050 931.050 ;
        RECT 236.400 925.050 237.450 928.950 ;
        RECT 238.950 925.950 244.050 928.050 ;
        RECT 244.950 925.950 250.050 928.050 ;
        RECT 251.400 925.050 252.450 928.950 ;
        RECT 260.400 925.050 261.450 940.950 ;
        RECT 263.400 937.050 264.450 952.950 ;
        RECT 275.400 946.050 276.450 962.100 ;
        RECT 287.400 961.350 288.600 962.100 ;
        RECT 293.400 961.350 294.600 962.100 ;
        RECT 304.950 961.950 307.050 964.050 ;
        RECT 313.950 962.100 316.050 964.200 ;
        RECT 319.950 962.100 322.050 964.200 ;
        RECT 334.950 962.100 337.050 964.200 ;
        RECT 340.950 962.100 343.050 964.200 ;
        RECT 283.950 958.950 286.050 961.050 ;
        RECT 286.950 958.950 289.050 961.050 ;
        RECT 289.950 958.950 292.050 961.050 ;
        RECT 292.950 958.950 295.050 961.050 ;
        RECT 301.950 958.950 304.050 961.050 ;
        RECT 284.400 957.000 285.600 958.650 ;
        RECT 290.400 957.900 291.600 958.650 ;
        RECT 283.950 952.950 286.050 957.000 ;
        RECT 289.950 955.800 292.050 957.900 ;
        RECT 295.950 952.950 298.050 957.900 ;
        RECT 302.400 952.050 303.450 958.950 ;
        RECT 289.950 949.950 292.050 952.050 ;
        RECT 301.950 949.950 304.050 952.050 ;
        RECT 265.950 943.950 268.050 946.050 ;
        RECT 274.950 943.950 277.050 946.050 ;
        RECT 262.950 934.950 265.050 937.050 ;
        RECT 229.950 922.950 232.050 925.050 ;
        RECT 235.950 922.950 238.050 925.050 ;
        RECT 249.000 924.900 252.450 925.050 ;
        RECT 230.400 918.600 231.450 922.950 ;
        RECT 241.950 922.800 244.050 924.900 ;
        RECT 247.950 923.400 252.450 924.900 ;
        RECT 247.950 922.950 252.000 923.400 ;
        RECT 259.950 922.950 262.050 925.050 ;
        RECT 247.950 922.800 250.050 922.950 ;
        RECT 230.400 916.350 231.600 918.600 ;
        RECT 235.950 917.100 238.050 919.200 ;
        RECT 236.400 916.350 237.600 917.100 ;
        RECT 226.950 913.950 229.050 916.050 ;
        RECT 229.950 913.950 232.050 916.050 ;
        RECT 232.950 913.950 235.050 916.050 ;
        RECT 235.950 913.950 238.050 916.050 ;
        RECT 220.950 910.950 223.050 913.050 ;
        RECT 227.400 911.400 228.600 913.650 ;
        RECT 233.400 912.900 234.600 913.650 ;
        RECT 227.400 901.050 228.450 911.400 ;
        RECT 232.950 910.800 235.050 912.900 ;
        RECT 226.950 898.950 229.050 901.050 ;
        RECT 211.950 889.950 217.050 892.050 ;
        RECT 217.950 889.950 220.050 892.050 ;
        RECT 220.950 886.950 223.050 892.050 ;
        RECT 188.400 884.400 192.450 885.450 ;
        RECT 178.950 880.950 181.050 883.050 ;
        RECT 181.950 880.950 184.050 883.050 ;
        RECT 184.950 880.950 187.050 883.050 ;
        RECT 182.400 879.900 183.600 880.650 ;
        RECT 181.950 877.800 184.050 879.900 ;
        RECT 160.950 868.950 163.050 871.050 ;
        RECT 172.950 868.950 175.050 871.050 ;
        RECT 191.400 855.450 192.450 884.400 ;
        RECT 193.950 883.950 196.050 886.050 ;
        RECT 202.950 884.100 205.050 886.200 ;
        RECT 210.000 885.600 214.050 886.050 ;
        RECT 194.400 877.050 195.450 883.950 ;
        RECT 203.400 883.350 204.600 884.100 ;
        RECT 209.400 883.950 214.050 885.600 ;
        RECT 209.400 883.350 210.600 883.950 ;
        RECT 220.950 883.800 223.050 885.900 ;
        RECT 199.950 880.950 202.050 883.050 ;
        RECT 202.950 880.950 205.050 883.050 ;
        RECT 205.950 880.950 208.050 883.050 ;
        RECT 208.950 880.950 211.050 883.050 ;
        RECT 200.400 878.400 201.600 880.650 ;
        RECT 206.400 879.900 207.600 880.650 ;
        RECT 193.950 874.950 196.050 877.050 ;
        RECT 200.400 871.050 201.450 878.400 ;
        RECT 205.950 877.800 208.050 879.900 ;
        RECT 221.400 871.050 222.450 883.800 ;
        RECT 227.400 880.050 228.450 898.950 ;
        RECT 242.400 898.050 243.450 922.800 ;
        RECT 250.950 917.100 253.050 919.200 ;
        RECT 251.400 916.350 252.600 917.100 ;
        RECT 250.950 913.950 253.050 916.050 ;
        RECT 253.950 913.950 256.050 916.050 ;
        RECT 254.400 911.400 255.600 913.650 ;
        RECT 260.400 913.050 261.450 922.950 ;
        RECT 262.950 916.950 265.050 919.050 ;
        RECT 241.950 895.950 244.050 898.050 ;
        RECT 254.400 895.050 255.450 911.400 ;
        RECT 259.950 910.950 262.050 913.050 ;
        RECT 263.400 910.050 264.450 916.950 ;
        RECT 266.400 913.050 267.450 943.950 ;
        RECT 274.950 917.100 277.050 919.200 ;
        RECT 281.400 918.450 282.600 918.600 ;
        RECT 281.400 917.400 288.450 918.450 ;
        RECT 275.400 916.350 276.600 917.100 ;
        RECT 281.400 916.350 282.600 917.400 ;
        RECT 271.950 913.950 274.050 916.050 ;
        RECT 274.950 913.950 277.050 916.050 ;
        RECT 277.950 913.950 280.050 916.050 ;
        RECT 280.950 913.950 283.050 916.050 ;
        RECT 265.950 910.950 268.050 913.050 ;
        RECT 272.400 912.900 273.600 913.650 ;
        RECT 271.950 910.800 274.050 912.900 ;
        RECT 278.400 912.000 279.600 913.650 ;
        RECT 262.950 907.950 265.050 910.050 ;
        RECT 277.950 907.950 280.050 912.000 ;
        RECT 287.400 901.050 288.450 917.400 ;
        RECT 290.400 913.050 291.450 949.950 ;
        RECT 305.400 949.050 306.450 961.950 ;
        RECT 314.400 961.350 315.600 962.100 ;
        RECT 320.400 961.350 321.600 962.100 ;
        RECT 335.400 961.350 336.600 962.100 ;
        RECT 341.400 961.350 342.600 962.100 ;
        RECT 310.950 958.950 313.050 961.050 ;
        RECT 313.950 958.950 316.050 961.050 ;
        RECT 316.950 958.950 319.050 961.050 ;
        RECT 319.950 958.950 322.050 961.050 ;
        RECT 334.950 958.950 337.050 961.050 ;
        RECT 337.950 958.950 340.050 961.050 ;
        RECT 340.950 958.950 343.050 961.050 ;
        RECT 343.950 958.950 346.050 961.050 ;
        RECT 311.400 956.400 312.600 958.650 ;
        RECT 317.400 957.900 318.600 958.650 ;
        RECT 338.400 957.900 339.600 958.650 ;
        RECT 344.400 957.900 345.600 958.650 ;
        RECT 304.950 946.950 307.050 949.050 ;
        RECT 311.400 925.050 312.450 956.400 ;
        RECT 316.950 955.800 319.050 957.900 ;
        RECT 325.950 955.800 328.050 957.900 ;
        RECT 331.950 955.800 334.050 957.900 ;
        RECT 337.950 955.800 340.050 957.900 ;
        RECT 343.800 955.800 345.900 957.900 ;
        RECT 316.950 954.300 319.050 954.750 ;
        RECT 322.950 954.300 325.050 954.750 ;
        RECT 316.950 953.250 325.050 954.300 ;
        RECT 316.950 952.650 319.050 953.250 ;
        RECT 322.950 952.650 325.050 953.250 ;
        RECT 326.400 943.050 327.450 955.800 ;
        RECT 332.400 949.050 333.450 955.800 ;
        RECT 337.950 954.300 340.050 954.750 ;
        RECT 346.950 954.300 349.050 958.050 ;
        RECT 350.400 955.050 351.450 973.950 ;
        RECT 403.950 970.950 406.050 973.050 ;
        RECT 427.950 970.950 430.050 973.050 ;
        RECT 433.950 970.950 436.050 973.050 ;
        RECT 478.950 970.950 481.050 973.050 ;
        RECT 514.950 970.950 517.050 973.050 ;
        RECT 526.950 970.950 529.050 973.050 ;
        RECT 404.400 964.200 405.450 970.950 ;
        RECT 409.950 967.950 412.050 970.050 ;
        RECT 352.950 962.100 355.050 964.200 ;
        RECT 358.950 962.100 361.050 964.200 ;
        RECT 337.950 954.000 349.050 954.300 ;
        RECT 337.950 953.250 348.450 954.000 ;
        RECT 337.950 952.650 340.050 953.250 ;
        RECT 349.950 952.950 352.050 955.050 ;
        RECT 331.950 946.950 334.050 949.050 ;
        RECT 353.400 943.050 354.450 962.100 ;
        RECT 359.400 961.350 360.600 962.100 ;
        RECT 367.950 961.950 370.050 964.050 ;
        RECT 379.950 962.100 382.050 964.200 ;
        RECT 394.950 962.100 397.050 964.200 ;
        RECT 403.950 962.100 406.050 964.200 ;
        RECT 410.400 963.600 411.450 967.950 ;
        RECT 428.400 963.600 429.450 970.950 ;
        RECT 434.400 963.600 435.450 970.950 ;
        RECT 479.400 964.200 480.450 970.950 ;
        RECT 490.950 967.950 493.050 970.050 ;
        RECT 358.950 958.950 361.050 961.050 ;
        RECT 361.950 958.950 364.050 961.050 ;
        RECT 362.400 957.900 363.600 958.650 ;
        RECT 361.950 955.800 364.050 957.900 ;
        RECT 368.400 949.050 369.450 961.950 ;
        RECT 380.400 961.350 381.600 962.100 ;
        RECT 376.950 958.950 379.050 961.050 ;
        RECT 379.950 958.950 382.050 961.050 ;
        RECT 382.950 958.950 385.050 961.050 ;
        RECT 377.400 956.400 378.600 958.650 ;
        RECT 383.400 957.900 384.600 958.650 ;
        RECT 377.400 952.050 378.450 956.400 ;
        RECT 382.950 955.800 385.050 957.900 ;
        RECT 395.400 952.050 396.450 962.100 ;
        RECT 404.400 961.350 405.600 962.100 ;
        RECT 410.400 961.350 411.600 963.600 ;
        RECT 428.400 961.350 429.600 963.600 ;
        RECT 434.400 961.350 435.600 963.600 ;
        RECT 454.950 962.100 457.050 964.200 ;
        RECT 473.400 963.450 474.600 963.600 ;
        RECT 467.400 962.400 474.600 963.450 ;
        RECT 455.400 961.350 456.600 962.100 ;
        RECT 400.950 958.950 403.050 961.050 ;
        RECT 403.950 958.950 406.050 961.050 ;
        RECT 406.950 958.950 409.050 961.050 ;
        RECT 409.950 958.950 412.050 961.050 ;
        RECT 424.950 958.950 427.050 961.050 ;
        RECT 427.950 958.950 430.050 961.050 ;
        RECT 430.950 958.950 433.050 961.050 ;
        RECT 433.950 958.950 436.050 961.050 ;
        RECT 451.950 958.950 454.050 961.050 ;
        RECT 454.950 958.950 457.050 961.050 ;
        RECT 457.950 958.950 460.050 961.050 ;
        RECT 401.400 957.900 402.600 958.650 ;
        RECT 400.950 955.800 403.050 957.900 ;
        RECT 407.400 956.400 408.600 958.650 ;
        RECT 425.400 957.900 426.600 958.650 ;
        RECT 376.950 949.950 379.050 952.050 ;
        RECT 394.950 949.950 397.050 952.050 ;
        RECT 367.950 946.950 370.050 949.050 ;
        RECT 316.950 940.950 319.050 943.050 ;
        RECT 325.950 940.950 328.050 943.050 ;
        RECT 352.950 940.950 355.050 943.050 ;
        RECT 317.400 934.050 318.450 940.950 ;
        RECT 316.950 931.950 319.050 934.050 ;
        RECT 319.950 928.950 322.050 931.050 ;
        RECT 310.950 922.950 313.050 925.050 ;
        RECT 298.950 917.100 301.050 919.200 ;
        RECT 320.400 918.600 321.450 928.950 ;
        RECT 331.950 925.950 334.050 928.050 ;
        RECT 305.400 918.450 306.600 918.600 ;
        RECT 305.400 917.400 312.450 918.450 ;
        RECT 299.400 916.350 300.600 917.100 ;
        RECT 305.400 916.350 306.600 917.400 ;
        RECT 295.950 913.950 298.050 916.050 ;
        RECT 298.950 913.950 301.050 916.050 ;
        RECT 301.950 913.950 304.050 916.050 ;
        RECT 304.950 913.950 307.050 916.050 ;
        RECT 289.950 910.950 292.050 913.050 ;
        RECT 296.400 912.900 297.600 913.650 ;
        RECT 295.950 910.800 298.050 912.900 ;
        RECT 302.400 911.400 303.600 913.650 ;
        RECT 302.400 901.050 303.450 911.400 ;
        RECT 286.950 898.950 289.050 901.050 ;
        RECT 301.950 898.950 304.050 901.050 ;
        RECT 286.950 895.800 289.050 897.900 ;
        RECT 253.950 892.950 256.050 895.050 ;
        RECT 229.950 886.950 235.050 889.050 ;
        RECT 256.950 886.950 262.050 889.050 ;
        RECT 235.950 884.100 238.050 886.200 ;
        RECT 246.000 885.600 250.050 886.050 ;
        RECT 236.400 883.350 237.600 884.100 ;
        RECT 245.400 883.950 250.050 885.600 ;
        RECT 262.950 884.100 265.050 886.200 ;
        RECT 268.950 885.000 271.050 889.050 ;
        RECT 245.400 883.350 246.600 883.950 ;
        RECT 263.400 883.350 264.600 884.100 ;
        RECT 269.400 883.350 270.600 885.000 ;
        RECT 280.950 884.100 283.050 886.200 ;
        RECT 287.400 885.600 288.450 895.800 ;
        RECT 311.400 895.050 312.450 917.400 ;
        RECT 320.400 916.350 321.600 918.600 ;
        RECT 325.950 917.100 328.050 919.200 ;
        RECT 326.400 916.350 327.600 917.100 ;
        RECT 313.950 913.950 316.050 916.050 ;
        RECT 319.950 913.950 322.050 916.050 ;
        RECT 322.950 913.950 325.050 916.050 ;
        RECT 325.950 913.950 328.050 916.050 ;
        RECT 310.950 892.950 313.050 895.050 ;
        RECT 301.950 886.950 304.050 889.050 ;
        RECT 230.400 880.950 232.500 883.050 ;
        RECT 235.950 880.950 238.050 883.050 ;
        RECT 238.950 880.950 241.050 883.050 ;
        RECT 245.100 880.950 247.200 883.050 ;
        RECT 262.950 880.950 265.050 883.050 ;
        RECT 265.950 880.950 268.050 883.050 ;
        RECT 268.950 880.950 271.050 883.050 ;
        RECT 271.950 880.950 274.050 883.050 ;
        RECT 226.950 877.950 229.050 880.050 ;
        RECT 230.400 879.900 231.600 880.650 ;
        RECT 229.950 877.800 232.050 879.900 ;
        RECT 239.400 879.000 240.600 880.650 ;
        RECT 238.950 874.950 241.050 879.000 ;
        RECT 266.400 878.400 267.600 880.650 ;
        RECT 272.400 878.400 273.600 880.650 ;
        RECT 266.400 877.050 267.450 878.400 ;
        RECT 265.950 876.450 268.050 877.050 ;
        RECT 265.950 875.400 270.450 876.450 ;
        RECT 265.950 874.950 268.050 875.400 ;
        RECT 199.950 868.950 202.050 871.050 ;
        RECT 220.950 868.950 223.050 871.050 ;
        RECT 200.400 861.450 201.450 868.950 ;
        RECT 265.950 865.950 268.050 868.050 ;
        RECT 200.400 860.400 204.450 861.450 ;
        RECT 188.400 854.400 192.450 855.450 ;
        RECT 169.950 850.950 172.050 853.050 ;
        RECT 184.950 850.950 187.050 853.050 ;
        RECT 146.400 839.400 150.450 840.450 ;
        RECT 133.950 835.950 136.050 838.050 ;
        RECT 136.950 835.950 139.050 838.050 ;
        RECT 139.950 835.950 142.050 838.050 ;
        RECT 142.950 835.950 145.050 838.050 ;
        RECT 119.400 833.400 126.450 834.450 ;
        RECT 134.400 834.000 135.600 835.650 ;
        RECT 133.950 831.450 136.050 834.000 ;
        RECT 131.400 830.400 136.050 831.450 ;
        RECT 118.950 817.950 121.050 820.050 ;
        RECT 119.400 811.050 120.450 817.950 ;
        RECT 118.950 807.000 121.050 811.050 ;
        RECT 119.400 805.350 120.600 807.000 ;
        RECT 124.950 806.100 127.050 808.200 ;
        RECT 125.400 805.350 126.600 806.100 ;
        RECT 115.950 802.950 118.050 805.050 ;
        RECT 118.950 802.950 121.050 805.050 ;
        RECT 121.950 802.950 124.050 805.050 ;
        RECT 124.950 802.950 127.050 805.050 ;
        RECT 116.400 801.900 117.600 802.650 ;
        RECT 122.400 801.900 123.600 802.650 ;
        RECT 131.400 801.900 132.450 830.400 ;
        RECT 133.950 829.950 136.050 830.400 ;
        RECT 140.400 833.400 141.600 835.650 ;
        RECT 140.400 811.050 141.450 833.400 ;
        RECT 149.400 829.050 150.450 839.400 ;
        RECT 160.950 839.100 163.050 841.200 ;
        RECT 170.400 840.600 171.450 850.950 ;
        RECT 176.250 847.500 178.350 848.400 ;
        RECT 174.150 846.300 178.350 847.500 ;
        RECT 161.400 838.350 162.600 839.100 ;
        RECT 170.400 838.350 171.600 840.600 ;
        RECT 160.950 835.950 163.050 838.050 ;
        RECT 163.950 835.950 166.050 838.050 ;
        RECT 169.950 835.950 172.050 838.050 ;
        RECT 164.400 833.400 165.600 835.650 ;
        RECT 148.950 826.950 151.050 829.050 ;
        RECT 164.400 820.050 165.450 833.400 ;
        RECT 166.950 832.950 169.050 835.050 ;
        RECT 163.950 817.950 166.050 820.050 ;
        RECT 167.400 816.450 168.450 832.950 ;
        RECT 174.150 827.700 175.350 846.300 ;
        RECT 178.950 839.100 181.050 841.200 ;
        RECT 179.400 838.350 180.600 839.100 ;
        RECT 179.100 835.950 181.200 838.050 ;
        RECT 185.400 832.050 186.450 850.950 ;
        RECT 188.400 850.050 189.450 854.400 ;
        RECT 187.950 847.950 190.050 850.050 ;
        RECT 191.550 849.300 193.650 851.400 ;
        RECT 191.550 842.700 192.750 849.300 ;
        RECT 191.550 840.600 193.650 842.700 ;
        RECT 178.950 829.950 181.050 832.050 ;
        RECT 184.950 829.950 187.050 832.050 ;
        RECT 173.850 825.600 175.950 827.700 ;
        RECT 164.400 815.400 168.450 816.450 ;
        RECT 133.950 808.950 136.050 811.050 ;
        RECT 139.950 808.950 142.050 811.050 ;
        RECT 134.400 801.900 135.450 808.950 ;
        RECT 142.950 806.100 145.050 808.200 ;
        RECT 143.400 805.350 144.600 806.100 ;
        RECT 151.950 805.950 154.050 808.050 ;
        RECT 164.400 807.600 165.450 815.400 ;
        RECT 169.950 811.950 172.050 814.050 ;
        RECT 170.400 807.600 171.450 811.950 ;
        RECT 139.950 802.950 142.050 805.050 ;
        RECT 142.950 802.950 145.050 805.050 ;
        RECT 145.950 802.950 148.050 805.050 ;
        RECT 140.400 801.900 141.600 802.650 ;
        RECT 109.950 799.800 112.050 801.900 ;
        RECT 115.950 799.800 118.050 801.900 ;
        RECT 121.950 799.800 124.050 801.900 ;
        RECT 130.800 799.800 132.900 801.900 ;
        RECT 133.950 799.800 136.050 801.900 ;
        RECT 139.950 799.800 142.050 801.900 ;
        RECT 146.400 800.400 147.600 802.650 ;
        RECT 146.400 796.050 147.450 800.400 ;
        RECT 77.400 794.400 81.450 795.450 ;
        RECT 49.950 784.950 52.050 787.050 ;
        RECT 44.400 760.350 45.600 762.600 ;
        RECT 40.950 757.950 43.050 760.050 ;
        RECT 43.950 757.950 46.050 760.050 ;
        RECT 41.400 755.400 42.600 757.650 ;
        RECT 34.950 751.950 37.050 754.050 ;
        RECT 41.400 751.050 42.450 755.400 ;
        RECT 46.950 754.950 49.050 757.050 ;
        RECT 43.950 751.950 46.050 754.050 ;
        RECT 40.950 748.950 43.050 751.050 ;
        RECT 34.950 724.950 37.050 727.050 ;
        RECT 37.950 724.950 40.050 727.050 ;
        RECT 38.400 722.400 39.600 724.650 ;
        RECT 38.400 717.450 39.450 722.400 ;
        RECT 38.400 716.400 42.450 717.450 ;
        RECT 28.950 712.950 31.050 715.050 ;
        RECT 37.950 712.950 40.050 715.050 ;
        RECT 31.950 697.950 34.050 700.050 ;
        RECT 10.350 693.300 12.450 695.400 ;
        RECT 16.950 694.950 19.050 697.050 ;
        RECT 25.950 694.950 28.050 697.050 ;
        RECT 11.250 686.700 12.450 693.300 ;
        RECT 10.350 684.600 12.450 686.700 ;
        RECT 4.950 679.950 7.050 682.050 ;
        RECT 5.400 678.900 6.600 679.650 ;
        RECT 4.950 676.800 7.050 678.900 ;
        RECT 11.250 671.700 12.450 684.600 ;
        RECT 10.350 669.600 12.450 671.700 ;
        RECT 17.400 655.050 18.450 694.950 ;
        RECT 25.650 691.500 27.750 692.400 ;
        RECT 25.650 690.300 29.850 691.500 ;
        RECT 22.950 683.100 25.050 685.200 ;
        RECT 23.400 682.350 24.600 683.100 ;
        RECT 22.800 679.950 24.900 682.050 ;
        RECT 22.950 673.950 25.050 676.050 ;
        RECT 4.950 652.950 7.050 655.050 ;
        RECT 16.950 652.950 19.050 655.050 ;
        RECT 5.400 610.050 6.450 652.950 ;
        RECT 13.950 646.950 16.050 649.050 ;
        RECT 16.950 646.950 19.050 649.050 ;
        RECT 17.400 644.400 18.600 646.650 ;
        RECT 13.950 640.950 16.050 643.050 ;
        RECT 10.350 615.300 12.450 617.400 ;
        RECT 4.950 607.950 7.050 610.050 ;
        RECT 11.250 608.700 12.450 615.300 ;
        RECT 10.350 606.600 12.450 608.700 ;
        RECT 4.950 601.950 7.050 604.050 ;
        RECT 5.400 600.900 6.600 601.650 ;
        RECT 4.950 598.800 7.050 600.900 ;
        RECT 11.250 593.700 12.450 606.600 ;
        RECT 14.400 601.050 15.450 640.950 ;
        RECT 17.400 637.050 18.450 644.400 ;
        RECT 23.400 643.050 24.450 673.950 ;
        RECT 28.650 671.700 29.850 690.300 ;
        RECT 32.400 684.600 33.450 697.950 ;
        RECT 32.400 682.350 33.600 684.600 ;
        RECT 31.950 679.950 34.050 682.050 ;
        RECT 38.400 676.050 39.450 712.950 ;
        RECT 37.950 673.950 40.050 676.050 ;
        RECT 41.400 673.050 42.450 716.400 ;
        RECT 44.400 700.050 45.450 751.950 ;
        RECT 43.950 697.950 46.050 700.050 ;
        RECT 47.400 694.050 48.450 754.950 ;
        RECT 50.400 754.050 51.450 784.950 ;
        RECT 52.950 761.100 55.050 763.200 ;
        RECT 58.950 761.100 61.050 763.200 ;
        RECT 64.950 761.100 67.050 763.200 ;
        RECT 53.400 757.050 54.450 761.100 ;
        RECT 59.400 760.350 60.600 761.100 ;
        RECT 65.400 760.350 66.600 761.100 ;
        RECT 58.950 757.950 61.050 760.050 ;
        RECT 61.950 757.950 64.050 760.050 ;
        RECT 64.950 757.950 67.050 760.050 ;
        RECT 52.950 754.950 55.050 757.050 ;
        RECT 62.400 755.400 63.600 757.650 ;
        RECT 49.950 751.950 52.050 754.050 ;
        RECT 62.400 739.050 63.450 755.400 ;
        RECT 77.400 751.050 78.450 794.400 ;
        RECT 103.950 793.950 106.050 796.050 ;
        RECT 145.950 793.950 148.050 796.050 ;
        RECT 152.400 793.050 153.450 805.950 ;
        RECT 164.400 805.350 165.600 807.600 ;
        RECT 170.400 805.350 171.600 807.600 ;
        RECT 154.950 802.950 157.050 805.050 ;
        RECT 160.950 802.950 163.050 805.050 ;
        RECT 163.950 802.950 166.050 805.050 ;
        RECT 166.950 802.950 169.050 805.050 ;
        RECT 169.950 802.950 172.050 805.050 ;
        RECT 151.950 790.950 154.050 793.050 ;
        RECT 83.100 766.500 85.200 768.600 ;
        RECT 80.100 757.950 82.200 760.050 ;
        RECT 83.100 759.900 84.000 766.500 ;
        RECT 92.100 766.200 94.200 768.300 ;
        RECT 86.400 763.350 87.600 765.600 ;
        RECT 85.800 760.950 87.900 763.050 ;
        RECT 90.000 759.900 92.100 760.200 ;
        RECT 83.100 759.000 92.100 759.900 ;
        RECT 80.400 756.900 81.600 757.650 ;
        RECT 79.950 754.800 82.050 756.900 ;
        RECT 83.100 753.900 84.000 759.000 ;
        RECT 90.000 758.100 92.100 759.000 ;
        RECT 84.900 757.200 87.000 758.100 ;
        RECT 84.900 756.000 92.100 757.200 ;
        RECT 90.000 755.100 92.100 756.000 ;
        RECT 82.500 751.800 84.600 753.900 ;
        RECT 85.800 752.100 87.900 754.200 ;
        RECT 93.000 753.600 93.900 766.200 ;
        RECT 94.950 762.450 97.050 763.200 ;
        RECT 94.950 761.400 99.450 762.450 ;
        RECT 94.950 761.100 97.050 761.400 ;
        RECT 95.400 760.350 96.600 761.100 ;
        RECT 94.800 757.950 96.900 760.050 ;
        RECT 86.400 751.050 87.600 751.800 ;
        RECT 92.400 751.500 94.500 753.600 ;
        RECT 98.400 751.050 99.450 761.400 ;
        RECT 100.950 760.950 103.050 763.050 ;
        RECT 113.400 762.450 114.600 762.600 ;
        RECT 110.400 761.400 114.600 762.450 ;
        RECT 76.950 748.950 79.050 751.050 ;
        RECT 85.950 748.950 88.050 751.050 ;
        RECT 97.950 748.950 100.050 751.050 ;
        RECT 61.950 736.950 64.050 739.050 ;
        RECT 55.950 728.100 58.050 730.200 ;
        RECT 62.400 729.450 63.450 736.950 ;
        RECT 101.400 736.050 102.450 760.950 ;
        RECT 106.950 739.950 109.050 742.050 ;
        RECT 85.950 733.950 88.050 736.050 ;
        RECT 100.950 733.950 103.050 736.050 ;
        RECT 62.400 728.400 66.450 729.450 ;
        RECT 56.400 727.350 57.600 728.100 ;
        RECT 52.950 724.950 55.050 727.050 ;
        RECT 55.950 724.950 58.050 727.050 ;
        RECT 58.950 724.950 61.050 727.050 ;
        RECT 53.400 722.400 54.600 724.650 ;
        RECT 59.400 723.450 60.600 724.650 ;
        RECT 65.400 723.450 66.450 728.400 ;
        RECT 67.950 727.950 70.050 730.050 ;
        RECT 76.950 728.100 79.050 730.200 ;
        RECT 68.400 723.900 69.450 727.950 ;
        RECT 77.400 727.350 78.600 728.100 ;
        RECT 73.950 724.950 76.050 727.050 ;
        RECT 76.950 724.950 79.050 727.050 ;
        RECT 79.950 724.950 82.050 727.050 ;
        RECT 74.400 723.900 75.600 724.650 ;
        RECT 80.400 723.900 81.600 724.650 ;
        RECT 86.400 723.900 87.450 733.950 ;
        RECT 102.000 732.450 106.050 733.050 ;
        RECT 101.400 730.950 106.050 732.450 ;
        RECT 91.950 727.950 94.050 730.050 ;
        RECT 101.400 729.600 102.450 730.950 ;
        RECT 107.400 730.050 108.450 739.950 ;
        RECT 110.400 739.050 111.450 761.400 ;
        RECT 113.400 760.350 114.600 761.400 ;
        RECT 121.950 761.100 124.050 763.200 ;
        RECT 139.950 761.100 142.050 763.200 ;
        RECT 145.950 761.100 148.050 763.200 ;
        RECT 122.400 760.350 123.600 761.100 ;
        RECT 140.400 760.350 141.600 761.100 ;
        RECT 146.400 760.350 147.600 761.100 ;
        RECT 113.100 757.950 115.200 760.050 ;
        RECT 116.400 757.950 118.500 760.050 ;
        RECT 121.800 757.950 123.900 760.050 ;
        RECT 139.950 757.950 142.050 760.050 ;
        RECT 142.950 757.950 145.050 760.050 ;
        RECT 145.950 757.950 148.050 760.050 ;
        RECT 148.950 757.950 151.050 760.050 ;
        RECT 116.400 756.900 117.600 757.650 ;
        RECT 115.950 754.800 118.050 756.900 ;
        RECT 143.400 755.400 144.600 757.650 ;
        RECT 149.400 755.400 150.600 757.650 ;
        RECT 116.400 753.450 117.450 754.800 ;
        RECT 113.400 752.400 117.450 753.450 ;
        RECT 109.950 736.950 112.050 739.050 ;
        RECT 109.950 730.950 112.050 733.050 ;
        RECT 59.400 722.400 66.450 723.450 ;
        RECT 53.400 715.050 54.450 722.400 ;
        RECT 67.950 721.800 70.050 723.900 ;
        RECT 73.950 721.800 76.050 723.900 ;
        RECT 79.950 721.800 82.050 723.900 ;
        RECT 85.950 721.800 88.050 723.900 ;
        RECT 92.400 721.050 93.450 727.950 ;
        RECT 101.400 727.350 102.600 729.600 ;
        RECT 106.950 727.950 109.050 730.050 ;
        RECT 97.950 724.950 100.050 727.050 ;
        RECT 100.950 724.950 103.050 727.050 ;
        RECT 103.950 724.950 106.050 727.050 ;
        RECT 98.400 723.000 99.600 724.650 ;
        RECT 104.400 723.900 105.600 724.650 ;
        RECT 91.950 718.950 94.050 721.050 ;
        RECT 97.950 718.950 100.050 723.000 ;
        RECT 103.950 721.800 106.050 723.900 ;
        RECT 110.400 721.050 111.450 730.950 ;
        RECT 113.400 721.050 114.450 752.400 ;
        RECT 127.950 739.950 130.050 742.050 ;
        RECT 121.950 728.100 124.050 730.200 ;
        RECT 128.400 729.600 129.450 739.950 ;
        RECT 143.400 733.050 144.450 755.400 ;
        RECT 149.400 742.050 150.450 755.400 ;
        RECT 148.950 739.950 151.050 742.050 ;
        RECT 148.950 736.800 151.050 738.900 ;
        RECT 142.950 730.950 145.050 733.050 ;
        RECT 122.400 727.350 123.600 728.100 ;
        RECT 128.400 727.350 129.600 729.600 ;
        RECT 139.950 727.950 142.050 730.050 ;
        RECT 149.400 729.600 150.450 736.800 ;
        RECT 155.400 730.200 156.450 802.950 ;
        RECT 161.400 800.400 162.600 802.650 ;
        RECT 167.400 801.900 168.600 802.650 ;
        RECT 161.400 781.050 162.450 800.400 ;
        RECT 166.950 799.800 169.050 801.900 ;
        RECT 160.950 778.950 163.050 781.050 ;
        RECT 163.950 771.450 166.050 772.050 ;
        RECT 167.400 771.450 168.450 799.800 ;
        RECT 179.400 787.050 180.450 829.950 ;
        RECT 191.550 827.700 192.750 840.600 ;
        RECT 196.950 835.950 199.050 838.050 ;
        RECT 197.400 834.900 198.600 835.650 ;
        RECT 196.950 832.800 199.050 834.900 ;
        RECT 191.550 825.600 193.650 827.700 ;
        RECT 196.950 820.950 199.050 823.050 ;
        RECT 190.950 806.100 193.050 808.200 ;
        RECT 197.400 807.600 198.450 820.950 ;
        RECT 203.400 820.050 204.450 860.400 ;
        RECT 256.950 859.950 259.050 862.050 ;
        RECT 229.950 856.950 232.050 859.050 ;
        RECT 211.950 844.950 214.050 847.050 ;
        RECT 220.950 844.950 223.050 847.050 ;
        RECT 202.950 817.950 205.050 820.050 ;
        RECT 206.850 813.300 208.950 815.400 ;
        RECT 212.400 814.050 213.450 844.950 ;
        RECT 221.400 840.600 222.450 844.950 ;
        RECT 221.400 838.350 222.600 840.600 ;
        RECT 217.950 835.950 220.050 838.050 ;
        RECT 220.950 835.950 223.050 838.050 ;
        RECT 218.400 834.900 219.600 835.650 ;
        RECT 217.950 832.800 220.050 834.900 ;
        RECT 230.400 832.050 231.450 856.950 ;
        RECT 244.950 850.950 247.050 853.050 ;
        RECT 232.950 839.100 235.050 841.200 ;
        RECT 238.950 839.100 241.050 841.200 ;
        RECT 245.400 840.600 246.450 850.950 ;
        RECT 233.400 835.050 234.450 839.100 ;
        RECT 239.400 838.350 240.600 839.100 ;
        RECT 245.400 838.350 246.600 840.600 ;
        RECT 238.950 835.950 241.050 838.050 ;
        RECT 241.950 835.950 244.050 838.050 ;
        RECT 244.950 835.950 247.050 838.050 ;
        RECT 232.950 832.950 235.050 835.050 ;
        RECT 242.400 834.000 243.600 835.650 ;
        RECT 257.400 834.900 258.450 859.950 ;
        RECT 266.400 840.600 267.450 865.950 ;
        RECT 269.400 862.050 270.450 875.400 ;
        RECT 272.400 874.050 273.450 878.400 ;
        RECT 271.950 871.950 274.050 874.050 ;
        RECT 281.400 868.050 282.450 884.100 ;
        RECT 287.400 883.350 288.600 885.600 ;
        RECT 292.950 884.100 295.050 886.200 ;
        RECT 293.400 883.350 294.600 884.100 ;
        RECT 286.950 880.950 289.050 883.050 ;
        RECT 289.950 880.950 292.050 883.050 ;
        RECT 292.950 880.950 295.050 883.050 ;
        RECT 295.950 880.950 298.050 883.050 ;
        RECT 290.400 879.000 291.600 880.650 ;
        RECT 296.400 879.900 297.600 880.650 ;
        RECT 289.950 874.950 292.050 879.000 ;
        RECT 295.950 877.800 298.050 879.900 ;
        RECT 296.400 874.050 297.450 877.800 ;
        RECT 302.400 877.050 303.450 886.950 ;
        RECT 314.400 885.600 315.450 913.950 ;
        RECT 323.400 911.400 324.600 913.650 ;
        RECT 332.400 913.050 333.450 925.950 ;
        RECT 343.950 917.100 346.050 919.200 ;
        RECT 344.400 916.350 345.600 917.100 ;
        RECT 343.950 913.950 346.050 916.050 ;
        RECT 346.950 913.950 349.050 916.050 ;
        RECT 323.400 907.050 324.450 911.400 ;
        RECT 331.950 910.950 334.050 913.050 ;
        RECT 347.400 912.900 348.600 913.650 ;
        RECT 346.950 910.800 349.050 912.900 ;
        RECT 322.950 904.950 325.050 907.050 ;
        RECT 346.950 898.950 349.050 901.050 ;
        RECT 314.400 883.350 315.600 885.600 ;
        RECT 319.950 885.000 322.050 889.050 ;
        RECT 320.400 883.350 321.600 885.000 ;
        RECT 334.950 884.100 337.050 886.200 ;
        RECT 340.950 884.100 343.050 886.200 ;
        RECT 347.400 885.600 348.450 898.950 ;
        RECT 353.400 898.050 354.450 940.950 ;
        RECT 361.950 937.950 364.050 940.050 ;
        RECT 362.400 918.600 363.450 937.950 ;
        RECT 368.400 918.600 369.450 946.950 ;
        RECT 407.400 931.050 408.450 956.400 ;
        RECT 424.950 955.800 427.050 957.900 ;
        RECT 431.400 956.400 432.600 958.650 ;
        RECT 452.400 956.400 453.600 958.650 ;
        RECT 458.400 956.400 459.600 958.650 ;
        RECT 431.400 952.050 432.450 956.400 ;
        RECT 430.950 949.950 433.050 952.050 ;
        RECT 452.400 931.050 453.450 956.400 ;
        RECT 458.400 949.050 459.450 956.400 ;
        RECT 457.950 946.950 460.050 949.050 ;
        RECT 376.950 928.950 379.050 931.050 ;
        RECT 406.950 928.950 409.050 931.050 ;
        RECT 451.950 928.950 454.050 931.050 ;
        RECT 362.400 916.350 363.600 918.600 ;
        RECT 368.400 916.350 369.600 918.600 ;
        RECT 361.950 913.950 364.050 916.050 ;
        RECT 364.950 913.950 367.050 916.050 ;
        RECT 367.950 913.950 370.050 916.050 ;
        RECT 370.950 913.950 373.050 916.050 ;
        RECT 365.400 912.900 366.600 913.650 ;
        RECT 364.950 910.800 367.050 912.900 ;
        RECT 371.400 912.450 372.600 913.650 ;
        RECT 377.400 912.450 378.450 928.950 ;
        RECT 458.400 928.050 459.450 946.950 ;
        RECT 467.400 946.050 468.450 962.400 ;
        RECT 473.400 961.350 474.600 962.400 ;
        RECT 478.950 962.100 481.050 964.200 ;
        RECT 479.400 961.350 480.600 962.100 ;
        RECT 472.950 958.950 475.050 961.050 ;
        RECT 475.950 958.950 478.050 961.050 ;
        RECT 478.950 958.950 481.050 961.050 ;
        RECT 481.950 958.950 484.050 961.050 ;
        RECT 476.400 957.900 477.600 958.650 ;
        RECT 475.950 952.950 478.050 957.900 ;
        RECT 482.400 957.000 483.600 958.650 ;
        RECT 481.950 952.950 484.050 957.000 ;
        RECT 491.400 952.050 492.450 967.950 ;
        RECT 499.950 962.100 502.050 964.200 ;
        RECT 505.950 962.100 508.050 964.200 ;
        RECT 500.400 961.350 501.600 962.100 ;
        RECT 506.400 961.350 507.600 962.100 ;
        RECT 496.950 958.950 499.050 961.050 ;
        RECT 499.950 958.950 502.050 961.050 ;
        RECT 502.950 958.950 505.050 961.050 ;
        RECT 505.950 958.950 508.050 961.050 ;
        RECT 497.400 957.000 498.600 958.650 ;
        RECT 503.400 957.000 504.600 958.650 ;
        RECT 496.950 952.950 499.050 957.000 ;
        RECT 502.950 952.950 505.050 957.000 ;
        RECT 490.950 949.950 493.050 952.050 ;
        RECT 466.950 943.950 469.050 946.050 ;
        RECT 467.400 940.050 468.450 943.950 ;
        RECT 466.950 937.950 469.050 940.050 ;
        RECT 490.950 937.950 493.050 940.050 ;
        RECT 412.950 925.950 415.050 928.050 ;
        RECT 448.950 925.950 451.050 928.050 ;
        RECT 457.950 925.950 460.050 928.050 ;
        RECT 385.950 917.100 388.050 919.200 ;
        RECT 391.950 917.100 394.050 919.200 ;
        RECT 413.400 918.600 414.450 925.950 ;
        RECT 430.950 922.950 433.050 925.050 ;
        RECT 436.950 922.950 439.050 925.050 ;
        RECT 386.400 916.350 387.600 917.100 ;
        RECT 392.400 916.350 393.600 917.100 ;
        RECT 413.400 916.350 414.600 918.600 ;
        RECT 421.950 917.100 424.050 919.200 ;
        RECT 431.400 918.600 432.450 922.950 ;
        RECT 385.950 913.950 388.050 916.050 ;
        RECT 388.950 913.950 391.050 916.050 ;
        RECT 391.950 913.950 394.050 916.050 ;
        RECT 394.950 913.950 397.050 916.050 ;
        RECT 409.950 913.950 412.050 916.050 ;
        RECT 412.950 913.950 415.050 916.050 ;
        RECT 371.400 911.400 378.450 912.450 ;
        RECT 382.950 910.950 385.050 913.050 ;
        RECT 389.400 911.400 390.600 913.650 ;
        RECT 395.400 912.000 396.600 913.650 ;
        RECT 410.400 912.000 411.600 913.650 ;
        RECT 379.950 904.950 382.050 907.050 ;
        RECT 352.950 895.950 355.050 898.050 ;
        RECT 358.950 892.950 361.050 895.050 ;
        RECT 355.950 886.950 358.050 889.050 ;
        RECT 313.950 880.950 316.050 883.050 ;
        RECT 316.950 880.950 319.050 883.050 ;
        RECT 319.950 880.950 322.050 883.050 ;
        RECT 322.950 880.950 325.050 883.050 ;
        RECT 317.400 879.900 318.600 880.650 ;
        RECT 316.950 877.800 319.050 879.900 ;
        RECT 323.400 878.400 324.600 880.650 ;
        RECT 301.950 874.950 304.050 877.050 ;
        RECT 295.950 871.950 298.050 874.050 ;
        RECT 280.950 865.950 283.050 868.050 ;
        RECT 268.950 859.950 271.050 862.050 ;
        RECT 283.800 850.950 285.900 853.050 ;
        RECT 286.950 850.950 289.050 853.050 ;
        RECT 284.400 844.050 285.450 850.950 ;
        RECT 283.950 841.950 286.050 844.050 ;
        RECT 266.400 838.350 267.600 840.600 ;
        RECT 280.950 839.100 283.050 841.200 ;
        RECT 287.400 840.600 288.450 850.950 ;
        RECT 281.400 838.350 282.600 839.100 ;
        RECT 287.400 838.350 288.600 840.600 ;
        RECT 262.950 835.950 265.050 838.050 ;
        RECT 265.950 835.950 268.050 838.050 ;
        RECT 280.950 835.950 283.050 838.050 ;
        RECT 283.950 835.950 286.050 838.050 ;
        RECT 286.950 835.950 289.050 838.050 ;
        RECT 263.400 834.900 264.600 835.650 ;
        RECT 284.400 834.900 285.600 835.650 ;
        RECT 296.400 835.050 297.450 871.950 ;
        RECT 323.400 868.050 324.450 878.400 ;
        RECT 325.950 877.800 328.050 879.900 ;
        RECT 326.400 871.050 327.450 877.800 ;
        RECT 325.950 868.950 328.050 871.050 ;
        RECT 322.950 865.950 325.050 868.050 ;
        RECT 301.950 862.950 304.050 865.050 ;
        RECT 307.950 862.950 310.050 865.050 ;
        RECT 302.400 859.050 303.450 862.950 ;
        RECT 308.400 859.050 309.450 862.950 ;
        RECT 301.950 856.950 304.050 859.050 ;
        RECT 307.950 856.950 310.050 859.050 ;
        RECT 304.800 850.950 306.900 853.050 ;
        RECT 307.950 850.950 310.050 853.050 ;
        RECT 305.400 840.600 306.450 850.950 ;
        RECT 308.400 844.050 309.450 850.950 ;
        RECT 307.950 841.950 310.050 844.050 ;
        RECT 326.400 840.600 327.450 868.950 ;
        RECT 335.400 862.050 336.450 884.100 ;
        RECT 341.400 883.350 342.600 884.100 ;
        RECT 347.400 883.350 348.600 885.600 ;
        RECT 340.950 880.950 343.050 883.050 ;
        RECT 343.950 880.950 346.050 883.050 ;
        RECT 346.950 880.950 349.050 883.050 ;
        RECT 349.950 880.950 352.050 883.050 ;
        RECT 344.400 879.900 345.600 880.650 ;
        RECT 350.400 879.900 351.600 880.650 ;
        RECT 356.400 880.050 357.450 886.950 ;
        RECT 343.950 877.800 346.050 879.900 ;
        RECT 349.950 877.800 352.050 879.900 ;
        RECT 355.950 877.950 358.050 880.050 ;
        RECT 337.950 865.950 340.050 868.050 ;
        RECT 334.950 859.950 337.050 862.050 ;
        RECT 305.400 838.350 306.600 840.600 ;
        RECT 326.400 838.350 327.600 840.600 ;
        RECT 298.950 835.950 301.050 838.050 ;
        RECT 304.950 835.950 307.050 838.050 ;
        RECT 307.950 835.950 310.050 838.050 ;
        RECT 322.950 835.950 325.050 838.050 ;
        RECT 325.950 835.950 328.050 838.050 ;
        RECT 328.950 835.950 331.050 838.050 ;
        RECT 229.950 829.950 232.050 832.050 ;
        RECT 241.950 829.950 244.050 834.000 ;
        RECT 256.950 832.800 259.050 834.900 ;
        RECT 262.950 832.800 265.050 834.900 ;
        RECT 283.950 832.800 286.050 834.900 ;
        RECT 295.950 832.950 298.050 835.050 ;
        RECT 247.950 826.950 250.050 829.050 ;
        RECT 191.400 805.350 192.600 806.100 ;
        RECT 197.400 805.350 198.600 807.600 ;
        RECT 187.950 802.950 190.050 805.050 ;
        RECT 190.950 802.950 193.050 805.050 ;
        RECT 193.950 802.950 196.050 805.050 ;
        RECT 196.950 802.950 199.050 805.050 ;
        RECT 202.950 802.950 205.050 805.050 ;
        RECT 188.400 800.400 189.600 802.650 ;
        RECT 194.400 801.900 195.600 802.650 ;
        RECT 178.950 784.950 181.050 787.050 ;
        RECT 188.400 775.050 189.450 800.400 ;
        RECT 193.950 799.800 196.050 801.900 ;
        RECT 203.400 800.400 204.600 802.650 ;
        RECT 203.400 787.050 204.450 800.400 ;
        RECT 207.150 794.700 208.350 813.300 ;
        RECT 211.950 811.950 214.050 814.050 ;
        RECT 224.550 813.300 226.650 815.400 ;
        RECT 217.950 805.950 220.050 808.050 ;
        RECT 212.100 802.950 214.200 805.050 ;
        RECT 212.400 801.900 213.600 802.650 ;
        RECT 218.400 801.900 219.450 805.950 ;
        RECT 211.950 799.800 214.050 801.900 ;
        RECT 217.950 799.800 220.050 801.900 ;
        RECT 224.550 800.400 225.750 813.300 ;
        RECT 229.950 806.100 232.050 808.200 ;
        RECT 235.950 806.100 238.050 808.200 ;
        RECT 230.400 805.350 231.600 806.100 ;
        RECT 229.950 802.950 232.050 805.050 ;
        RECT 224.550 798.300 226.650 800.400 ;
        RECT 207.150 793.500 211.350 794.700 ;
        RECT 209.250 792.600 211.350 793.500 ;
        RECT 224.550 791.700 225.750 798.300 ;
        RECT 224.550 789.600 226.650 791.700 ;
        RECT 202.950 784.950 205.050 787.050 ;
        RECT 236.400 775.050 237.450 806.100 ;
        RECT 241.950 805.950 244.050 808.050 ;
        RECT 248.400 807.600 249.450 826.950 ;
        RECT 280.950 817.950 283.050 820.050 ;
        RECT 281.400 813.450 282.450 817.950 ;
        RECT 274.500 809.400 276.600 811.500 ;
        RECT 281.400 811.200 282.600 813.450 ;
        RECT 175.950 772.950 178.050 775.050 ;
        RECT 187.950 772.950 190.050 775.050 ;
        RECT 235.950 772.950 238.050 775.050 ;
        RECT 163.950 770.400 168.450 771.450 ;
        RECT 163.950 769.950 166.050 770.400 ;
        RECT 164.400 762.600 165.450 769.950 ;
        RECT 164.400 760.350 165.600 762.600 ;
        RECT 163.950 757.950 166.050 760.050 ;
        RECT 166.950 757.950 169.050 760.050 ;
        RECT 169.950 757.950 172.050 760.050 ;
        RECT 167.400 756.900 168.600 757.650 ;
        RECT 176.400 757.050 177.450 772.950 ;
        RECT 242.400 769.050 243.450 805.950 ;
        RECT 248.400 805.350 249.600 807.600 ;
        RECT 253.950 806.100 256.050 808.200 ;
        RECT 254.400 805.350 255.600 806.100 ;
        RECT 247.950 802.950 250.050 805.050 ;
        RECT 250.950 802.950 253.050 805.050 ;
        RECT 253.950 802.950 256.050 805.050 ;
        RECT 256.950 802.950 259.050 805.050 ;
        RECT 272.100 802.950 274.200 805.050 ;
        RECT 251.400 800.400 252.600 802.650 ;
        RECT 257.400 800.400 258.600 802.650 ;
        RECT 272.400 801.900 273.600 802.650 ;
        RECT 251.400 793.050 252.450 800.400 ;
        RECT 250.950 790.950 253.050 793.050 ;
        RECT 257.400 784.050 258.450 800.400 ;
        RECT 262.950 799.800 265.050 801.900 ;
        RECT 271.950 799.800 274.050 801.900 ;
        RECT 256.950 781.950 259.050 784.050 ;
        RECT 211.800 766.500 213.900 768.600 ;
        RECT 184.950 761.100 187.050 763.200 ;
        RECT 190.950 762.000 193.050 766.050 ;
        RECT 205.950 763.950 208.050 766.050 ;
        RECT 185.400 760.350 186.600 761.100 ;
        RECT 191.400 760.350 192.600 762.000 ;
        RECT 184.950 757.950 187.050 760.050 ;
        RECT 187.950 757.950 190.050 760.050 ;
        RECT 190.950 757.950 193.050 760.050 ;
        RECT 166.950 754.800 169.050 756.900 ;
        RECT 175.950 754.950 178.050 757.050 ;
        RECT 188.400 755.400 189.600 757.650 ;
        RECT 206.400 756.450 207.450 763.950 ;
        RECT 209.100 757.950 211.200 760.050 ;
        RECT 212.100 759.300 213.300 766.500 ;
        RECT 215.400 763.350 216.600 765.600 ;
        RECT 221.400 765.300 223.500 767.400 ;
        RECT 241.950 766.950 244.050 769.050 ;
        RECT 253.950 766.950 256.050 769.050 ;
        RECT 215.100 760.950 217.200 763.050 ;
        RECT 218.100 761.700 220.200 763.800 ;
        RECT 218.100 759.300 219.000 761.700 ;
        RECT 212.100 758.100 219.000 759.300 ;
        RECT 209.400 756.450 210.600 757.650 ;
        RECT 206.400 755.400 210.600 756.450 ;
        RECT 188.400 742.050 189.450 755.400 ;
        RECT 212.100 752.700 213.000 758.100 ;
        RECT 213.900 756.300 216.000 757.200 ;
        RECT 221.700 756.300 222.600 765.300 ;
        RECT 224.400 762.450 225.600 762.600 ;
        RECT 224.400 761.400 228.450 762.450 ;
        RECT 224.400 760.350 225.600 761.400 ;
        RECT 227.400 760.050 228.450 761.400 ;
        RECT 241.950 761.100 244.050 763.200 ;
        RECT 242.400 760.350 243.600 761.100 ;
        RECT 250.950 760.950 253.050 763.050 ;
        RECT 223.800 757.950 225.900 760.050 ;
        RECT 226.950 757.950 229.050 760.050 ;
        RECT 238.950 757.950 241.050 760.050 ;
        RECT 241.950 757.950 244.050 760.050 ;
        RECT 244.950 757.950 247.050 760.050 ;
        RECT 213.900 755.100 222.600 756.300 ;
        RECT 211.800 750.600 213.900 752.700 ;
        RECT 215.100 752.100 217.200 754.200 ;
        RECT 219.000 753.300 221.100 755.100 ;
        RECT 215.400 751.050 216.600 751.800 ;
        RECT 214.950 748.950 217.050 751.050 ;
        RECT 227.400 742.050 228.450 757.950 ;
        RECT 239.400 756.900 240.600 757.650 ;
        RECT 238.950 754.800 241.050 756.900 ;
        RECT 245.400 755.400 246.600 757.650 ;
        RECT 187.950 739.950 190.050 742.050 ;
        RECT 226.950 739.950 229.050 742.050 ;
        RECT 220.950 736.950 223.050 739.050 ;
        RECT 184.950 733.950 187.050 736.050 ;
        RECT 196.950 733.950 199.050 736.050 ;
        RECT 157.950 730.950 160.050 733.050 ;
        RECT 118.950 724.950 121.050 727.050 ;
        RECT 121.950 724.950 124.050 727.050 ;
        RECT 124.950 724.950 127.050 727.050 ;
        RECT 127.950 724.950 130.050 727.050 ;
        RECT 119.400 723.000 120.600 724.650 ;
        RECT 109.950 718.950 112.050 721.050 ;
        RECT 112.950 718.950 115.050 721.050 ;
        RECT 118.950 718.950 121.050 723.000 ;
        RECT 125.400 722.400 126.600 724.650 ;
        RECT 125.400 721.050 126.450 722.400 ;
        RECT 124.950 718.950 127.050 721.050 ;
        RECT 113.400 715.050 114.450 718.950 ;
        RECT 52.950 712.950 55.050 715.050 ;
        RECT 112.950 712.950 115.050 715.050 ;
        RECT 67.950 703.950 70.050 706.050 ;
        RECT 46.950 693.450 49.050 694.050 ;
        RECT 44.400 692.400 49.050 693.450 ;
        RECT 44.400 678.900 45.450 692.400 ;
        RECT 46.950 691.950 49.050 692.400 ;
        RECT 52.950 684.000 55.050 688.050 ;
        RECT 53.400 682.350 54.600 684.000 ;
        RECT 58.950 683.100 61.050 685.200 ;
        RECT 64.950 683.100 67.050 685.200 ;
        RECT 59.400 682.350 60.600 683.100 ;
        RECT 49.950 679.950 52.050 682.050 ;
        RECT 52.950 679.950 55.050 682.050 ;
        RECT 55.950 679.950 58.050 682.050 ;
        RECT 58.950 679.950 61.050 682.050 ;
        RECT 43.950 676.800 46.050 678.900 ;
        RECT 50.400 677.400 51.600 679.650 ;
        RECT 56.400 678.900 57.600 679.650 ;
        RECT 65.400 679.050 66.450 683.100 ;
        RECT 50.400 673.050 51.450 677.400 ;
        RECT 55.950 676.800 58.050 678.900 ;
        RECT 64.950 676.950 67.050 679.050 ;
        RECT 68.400 673.050 69.450 703.950 ;
        RECT 125.400 703.050 126.450 718.950 ;
        RECT 140.400 718.050 141.450 727.950 ;
        RECT 149.400 727.350 150.600 729.600 ;
        RECT 154.950 728.100 157.050 730.200 ;
        RECT 145.950 724.950 148.050 727.050 ;
        RECT 148.950 724.950 151.050 727.050 ;
        RECT 151.950 724.950 154.050 727.050 ;
        RECT 146.400 723.900 147.600 724.650 ;
        RECT 145.950 721.800 148.050 723.900 ;
        RECT 152.400 722.400 153.600 724.650 ;
        RECT 152.400 718.050 153.450 722.400 ;
        RECT 139.950 715.950 142.050 718.050 ;
        RECT 151.950 715.950 154.050 718.050 ;
        RECT 124.950 700.950 127.050 703.050 ;
        RECT 88.950 697.950 91.050 700.050 ;
        RECT 76.950 691.950 79.050 694.050 ;
        RECT 70.950 683.100 73.050 685.200 ;
        RECT 77.400 684.600 78.450 691.950 ;
        RECT 28.050 669.600 30.150 671.700 ;
        RECT 40.950 670.950 43.050 673.050 ;
        RECT 49.950 670.950 52.050 673.050 ;
        RECT 58.950 670.950 61.050 673.050 ;
        RECT 67.950 670.950 70.050 673.050 ;
        RECT 50.400 667.050 51.450 670.950 ;
        RECT 49.950 664.950 52.050 667.050 ;
        RECT 49.950 658.950 52.050 661.050 ;
        RECT 28.950 652.950 31.050 655.050 ;
        RECT 29.400 645.900 30.450 652.950 ;
        RECT 37.950 650.100 40.050 652.200 ;
        RECT 38.400 649.350 39.600 650.100 ;
        RECT 46.950 649.950 49.050 652.050 ;
        RECT 34.950 646.950 37.050 649.050 ;
        RECT 37.950 646.950 40.050 649.050 ;
        RECT 40.950 646.950 43.050 649.050 ;
        RECT 35.400 645.900 36.600 646.650 ;
        RECT 41.400 645.900 42.600 646.650 ;
        RECT 28.950 643.800 31.050 645.900 ;
        RECT 34.950 643.800 37.050 645.900 ;
        RECT 40.950 643.800 43.050 645.900 ;
        RECT 22.950 640.950 25.050 643.050 ;
        RECT 16.950 634.950 19.050 637.050 ;
        RECT 41.400 619.050 42.450 643.800 ;
        RECT 43.950 631.950 46.050 634.050 ;
        RECT 40.950 616.950 43.050 619.050 ;
        RECT 25.650 613.500 27.750 614.400 ;
        RECT 25.650 612.300 29.850 613.500 ;
        RECT 16.950 605.100 19.050 607.200 ;
        RECT 22.950 605.100 25.050 607.200 ;
        RECT 13.950 598.950 16.050 601.050 ;
        RECT 17.400 595.050 18.450 605.100 ;
        RECT 23.400 604.350 24.600 605.100 ;
        RECT 22.800 601.950 24.900 604.050 ;
        RECT 19.950 598.950 22.050 601.050 ;
        RECT 10.350 591.600 12.450 593.700 ;
        RECT 16.950 592.950 19.050 595.050 ;
        RECT 20.400 573.600 21.450 598.950 ;
        RECT 28.650 593.700 29.850 612.300 ;
        RECT 31.950 605.100 34.050 607.200 ;
        RECT 37.950 605.100 40.050 607.200 ;
        RECT 32.400 604.350 33.600 605.100 ;
        RECT 31.950 601.950 34.050 604.050 ;
        RECT 28.050 591.600 30.150 593.700 ;
        RECT 20.400 571.350 21.600 573.600 ;
        RECT 16.950 568.950 19.050 571.050 ;
        RECT 19.950 568.950 22.050 571.050 ;
        RECT 22.950 568.950 25.050 571.050 ;
        RECT 23.400 567.900 24.600 568.650 ;
        RECT 22.950 565.800 25.050 567.900 ;
        RECT 28.950 565.800 31.050 567.900 ;
        RECT 29.400 559.050 30.450 565.800 ;
        RECT 38.400 565.050 39.450 605.100 ;
        RECT 44.400 601.050 45.450 631.950 ;
        RECT 47.400 613.050 48.450 649.950 ;
        RECT 50.400 646.050 51.450 658.950 ;
        RECT 59.400 652.200 60.450 670.950 ;
        RECT 71.400 661.050 72.450 683.100 ;
        RECT 77.400 682.350 78.600 684.600 ;
        RECT 82.950 683.100 85.050 685.200 ;
        RECT 83.400 682.350 84.600 683.100 ;
        RECT 76.950 679.950 79.050 682.050 ;
        RECT 79.950 679.950 82.050 682.050 ;
        RECT 82.950 679.950 85.050 682.050 ;
        RECT 80.400 678.900 81.600 679.650 ;
        RECT 79.950 676.800 82.050 678.900 ;
        RECT 70.950 658.950 73.050 661.050 ;
        RECT 74.850 657.300 76.950 659.400 ;
        RECT 58.950 650.100 61.050 652.200 ;
        RECT 64.950 650.100 67.050 652.200 ;
        RECT 59.400 649.350 60.600 650.100 ;
        RECT 65.400 649.350 66.600 650.100 ;
        RECT 55.950 646.950 58.050 649.050 ;
        RECT 58.950 646.950 61.050 649.050 ;
        RECT 61.950 646.950 64.050 649.050 ;
        RECT 64.950 646.950 67.050 649.050 ;
        RECT 70.950 646.950 73.050 649.050 ;
        RECT 49.950 643.950 52.050 646.050 ;
        RECT 56.400 644.400 57.600 646.650 ;
        RECT 62.400 645.000 63.600 646.650 ;
        RECT 56.400 634.050 57.450 644.400 ;
        RECT 61.950 640.950 64.050 645.000 ;
        RECT 71.400 644.400 72.600 646.650 ;
        RECT 71.400 634.050 72.450 644.400 ;
        RECT 75.150 638.700 76.350 657.300 ;
        RECT 85.950 649.950 88.050 652.050 ;
        RECT 80.100 646.950 82.200 649.050 ;
        RECT 80.400 645.900 81.600 646.650 ;
        RECT 86.400 645.900 87.450 649.950 ;
        RECT 79.950 643.800 82.050 645.900 ;
        RECT 85.950 643.800 88.050 645.900 ;
        RECT 75.150 637.500 79.350 638.700 ;
        RECT 77.250 636.600 79.350 637.500 ;
        RECT 89.400 634.050 90.450 697.950 ;
        RECT 103.800 688.200 105.900 690.300 ;
        RECT 112.800 688.500 114.900 690.600 ;
        RECT 133.800 688.500 135.900 690.600 ;
        RECT 100.950 683.100 103.050 685.200 ;
        RECT 101.400 682.350 102.600 683.100 ;
        RECT 101.100 679.950 103.200 682.050 ;
        RECT 104.100 675.600 105.000 688.200 ;
        RECT 110.400 685.350 111.600 687.600 ;
        RECT 110.100 682.950 112.200 685.050 ;
        RECT 105.900 681.900 108.000 682.200 ;
        RECT 114.000 681.900 114.900 688.500 ;
        RECT 105.900 681.000 114.900 681.900 ;
        RECT 105.900 680.100 108.000 681.000 ;
        RECT 111.000 679.200 113.100 680.100 ;
        RECT 105.900 678.000 113.100 679.200 ;
        RECT 105.900 677.100 108.000 678.000 ;
        RECT 103.500 673.500 105.600 675.600 ;
        RECT 110.100 674.100 112.200 676.200 ;
        RECT 114.000 675.900 114.900 681.000 ;
        RECT 115.800 679.950 117.900 682.050 ;
        RECT 131.100 679.950 133.200 682.050 ;
        RECT 134.100 681.300 135.300 688.500 ;
        RECT 137.400 685.350 138.600 687.600 ;
        RECT 143.400 687.300 145.500 689.400 ;
        RECT 137.100 682.950 139.200 685.050 ;
        RECT 140.100 683.700 142.200 685.800 ;
        RECT 140.100 681.300 141.000 683.700 ;
        RECT 134.100 680.100 141.000 681.300 ;
        RECT 116.400 678.450 117.600 679.650 ;
        RECT 131.400 678.450 132.600 679.650 ;
        RECT 116.400 677.400 120.450 678.450 ;
        RECT 113.400 673.800 115.500 675.900 ;
        RECT 110.400 672.000 111.600 673.800 ;
        RECT 119.400 673.050 120.450 677.400 ;
        RECT 128.400 677.400 132.600 678.450 ;
        RECT 109.950 667.950 112.050 672.000 ;
        RECT 118.950 670.950 121.050 673.050 ;
        RECT 103.950 664.950 106.050 667.050 ;
        RECT 97.950 661.950 100.050 664.050 ;
        RECT 92.550 657.300 94.650 659.400 ;
        RECT 92.550 644.400 93.750 657.300 ;
        RECT 98.400 651.600 99.450 661.950 ;
        RECT 98.400 649.350 99.600 651.600 ;
        RECT 97.950 646.950 100.050 649.050 ;
        RECT 92.550 642.300 94.650 644.400 ;
        RECT 92.550 635.700 93.750 642.300 ;
        RECT 55.950 631.950 58.050 634.050 ;
        RECT 70.950 631.950 73.050 634.050 ;
        RECT 88.950 631.950 91.050 634.050 ;
        RECT 92.550 633.600 94.650 635.700 ;
        RECT 64.950 619.950 67.050 622.050 ;
        RECT 52.950 616.950 55.050 619.050 ;
        RECT 46.950 610.950 49.050 613.050 ;
        RECT 53.400 607.200 54.450 616.950 ;
        RECT 58.950 610.950 61.050 613.050 ;
        RECT 52.950 605.100 55.050 607.200 ;
        RECT 59.400 606.600 60.450 610.950 ;
        RECT 53.400 604.350 54.600 605.100 ;
        RECT 59.400 604.350 60.600 606.600 ;
        RECT 49.950 601.950 52.050 604.050 ;
        RECT 52.950 601.950 55.050 604.050 ;
        RECT 55.950 601.950 58.050 604.050 ;
        RECT 58.950 601.950 61.050 604.050 ;
        RECT 43.950 598.950 46.050 601.050 ;
        RECT 50.400 600.900 51.600 601.650 ;
        RECT 49.950 598.800 52.050 600.900 ;
        RECT 56.400 599.400 57.600 601.650 ;
        RECT 44.100 568.950 46.200 571.050 ;
        RECT 44.400 567.000 45.600 568.650 ;
        RECT 50.400 567.450 51.450 598.800 ;
        RECT 56.400 595.050 57.450 599.400 ;
        RECT 55.950 592.950 58.050 595.050 ;
        RECT 58.950 589.950 61.050 592.050 ;
        RECT 52.950 574.950 55.050 577.050 ;
        RECT 37.950 562.950 40.050 565.050 ;
        RECT 43.950 562.950 46.050 567.000 ;
        RECT 47.400 566.400 51.450 567.450 ;
        RECT 28.950 556.950 31.050 559.050 ;
        RECT 37.950 532.950 40.050 535.050 ;
        RECT 38.400 528.600 39.450 532.950 ;
        RECT 38.400 526.350 39.600 528.600 ;
        RECT 14.100 523.950 16.200 526.050 ;
        RECT 19.500 523.950 21.600 526.050 ;
        RECT 34.950 523.950 37.050 526.050 ;
        RECT 37.950 523.950 40.050 526.050 ;
        RECT 20.400 522.900 21.600 523.650 ;
        RECT 19.950 520.800 22.050 522.900 ;
        RECT 43.950 520.950 46.050 523.050 ;
        RECT 44.400 517.050 45.450 520.950 ;
        RECT 43.950 514.950 46.050 517.050 ;
        RECT 19.950 505.950 22.050 508.050 ;
        RECT 20.400 495.600 21.450 505.950 ;
        RECT 20.400 493.350 21.600 495.600 ;
        RECT 14.100 490.950 16.200 493.050 ;
        RECT 19.500 490.950 21.600 493.050 ;
        RECT 37.800 490.950 39.900 493.050 ;
        RECT 17.100 445.950 19.200 448.050 ;
        RECT 22.500 445.950 24.600 448.050 ;
        RECT 38.100 445.950 40.200 448.050 ;
        RECT 43.500 445.950 45.600 448.050 ;
        RECT 23.400 444.900 24.600 445.650 ;
        RECT 44.400 444.900 45.600 445.650 ;
        RECT 22.950 442.800 25.050 444.900 ;
        RECT 43.950 442.800 46.050 444.900 ;
        RECT 31.950 433.950 34.050 436.050 ;
        RECT 19.950 427.950 22.050 430.050 ;
        RECT 8.850 423.300 10.950 425.400 ;
        RECT 4.950 412.950 7.050 415.050 ;
        RECT 5.400 410.400 6.600 412.650 ;
        RECT 5.400 403.050 6.450 410.400 ;
        RECT 9.150 404.700 10.350 423.300 ;
        RECT 14.100 412.950 16.200 415.050 ;
        RECT 9.150 403.500 13.350 404.700 ;
        RECT 4.950 400.950 7.050 403.050 ;
        RECT 11.250 402.600 13.350 403.500 ;
        RECT 1.950 394.950 4.050 397.050 ;
        RECT 2.400 327.450 3.450 394.950 ;
        RECT 5.400 352.050 6.450 400.950 ;
        RECT 20.400 372.600 21.450 427.950 ;
        RECT 26.550 423.300 28.650 425.400 ;
        RECT 26.550 410.400 27.750 423.300 ;
        RECT 32.400 418.200 33.450 433.950 ;
        RECT 47.400 430.050 48.450 566.400 ;
        RECT 53.400 529.200 54.450 574.950 ;
        RECT 59.400 535.050 60.450 589.950 ;
        RECT 65.400 577.050 66.450 619.950 ;
        RECT 71.400 610.050 72.450 631.950 ;
        RECT 82.950 613.950 85.050 616.050 ;
        RECT 70.950 607.950 73.050 610.050 ;
        RECT 76.950 605.100 79.050 607.200 ;
        RECT 83.400 606.600 84.450 613.950 ;
        RECT 95.250 613.500 97.350 614.400 ;
        RECT 93.150 612.300 97.350 613.500 ;
        RECT 77.400 604.350 78.600 605.100 ;
        RECT 83.400 604.350 84.600 606.600 ;
        RECT 88.950 606.000 91.050 610.050 ;
        RECT 89.400 604.350 90.600 606.000 ;
        RECT 73.950 601.950 76.050 604.050 ;
        RECT 76.950 601.950 79.050 604.050 ;
        RECT 79.950 601.950 82.050 604.050 ;
        RECT 82.950 601.950 85.050 604.050 ;
        RECT 88.950 601.950 91.050 604.050 ;
        RECT 74.400 599.400 75.600 601.650 ;
        RECT 80.400 600.900 81.600 601.650 ;
        RECT 74.400 592.050 75.450 599.400 ;
        RECT 79.950 598.800 82.050 600.900 ;
        RECT 88.950 595.950 91.050 598.050 ;
        RECT 73.950 589.950 76.050 592.050 ;
        RECT 74.850 579.300 76.950 581.400 ;
        RECT 64.950 574.950 67.050 577.050 ;
        RECT 62.100 568.950 64.200 571.050 ;
        RECT 70.950 568.950 73.050 571.050 ;
        RECT 71.400 567.000 72.600 568.650 ;
        RECT 70.950 562.950 73.050 567.000 ;
        RECT 75.150 560.700 76.350 579.300 ;
        RECT 80.100 568.950 82.200 571.050 ;
        RECT 80.400 567.450 81.600 568.650 ;
        RECT 80.400 566.400 84.450 567.450 ;
        RECT 75.150 559.500 79.350 560.700 ;
        RECT 77.250 558.600 79.350 559.500 ;
        RECT 58.950 532.950 61.050 535.050 ;
        RECT 67.950 532.950 70.050 535.050 ;
        RECT 52.950 527.100 55.050 529.200 ;
        RECT 58.950 527.100 61.050 529.200 ;
        RECT 53.400 526.350 54.600 527.100 ;
        RECT 59.400 526.350 60.600 527.100 ;
        RECT 52.950 523.950 55.050 526.050 ;
        RECT 55.950 523.950 58.050 526.050 ;
        RECT 58.950 523.950 61.050 526.050 ;
        RECT 64.950 523.950 67.050 529.200 ;
        RECT 49.950 520.950 52.050 523.050 ;
        RECT 56.400 522.900 57.600 523.650 ;
        RECT 50.400 514.050 51.450 520.950 ;
        RECT 55.950 520.800 58.050 522.900 ;
        RECT 61.950 517.950 64.050 523.050 ;
        RECT 64.950 520.800 67.050 522.900 ;
        RECT 65.400 517.050 66.450 520.800 ;
        RECT 68.400 517.050 69.450 532.950 ;
        RECT 83.400 532.050 84.450 566.400 ;
        RECT 89.400 559.050 90.450 595.950 ;
        RECT 93.150 593.700 94.350 612.300 ;
        RECT 97.950 605.100 100.050 607.200 ;
        RECT 98.400 604.350 99.600 605.100 ;
        RECT 98.100 601.950 100.200 604.050 ;
        RECT 92.850 591.600 94.950 593.700 ;
        RECT 92.550 579.300 94.650 581.400 ;
        RECT 92.550 566.400 93.750 579.300 ;
        RECT 97.950 572.100 100.050 574.200 ;
        RECT 104.400 574.050 105.450 664.950 ;
        RECT 124.950 661.950 127.050 664.050 ;
        RECT 125.400 652.200 126.450 661.950 ;
        RECT 106.950 650.100 109.050 652.200 ;
        RECT 118.950 650.100 121.050 652.200 ;
        RECT 124.950 650.100 127.050 652.200 ;
        RECT 128.400 652.050 129.450 677.400 ;
        RECT 134.100 674.700 135.000 680.100 ;
        RECT 135.900 678.300 138.000 679.200 ;
        RECT 143.700 678.300 144.600 687.300 ;
        RECT 158.400 685.200 159.450 730.950 ;
        RECT 160.950 727.950 163.050 730.050 ;
        RECT 169.950 728.100 172.050 730.200 ;
        RECT 161.400 723.900 162.450 727.950 ;
        RECT 170.400 727.350 171.600 728.100 ;
        RECT 167.100 724.950 169.200 727.050 ;
        RECT 170.400 724.950 172.500 727.050 ;
        RECT 175.800 724.950 177.900 727.050 ;
        RECT 167.400 723.900 168.600 724.650 ;
        RECT 160.950 721.800 163.050 723.900 ;
        RECT 166.950 721.800 169.050 723.900 ;
        RECT 176.400 722.400 177.600 724.650 ;
        RECT 167.400 718.050 168.450 721.800 ;
        RECT 176.400 718.050 177.450 722.400 ;
        RECT 166.950 715.950 169.050 718.050 ;
        RECT 175.950 715.950 178.050 718.050 ;
        RECT 146.400 684.450 147.600 684.600 ;
        RECT 146.400 684.000 150.450 684.450 ;
        RECT 146.400 683.400 151.050 684.000 ;
        RECT 146.400 682.350 147.600 683.400 ;
        RECT 145.800 679.950 147.900 682.050 ;
        RECT 148.950 679.950 151.050 683.400 ;
        RECT 157.950 683.100 160.050 685.200 ;
        RECT 163.950 683.100 166.050 685.200 ;
        RECT 178.950 683.100 181.050 685.200 ;
        RECT 185.400 684.600 186.450 733.950 ;
        RECT 190.950 728.100 193.050 730.200 ;
        RECT 197.400 729.600 198.450 733.950 ;
        RECT 191.400 727.350 192.600 728.100 ;
        RECT 197.400 727.350 198.600 729.600 ;
        RECT 208.950 727.950 211.050 730.050 ;
        RECT 221.400 729.600 222.450 736.950 ;
        RECT 245.400 733.050 246.450 755.400 ;
        RECT 247.950 754.950 250.050 757.050 ;
        RECT 244.950 730.950 247.050 733.050 ;
        RECT 190.950 724.950 193.050 727.050 ;
        RECT 193.950 724.950 196.050 727.050 ;
        RECT 196.950 724.950 199.050 727.050 ;
        RECT 199.950 724.950 202.050 727.050 ;
        RECT 194.400 723.900 195.600 724.650 ;
        RECT 200.400 723.900 201.600 724.650 ;
        RECT 209.400 723.900 210.450 727.950 ;
        RECT 221.400 727.350 222.600 729.600 ;
        RECT 241.950 728.100 244.050 730.200 ;
        RECT 248.400 729.600 249.450 754.950 ;
        RECT 242.400 727.350 243.600 728.100 ;
        RECT 248.400 727.350 249.600 729.600 ;
        RECT 251.400 729.450 252.450 760.950 ;
        RECT 254.400 756.900 255.450 766.950 ;
        RECT 263.400 762.600 264.450 799.800 ;
        RECT 275.100 796.800 276.000 809.400 ;
        RECT 281.100 808.800 283.200 810.900 ;
        RECT 284.400 809.100 286.500 811.200 ;
        RECT 276.900 807.000 279.000 807.900 ;
        RECT 276.900 805.800 284.100 807.000 ;
        RECT 282.000 804.900 284.100 805.800 ;
        RECT 276.900 804.000 279.000 804.900 ;
        RECT 285.000 804.000 285.900 809.100 ;
        RECT 287.400 807.450 288.600 807.600 ;
        RECT 287.400 806.400 291.450 807.450 ;
        RECT 287.400 805.350 288.600 806.400 ;
        RECT 276.900 803.100 285.900 804.000 ;
        RECT 276.900 802.800 279.000 803.100 ;
        RECT 281.100 799.950 283.200 802.050 ;
        RECT 281.400 797.400 282.600 799.650 ;
        RECT 274.800 794.700 276.900 796.800 ;
        RECT 285.000 796.500 285.900 803.100 ;
        RECT 286.800 802.950 288.900 805.050 ;
        RECT 283.800 794.400 285.900 796.500 ;
        RECT 290.400 778.050 291.450 806.400 ;
        RECT 289.950 775.950 292.050 778.050 ;
        RECT 299.400 777.450 300.450 835.950 ;
        RECT 308.400 834.900 309.600 835.650 ;
        RECT 323.400 834.900 324.600 835.650 ;
        RECT 329.400 834.900 330.600 835.650 ;
        RECT 307.950 832.800 310.050 834.900 ;
        RECT 322.950 832.800 325.050 834.900 ;
        RECT 328.950 832.800 331.050 834.900 ;
        RECT 323.400 823.050 324.450 832.800 ;
        RECT 325.950 826.950 328.050 829.050 ;
        RECT 331.950 826.950 334.050 829.050 ;
        RECT 319.800 822.000 321.900 823.050 ;
        RECT 319.800 820.950 322.050 822.000 ;
        RECT 322.950 820.950 325.050 823.050 ;
        RECT 319.950 819.450 322.050 820.950 ;
        RECT 319.950 819.000 324.450 819.450 ;
        RECT 320.400 818.400 325.050 819.000 ;
        RECT 322.950 814.950 325.050 818.400 ;
        RECT 313.950 811.950 316.050 814.050 ;
        RECT 314.400 811.200 315.600 811.950 ;
        RECT 309.900 807.900 312.000 809.700 ;
        RECT 313.800 808.800 315.900 810.900 ;
        RECT 317.100 810.300 319.200 812.400 ;
        RECT 308.400 806.700 317.100 807.900 ;
        RECT 305.100 802.950 307.200 805.050 ;
        RECT 305.400 801.450 306.600 802.650 ;
        RECT 302.400 800.400 306.600 801.450 ;
        RECT 302.400 793.050 303.450 800.400 ;
        RECT 308.400 797.700 309.300 806.700 ;
        RECT 315.000 805.800 317.100 806.700 ;
        RECT 318.000 804.900 318.900 810.300 ;
        RECT 326.400 808.200 327.450 826.950 ;
        RECT 332.400 817.050 333.450 826.950 ;
        RECT 331.950 814.950 334.050 817.050 ;
        RECT 335.400 814.050 336.450 859.950 ;
        RECT 338.400 859.050 339.450 865.950 ;
        RECT 359.400 862.050 360.450 892.950 ;
        RECT 367.950 884.100 370.050 886.200 ;
        RECT 368.400 883.350 369.600 884.100 ;
        RECT 364.950 880.950 367.050 883.050 ;
        RECT 367.950 880.950 370.050 883.050 ;
        RECT 365.400 879.900 366.600 880.650 ;
        RECT 364.950 877.800 367.050 879.900 ;
        RECT 358.950 859.950 361.050 862.050 ;
        RECT 370.950 859.950 373.050 862.050 ;
        RECT 337.950 856.950 340.050 859.050 ;
        RECT 355.950 850.950 358.050 853.050 ;
        RECT 349.950 839.100 352.050 841.200 ;
        RECT 350.400 838.350 351.600 839.100 ;
        RECT 343.950 835.950 346.050 838.050 ;
        RECT 346.950 835.950 349.050 838.050 ;
        RECT 349.950 835.950 352.050 838.050 ;
        RECT 347.400 834.900 348.600 835.650 ;
        RECT 346.950 832.800 349.050 834.900 ;
        RECT 356.400 829.050 357.450 850.950 ;
        RECT 364.950 844.950 367.050 847.050 ;
        RECT 358.950 839.100 361.050 841.200 ;
        RECT 365.400 840.600 366.450 844.950 ;
        RECT 371.400 840.600 372.450 859.950 ;
        RECT 359.400 834.450 360.450 839.100 ;
        RECT 365.400 838.350 366.600 840.600 ;
        RECT 371.400 838.350 372.600 840.600 ;
        RECT 364.950 835.950 367.050 838.050 ;
        RECT 367.950 835.950 370.050 838.050 ;
        RECT 370.950 835.950 373.050 838.050 ;
        RECT 373.950 835.950 376.050 838.050 ;
        RECT 368.400 834.900 369.600 835.650 ;
        RECT 359.400 833.400 363.450 834.450 ;
        RECT 349.950 826.950 352.050 829.050 ;
        RECT 355.950 826.950 358.050 829.050 ;
        RECT 350.400 820.050 351.450 826.950 ;
        RECT 349.950 817.950 352.050 820.050 ;
        RECT 328.950 811.950 331.050 814.050 ;
        RECT 334.950 811.950 337.050 814.050 ;
        RECT 319.950 806.100 322.050 808.200 ;
        RECT 325.950 806.100 328.050 808.200 ;
        RECT 320.400 805.350 321.600 806.100 ;
        RECT 312.000 803.700 318.900 804.900 ;
        RECT 312.000 801.300 312.900 803.700 ;
        RECT 310.800 799.200 312.900 801.300 ;
        RECT 313.800 799.950 315.900 802.050 ;
        RECT 307.500 795.600 309.600 797.700 ;
        RECT 314.400 797.400 315.600 799.650 ;
        RECT 317.700 796.500 318.900 803.700 ;
        RECT 319.800 802.950 321.900 805.050 ;
        RECT 322.950 802.950 325.050 805.050 ;
        RECT 317.100 794.400 319.200 796.500 ;
        RECT 301.950 790.950 304.050 793.050 ;
        RECT 307.950 787.950 310.050 790.050 ;
        RECT 299.400 776.400 303.450 777.450 ;
        RECT 271.950 763.950 274.050 766.050 ;
        RECT 263.400 760.350 264.600 762.600 ;
        RECT 259.950 757.950 262.050 760.050 ;
        RECT 262.950 757.950 265.050 760.050 ;
        RECT 265.950 757.950 268.050 760.050 ;
        RECT 253.950 754.800 256.050 756.900 ;
        RECT 260.400 755.400 261.600 757.650 ;
        RECT 266.400 755.400 267.600 757.650 ;
        RECT 260.400 739.050 261.450 755.400 ;
        RECT 266.400 751.050 267.450 755.400 ;
        RECT 265.950 748.950 268.050 751.050 ;
        RECT 272.400 748.050 273.450 763.950 ;
        RECT 277.950 761.100 280.050 763.200 ;
        RECT 286.950 761.100 289.050 763.200 ;
        RECT 292.950 761.100 295.050 763.200 ;
        RECT 298.950 761.100 301.050 766.050 ;
        RECT 278.400 751.050 279.450 761.100 ;
        RECT 287.400 760.350 288.600 761.100 ;
        RECT 293.400 760.350 294.600 761.100 ;
        RECT 283.950 757.950 286.050 760.050 ;
        RECT 286.950 757.950 289.050 760.050 ;
        RECT 289.950 757.950 292.050 760.050 ;
        RECT 292.950 757.950 295.050 760.050 ;
        RECT 295.950 757.950 298.050 760.050 ;
        RECT 284.400 756.900 285.600 757.650 ;
        RECT 283.950 754.800 286.050 756.900 ;
        RECT 290.400 755.400 291.600 757.650 ;
        RECT 296.400 755.400 297.600 757.650 ;
        RECT 277.950 748.950 280.050 751.050 ;
        RECT 290.400 748.050 291.450 755.400 ;
        RECT 271.950 745.950 274.050 748.050 ;
        RECT 289.950 745.950 292.050 748.050 ;
        RECT 280.950 739.950 283.050 742.050 ;
        RECT 259.950 736.950 262.050 739.050 ;
        RECT 259.950 730.950 262.050 735.900 ;
        RECT 271.950 733.950 274.050 736.050 ;
        RECT 272.400 733.200 273.600 733.950 ;
        RECT 267.900 729.900 270.000 731.700 ;
        RECT 271.800 730.800 273.900 732.900 ;
        RECT 275.100 732.300 277.200 734.400 ;
        RECT 251.400 728.400 255.450 729.450 ;
        RECT 215.100 724.950 217.200 727.050 ;
        RECT 220.500 724.950 222.600 727.050 ;
        RECT 223.800 724.950 225.900 727.050 ;
        RECT 238.950 724.950 241.050 727.050 ;
        RECT 241.950 724.950 244.050 727.050 ;
        RECT 244.950 724.950 247.050 727.050 ;
        RECT 247.950 724.950 250.050 727.050 ;
        RECT 193.950 721.800 196.050 723.900 ;
        RECT 199.950 721.800 202.050 723.900 ;
        RECT 208.950 721.800 211.050 723.900 ;
        RECT 215.400 722.400 216.600 724.650 ;
        RECT 224.400 723.900 225.600 724.650 ;
        RECT 239.400 723.900 240.600 724.650 ;
        RECT 245.400 723.900 246.600 724.650 ;
        RECT 254.400 723.900 255.450 728.400 ;
        RECT 259.950 727.800 262.050 729.900 ;
        RECT 266.400 728.700 275.100 729.900 ;
        RECT 202.950 715.950 205.050 718.050 ;
        RECT 196.950 694.950 199.050 697.050 ;
        RECT 164.400 682.350 165.600 683.100 ;
        RECT 179.400 682.350 180.600 683.100 ;
        RECT 185.400 682.350 186.600 684.600 ;
        RECT 160.950 679.950 163.050 682.050 ;
        RECT 163.950 679.950 166.050 682.050 ;
        RECT 178.950 679.950 181.050 682.050 ;
        RECT 181.950 679.950 184.050 682.050 ;
        RECT 184.950 679.950 187.050 682.050 ;
        RECT 135.900 677.100 144.600 678.300 ;
        RECT 161.400 677.400 162.600 679.650 ;
        RECT 182.400 677.400 183.600 679.650 ;
        RECT 133.800 672.600 135.900 674.700 ;
        RECT 137.100 674.100 139.200 676.200 ;
        RECT 141.000 675.300 143.100 677.100 ;
        RECT 137.400 673.050 138.600 673.800 ;
        RECT 136.950 670.950 139.050 673.050 ;
        RECT 161.400 670.050 162.450 677.400 ;
        RECT 160.950 667.950 163.050 670.050 ;
        RECT 182.400 664.050 183.450 677.400 ;
        RECT 181.950 661.950 184.050 664.050 ;
        RECT 145.950 655.950 148.050 658.050 ;
        RECT 182.850 657.300 184.950 659.400 ;
        RECT 133.950 652.950 136.050 655.050 ;
        RECT 107.400 598.050 108.450 650.100 ;
        RECT 119.400 649.350 120.600 650.100 ;
        RECT 125.400 649.350 126.600 650.100 ;
        RECT 127.950 649.950 130.050 652.050 ;
        RECT 130.950 650.100 133.050 652.200 ;
        RECT 118.950 646.950 121.050 649.050 ;
        RECT 121.950 646.950 124.050 649.050 ;
        RECT 124.950 646.950 127.050 649.050 ;
        RECT 122.400 645.900 123.600 646.650 ;
        RECT 121.950 643.800 124.050 645.900 ;
        RECT 124.950 640.950 127.050 643.050 ;
        RECT 125.400 637.050 126.450 640.950 ;
        RECT 131.400 637.050 132.450 650.100 ;
        RECT 134.400 643.050 135.450 652.950 ;
        RECT 139.950 651.000 142.050 655.050 ;
        RECT 146.400 651.600 147.450 655.950 ;
        RECT 140.400 649.350 141.600 651.000 ;
        RECT 146.400 649.350 147.600 651.600 ;
        RECT 154.950 649.950 157.050 652.050 ;
        RECT 169.950 650.100 172.050 652.200 ;
        RECT 139.950 646.950 142.050 649.050 ;
        RECT 142.950 646.950 145.050 649.050 ;
        RECT 145.950 646.950 148.050 649.050 ;
        RECT 148.950 646.950 151.050 649.050 ;
        RECT 136.950 643.950 139.050 646.050 ;
        RECT 143.400 644.400 144.600 646.650 ;
        RECT 149.400 645.900 150.600 646.650 ;
        RECT 155.400 645.900 156.450 649.950 ;
        RECT 170.400 649.350 171.600 650.100 ;
        RECT 166.950 646.950 169.050 649.050 ;
        RECT 169.950 646.950 172.050 649.050 ;
        RECT 172.950 646.950 175.050 649.050 ;
        RECT 178.950 646.950 181.050 649.050 ;
        RECT 133.950 640.950 136.050 643.050 ;
        RECT 124.950 636.450 127.050 637.050 ;
        RECT 122.400 635.400 127.050 636.450 ;
        RECT 110.550 615.300 112.650 617.400 ;
        RECT 110.550 608.700 111.750 615.300 ;
        RECT 110.550 606.600 112.650 608.700 ;
        RECT 106.950 595.950 109.050 598.050 ;
        RECT 110.550 593.700 111.750 606.600 ;
        RECT 115.950 601.950 118.050 604.050 ;
        RECT 116.400 600.900 117.600 601.650 ;
        RECT 115.950 598.800 118.050 600.900 ;
        RECT 110.550 591.600 112.650 593.700 ;
        RECT 106.950 586.950 109.050 589.050 ;
        RECT 98.400 571.350 99.600 572.100 ;
        RECT 103.950 571.950 106.050 574.050 ;
        RECT 107.400 573.600 108.450 586.950 ;
        RECT 112.350 579.300 114.450 581.400 ;
        RECT 107.400 571.350 108.600 573.600 ;
        RECT 97.950 568.950 100.050 571.050 ;
        RECT 106.950 568.950 109.050 571.050 ;
        RECT 92.550 564.300 94.650 566.400 ;
        RECT 103.950 565.950 106.050 568.050 ;
        RECT 113.250 566.400 114.450 579.300 ;
        RECT 115.950 571.950 118.050 574.050 ;
        RECT 122.400 573.450 123.450 635.400 ;
        RECT 124.950 634.950 127.050 635.400 ;
        RECT 130.950 634.950 133.050 637.050 ;
        RECT 130.950 613.950 133.050 616.050 ;
        RECT 124.950 604.950 127.050 607.050 ;
        RECT 125.400 600.900 126.450 604.950 ;
        RECT 131.400 601.050 132.450 613.950 ;
        RECT 137.400 607.200 138.450 643.950 ;
        RECT 143.400 643.050 144.450 644.400 ;
        RECT 148.950 643.800 151.050 645.900 ;
        RECT 154.950 643.800 157.050 645.900 ;
        RECT 167.400 645.000 168.600 646.650 ;
        RECT 173.400 645.900 174.600 646.650 ;
        RECT 142.950 640.950 145.050 643.050 ;
        RECT 166.950 640.950 169.050 645.000 ;
        RECT 172.950 643.800 175.050 645.900 ;
        RECT 179.400 644.400 180.600 646.650 ;
        RECT 143.400 607.200 144.450 640.950 ;
        RECT 179.400 634.050 180.450 644.400 ;
        RECT 183.150 638.700 184.350 657.300 ;
        RECT 193.950 655.950 196.050 658.050 ;
        RECT 188.100 646.950 190.200 649.050 ;
        RECT 188.400 645.900 189.600 646.650 ;
        RECT 194.400 645.900 195.450 655.950 ;
        RECT 187.950 643.800 190.050 645.900 ;
        RECT 193.950 643.800 196.050 645.900 ;
        RECT 183.150 637.500 187.350 638.700 ;
        RECT 190.950 637.950 193.050 640.050 ;
        RECT 185.250 636.600 187.350 637.500 ;
        RECT 178.950 631.950 181.050 634.050 ;
        RECT 191.400 607.200 192.450 637.950 ;
        RECT 197.400 622.050 198.450 694.950 ;
        RECT 203.400 684.600 204.450 715.950 ;
        RECT 209.400 684.600 210.450 721.800 ;
        RECT 215.400 718.050 216.450 722.400 ;
        RECT 223.950 721.800 226.050 723.900 ;
        RECT 238.950 721.800 241.050 723.900 ;
        RECT 244.950 721.800 247.050 723.900 ;
        RECT 253.950 721.800 256.050 723.900 ;
        RECT 239.400 718.050 240.450 721.800 ;
        RECT 260.400 718.050 261.450 727.800 ;
        RECT 263.100 724.950 265.200 727.050 ;
        RECT 263.400 723.900 264.600 724.650 ;
        RECT 262.950 721.800 265.050 723.900 ;
        RECT 266.400 719.700 267.300 728.700 ;
        RECT 273.000 727.800 275.100 728.700 ;
        RECT 276.000 726.900 276.900 732.300 ;
        RECT 277.950 728.100 280.050 730.200 ;
        RECT 278.400 727.350 279.600 728.100 ;
        RECT 270.000 725.700 276.900 726.900 ;
        RECT 270.000 723.300 270.900 725.700 ;
        RECT 268.800 721.200 270.900 723.300 ;
        RECT 271.800 721.950 273.900 724.050 ;
        RECT 214.950 715.950 217.050 718.050 ;
        RECT 238.950 715.950 241.050 718.050 ;
        RECT 259.950 715.950 262.050 718.050 ;
        RECT 265.500 717.600 267.600 719.700 ;
        RECT 272.400 719.400 273.600 721.650 ;
        RECT 275.700 718.500 276.900 725.700 ;
        RECT 277.800 724.950 279.900 727.050 ;
        RECT 275.100 716.400 277.200 718.500 ;
        RECT 259.950 712.800 262.050 714.900 ;
        RECT 226.950 706.950 229.050 709.050 ;
        RECT 220.950 703.950 223.050 706.050 ;
        RECT 217.950 700.950 220.050 703.050 ;
        RECT 203.400 682.350 204.600 684.600 ;
        RECT 209.400 682.350 210.600 684.600 ;
        RECT 202.950 679.950 205.050 682.050 ;
        RECT 205.950 679.950 208.050 682.050 ;
        RECT 208.950 679.950 211.050 682.050 ;
        RECT 211.950 679.950 214.050 682.050 ;
        RECT 206.400 677.400 207.600 679.650 ;
        RECT 212.400 677.400 213.600 679.650 ;
        RECT 206.400 670.050 207.450 677.400 ;
        RECT 205.950 667.950 208.050 670.050 ;
        RECT 212.400 666.450 213.450 677.400 ;
        RECT 218.400 676.050 219.450 700.950 ;
        RECT 217.950 673.950 220.050 676.050 ;
        RECT 217.950 667.950 220.050 670.050 ;
        RECT 212.400 665.400 216.450 666.450 ;
        RECT 211.950 661.950 214.050 664.050 ;
        RECT 200.550 657.300 202.650 659.400 ;
        RECT 200.550 644.400 201.750 657.300 ;
        RECT 205.950 650.100 208.050 652.200 ;
        RECT 206.400 649.350 207.600 650.100 ;
        RECT 205.950 646.950 208.050 649.050 ;
        RECT 200.550 642.300 202.650 644.400 ;
        RECT 200.550 635.700 201.750 642.300 ;
        RECT 200.550 633.600 202.650 635.700 ;
        RECT 212.400 634.050 213.450 661.950 ;
        RECT 211.950 631.950 214.050 634.050 ;
        RECT 196.950 619.950 199.050 622.050 ;
        RECT 215.400 621.450 216.450 665.400 ;
        RECT 218.400 652.050 219.450 667.950 ;
        RECT 217.950 649.950 220.050 652.050 ;
        RECT 215.400 620.400 219.450 621.450 ;
        RECT 202.950 616.950 205.050 619.050 ;
        RECT 197.250 613.500 199.350 614.400 ;
        RECT 195.150 612.300 199.350 613.500 ;
        RECT 136.950 605.100 139.050 607.200 ;
        RECT 142.950 605.100 145.050 607.200 ;
        RECT 148.950 605.100 151.050 607.200 ;
        RECT 137.400 604.350 138.600 605.100 ;
        RECT 143.400 604.350 144.600 605.100 ;
        RECT 136.950 601.950 139.050 604.050 ;
        RECT 139.950 601.950 142.050 604.050 ;
        RECT 142.950 601.950 145.050 604.050 ;
        RECT 124.950 598.800 127.050 600.900 ;
        RECT 130.950 598.950 133.050 601.050 ;
        RECT 140.400 600.900 141.600 601.650 ;
        RECT 139.950 598.800 142.050 600.900 ;
        RECT 149.400 595.050 150.450 605.100 ;
        RECT 154.950 604.950 157.050 607.050 ;
        RECT 163.950 605.100 166.050 607.200 ;
        RECT 190.950 605.100 193.050 607.200 ;
        RECT 142.950 592.950 145.050 595.050 ;
        RECT 148.950 592.950 151.050 595.050 ;
        RECT 139.950 583.950 142.050 586.050 ;
        RECT 130.050 579.300 132.150 581.400 ;
        RECT 119.400 572.400 123.450 573.450 ;
        RECT 88.950 556.950 91.050 559.050 ;
        RECT 92.550 557.700 93.750 564.300 ;
        RECT 92.550 555.600 94.650 557.700 ;
        RECT 104.400 547.050 105.450 565.950 ;
        RECT 112.350 564.300 114.450 566.400 ;
        RECT 113.250 557.700 114.450 564.300 ;
        RECT 112.350 555.600 114.450 557.700 ;
        RECT 103.950 544.950 106.050 547.050 ;
        RECT 85.950 532.950 88.050 535.050 ;
        RECT 82.950 529.950 85.050 532.050 ;
        RECT 86.400 529.200 87.450 532.950 ;
        RECT 88.950 529.950 91.050 532.050 ;
        RECT 116.400 531.450 117.450 571.950 ;
        RECT 113.400 530.400 117.450 531.450 ;
        RECT 73.950 527.100 76.050 529.200 ;
        RECT 79.950 527.100 82.050 529.200 ;
        RECT 85.950 527.100 88.050 529.200 ;
        RECT 74.400 526.350 75.600 527.100 ;
        RECT 80.400 526.350 81.600 527.100 ;
        RECT 73.950 523.950 76.050 526.050 ;
        RECT 76.950 523.950 79.050 526.050 ;
        RECT 79.950 523.950 82.050 526.050 ;
        RECT 82.950 523.950 85.050 526.050 ;
        RECT 77.400 522.900 78.600 523.650 ;
        RECT 83.400 522.900 84.600 523.650 ;
        RECT 89.400 523.050 90.450 529.950 ;
        RECT 91.950 527.100 94.050 529.200 ;
        RECT 100.950 527.100 103.050 529.200 ;
        RECT 106.950 527.100 109.050 529.200 ;
        RECT 76.950 520.800 79.050 522.900 ;
        RECT 82.950 520.800 85.050 522.900 ;
        RECT 88.950 520.950 91.050 523.050 ;
        RECT 64.800 514.950 66.900 517.050 ;
        RECT 67.950 514.950 70.050 517.050 ;
        RECT 49.950 511.950 52.050 514.050 ;
        RECT 58.950 511.950 61.050 514.050 ;
        RECT 79.950 511.950 82.050 514.050 ;
        RECT 55.800 490.950 57.900 493.050 ;
        RECT 56.400 489.000 57.600 490.650 ;
        RECT 55.950 484.950 58.050 489.000 ;
        RECT 46.950 427.950 49.050 430.050 ;
        RECT 44.850 423.300 46.950 425.400 ;
        RECT 31.950 416.100 34.050 418.200 ;
        RECT 32.400 415.350 33.600 416.100 ;
        RECT 31.950 412.950 34.050 415.050 ;
        RECT 40.950 412.950 43.050 415.050 ;
        RECT 41.400 410.400 42.600 412.650 ;
        RECT 26.550 408.300 28.650 410.400 ;
        RECT 26.550 401.700 27.750 408.300 ;
        RECT 31.950 406.950 34.050 409.050 ;
        RECT 26.550 399.600 28.650 401.700 ;
        RECT 32.400 396.450 33.450 406.950 ;
        RECT 41.400 403.050 42.450 410.400 ;
        RECT 45.150 404.700 46.350 423.300 ;
        RECT 50.100 412.950 52.200 415.050 ;
        RECT 50.400 411.000 51.600 412.650 ;
        RECT 49.950 406.950 52.050 411.000 ;
        RECT 52.950 409.950 55.050 412.050 ;
        RECT 45.150 403.500 49.350 404.700 ;
        RECT 40.950 400.950 43.050 403.050 ;
        RECT 47.250 402.600 49.350 403.500 ;
        RECT 29.400 395.400 33.450 396.450 ;
        RECT 20.400 370.350 21.600 372.600 ;
        RECT 16.950 367.950 19.050 370.050 ;
        RECT 19.950 367.950 22.050 370.050 ;
        RECT 29.400 367.050 30.450 395.400 ;
        RECT 37.950 379.950 40.050 382.050 ;
        RECT 49.950 379.950 52.050 382.050 ;
        RECT 38.400 372.600 39.450 379.950 ;
        RECT 38.400 370.350 39.600 372.600 ;
        RECT 43.950 371.100 46.050 373.200 ;
        RECT 44.400 370.350 45.600 371.100 ;
        RECT 34.950 367.950 37.050 370.050 ;
        RECT 37.950 367.950 40.050 370.050 ;
        RECT 40.950 367.950 43.050 370.050 ;
        RECT 43.950 367.950 46.050 370.050 ;
        RECT 28.950 364.950 31.050 367.050 ;
        RECT 35.400 366.450 36.600 367.650 ;
        RECT 41.400 366.900 42.600 367.650 ;
        RECT 32.400 365.400 36.600 366.450 ;
        RECT 4.950 349.950 7.050 352.050 ;
        RECT 25.950 349.950 28.050 352.050 ;
        RECT 16.950 338.100 19.050 340.200 ;
        RECT 17.400 337.350 18.600 338.100 ;
        RECT 13.950 334.950 16.050 337.050 ;
        RECT 16.950 334.950 19.050 337.050 ;
        RECT 19.950 334.950 22.050 337.050 ;
        RECT 20.400 333.900 21.600 334.650 ;
        RECT 19.950 331.800 22.050 333.900 ;
        RECT 2.400 326.400 6.450 327.450 ;
        RECT 5.400 226.050 6.450 326.400 ;
        RECT 20.400 294.600 21.450 331.800 ;
        RECT 26.400 316.050 27.450 349.950 ;
        RECT 32.400 333.450 33.450 365.400 ;
        RECT 40.950 364.800 43.050 366.900 ;
        RECT 40.950 343.950 43.050 346.050 ;
        RECT 41.400 339.600 42.450 343.950 ;
        RECT 43.950 340.950 46.050 343.050 ;
        RECT 41.400 337.350 42.600 339.600 ;
        RECT 35.100 334.950 37.200 337.050 ;
        RECT 40.500 334.950 42.600 337.050 ;
        RECT 35.400 333.900 36.600 334.650 ;
        RECT 34.950 333.450 37.050 333.900 ;
        RECT 32.400 332.400 37.050 333.450 ;
        RECT 34.950 331.800 37.050 332.400 ;
        RECT 25.950 313.950 28.050 316.050 ;
        RECT 26.400 294.600 27.450 313.950 ;
        RECT 32.250 301.500 34.350 302.400 ;
        RECT 30.150 300.300 34.350 301.500 ;
        RECT 20.400 292.350 21.600 294.600 ;
        RECT 26.400 292.350 27.600 294.600 ;
        RECT 13.950 289.950 16.050 292.050 ;
        RECT 16.950 289.950 19.050 292.050 ;
        RECT 19.950 289.950 22.050 292.050 ;
        RECT 25.950 289.950 28.050 292.050 ;
        RECT 17.400 287.400 18.600 289.650 ;
        RECT 17.400 265.050 18.450 287.400 ;
        RECT 30.150 281.700 31.350 300.300 ;
        RECT 44.400 295.200 45.450 340.950 ;
        RECT 50.400 328.050 51.450 379.950 ;
        RECT 53.400 346.050 54.450 409.950 ;
        RECT 56.400 403.050 57.450 484.950 ;
        RECT 59.400 418.200 60.450 511.950 ;
        RECT 68.850 501.300 70.950 503.400 ;
        RECT 64.950 490.950 67.050 493.050 ;
        RECT 65.400 489.000 66.600 490.650 ;
        RECT 64.950 484.950 67.050 489.000 ;
        RECT 65.400 481.050 66.450 484.950 ;
        RECT 69.150 482.700 70.350 501.300 ;
        RECT 74.100 490.950 76.200 493.050 ;
        RECT 74.400 489.900 75.600 490.650 ;
        RECT 73.950 487.800 76.050 489.900 ;
        RECT 69.150 481.500 73.350 482.700 ;
        RECT 64.950 478.950 67.050 481.050 ;
        RECT 71.250 480.600 73.350 481.500 ;
        RECT 80.400 472.050 81.450 511.950 ;
        RECT 83.400 511.050 84.450 520.800 ;
        RECT 92.400 514.050 93.450 527.100 ;
        RECT 101.400 526.350 102.600 527.100 ;
        RECT 107.400 526.350 108.600 527.100 ;
        RECT 97.950 523.950 100.050 526.050 ;
        RECT 100.950 523.950 103.050 526.050 ;
        RECT 103.950 523.950 106.050 526.050 ;
        RECT 106.950 523.950 109.050 526.050 ;
        RECT 98.400 521.400 99.600 523.650 ;
        RECT 104.400 522.900 105.600 523.650 ;
        RECT 98.400 517.050 99.450 521.400 ;
        RECT 103.950 520.800 106.050 522.900 ;
        RECT 97.950 514.950 100.050 517.050 ;
        RECT 91.950 511.950 94.050 514.050 ;
        RECT 82.950 508.950 85.050 511.050 ;
        RECT 83.400 489.900 84.450 508.950 ;
        RECT 86.550 501.300 88.650 503.400 ;
        RECT 104.850 501.300 106.950 503.400 ;
        RECT 82.950 487.800 85.050 489.900 ;
        RECT 86.550 488.400 87.750 501.300 ;
        RECT 91.950 494.100 94.050 496.200 ;
        RECT 92.400 493.350 93.600 494.100 ;
        RECT 91.950 490.950 94.050 493.050 ;
        RECT 100.950 490.950 103.050 493.050 ;
        RECT 101.400 488.400 102.600 490.650 ;
        RECT 79.950 469.950 82.050 472.050 ;
        RECT 83.400 463.050 84.450 487.800 ;
        RECT 86.550 486.300 88.650 488.400 ;
        RECT 86.550 479.700 87.750 486.300 ;
        RECT 101.400 481.050 102.450 488.400 ;
        RECT 105.150 482.700 106.350 501.300 ;
        RECT 113.400 495.450 114.450 530.400 ;
        RECT 115.950 527.100 118.050 529.200 ;
        RECT 116.400 523.050 117.450 527.100 ;
        RECT 115.950 520.950 118.050 523.050 ;
        RECT 113.400 494.400 117.450 495.450 ;
        RECT 110.100 490.950 112.200 493.050 ;
        RECT 110.400 489.900 111.600 490.650 ;
        RECT 109.950 489.450 112.050 489.900 ;
        RECT 109.950 488.400 114.450 489.450 ;
        RECT 109.950 487.800 112.050 488.400 ;
        RECT 113.400 484.050 114.450 488.400 ;
        RECT 105.150 481.500 109.350 482.700 ;
        RECT 112.950 481.950 115.050 484.050 ;
        RECT 86.550 477.600 88.650 479.700 ;
        RECT 100.950 478.950 103.050 481.050 ;
        RECT 107.250 480.600 109.350 481.500 ;
        RECT 97.950 463.950 100.050 466.050 ;
        RECT 82.950 460.950 85.050 463.050 ;
        RECT 83.400 457.050 84.450 460.950 ;
        RECT 61.950 454.950 64.050 457.050 ;
        RECT 82.950 454.950 85.050 457.050 ;
        RECT 62.400 450.600 63.450 454.950 ;
        RECT 76.950 451.950 79.050 454.050 ;
        RECT 62.400 448.350 63.600 450.600 ;
        RECT 62.100 445.950 64.200 448.050 ;
        RECT 67.500 445.950 69.600 448.050 ;
        RECT 68.400 443.400 69.600 445.650 ;
        RECT 68.400 436.050 69.450 443.400 ;
        RECT 77.400 442.050 78.450 451.950 ;
        RECT 83.400 450.600 84.450 454.950 ;
        RECT 83.400 448.350 84.600 450.600 ;
        RECT 88.950 449.100 91.050 451.200 ;
        RECT 94.950 449.100 97.050 451.200 ;
        RECT 89.400 448.350 90.600 449.100 ;
        RECT 82.950 445.950 85.050 448.050 ;
        RECT 85.950 445.950 88.050 448.050 ;
        RECT 88.950 445.950 91.050 448.050 ;
        RECT 86.400 444.000 87.600 445.650 ;
        RECT 76.950 439.950 79.050 442.050 ;
        RECT 85.950 439.950 88.050 444.000 ;
        RECT 67.950 433.950 70.050 436.050 ;
        RECT 85.950 427.950 88.050 430.050 ;
        RECT 62.550 423.300 64.650 425.400 ;
        RECT 58.950 416.100 61.050 418.200 ;
        RECT 55.950 400.950 58.050 403.050 ;
        RECT 56.400 379.050 57.450 400.950 ;
        RECT 59.400 397.050 60.450 416.100 ;
        RECT 62.550 410.400 63.750 423.300 ;
        RECT 76.950 421.950 79.050 424.050 ;
        RECT 67.950 416.100 70.050 418.200 ;
        RECT 68.400 415.350 69.600 416.100 ;
        RECT 73.950 415.950 76.050 418.050 ;
        RECT 67.950 412.950 70.050 415.050 ;
        RECT 62.550 408.300 64.650 410.400 ;
        RECT 62.550 401.700 63.750 408.300 ;
        RECT 74.400 406.050 75.450 415.950 ;
        RECT 73.950 403.950 76.050 406.050 ;
        RECT 62.550 399.600 64.650 401.700 ;
        RECT 77.400 400.050 78.450 421.950 ;
        RECT 86.400 417.600 87.450 427.950 ;
        RECT 95.400 424.050 96.450 449.100 ;
        RECT 98.400 445.050 99.450 463.950 ;
        RECT 109.950 457.950 112.050 460.050 ;
        RECT 103.950 450.000 106.050 454.050 ;
        RECT 110.400 450.600 111.450 457.950 ;
        RECT 116.400 451.050 117.450 494.400 ;
        RECT 104.400 448.350 105.600 450.000 ;
        RECT 110.400 448.350 111.600 450.600 ;
        RECT 115.950 448.950 118.050 451.050 ;
        RECT 103.950 445.950 106.050 448.050 ;
        RECT 106.950 445.950 109.050 448.050 ;
        RECT 109.950 445.950 112.050 448.050 ;
        RECT 112.950 445.950 115.050 448.050 ;
        RECT 97.950 442.950 100.050 445.050 ;
        RECT 107.400 444.900 108.600 445.650 ;
        RECT 113.400 445.050 114.600 445.650 ;
        RECT 106.950 442.800 109.050 444.900 ;
        RECT 113.400 443.400 118.050 445.050 ;
        RECT 119.400 444.900 120.450 572.400 ;
        RECT 124.800 568.950 126.900 571.050 ;
        RECT 125.400 567.900 126.600 568.650 ;
        RECT 124.950 565.800 127.050 567.900 ;
        RECT 130.650 560.700 131.850 579.300 ;
        RECT 133.950 568.950 136.050 571.050 ;
        RECT 134.400 567.450 135.600 568.650 ;
        RECT 140.400 567.450 141.450 583.950 ;
        RECT 134.400 566.400 141.450 567.450 ;
        RECT 127.650 559.500 131.850 560.700 ;
        RECT 127.650 558.600 129.750 559.500 ;
        RECT 139.950 547.950 142.050 550.050 ;
        RECT 124.950 544.950 127.050 547.050 ;
        RECT 125.400 528.600 126.450 544.950 ;
        RECT 125.400 526.350 126.600 528.600 ;
        RECT 130.950 527.100 133.050 529.200 ;
        RECT 131.400 526.350 132.600 527.100 ;
        RECT 124.950 523.950 127.050 526.050 ;
        RECT 127.950 523.950 130.050 526.050 ;
        RECT 130.950 523.950 133.050 526.050 ;
        RECT 133.950 523.950 136.050 526.050 ;
        RECT 128.400 522.900 129.600 523.650 ;
        RECT 127.950 520.800 130.050 522.900 ;
        RECT 134.400 521.400 135.600 523.650 ;
        RECT 134.400 511.050 135.450 521.400 ;
        RECT 133.950 508.950 136.050 511.050 ;
        RECT 122.550 501.300 124.650 503.400 ;
        RECT 122.550 488.400 123.750 501.300 ;
        RECT 127.950 499.950 130.050 502.050 ;
        RECT 128.400 495.600 129.450 499.950 ;
        RECT 134.400 496.200 135.450 508.950 ;
        RECT 128.400 493.350 129.600 495.600 ;
        RECT 133.950 494.100 136.050 496.200 ;
        RECT 127.950 490.950 130.050 493.050 ;
        RECT 122.550 486.300 124.650 488.400 ;
        RECT 122.550 479.700 123.750 486.300 ;
        RECT 122.550 477.600 124.650 479.700 ;
        RECT 124.950 469.950 127.050 472.050 ;
        RECT 121.950 460.950 124.050 463.050 ;
        RECT 122.400 445.050 123.450 460.950 ;
        RECT 125.400 454.050 126.450 469.950 ;
        RECT 140.400 460.050 141.450 547.950 ;
        RECT 143.400 523.050 144.450 592.950 ;
        RECT 155.400 586.050 156.450 604.950 ;
        RECT 164.400 604.350 165.600 605.100 ;
        RECT 191.400 604.350 192.600 605.100 ;
        RECT 164.100 601.950 166.200 604.050 ;
        RECT 182.100 601.950 184.200 604.050 ;
        RECT 190.950 601.950 193.050 604.050 ;
        RECT 195.150 593.700 196.350 612.300 ;
        RECT 200.400 606.450 201.600 606.600 ;
        RECT 203.400 606.450 204.450 616.950 ;
        RECT 200.400 605.400 204.450 606.450 ;
        RECT 212.550 615.300 214.650 617.400 ;
        RECT 212.550 608.700 213.750 615.300 ;
        RECT 218.400 613.050 219.450 620.400 ;
        RECT 217.950 610.950 220.050 613.050 ;
        RECT 212.550 606.600 214.650 608.700 ;
        RECT 200.400 604.350 201.600 605.400 ;
        RECT 200.100 601.950 202.200 604.050 ;
        RECT 194.850 591.600 196.950 593.700 ;
        RECT 205.950 592.950 208.050 595.050 ;
        RECT 212.550 593.700 213.750 606.600 ;
        RECT 221.400 606.450 222.450 703.950 ;
        RECT 227.400 697.050 228.450 706.950 ;
        RECT 229.950 697.950 232.050 700.050 ;
        RECT 256.950 697.950 259.050 700.050 ;
        RECT 226.950 694.950 229.050 697.050 ;
        RECT 230.400 684.600 231.450 697.950 ;
        RECT 230.400 682.350 231.600 684.600 ;
        RECT 235.950 683.100 238.050 685.200 ;
        RECT 244.950 683.100 247.050 685.200 ;
        RECT 250.950 683.100 253.050 685.200 ;
        RECT 257.400 684.600 258.450 697.950 ;
        RECT 260.400 694.050 261.450 712.800 ;
        RECT 259.950 691.950 262.050 694.050 ;
        RECT 281.400 684.600 282.450 739.950 ;
        RECT 283.950 736.950 286.050 739.050 ;
        RECT 284.400 724.050 285.450 736.950 ;
        RECT 296.400 736.050 297.450 755.400 ;
        RECT 302.400 748.050 303.450 776.400 ;
        RECT 304.950 775.950 307.050 778.050 ;
        RECT 305.400 756.900 306.450 775.950 ;
        RECT 308.400 762.450 309.450 787.950 ;
        RECT 323.400 781.050 324.450 802.950 ;
        RECT 329.400 802.050 330.450 811.950 ;
        RECT 362.400 808.050 363.450 833.400 ;
        RECT 367.950 832.800 370.050 834.900 ;
        RECT 374.400 833.400 375.600 835.650 ;
        RECT 374.400 817.050 375.450 833.400 ;
        RECT 376.950 817.950 379.050 820.050 ;
        RECT 373.950 814.950 376.050 817.050 ;
        RECT 355.950 805.950 358.050 808.050 ;
        RECT 361.950 805.950 364.050 808.050 ;
        RECT 367.950 806.100 370.050 808.200 ;
        RECT 334.950 802.950 337.050 805.050 ;
        RECT 337.950 802.950 340.050 805.050 ;
        RECT 340.950 802.950 343.050 805.050 ;
        RECT 343.950 802.950 346.050 805.050 ;
        RECT 346.950 802.950 349.050 805.050 ;
        RECT 328.950 799.950 331.050 802.050 ;
        RECT 335.400 801.000 336.600 802.650 ;
        RECT 341.400 801.900 342.600 802.650 ;
        RECT 328.950 796.800 331.050 798.900 ;
        RECT 334.950 796.950 337.050 801.000 ;
        RECT 340.950 799.800 343.050 801.900 ;
        RECT 347.400 800.400 348.600 802.650 ;
        RECT 325.950 787.950 328.050 790.050 ;
        RECT 322.950 778.950 325.050 781.050 ;
        RECT 326.400 769.050 327.450 787.950 ;
        RECT 329.400 787.050 330.450 796.800 ;
        RECT 347.400 793.050 348.450 800.400 ;
        RECT 349.950 799.950 352.050 802.050 ;
        RECT 346.950 790.950 349.050 793.050 ;
        RECT 350.400 787.050 351.450 799.950 ;
        RECT 328.950 784.950 331.050 787.050 ;
        RECT 349.950 784.950 352.050 787.050 ;
        RECT 325.950 766.950 328.050 769.050 ;
        RECT 311.400 762.450 312.600 762.600 ;
        RECT 308.400 761.400 312.600 762.450 ;
        RECT 311.400 760.350 312.600 761.400 ;
        RECT 310.950 757.950 313.050 760.050 ;
        RECT 313.950 757.950 316.050 760.050 ;
        RECT 316.950 757.950 319.050 760.050 ;
        RECT 304.800 754.800 306.900 756.900 ;
        RECT 307.950 751.950 310.050 757.050 ;
        RECT 314.400 756.900 315.600 757.650 ;
        RECT 313.950 754.800 316.050 756.900 ;
        RECT 301.950 745.950 304.050 748.050 ;
        RECT 298.950 739.950 301.050 742.050 ;
        RECT 295.950 733.950 298.050 736.050 ;
        RECT 296.400 729.600 297.450 733.950 ;
        RECT 299.400 733.050 300.450 739.950 ;
        RECT 298.950 730.950 301.050 733.050 ;
        RECT 314.400 730.200 315.450 754.800 ;
        RECT 296.400 727.350 297.600 729.600 ;
        RECT 301.950 728.100 304.050 730.200 ;
        RECT 313.950 728.100 316.050 730.200 ;
        RECT 302.400 727.350 303.600 728.100 ;
        RECT 295.950 724.950 298.050 727.050 ;
        RECT 298.950 724.950 301.050 727.050 ;
        RECT 301.950 724.950 304.050 727.050 ;
        RECT 283.950 721.950 286.050 724.050 ;
        RECT 299.400 723.900 300.600 724.650 ;
        RECT 298.950 721.800 301.050 723.900 ;
        RECT 314.400 688.050 315.450 728.100 ;
        RECT 317.100 724.950 319.200 727.050 ;
        RECT 320.400 724.950 322.500 727.050 ;
        RECT 325.800 724.950 327.900 727.050 ;
        RECT 317.400 722.400 318.600 724.650 ;
        RECT 326.400 724.050 327.600 724.650 ;
        RECT 329.400 724.050 330.450 784.950 ;
        RECT 356.400 784.050 357.450 805.950 ;
        RECT 368.400 805.350 369.600 806.100 ;
        RECT 364.950 802.950 367.050 805.050 ;
        RECT 367.950 802.950 370.050 805.050 ;
        RECT 370.950 802.950 373.050 805.050 ;
        RECT 365.400 800.400 366.600 802.650 ;
        RECT 371.400 801.900 372.600 802.650 ;
        RECT 370.950 801.450 373.050 801.900 ;
        RECT 370.950 800.400 375.450 801.450 ;
        RECT 358.950 790.800 361.050 792.900 ;
        RECT 355.950 781.950 358.050 784.050 ;
        RECT 349.950 775.950 352.050 778.050 ;
        RECT 337.950 764.100 340.050 769.050 ;
        RECT 337.950 760.950 340.050 763.050 ;
        RECT 343.950 761.100 346.050 766.050 ;
        RECT 338.400 760.350 339.600 760.950 ;
        RECT 344.400 760.350 345.600 761.100 ;
        RECT 334.950 757.950 337.050 760.050 ;
        RECT 337.950 757.950 340.050 760.050 ;
        RECT 340.950 757.950 343.050 760.050 ;
        RECT 343.950 757.950 346.050 760.050 ;
        RECT 331.950 754.950 334.050 757.050 ;
        RECT 335.400 755.400 336.600 757.650 ;
        RECT 350.400 757.050 351.450 775.950 ;
        RECT 352.950 761.100 355.050 763.200 ;
        RECT 359.400 762.600 360.450 790.800 ;
        RECT 365.400 781.050 366.450 800.400 ;
        RECT 370.950 799.800 373.050 800.400 ;
        RECT 364.950 778.950 367.050 781.050 ;
        RECT 332.400 748.050 333.450 754.950 ;
        RECT 335.400 751.050 336.450 755.400 ;
        RECT 349.950 754.950 352.050 757.050 ;
        RECT 353.400 756.450 354.450 761.100 ;
        RECT 359.400 760.350 360.600 762.600 ;
        RECT 358.950 757.950 361.050 760.050 ;
        RECT 361.950 757.950 364.050 760.050 ;
        RECT 364.950 757.950 367.050 760.050 ;
        RECT 362.400 756.900 363.600 757.650 ;
        RECT 374.400 756.900 375.450 800.400 ;
        RECT 377.400 790.050 378.450 817.950 ;
        RECT 380.400 796.050 381.450 904.950 ;
        RECT 383.400 904.050 384.450 910.950 ;
        RECT 382.950 901.950 385.050 904.050 ;
        RECT 389.400 898.050 390.450 911.400 ;
        RECT 394.950 907.950 397.050 912.000 ;
        RECT 409.950 907.950 412.050 912.000 ;
        RECT 422.400 907.050 423.450 917.100 ;
        RECT 431.400 916.350 432.600 918.600 ;
        RECT 427.950 913.950 430.050 916.050 ;
        RECT 430.950 913.950 433.050 916.050 ;
        RECT 428.400 911.400 429.600 913.650 ;
        RECT 437.400 912.900 438.450 922.950 ;
        RECT 449.400 921.450 450.450 925.950 ;
        RECT 472.950 922.950 475.050 925.050 ;
        RECT 449.400 920.400 453.450 921.450 ;
        RECT 452.400 919.200 453.450 920.400 ;
        RECT 460.950 919.950 463.050 922.050 ;
        RECT 446.400 918.450 447.600 918.600 ;
        RECT 440.400 917.400 447.600 918.450 ;
        RECT 428.400 907.050 429.450 911.400 ;
        RECT 436.950 910.800 439.050 912.900 ;
        RECT 421.950 904.950 424.050 907.050 ;
        RECT 427.950 904.950 430.050 907.050 ;
        RECT 440.400 901.050 441.450 917.400 ;
        RECT 446.400 916.350 447.600 917.400 ;
        RECT 451.950 917.100 454.050 919.200 ;
        RECT 452.400 916.350 453.600 917.100 ;
        RECT 445.950 913.950 448.050 916.050 ;
        RECT 448.950 913.950 451.050 916.050 ;
        RECT 451.950 913.950 454.050 916.050 ;
        RECT 454.950 913.950 457.050 916.050 ;
        RECT 449.400 912.900 450.600 913.650 ;
        RECT 448.950 910.800 451.050 912.900 ;
        RECT 455.400 911.400 456.600 913.650 ;
        RECT 448.950 907.650 451.050 909.750 ;
        RECT 409.950 898.950 412.050 901.050 ;
        RECT 439.950 898.950 442.050 901.050 ;
        RECT 388.950 895.950 391.050 898.050 ;
        RECT 388.950 884.100 391.050 886.200 ;
        RECT 410.400 885.600 411.450 898.950 ;
        RECT 389.400 883.350 390.600 884.100 ;
        RECT 410.400 883.350 411.600 885.600 ;
        RECT 385.950 880.950 388.050 883.050 ;
        RECT 388.950 880.950 391.050 883.050 ;
        RECT 391.950 880.950 394.050 883.050 ;
        RECT 406.950 880.950 409.050 883.050 ;
        RECT 409.950 880.950 412.050 883.050 ;
        RECT 412.950 880.950 415.050 883.050 ;
        RECT 430.950 880.950 433.050 883.050 ;
        RECT 433.950 880.950 436.050 883.050 ;
        RECT 436.950 880.950 439.050 883.050 ;
        RECT 439.950 880.950 442.050 883.050 ;
        RECT 442.950 880.950 445.050 883.050 ;
        RECT 386.400 878.400 387.600 880.650 ;
        RECT 407.400 878.400 408.600 880.650 ;
        RECT 413.400 878.400 414.600 880.650 ;
        RECT 431.400 879.900 432.600 880.650 ;
        RECT 437.400 879.900 438.600 880.650 ;
        RECT 386.400 874.050 387.450 878.400 ;
        RECT 385.950 871.950 388.050 874.050 ;
        RECT 407.400 856.050 408.450 878.400 ;
        RECT 413.400 865.050 414.450 878.400 ;
        RECT 418.950 877.800 421.050 879.900 ;
        RECT 430.950 877.800 433.050 879.900 ;
        RECT 436.950 877.800 439.050 879.900 ;
        RECT 443.400 879.000 444.600 880.650 ;
        RECT 449.400 879.900 450.450 907.650 ;
        RECT 455.400 892.050 456.450 911.400 ;
        RECT 457.950 904.950 460.050 907.050 ;
        RECT 458.400 895.050 459.450 904.950 ;
        RECT 461.400 901.050 462.450 919.950 ;
        RECT 466.950 916.950 469.050 919.050 ;
        RECT 473.400 918.600 474.450 922.950 ;
        RECT 475.950 919.950 478.050 925.050 ;
        RECT 467.400 912.900 468.450 916.950 ;
        RECT 473.400 916.350 474.600 918.600 ;
        RECT 478.950 917.100 481.050 919.200 ;
        RECT 479.400 916.350 480.600 917.100 ;
        RECT 472.950 913.950 475.050 916.050 ;
        RECT 475.950 913.950 478.050 916.050 ;
        RECT 478.950 913.950 481.050 916.050 ;
        RECT 481.950 913.950 484.050 916.050 ;
        RECT 476.400 912.900 477.600 913.650 ;
        RECT 466.950 910.800 469.050 912.900 ;
        RECT 475.950 910.800 478.050 912.900 ;
        RECT 482.400 911.400 483.600 913.650 ;
        RECT 491.400 913.050 492.450 937.950 ;
        RECT 502.950 934.950 505.050 937.050 ;
        RECT 496.950 925.950 499.050 928.050 ;
        RECT 497.400 918.600 498.450 925.950 ;
        RECT 503.400 918.600 504.450 934.950 ;
        RECT 511.950 922.950 514.050 925.050 ;
        RECT 497.400 916.350 498.600 918.600 ;
        RECT 503.400 916.350 504.600 918.600 ;
        RECT 496.950 913.950 499.050 916.050 ;
        RECT 499.950 913.950 502.050 916.050 ;
        RECT 502.950 913.950 505.050 916.050 ;
        RECT 505.950 913.950 508.050 916.050 ;
        RECT 460.950 898.950 463.050 901.050 ;
        RECT 482.400 898.050 483.450 911.400 ;
        RECT 490.950 910.950 493.050 913.050 ;
        RECT 500.400 912.900 501.600 913.650 ;
        RECT 506.400 912.900 507.600 913.650 ;
        RECT 512.400 912.900 513.450 922.950 ;
        RECT 499.950 910.800 502.050 912.900 ;
        RECT 505.950 910.800 508.050 912.900 ;
        RECT 511.950 910.800 514.050 912.900 ;
        RECT 482.400 896.400 487.050 898.050 ;
        RECT 483.000 895.950 487.050 896.400 ;
        RECT 457.950 892.950 460.050 895.050 ;
        RECT 481.950 892.950 484.050 895.050 ;
        RECT 454.950 889.950 457.050 892.050 ;
        RECT 458.400 886.200 459.450 892.950 ;
        RECT 478.950 889.950 481.050 892.050 ;
        RECT 472.950 886.950 475.050 889.050 ;
        RECT 457.950 884.100 460.050 886.200 ;
        RECT 458.400 883.350 459.600 884.100 ;
        RECT 463.950 883.950 466.050 886.050 ;
        RECT 464.400 883.350 465.600 883.950 ;
        RECT 457.950 880.950 460.050 883.050 ;
        RECT 460.950 880.950 463.050 883.050 ;
        RECT 463.950 880.950 466.050 883.050 ;
        RECT 466.950 880.950 469.050 883.050 ;
        RECT 412.950 862.950 415.050 865.050 ;
        RECT 412.950 859.800 415.050 861.900 ;
        RECT 406.950 853.950 409.050 856.050 ;
        RECT 403.950 847.950 406.050 850.050 ;
        RECT 382.950 844.950 385.050 847.050 ;
        RECT 383.400 835.050 384.450 844.950 ;
        RECT 391.950 839.100 394.050 841.200 ;
        RECT 397.950 839.100 400.050 841.200 ;
        RECT 392.400 838.350 393.600 839.100 ;
        RECT 398.400 838.350 399.600 839.100 ;
        RECT 388.950 835.950 391.050 838.050 ;
        RECT 391.950 835.950 394.050 838.050 ;
        RECT 394.950 835.950 397.050 838.050 ;
        RECT 397.950 835.950 400.050 838.050 ;
        RECT 382.950 832.950 385.050 835.050 ;
        RECT 389.400 833.400 390.600 835.650 ;
        RECT 395.400 833.400 396.600 835.650 ;
        RECT 389.400 829.050 390.450 833.400 ;
        RECT 395.400 829.050 396.450 833.400 ;
        RECT 388.950 826.950 391.050 829.050 ;
        RECT 394.950 826.950 397.050 829.050 ;
        RECT 391.950 822.450 394.050 823.050 ;
        RECT 397.950 822.450 400.050 823.050 ;
        RECT 391.950 821.400 400.050 822.450 ;
        RECT 391.950 820.950 394.050 821.400 ;
        RECT 397.950 820.950 400.050 821.400 ;
        RECT 397.950 811.950 400.050 814.050 ;
        RECT 391.950 806.100 394.050 808.200 ;
        RECT 392.400 805.350 393.600 806.100 ;
        RECT 388.950 802.950 391.050 805.050 ;
        RECT 391.950 802.950 394.050 805.050 ;
        RECT 389.400 801.900 390.600 802.650 ;
        RECT 388.950 799.800 391.050 801.900 ;
        RECT 398.400 801.450 399.450 811.950 ;
        RECT 404.400 808.200 405.450 847.950 ;
        RECT 413.400 840.600 414.450 859.800 ;
        RECT 419.400 853.050 420.450 877.800 ;
        RECT 442.950 871.950 445.050 879.000 ;
        RECT 448.950 877.800 451.050 879.900 ;
        RECT 461.400 878.400 462.600 880.650 ;
        RECT 467.400 879.900 468.600 880.650 ;
        RECT 418.950 850.950 421.050 853.050 ;
        RECT 442.950 850.950 445.050 853.050 ;
        RECT 413.400 838.350 414.600 840.600 ;
        RECT 421.950 840.450 424.050 841.200 ;
        RECT 443.400 840.600 444.450 850.950 ;
        RECT 421.950 839.400 426.450 840.450 ;
        RECT 421.950 839.100 424.050 839.400 ;
        RECT 422.400 838.350 423.600 839.100 ;
        RECT 406.950 835.950 409.050 838.050 ;
        RECT 413.100 835.950 415.200 838.050 ;
        RECT 416.400 835.950 418.500 838.050 ;
        RECT 421.800 835.950 423.900 838.050 ;
        RECT 407.400 817.050 408.450 835.950 ;
        RECT 416.400 833.400 417.600 835.650 ;
        RECT 416.400 829.050 417.450 833.400 ;
        RECT 415.950 826.950 418.050 829.050 ;
        RECT 406.950 814.950 409.050 817.050 ;
        RECT 409.950 811.950 412.050 814.050 ;
        RECT 403.950 807.450 406.050 808.200 ;
        RECT 401.400 806.400 406.050 807.450 ;
        RECT 401.400 801.900 402.450 806.400 ;
        RECT 403.950 806.100 406.050 806.400 ;
        RECT 410.400 807.600 411.450 811.950 ;
        RECT 410.400 805.350 411.600 807.600 ;
        RECT 415.950 806.100 418.050 808.200 ;
        RECT 416.400 805.350 417.600 806.100 ;
        RECT 421.950 805.950 424.050 808.050 ;
        RECT 406.950 802.950 409.050 805.050 ;
        RECT 409.950 802.950 412.050 805.050 ;
        RECT 412.950 802.950 415.050 805.050 ;
        RECT 415.950 802.950 418.050 805.050 ;
        RECT 407.400 801.900 408.600 802.650 ;
        RECT 395.400 800.400 399.450 801.450 ;
        RECT 379.950 793.950 382.050 796.050 ;
        RECT 376.950 787.950 379.050 790.050 ;
        RECT 395.400 781.050 396.450 800.400 ;
        RECT 400.950 799.800 403.050 801.900 ;
        RECT 406.950 799.800 409.050 801.900 ;
        RECT 413.400 800.400 414.600 802.650 ;
        RECT 413.400 796.050 414.450 800.400 ;
        RECT 412.950 793.950 415.050 796.050 ;
        RECT 400.950 781.950 403.050 784.050 ;
        RECT 394.950 778.950 397.050 781.050 ;
        RECT 382.950 761.100 385.050 763.200 ;
        RECT 388.950 761.100 391.050 763.200 ;
        RECT 383.400 760.350 384.600 761.100 ;
        RECT 389.400 760.350 390.600 761.100 ;
        RECT 379.950 757.950 382.050 760.050 ;
        RECT 382.950 757.950 385.050 760.050 ;
        RECT 385.950 757.950 388.050 760.050 ;
        RECT 388.950 757.950 391.050 760.050 ;
        RECT 380.400 756.900 381.600 757.650 ;
        RECT 353.400 755.400 357.450 756.450 ;
        RECT 334.950 748.950 337.050 751.050 ;
        RECT 331.950 745.950 334.050 748.050 ;
        RECT 326.400 722.400 331.050 724.050 ;
        RECT 317.400 718.050 318.450 722.400 ;
        RECT 327.000 721.950 331.050 722.400 ;
        RECT 332.400 718.050 333.450 745.950 ;
        RECT 346.950 739.950 349.050 742.050 ;
        RECT 347.400 736.050 348.450 739.950 ;
        RECT 343.800 733.950 345.900 736.050 ;
        RECT 346.950 733.950 349.050 736.050 ;
        RECT 344.400 729.600 345.450 733.950 ;
        RECT 344.400 727.350 345.600 729.600 ;
        RECT 340.950 724.950 343.050 727.050 ;
        RECT 343.950 724.950 346.050 727.050 ;
        RECT 346.950 724.950 349.050 727.050 ;
        RECT 347.400 723.900 348.600 724.650 ;
        RECT 346.950 721.800 349.050 723.900 ;
        RECT 356.400 721.050 357.450 755.400 ;
        RECT 361.950 754.800 364.050 756.900 ;
        RECT 373.950 754.800 376.050 756.900 ;
        RECT 379.950 754.800 382.050 756.900 ;
        RECT 386.400 755.400 387.600 757.650 ;
        RECT 395.400 756.900 396.450 778.950 ;
        RECT 401.400 775.050 402.450 781.950 ;
        RECT 412.950 778.950 415.050 781.050 ;
        RECT 400.950 772.950 403.050 775.050 ;
        RECT 403.950 761.100 406.050 763.200 ;
        RECT 404.400 760.350 405.600 761.100 ;
        RECT 403.950 757.950 406.050 760.050 ;
        RECT 406.950 757.950 409.050 760.050 ;
        RECT 407.400 756.900 408.600 757.650 ;
        RECT 394.950 756.450 397.050 756.900 ;
        RECT 392.400 755.400 397.050 756.450 ;
        RECT 367.950 736.950 370.050 739.050 ;
        RECT 358.950 729.600 363.000 730.050 ;
        RECT 368.400 729.600 369.450 736.950 ;
        RECT 376.950 733.950 379.050 736.050 ;
        RECT 358.950 727.950 363.600 729.600 ;
        RECT 362.400 727.350 363.600 727.950 ;
        RECT 368.400 727.350 369.600 729.600 ;
        RECT 361.950 724.950 364.050 727.050 ;
        RECT 364.950 724.950 367.050 727.050 ;
        RECT 367.950 724.950 370.050 727.050 ;
        RECT 370.950 724.950 373.050 727.050 ;
        RECT 358.950 721.950 361.050 724.050 ;
        RECT 365.400 722.400 366.600 724.650 ;
        RECT 371.400 723.900 372.600 724.650 ;
        RECT 355.950 718.950 358.050 721.050 ;
        RECT 316.950 715.950 319.050 718.050 ;
        RECT 331.950 715.950 334.050 718.050 ;
        RECT 317.400 700.050 318.450 715.950 ;
        RECT 352.950 706.950 355.050 709.050 ;
        RECT 316.950 697.950 319.050 700.050 ;
        RECT 353.400 697.050 354.450 706.950 ;
        RECT 356.400 706.050 357.450 718.950 ;
        RECT 355.950 703.950 358.050 706.050 ;
        RECT 355.950 697.950 358.050 700.050 ;
        RECT 352.950 694.950 355.050 697.050 ;
        RECT 346.950 691.950 349.050 694.050 ;
        RECT 236.400 682.350 237.600 683.100 ;
        RECT 226.950 679.950 229.050 682.050 ;
        RECT 229.950 679.950 232.050 682.050 ;
        RECT 232.950 679.950 235.050 682.050 ;
        RECT 235.950 679.950 238.050 682.050 ;
        RECT 227.400 677.400 228.600 679.650 ;
        RECT 233.400 678.900 234.600 679.650 ;
        RECT 227.400 670.050 228.450 677.400 ;
        RECT 232.950 676.800 235.050 678.900 ;
        RECT 229.950 673.950 232.050 676.050 ;
        RECT 226.950 667.950 229.050 670.050 ;
        RECT 230.400 657.450 231.450 673.950 ;
        RECT 245.400 661.050 246.450 683.100 ;
        RECT 251.400 682.350 252.600 683.100 ;
        RECT 257.400 682.350 258.600 684.600 ;
        RECT 272.400 684.450 273.600 684.600 ;
        RECT 269.400 683.400 273.600 684.450 ;
        RECT 250.950 679.950 253.050 682.050 ;
        RECT 253.950 679.950 256.050 682.050 ;
        RECT 256.950 679.950 259.050 682.050 ;
        RECT 254.400 678.900 255.600 679.650 ;
        RECT 269.400 679.050 270.450 683.400 ;
        RECT 272.400 682.350 273.600 683.400 ;
        RECT 281.400 682.350 282.600 684.600 ;
        RECT 289.950 682.950 292.050 685.050 ;
        RECT 295.950 684.000 298.050 688.050 ;
        RECT 313.950 685.950 316.050 688.050 ;
        RECT 272.100 679.950 274.200 682.050 ;
        RECT 277.500 679.950 279.600 682.050 ;
        RECT 280.800 679.950 282.900 682.050 ;
        RECT 253.950 676.800 256.050 678.900 ;
        RECT 268.950 676.950 271.050 679.050 ;
        RECT 278.400 678.900 279.600 679.650 ;
        RECT 277.950 676.800 280.050 678.900 ;
        RECT 265.950 664.950 268.050 667.050 ;
        RECT 244.950 658.950 247.050 661.050 ;
        RECT 250.950 658.950 253.050 661.050 ;
        RECT 226.800 654.300 228.900 656.400 ;
        RECT 230.400 655.200 231.600 657.450 ;
        RECT 223.950 650.100 226.050 652.200 ;
        RECT 224.400 649.350 225.600 650.100 ;
        RECT 224.100 646.950 226.200 649.050 ;
        RECT 227.100 648.900 228.000 654.300 ;
        RECT 230.100 652.800 232.200 654.900 ;
        RECT 234.000 651.900 236.100 653.700 ;
        RECT 228.900 650.700 237.600 651.900 ;
        RECT 228.900 649.800 231.000 650.700 ;
        RECT 227.100 647.700 234.000 648.900 ;
        RECT 227.100 640.500 228.300 647.700 ;
        RECT 230.100 643.950 232.200 646.050 ;
        RECT 233.100 645.300 234.000 647.700 ;
        RECT 230.400 641.400 231.600 643.650 ;
        RECT 233.100 643.200 235.200 645.300 ;
        RECT 236.700 641.700 237.600 650.700 ;
        RECT 241.950 649.950 244.050 652.050 ;
        RECT 238.800 646.950 240.900 649.050 ;
        RECT 239.400 645.450 240.600 646.650 ;
        RECT 242.400 645.450 243.450 649.950 ;
        RECT 251.400 645.900 252.450 658.950 ;
        RECT 259.950 650.100 262.050 652.200 ;
        RECT 266.400 651.600 267.450 664.950 ;
        RECT 274.950 658.950 277.050 661.050 ;
        RECT 271.950 652.950 274.050 655.050 ;
        RECT 260.400 649.350 261.600 650.100 ;
        RECT 266.400 649.350 267.600 651.600 ;
        RECT 256.950 646.950 259.050 649.050 ;
        RECT 259.950 646.950 262.050 649.050 ;
        RECT 262.950 646.950 265.050 649.050 ;
        RECT 265.950 646.950 268.050 649.050 ;
        RECT 257.400 645.900 258.600 646.650 ;
        RECT 239.400 644.400 243.450 645.450 ;
        RECT 250.950 643.800 253.050 645.900 ;
        RECT 256.950 643.800 259.050 645.900 ;
        RECT 263.400 644.400 264.600 646.650 ;
        RECT 226.800 638.400 228.900 640.500 ;
        RECT 236.400 639.600 238.500 641.700 ;
        RECT 263.400 628.050 264.450 644.400 ;
        RECT 262.950 625.950 265.050 628.050 ;
        RECT 259.950 616.950 262.050 619.050 ;
        RECT 221.400 605.400 225.450 606.450 ;
        RECT 217.950 601.950 220.050 604.050 ;
        RECT 218.400 600.900 219.600 601.650 ;
        RECT 217.950 598.800 220.050 600.900 ;
        RECT 163.950 586.950 166.050 589.050 ;
        RECT 154.950 583.950 157.050 586.050 ;
        RECT 145.950 580.950 148.050 583.050 ;
        RECT 146.400 567.900 147.450 580.950 ;
        RECT 151.950 572.100 154.050 574.200 ;
        RECT 157.950 572.100 160.050 574.200 ;
        RECT 152.400 571.350 153.600 572.100 ;
        RECT 158.400 571.350 159.600 572.100 ;
        RECT 151.950 568.950 154.050 571.050 ;
        RECT 154.950 568.950 157.050 571.050 ;
        RECT 157.950 568.950 160.050 571.050 ;
        RECT 145.950 565.800 148.050 567.900 ;
        RECT 155.400 566.400 156.600 568.650 ;
        RECT 151.950 562.950 154.050 565.050 ;
        RECT 152.400 529.200 153.450 562.950 ;
        RECT 155.400 559.050 156.450 566.400 ;
        RECT 154.950 556.950 157.050 559.050 ;
        RECT 164.400 553.050 165.450 586.950 ;
        RECT 199.950 580.950 202.050 583.050 ;
        RECT 187.950 574.950 190.050 577.050 ;
        RECT 169.950 571.950 172.050 574.050 ;
        RECT 178.950 572.100 181.050 574.200 ;
        RECT 163.950 550.950 166.050 553.050 ;
        RECT 170.400 538.050 171.450 571.950 ;
        RECT 179.400 571.350 180.600 572.100 ;
        RECT 175.950 568.950 178.050 571.050 ;
        RECT 178.950 568.950 181.050 571.050 ;
        RECT 181.950 568.950 184.050 571.050 ;
        RECT 176.400 566.400 177.600 568.650 ;
        RECT 182.400 567.000 183.600 568.650 ;
        RECT 176.400 553.050 177.450 566.400 ;
        RECT 181.950 562.950 184.050 567.000 ;
        RECT 188.400 565.050 189.450 574.950 ;
        RECT 190.950 571.950 193.050 574.050 ;
        RECT 200.400 573.600 201.450 580.950 ;
        RECT 206.400 577.050 207.450 592.950 ;
        RECT 212.550 591.600 214.650 593.700 ;
        RECT 211.950 586.950 214.050 589.050 ;
        RECT 205.950 574.950 208.050 577.050 ;
        RECT 206.400 573.600 207.450 574.950 ;
        RECT 191.400 567.900 192.450 571.950 ;
        RECT 200.400 571.350 201.600 573.600 ;
        RECT 206.400 571.350 207.600 573.600 ;
        RECT 196.950 568.950 199.050 571.050 ;
        RECT 199.950 568.950 202.050 571.050 ;
        RECT 202.950 568.950 205.050 571.050 ;
        RECT 205.950 568.950 208.050 571.050 ;
        RECT 197.400 567.900 198.600 568.650 ;
        RECT 203.400 567.900 204.600 568.650 ;
        RECT 212.400 567.900 213.450 586.950 ;
        RECT 220.950 583.950 223.050 586.050 ;
        RECT 214.950 574.950 217.050 577.050 ;
        RECT 190.950 565.800 193.050 567.900 ;
        RECT 196.950 565.800 199.050 567.900 ;
        RECT 202.950 565.800 205.050 567.900 ;
        RECT 211.950 565.800 214.050 567.900 ;
        RECT 187.950 562.950 190.050 565.050 ;
        RECT 175.950 550.950 178.050 553.050 ;
        RECT 188.400 541.050 189.450 562.950 ;
        RECT 187.950 538.950 190.050 541.050 ;
        RECT 169.950 535.950 172.050 538.050 ;
        RECT 188.250 535.500 190.350 536.400 ;
        RECT 196.950 535.950 199.050 538.050 ;
        RECT 203.550 537.300 205.650 539.400 ;
        RECT 186.150 534.300 190.350 535.500 ;
        RECT 151.950 527.100 154.050 529.200 ;
        RECT 152.400 526.350 153.600 527.100 ;
        RECT 157.950 526.950 160.050 529.050 ;
        RECT 160.950 526.950 166.050 529.050 ;
        RECT 169.950 527.100 172.050 529.200 ;
        RECT 175.950 527.100 178.050 529.200 ;
        RECT 181.950 527.100 184.050 529.200 ;
        RECT 148.950 523.950 151.050 526.050 ;
        RECT 151.950 523.950 154.050 526.050 ;
        RECT 142.950 520.950 145.050 523.050 ;
        RECT 149.400 521.400 150.600 523.650 ;
        RECT 149.400 517.050 150.450 521.400 ;
        RECT 154.950 520.950 157.050 523.050 ;
        RECT 148.950 514.950 151.050 517.050 ;
        RECT 149.400 502.050 150.450 514.950 ;
        RECT 155.400 502.050 156.450 520.950 ;
        RECT 158.400 520.050 159.450 526.950 ;
        RECT 170.400 526.350 171.600 527.100 ;
        RECT 176.400 526.350 177.600 527.100 ;
        RECT 182.400 526.350 183.600 527.100 ;
        RECT 160.950 523.800 163.050 525.900 ;
        RECT 166.950 523.950 169.050 526.050 ;
        RECT 169.950 523.950 172.050 526.050 ;
        RECT 172.950 523.950 175.050 526.050 ;
        RECT 175.950 523.950 178.050 526.050 ;
        RECT 181.950 523.950 184.050 526.050 ;
        RECT 157.950 517.950 160.050 520.050 ;
        RECT 148.950 499.950 151.050 502.050 ;
        RECT 154.950 501.450 157.050 502.050 ;
        RECT 154.950 500.400 159.450 501.450 ;
        RECT 154.950 499.950 157.050 500.400 ;
        RECT 148.950 494.100 151.050 496.200 ;
        RECT 154.950 494.100 157.050 496.200 ;
        RECT 158.400 496.050 159.450 500.400 ;
        RECT 149.400 493.350 150.600 494.100 ;
        RECT 155.400 493.350 156.600 494.100 ;
        RECT 157.950 493.950 160.050 496.050 ;
        RECT 161.400 495.450 162.450 523.800 ;
        RECT 167.400 522.900 168.600 523.650 ;
        RECT 166.950 520.800 169.050 522.900 ;
        RECT 173.400 521.400 174.600 523.650 ;
        RECT 163.950 519.450 166.050 520.050 ;
        RECT 173.400 519.450 174.450 521.400 ;
        RECT 178.950 520.950 181.050 523.050 ;
        RECT 163.950 518.400 174.450 519.450 ;
        RECT 163.950 517.950 166.050 518.400 ;
        RECT 163.950 495.450 166.050 496.200 ;
        RECT 161.400 494.400 166.050 495.450 ;
        RECT 163.950 494.100 166.050 494.400 ;
        RECT 169.950 494.100 172.050 496.200 ;
        RECT 148.950 490.950 151.050 493.050 ;
        RECT 151.950 490.950 154.050 493.050 ;
        RECT 154.950 490.950 157.050 493.050 ;
        RECT 160.950 490.800 163.050 492.900 ;
        RECT 152.400 489.000 153.600 490.650 ;
        RECT 151.950 484.950 154.050 489.000 ;
        RECT 161.400 487.050 162.450 490.800 ;
        RECT 164.400 489.450 165.450 494.100 ;
        RECT 170.400 493.350 171.600 494.100 ;
        RECT 169.950 490.950 172.050 493.050 ;
        RECT 172.950 490.950 175.050 493.050 ;
        RECT 173.400 489.900 174.600 490.650 ;
        RECT 164.400 488.400 168.450 489.450 ;
        RECT 160.950 484.950 163.050 487.050 ;
        RECT 157.950 463.950 163.050 466.050 ;
        RECT 139.950 457.950 142.050 460.050 ;
        RECT 124.950 451.950 127.050 454.050 ;
        RECT 114.000 442.950 118.050 443.400 ;
        RECT 118.950 442.800 121.050 444.900 ;
        RECT 121.950 442.950 124.050 445.050 ;
        RECT 115.950 427.950 118.050 430.050 ;
        RECT 94.950 421.950 97.050 424.050 ;
        RECT 104.850 423.300 106.950 425.400 ;
        RECT 86.400 415.350 87.600 417.600 ;
        RECT 91.950 416.100 94.050 418.200 ;
        RECT 92.400 415.350 93.600 416.100 ;
        RECT 85.950 412.950 88.050 415.050 ;
        RECT 88.950 412.950 91.050 415.050 ;
        RECT 91.950 412.950 94.050 415.050 ;
        RECT 94.950 412.950 97.050 415.050 ;
        RECT 100.950 412.950 103.050 415.050 ;
        RECT 89.400 411.900 90.600 412.650 ;
        RECT 88.950 409.800 91.050 411.900 ;
        RECT 95.400 410.400 96.600 412.650 ;
        RECT 101.400 410.400 102.600 412.650 ;
        RECT 76.950 397.950 79.050 400.050 ;
        RECT 95.400 397.050 96.450 410.400 ;
        RECT 58.950 394.950 61.050 397.050 ;
        RECT 94.950 394.950 97.050 397.050 ;
        RECT 64.950 391.950 67.050 394.050 ;
        RECT 88.950 391.950 91.050 394.050 ;
        RECT 55.950 376.950 58.050 379.050 ;
        RECT 65.400 372.600 66.450 391.950 ;
        RECT 85.950 382.950 88.050 385.050 ;
        RECT 77.250 379.500 79.350 380.400 ;
        RECT 70.950 376.950 73.050 379.050 ;
        RECT 75.150 378.300 79.350 379.500 ;
        RECT 71.400 372.600 72.450 376.950 ;
        RECT 65.400 370.350 66.600 372.600 ;
        RECT 71.400 370.350 72.600 372.600 ;
        RECT 58.950 367.950 61.050 370.050 ;
        RECT 61.950 367.950 64.050 370.050 ;
        RECT 64.950 367.950 67.050 370.050 ;
        RECT 70.950 367.950 73.050 370.050 ;
        RECT 62.400 366.900 63.600 367.650 ;
        RECT 61.950 364.800 64.050 366.900 ;
        RECT 75.150 359.700 76.350 378.300 ;
        RECT 79.950 371.100 82.050 373.200 ;
        RECT 80.400 370.350 81.600 371.100 ;
        RECT 80.100 367.950 82.200 370.050 ;
        RECT 74.850 357.600 76.950 359.700 ;
        RECT 73.950 352.950 76.050 355.050 ;
        RECT 52.950 343.950 55.050 346.050 ;
        RECT 61.950 343.950 64.050 346.050 ;
        RECT 55.950 339.000 58.050 343.050 ;
        RECT 62.400 339.600 63.450 343.950 ;
        RECT 56.400 337.350 57.600 339.000 ;
        RECT 62.400 337.350 63.600 339.600 ;
        RECT 70.950 337.950 73.050 340.050 ;
        RECT 55.950 334.950 58.050 337.050 ;
        RECT 58.950 334.950 61.050 337.050 ;
        RECT 61.950 334.950 64.050 337.050 ;
        RECT 64.950 334.950 67.050 337.050 ;
        RECT 59.400 333.000 60.600 334.650 ;
        RECT 65.400 333.000 66.600 334.650 ;
        RECT 71.400 333.900 72.450 337.950 ;
        RECT 58.950 328.950 61.050 333.000 ;
        RECT 64.950 330.450 67.050 333.000 ;
        RECT 70.950 331.800 73.050 333.900 ;
        RECT 64.950 329.400 69.450 330.450 ;
        RECT 64.950 328.950 67.050 329.400 ;
        RECT 49.950 325.950 52.050 328.050 ;
        RECT 58.950 325.800 61.050 327.900 ;
        RECT 47.550 303.300 49.650 305.400 ;
        RECT 47.550 296.700 48.750 303.300 ;
        RECT 34.950 293.100 37.050 295.200 ;
        RECT 43.950 293.100 46.050 295.200 ;
        RECT 47.550 294.600 49.650 296.700 ;
        RECT 35.400 292.350 36.600 293.100 ;
        RECT 35.100 289.950 37.200 292.050 ;
        RECT 47.550 281.700 48.750 294.600 ;
        RECT 52.950 289.950 55.050 292.050 ;
        RECT 53.400 287.400 54.600 289.650 ;
        RECT 59.400 289.050 60.450 325.800 ;
        RECT 64.950 313.950 67.050 316.050 ;
        RECT 29.850 279.600 31.950 281.700 ;
        RECT 47.550 279.600 49.650 281.700 ;
        RECT 53.400 280.050 54.450 287.400 ;
        RECT 58.950 286.950 61.050 289.050 ;
        RECT 61.950 286.950 64.050 289.050 ;
        RECT 52.950 277.950 55.050 280.050 ;
        RECT 40.950 271.950 43.050 274.050 ;
        RECT 16.950 262.950 19.050 265.050 ;
        RECT 31.950 262.950 34.050 265.050 ;
        RECT 20.400 261.450 21.600 261.600 ;
        RECT 20.400 260.400 24.450 261.450 ;
        RECT 20.400 259.350 21.600 260.400 ;
        RECT 14.100 256.950 16.200 259.050 ;
        RECT 19.500 256.950 21.600 259.050 ;
        RECT 23.400 244.050 24.450 260.400 ;
        RECT 32.400 253.050 33.450 262.950 ;
        RECT 41.400 261.600 42.450 271.950 ;
        RECT 62.400 271.050 63.450 286.950 ;
        RECT 56.850 267.300 58.950 269.400 ;
        RECT 61.950 268.950 64.050 271.050 ;
        RECT 41.400 259.350 42.600 261.600 ;
        RECT 46.950 261.000 49.050 265.050 ;
        RECT 47.400 259.350 48.600 261.000 ;
        RECT 37.950 256.950 40.050 259.050 ;
        RECT 40.950 256.950 43.050 259.050 ;
        RECT 43.950 256.950 46.050 259.050 ;
        RECT 46.950 256.950 49.050 259.050 ;
        RECT 52.950 256.950 55.050 259.050 ;
        RECT 38.400 255.000 39.600 256.650 ;
        RECT 31.950 250.950 34.050 253.050 ;
        RECT 37.950 250.950 40.050 255.000 ;
        RECT 44.400 254.400 45.600 256.650 ;
        RECT 53.400 255.900 54.600 256.650 ;
        RECT 22.950 241.950 25.050 244.050 ;
        RECT 4.950 223.950 7.050 226.050 ;
        RECT 25.950 223.950 28.050 226.050 ;
        RECT 20.400 216.450 21.600 216.600 ;
        RECT 20.400 215.400 24.450 216.450 ;
        RECT 20.400 214.350 21.600 215.400 ;
        RECT 14.400 211.950 16.500 214.050 ;
        RECT 19.800 211.950 21.900 214.050 ;
        RECT 23.400 205.050 24.450 215.400 ;
        RECT 22.950 202.950 25.050 205.050 ;
        RECT 16.950 182.100 19.050 184.200 ;
        RECT 17.400 181.350 18.600 182.100 ;
        RECT 13.950 178.950 16.050 181.050 ;
        RECT 16.950 178.950 19.050 181.050 ;
        RECT 19.950 178.950 22.050 181.050 ;
        RECT 20.400 176.400 21.600 178.650 ;
        RECT 20.400 157.050 21.450 176.400 ;
        RECT 26.400 157.050 27.450 223.950 ;
        RECT 40.950 215.100 43.050 217.200 ;
        RECT 44.400 217.050 45.450 254.400 ;
        RECT 52.950 253.800 55.050 255.900 ;
        RECT 57.150 248.700 58.350 267.300 ;
        RECT 62.400 265.050 63.450 268.950 ;
        RECT 61.950 262.950 64.050 265.050 ;
        RECT 65.400 262.050 66.450 313.950 ;
        RECT 68.400 288.900 69.450 329.400 ;
        RECT 74.400 328.050 75.450 352.950 ;
        RECT 86.400 346.050 87.450 382.950 ;
        RECT 89.400 367.050 90.450 391.950 ;
        RECT 92.550 381.300 94.650 383.400 ;
        RECT 92.550 374.700 93.750 381.300 ;
        RECT 101.400 379.050 102.450 410.400 ;
        RECT 105.150 404.700 106.350 423.300 ;
        RECT 110.100 412.950 112.200 415.050 ;
        RECT 110.400 411.000 111.600 412.650 ;
        RECT 116.400 411.900 117.450 427.950 ;
        RECT 109.950 406.950 112.050 411.000 ;
        RECT 115.950 409.800 118.050 411.900 ;
        RECT 105.150 403.500 109.350 404.700 ;
        RECT 107.250 402.600 109.350 403.500 ;
        RECT 109.950 397.950 112.050 400.050 ;
        RECT 100.950 376.950 103.050 379.050 ;
        RECT 92.550 372.600 94.650 374.700 ;
        RECT 88.950 364.950 91.050 367.050 ;
        RECT 85.950 343.950 88.050 346.050 ;
        RECT 89.400 342.450 90.450 364.950 ;
        RECT 92.550 359.700 93.750 372.600 ;
        RECT 103.950 371.100 106.050 373.200 ;
        RECT 97.950 367.950 100.050 370.050 ;
        RECT 98.400 366.000 99.600 367.650 ;
        RECT 97.950 361.950 100.050 366.000 ;
        RECT 104.400 361.050 105.450 371.100 ;
        RECT 92.550 357.600 94.650 359.700 ;
        RECT 103.950 358.950 106.050 361.050 ;
        RECT 110.400 355.050 111.450 397.950 ;
        RECT 119.400 385.050 120.450 442.800 ;
        RECT 125.400 430.050 126.450 451.950 ;
        RECT 134.400 450.450 135.600 450.600 ;
        RECT 134.400 449.400 138.450 450.450 ;
        RECT 134.400 448.350 135.600 449.400 ;
        RECT 128.400 445.950 130.500 448.050 ;
        RECT 133.800 445.950 135.900 448.050 ;
        RECT 128.400 443.400 129.600 445.650 ;
        RECT 128.400 439.050 129.450 443.400 ;
        RECT 127.950 436.950 130.050 439.050 ;
        RECT 124.950 427.950 127.050 430.050 ;
        RECT 122.550 423.300 124.650 425.400 ;
        RECT 137.400 424.050 138.450 449.400 ;
        RECT 139.950 448.950 142.050 451.050 ;
        RECT 151.950 450.000 154.050 454.050 ;
        RECT 122.550 410.400 123.750 423.300 ;
        RECT 136.950 421.950 139.050 424.050 ;
        RECT 140.400 420.450 141.450 448.950 ;
        RECT 152.400 448.350 153.600 450.000 ;
        RECT 157.950 449.100 160.050 451.200 ;
        RECT 158.400 448.350 159.600 449.100 ;
        RECT 148.950 445.950 151.050 448.050 ;
        RECT 151.950 445.950 154.050 448.050 ;
        RECT 154.950 445.950 157.050 448.050 ;
        RECT 157.950 445.950 160.050 448.050 ;
        RECT 149.400 444.900 150.600 445.650 ;
        RECT 148.950 442.800 151.050 444.900 ;
        RECT 155.400 443.400 156.600 445.650 ;
        RECT 148.950 436.950 151.050 439.050 ;
        RECT 149.400 427.050 150.450 436.950 ;
        RECT 155.400 433.050 156.450 443.400 ;
        RECT 154.950 430.950 157.050 433.050 ;
        RECT 167.400 430.050 168.450 488.400 ;
        RECT 172.950 487.800 175.050 489.900 ;
        RECT 173.400 484.050 174.450 487.800 ;
        RECT 172.950 481.950 175.050 484.050 ;
        RECT 179.400 468.450 180.450 520.950 ;
        RECT 186.150 515.700 187.350 534.300 ;
        RECT 190.950 527.100 193.050 529.200 ;
        RECT 191.400 526.350 192.600 527.100 ;
        RECT 191.100 523.950 193.200 526.050 ;
        RECT 193.950 520.950 196.050 523.050 ;
        RECT 185.850 513.600 187.950 515.700 ;
        RECT 190.950 502.950 193.050 505.050 ;
        RECT 181.950 499.950 184.050 502.050 ;
        RECT 182.400 489.900 183.450 499.950 ;
        RECT 191.400 495.600 192.450 502.950 ;
        RECT 194.400 499.050 195.450 520.950 ;
        RECT 197.400 505.050 198.450 535.950 ;
        RECT 203.550 530.700 204.750 537.300 ;
        RECT 203.550 528.600 205.650 530.700 ;
        RECT 199.950 517.950 202.050 520.050 ;
        RECT 196.950 502.950 199.050 505.050 ;
        RECT 200.400 502.050 201.450 517.950 ;
        RECT 203.550 515.700 204.750 528.600 ;
        RECT 208.950 523.950 211.050 526.050 ;
        RECT 209.400 522.450 210.600 523.650 ;
        RECT 215.400 522.450 216.450 574.950 ;
        RECT 221.400 573.600 222.450 583.950 ;
        RECT 224.400 577.050 225.450 605.400 ;
        RECT 238.950 605.100 241.050 607.200 ;
        RECT 239.400 604.350 240.600 605.100 ;
        RECT 244.800 604.950 246.900 607.050 ;
        RECT 247.950 605.100 250.050 607.200 ;
        RECT 253.950 605.100 256.050 607.200 ;
        RECT 260.400 606.600 261.450 616.950 ;
        RECT 235.950 601.950 238.050 604.050 ;
        RECT 238.950 601.950 241.050 604.050 ;
        RECT 236.400 600.900 237.600 601.650 ;
        RECT 245.400 600.900 246.450 604.950 ;
        RECT 235.950 598.800 238.050 600.900 ;
        RECT 244.950 598.800 247.050 600.900 ;
        RECT 245.400 589.050 246.450 598.800 ;
        RECT 248.400 595.050 249.450 605.100 ;
        RECT 254.400 604.350 255.600 605.100 ;
        RECT 260.400 604.350 261.600 606.600 ;
        RECT 265.950 605.100 268.050 607.200 ;
        RECT 266.400 604.350 267.600 605.100 ;
        RECT 253.950 601.950 256.050 604.050 ;
        RECT 256.950 601.950 259.050 604.050 ;
        RECT 259.950 601.950 262.050 604.050 ;
        RECT 262.950 601.950 265.050 604.050 ;
        RECT 265.950 601.950 268.050 604.050 ;
        RECT 257.400 600.900 258.600 601.650 ;
        RECT 263.400 600.900 264.600 601.650 ;
        RECT 256.950 598.800 259.050 600.900 ;
        RECT 262.950 598.800 265.050 600.900 ;
        RECT 247.950 592.950 250.050 595.050 ;
        RECT 247.950 589.800 250.050 591.900 ;
        RECT 244.950 586.950 247.050 589.050 ;
        RECT 229.950 577.950 232.050 580.050 ;
        RECT 223.950 574.950 226.050 577.050 ;
        RECT 221.400 571.350 222.600 573.600 ;
        RECT 220.950 568.950 223.050 571.050 ;
        RECT 223.950 568.950 226.050 571.050 ;
        RECT 224.400 567.900 225.600 568.650 ;
        RECT 223.950 565.800 226.050 567.900 ;
        RECT 223.950 538.950 226.050 541.050 ;
        RECT 217.950 529.950 220.050 532.050 ;
        RECT 209.400 521.400 216.450 522.450 ;
        RECT 203.550 513.600 205.650 515.700 ;
        RECT 199.950 499.950 202.050 502.050 ;
        RECT 193.950 496.950 196.050 499.050 ;
        RECT 191.400 493.350 192.600 495.600 ;
        RECT 208.950 495.000 211.050 499.050 ;
        RECT 215.400 495.450 216.600 495.600 ;
        RECT 218.400 495.450 219.450 529.950 ;
        RECT 220.950 502.950 223.050 505.050 ;
        RECT 209.400 493.350 210.600 495.000 ;
        RECT 215.400 494.400 219.450 495.450 ;
        RECT 215.400 493.350 216.600 494.400 ;
        RECT 187.950 490.950 190.050 493.050 ;
        RECT 190.950 490.950 193.050 493.050 ;
        RECT 205.950 490.950 208.050 493.050 ;
        RECT 208.950 490.950 211.050 493.050 ;
        RECT 211.950 490.950 214.050 493.050 ;
        RECT 214.950 490.950 217.050 493.050 ;
        RECT 188.400 489.900 189.600 490.650 ;
        RECT 181.950 487.800 184.050 489.900 ;
        RECT 187.950 487.800 190.050 489.900 ;
        RECT 206.400 488.400 207.600 490.650 ;
        RECT 212.400 488.400 213.600 490.650 ;
        RECT 206.400 486.450 207.450 488.400 ;
        RECT 206.400 485.400 210.450 486.450 ;
        RECT 181.950 468.450 184.050 469.050 ;
        RECT 179.400 467.400 184.050 468.450 ;
        RECT 181.950 466.950 184.050 467.400 ;
        RECT 169.950 460.950 172.050 466.050 ;
        RECT 172.950 457.950 175.050 460.050 ;
        RECT 173.400 454.050 174.450 457.950 ;
        RECT 172.950 450.000 175.050 454.050 ;
        RECT 182.400 450.600 183.450 466.950 ;
        RECT 203.550 459.300 205.650 461.400 ;
        RECT 188.250 457.500 190.350 458.400 ;
        RECT 186.150 456.300 190.350 457.500 ;
        RECT 173.400 448.350 174.600 450.000 ;
        RECT 182.400 448.350 183.600 450.600 ;
        RECT 172.950 445.950 175.050 448.050 ;
        RECT 175.950 445.950 178.050 448.050 ;
        RECT 181.950 445.950 184.050 448.050 ;
        RECT 176.400 443.400 177.600 445.650 ;
        RECT 176.400 436.050 177.450 443.400 ;
        RECT 178.950 442.950 181.050 445.050 ;
        RECT 175.950 433.950 178.050 436.050 ;
        RECT 166.950 427.950 169.050 430.050 ;
        RECT 148.950 424.950 151.050 427.050 ;
        RECT 137.400 419.400 141.450 420.450 ;
        RECT 127.950 416.100 130.050 418.200 ;
        RECT 133.950 416.100 136.050 418.200 ;
        RECT 128.400 415.350 129.600 416.100 ;
        RECT 127.950 412.950 130.050 415.050 ;
        RECT 134.400 411.900 135.450 416.100 ;
        RECT 122.550 408.300 124.650 410.400 ;
        RECT 133.950 409.800 136.050 411.900 ;
        RECT 122.550 401.700 123.750 408.300 ;
        RECT 122.550 399.600 124.650 401.700 ;
        RECT 118.950 382.950 121.050 385.050 ;
        RECT 118.950 372.000 121.050 376.050 ;
        RECT 119.400 370.350 120.600 372.000 ;
        RECT 124.950 371.100 127.050 373.200 ;
        RECT 125.400 370.350 126.600 371.100 ;
        RECT 130.950 370.950 133.050 373.050 ;
        RECT 115.950 367.950 118.050 370.050 ;
        RECT 118.950 367.950 121.050 370.050 ;
        RECT 121.950 367.950 124.050 370.050 ;
        RECT 124.950 367.950 127.050 370.050 ;
        RECT 116.400 365.400 117.600 367.650 ;
        RECT 122.400 366.000 123.600 367.650 ;
        RECT 116.400 361.050 117.450 365.400 ;
        RECT 121.950 361.950 124.050 366.000 ;
        RECT 131.400 364.050 132.450 370.950 ;
        RECT 130.950 361.950 133.050 364.050 ;
        RECT 115.950 358.950 118.050 361.050 ;
        RECT 109.950 352.950 112.050 355.050 ;
        RECT 101.850 345.300 103.950 347.400 ;
        RECT 115.950 346.950 118.050 349.050 ;
        RECT 89.400 341.400 93.450 342.450 ;
        RECT 85.950 338.100 88.050 340.200 ;
        RECT 92.400 339.600 93.450 341.400 ;
        RECT 86.400 337.350 87.600 338.100 ;
        RECT 92.400 337.350 93.600 339.600 ;
        RECT 82.950 334.950 85.050 337.050 ;
        RECT 85.950 334.950 88.050 337.050 ;
        RECT 88.950 334.950 91.050 337.050 ;
        RECT 91.950 334.950 94.050 337.050 ;
        RECT 97.950 334.950 100.050 337.050 ;
        RECT 83.400 333.900 84.600 334.650 ;
        RECT 82.950 331.800 85.050 333.900 ;
        RECT 89.400 332.400 90.600 334.650 ;
        RECT 98.400 332.400 99.600 334.650 ;
        RECT 76.950 328.950 79.050 331.050 ;
        RECT 73.950 325.950 76.050 328.050 ;
        RECT 77.400 294.600 78.450 328.950 ;
        RECT 89.400 328.050 90.450 332.400 ;
        RECT 85.800 325.950 87.900 328.050 ;
        RECT 88.950 325.950 91.050 328.050 ;
        RECT 86.400 322.050 87.450 325.950 ;
        RECT 85.950 319.950 88.050 322.050 ;
        RECT 77.400 292.350 78.600 294.600 ;
        RECT 73.950 289.950 76.050 292.050 ;
        RECT 76.950 289.950 79.050 292.050 ;
        RECT 79.950 289.950 82.050 292.050 ;
        RECT 67.950 286.800 70.050 288.900 ;
        RECT 70.950 286.950 73.050 289.050 ;
        RECT 74.400 288.900 75.600 289.650 ;
        RECT 67.950 271.950 70.050 274.050 ;
        RECT 64.950 259.950 67.050 262.050 ;
        RECT 62.100 256.950 64.200 259.050 ;
        RECT 62.400 255.000 63.600 256.650 ;
        RECT 61.950 250.950 64.050 255.000 ;
        RECT 68.400 253.050 69.450 271.950 ;
        RECT 67.950 250.950 70.050 253.050 ;
        RECT 57.150 247.500 61.350 248.700 ;
        RECT 59.250 246.600 61.350 247.500 ;
        RECT 55.950 223.950 58.050 226.050 ;
        RECT 41.400 214.350 42.600 215.100 ;
        RECT 43.950 214.950 46.050 217.050 ;
        RECT 56.400 216.600 57.450 223.950 ;
        RECT 56.400 214.350 57.600 216.600 ;
        RECT 61.950 215.100 64.050 217.200 ;
        RECT 62.400 214.350 63.600 215.100 ;
        RECT 37.950 211.950 40.050 214.050 ;
        RECT 40.950 211.950 43.050 214.050 ;
        RECT 55.950 211.950 58.050 214.050 ;
        RECT 58.950 211.950 61.050 214.050 ;
        RECT 61.950 211.950 64.050 214.050 ;
        RECT 64.950 211.950 67.050 214.050 ;
        RECT 38.400 210.000 39.600 211.650 ;
        RECT 37.950 205.950 40.050 210.000 ;
        RECT 59.400 209.400 60.600 211.650 ;
        RECT 65.400 209.400 66.600 211.650 ;
        RECT 52.950 205.950 55.050 208.050 ;
        RECT 28.950 181.950 31.050 184.050 ;
        RECT 40.950 182.100 43.050 184.200 ;
        RECT 29.400 163.050 30.450 181.950 ;
        RECT 41.400 181.350 42.600 182.100 ;
        RECT 49.950 181.950 52.050 184.050 ;
        RECT 37.950 178.950 40.050 181.050 ;
        RECT 40.950 178.950 43.050 181.050 ;
        RECT 43.950 178.950 46.050 181.050 ;
        RECT 44.400 176.400 45.600 178.650 ;
        RECT 44.400 172.050 45.450 176.400 ;
        RECT 43.950 169.950 46.050 172.050 ;
        RECT 28.950 160.950 31.050 163.050 ;
        RECT 19.950 154.950 22.050 157.050 ;
        RECT 25.950 154.950 28.050 157.050 ;
        RECT 19.950 145.950 22.050 148.050 ;
        RECT 20.400 138.600 21.450 145.950 ;
        RECT 26.400 138.600 27.450 154.950 ;
        RECT 50.400 151.050 51.450 181.950 ;
        RECT 49.950 148.950 52.050 151.050 ;
        RECT 46.950 145.950 49.050 148.050 ;
        RECT 20.400 136.350 21.600 138.600 ;
        RECT 26.400 136.350 27.600 138.600 ;
        RECT 34.950 136.950 37.050 139.050 ;
        RECT 40.950 137.100 43.050 139.200 ;
        RECT 47.400 139.050 48.450 145.950 ;
        RECT 49.950 142.950 52.050 145.050 ;
        RECT 16.950 133.950 19.050 136.050 ;
        RECT 19.950 133.950 22.050 136.050 ;
        RECT 22.950 133.950 25.050 136.050 ;
        RECT 25.950 133.950 28.050 136.050 ;
        RECT 17.400 131.400 18.600 133.650 ;
        RECT 23.400 132.000 24.600 133.650 ;
        RECT 17.400 106.200 18.450 131.400 ;
        RECT 22.950 127.950 25.050 132.000 ;
        RECT 35.400 127.050 36.450 136.950 ;
        RECT 41.400 136.350 42.600 137.100 ;
        RECT 46.950 136.950 49.050 139.050 ;
        RECT 40.950 133.950 43.050 136.050 ;
        RECT 43.950 133.950 46.050 136.050 ;
        RECT 44.400 132.900 45.600 133.650 ;
        RECT 50.400 132.900 51.450 142.950 ;
        RECT 53.400 139.050 54.450 205.950 ;
        RECT 59.400 205.050 60.450 209.400 ;
        RECT 58.950 202.950 61.050 205.050 ;
        RECT 59.400 187.050 60.450 202.950 ;
        RECT 58.950 184.950 61.050 187.050 ;
        RECT 55.950 183.600 60.000 184.050 ;
        RECT 65.400 183.600 66.450 209.400 ;
        RECT 71.400 196.050 72.450 286.950 ;
        RECT 73.950 286.800 76.050 288.900 ;
        RECT 80.400 287.400 81.600 289.650 ;
        RECT 80.400 280.050 81.450 287.400 ;
        RECT 79.950 277.950 82.050 280.050 ;
        RECT 74.550 267.300 76.650 269.400 ;
        RECT 74.550 254.400 75.750 267.300 ;
        RECT 79.950 260.100 82.050 262.200 ;
        RECT 80.400 259.350 81.600 260.100 ;
        RECT 79.950 256.950 82.050 259.050 ;
        RECT 74.550 252.300 76.650 254.400 ;
        RECT 82.950 253.950 85.050 256.050 ;
        RECT 74.550 245.700 75.750 252.300 ;
        RECT 74.550 243.600 76.650 245.700 ;
        RECT 76.950 232.950 79.050 235.050 ;
        RECT 73.950 215.100 76.050 217.200 ;
        RECT 74.400 208.050 75.450 215.100 ;
        RECT 73.950 205.950 76.050 208.050 ;
        RECT 73.950 196.950 76.050 199.050 ;
        RECT 70.950 193.950 73.050 196.050 ;
        RECT 55.950 181.950 60.600 183.600 ;
        RECT 59.400 181.350 60.600 181.950 ;
        RECT 65.400 181.350 66.600 183.600 ;
        RECT 58.950 178.950 61.050 181.050 ;
        RECT 61.950 178.950 64.050 181.050 ;
        RECT 64.950 178.950 67.050 181.050 ;
        RECT 67.950 178.950 70.050 181.050 ;
        RECT 62.400 177.900 63.600 178.650 ;
        RECT 68.400 177.900 69.600 178.650 ;
        RECT 74.400 177.900 75.450 196.950 ;
        RECT 61.950 175.800 64.050 177.900 ;
        RECT 67.950 175.800 70.050 177.900 ;
        RECT 73.950 175.800 76.050 177.900 ;
        RECT 62.400 145.050 63.450 175.800 ;
        RECT 77.400 175.050 78.450 232.950 ;
        RECT 83.400 217.200 84.450 253.950 ;
        RECT 86.400 253.050 87.450 319.950 ;
        RECT 98.400 316.050 99.450 332.400 ;
        RECT 102.150 326.700 103.350 345.300 ;
        RECT 112.950 340.950 115.050 343.050 ;
        RECT 107.100 334.950 109.200 337.050 ;
        RECT 107.400 333.900 108.600 334.650 ;
        RECT 106.950 331.800 109.050 333.900 ;
        RECT 102.150 325.500 106.350 326.700 ;
        RECT 104.250 324.600 106.350 325.500 ;
        RECT 97.950 313.950 100.050 316.050 ;
        RECT 88.950 304.950 91.050 307.050 ;
        RECT 85.950 250.950 88.050 253.050 ;
        RECT 82.950 215.100 85.050 217.200 ;
        RECT 89.400 216.600 90.450 304.950 ;
        RECT 104.400 294.450 105.600 294.600 ;
        RECT 104.400 293.400 108.450 294.450 ;
        RECT 104.400 292.350 105.600 293.400 ;
        RECT 98.400 289.950 100.500 292.050 ;
        RECT 103.800 289.950 105.900 292.050 ;
        RECT 107.400 288.900 108.450 293.400 ;
        RECT 113.400 289.050 114.450 340.950 ;
        RECT 116.400 304.050 117.450 346.950 ;
        RECT 119.550 345.300 121.650 347.400 ;
        RECT 119.550 332.400 120.750 345.300 ;
        RECT 124.950 338.100 127.050 340.200 ;
        RECT 125.400 337.350 126.600 338.100 ;
        RECT 124.950 334.950 127.050 337.050 ;
        RECT 119.550 330.300 121.650 332.400 ;
        RECT 119.550 323.700 120.750 330.300 ;
        RECT 119.550 321.600 121.650 323.700 ;
        RECT 115.950 301.950 118.050 304.050 ;
        RECT 121.950 294.000 124.050 298.050 ;
        RECT 122.400 292.350 123.600 294.000 ;
        RECT 127.950 293.100 130.050 295.200 ;
        RECT 128.400 292.350 129.600 293.100 ;
        RECT 118.950 289.950 121.050 292.050 ;
        RECT 121.950 289.950 124.050 292.050 ;
        RECT 124.950 289.950 127.050 292.050 ;
        RECT 127.950 289.950 130.050 292.050 ;
        RECT 106.950 286.800 109.050 288.900 ;
        RECT 112.950 286.950 115.050 289.050 ;
        RECT 119.400 287.400 120.600 289.650 ;
        RECT 125.400 288.900 126.600 289.650 ;
        RECT 91.950 277.950 94.050 280.050 ;
        RECT 92.400 235.050 93.450 277.950 ;
        RECT 119.400 271.050 120.450 287.400 ;
        RECT 124.950 286.800 127.050 288.900 ;
        RECT 125.400 283.050 126.450 286.800 ;
        RECT 124.950 280.950 127.050 283.050 ;
        RECT 97.950 268.950 100.050 271.050 ;
        RECT 118.950 268.950 121.050 271.050 ;
        RECT 98.400 261.600 99.450 268.950 ;
        RECT 121.950 264.450 124.050 268.050 ;
        RECT 119.400 264.000 124.050 264.450 ;
        RECT 125.400 264.450 126.450 280.950 ;
        RECT 119.400 263.400 123.450 264.000 ;
        RECT 125.400 263.400 129.450 264.450 ;
        RECT 98.400 259.350 99.600 261.600 ;
        RECT 103.950 260.100 106.050 262.200 ;
        RECT 112.950 260.100 115.050 262.200 ;
        RECT 119.400 261.450 120.450 263.400 ;
        RECT 116.400 260.400 120.450 261.450 ;
        RECT 104.400 259.350 105.600 260.100 ;
        RECT 97.950 256.950 100.050 259.050 ;
        RECT 100.950 256.950 103.050 259.050 ;
        RECT 103.950 256.950 106.050 259.050 ;
        RECT 106.950 256.950 109.050 259.050 ;
        RECT 101.400 254.400 102.600 256.650 ;
        RECT 107.400 255.900 108.600 256.650 ;
        RECT 97.950 250.950 100.050 253.050 ;
        RECT 91.950 232.950 94.050 235.050 ;
        RECT 98.400 217.050 99.450 250.950 ;
        RECT 101.400 238.050 102.450 254.400 ;
        RECT 106.950 253.800 109.050 255.900 ;
        RECT 113.400 244.050 114.450 260.100 ;
        RECT 116.400 255.900 117.450 260.400 ;
        RECT 121.950 260.100 124.050 262.200 ;
        RECT 128.400 261.600 129.450 263.400 ;
        RECT 134.400 262.050 135.450 409.800 ;
        RECT 137.400 406.050 138.450 419.400 ;
        RECT 139.950 415.950 142.050 418.050 ;
        RECT 151.950 416.100 154.050 418.200 ;
        RECT 157.950 416.100 160.050 418.200 ;
        RECT 136.950 403.950 139.050 406.050 ;
        RECT 137.400 373.050 138.450 403.950 ;
        RECT 140.400 397.050 141.450 415.950 ;
        RECT 152.400 415.350 153.600 416.100 ;
        RECT 158.400 415.350 159.600 416.100 ;
        RECT 148.950 412.950 151.050 415.050 ;
        RECT 151.950 412.950 154.050 415.050 ;
        RECT 154.950 412.950 157.050 415.050 ;
        RECT 157.950 412.950 160.050 415.050 ;
        RECT 149.400 411.900 150.600 412.650 ;
        RECT 148.950 409.800 151.050 411.900 ;
        RECT 155.400 411.000 156.600 412.650 ;
        RECT 154.950 406.950 157.050 411.000 ;
        RECT 160.950 409.950 163.050 412.050 ;
        RECT 139.950 394.950 142.050 397.050 ;
        RECT 139.950 375.450 144.000 376.050 ;
        RECT 139.950 373.950 144.450 375.450 ;
        RECT 136.950 370.950 139.050 373.050 ;
        RECT 143.400 372.600 144.450 373.950 ;
        RECT 161.400 373.200 162.450 409.950 ;
        RECT 167.400 409.050 168.450 427.950 ;
        RECT 179.400 427.050 180.450 442.950 ;
        RECT 186.150 437.700 187.350 456.300 ;
        RECT 203.550 452.700 204.750 459.300 ;
        RECT 209.400 454.050 210.450 485.400 ;
        RECT 190.950 449.100 193.050 451.200 ;
        RECT 196.950 449.100 199.050 451.200 ;
        RECT 203.550 450.600 205.650 452.700 ;
        RECT 208.950 451.950 211.050 454.050 ;
        RECT 212.400 451.050 213.450 488.400 ;
        RECT 221.400 481.050 222.450 502.950 ;
        RECT 220.950 478.950 223.050 481.050 ;
        RECT 217.950 475.950 220.050 478.050 ;
        RECT 218.400 469.050 219.450 475.950 ;
        RECT 224.400 472.050 225.450 538.950 ;
        RECT 230.400 532.050 231.450 577.950 ;
        RECT 248.400 576.450 249.450 589.800 ;
        RECT 272.400 580.050 273.450 652.950 ;
        RECT 275.400 646.050 276.450 658.950 ;
        RECT 283.950 651.000 286.050 655.050 ;
        RECT 290.400 651.600 291.450 682.950 ;
        RECT 296.400 682.350 297.600 684.000 ;
        RECT 301.950 683.100 304.050 685.200 ;
        RECT 319.950 683.100 322.050 685.200 ;
        RECT 340.950 683.100 343.050 685.200 ;
        RECT 347.400 684.600 348.450 691.950 ;
        RECT 302.400 682.350 303.600 683.100 ;
        RECT 320.400 682.350 321.600 683.100 ;
        RECT 341.400 682.350 342.600 683.100 ;
        RECT 347.400 682.350 348.600 684.600 ;
        RECT 352.950 682.950 355.050 688.050 ;
        RECT 356.400 685.200 357.450 697.950 ;
        RECT 359.400 693.450 360.450 721.950 ;
        RECT 365.400 700.050 366.450 722.400 ;
        RECT 370.950 721.800 373.050 723.900 ;
        RECT 364.950 697.950 367.050 700.050 ;
        RECT 359.400 692.400 363.450 693.450 ;
        RECT 358.950 688.950 361.050 691.050 ;
        RECT 355.950 683.100 358.050 685.200 ;
        RECT 295.950 679.950 298.050 682.050 ;
        RECT 298.950 679.950 301.050 682.050 ;
        RECT 301.950 679.950 304.050 682.050 ;
        RECT 304.950 679.950 307.050 682.050 ;
        RECT 319.950 679.950 322.050 682.050 ;
        RECT 322.950 679.950 325.050 682.050 ;
        RECT 340.950 679.950 343.050 682.050 ;
        RECT 343.950 679.950 346.050 682.050 ;
        RECT 346.950 679.950 349.050 682.050 ;
        RECT 349.950 679.950 352.050 682.050 ;
        RECT 299.400 678.900 300.600 679.650 ;
        RECT 298.950 676.800 301.050 678.900 ;
        RECT 305.400 677.400 306.600 679.650 ;
        RECT 305.400 667.050 306.450 677.400 ;
        RECT 337.950 676.950 340.050 679.050 ;
        RECT 344.400 677.400 345.600 679.650 ;
        RECT 350.400 677.400 351.600 679.650 ;
        RECT 338.400 670.050 339.450 676.950 ;
        RECT 337.950 667.950 340.050 670.050 ;
        RECT 304.950 664.950 307.050 667.050 ;
        RECT 334.950 664.950 337.050 667.050 ;
        RECT 301.350 657.300 303.450 659.400 ;
        RECT 319.050 657.300 321.150 659.400 ;
        RECT 284.400 649.350 285.600 651.000 ;
        RECT 290.400 649.350 291.600 651.600 ;
        RECT 295.950 650.100 298.050 652.200 ;
        RECT 296.400 649.350 297.600 650.100 ;
        RECT 283.950 646.950 286.050 649.050 ;
        RECT 286.950 646.950 289.050 649.050 ;
        RECT 289.950 646.950 292.050 649.050 ;
        RECT 295.950 646.950 298.050 649.050 ;
        RECT 274.950 643.950 277.050 646.050 ;
        RECT 287.400 645.900 288.600 646.650 ;
        RECT 286.950 643.800 289.050 645.900 ;
        RECT 302.250 644.400 303.450 657.300 ;
        RECT 313.800 646.950 315.900 649.050 ;
        RECT 314.400 645.900 315.600 646.650 ;
        RECT 301.350 642.300 303.450 644.400 ;
        RECT 313.950 643.800 316.050 645.900 ;
        RECT 302.250 635.700 303.450 642.300 ;
        RECT 304.950 637.950 307.050 640.050 ;
        RECT 319.650 638.700 320.850 657.300 ;
        RECT 328.950 652.950 331.050 655.050 ;
        RECT 329.400 649.050 330.450 652.950 ;
        RECT 331.950 650.100 334.050 652.200 ;
        RECT 322.950 646.950 325.050 649.050 ;
        RECT 328.950 646.950 331.050 649.050 ;
        RECT 323.400 644.400 324.600 646.650 ;
        RECT 332.400 645.900 333.450 650.100 ;
        RECT 323.400 640.050 324.450 644.400 ;
        RECT 331.950 643.800 334.050 645.900 ;
        RECT 274.950 631.950 277.050 634.050 ;
        RECT 301.350 633.600 303.450 635.700 ;
        RECT 275.400 600.900 276.450 631.950 ;
        RECT 301.350 615.300 303.450 617.400 ;
        RECT 289.950 610.950 292.050 613.050 ;
        RECT 280.950 605.100 283.050 607.200 ;
        RECT 290.400 606.600 291.450 610.950 ;
        RECT 302.250 608.700 303.450 615.300 ;
        RECT 301.350 606.600 303.450 608.700 ;
        RECT 281.400 604.350 282.600 605.100 ;
        RECT 290.400 604.350 291.600 606.600 ;
        RECT 281.100 601.950 283.200 604.050 ;
        RECT 284.400 601.950 286.500 604.050 ;
        RECT 289.800 601.950 291.900 604.050 ;
        RECT 295.950 601.950 298.050 604.050 ;
        RECT 274.950 598.800 277.050 600.900 ;
        RECT 284.400 599.400 285.600 601.650 ;
        RECT 296.400 599.400 297.600 601.650 ;
        RECT 271.950 577.950 274.050 580.050 ;
        RECT 277.950 577.950 280.050 580.050 ;
        RECT 245.400 575.400 249.450 576.450 ;
        RECT 238.950 572.100 241.050 574.200 ;
        RECT 245.400 573.600 246.450 575.400 ;
        RECT 239.400 571.350 240.600 572.100 ;
        RECT 245.400 571.350 246.600 573.600 ;
        RECT 253.800 572.100 255.900 574.200 ;
        RECT 238.950 568.950 241.050 571.050 ;
        RECT 241.950 568.950 244.050 571.050 ;
        RECT 244.950 568.950 247.050 571.050 ;
        RECT 247.950 568.950 250.050 571.050 ;
        RECT 242.400 567.900 243.600 568.650 ;
        RECT 248.400 567.900 249.600 568.650 ;
        RECT 241.950 565.800 244.050 567.900 ;
        RECT 247.950 565.800 250.050 567.900 ;
        RECT 232.950 550.950 235.050 553.050 ;
        RECT 229.950 529.950 232.050 532.050 ;
        RECT 233.400 528.600 234.450 550.950 ;
        RECT 233.400 526.350 234.600 528.600 ;
        RECT 238.950 528.000 241.050 532.050 ;
        RECT 242.400 529.200 243.450 565.800 ;
        RECT 254.400 565.050 255.450 572.100 ;
        RECT 256.950 571.950 259.050 574.050 ;
        RECT 268.950 572.100 271.050 574.200 ;
        RECT 257.400 567.900 258.450 571.950 ;
        RECT 269.400 571.350 270.600 572.100 ;
        RECT 265.950 568.950 268.050 571.050 ;
        RECT 268.950 568.950 271.050 571.050 ;
        RECT 271.950 568.950 274.050 571.050 ;
        RECT 256.950 565.800 259.050 567.900 ;
        RECT 266.400 567.000 267.600 568.650 ;
        RECT 272.400 567.900 273.600 568.650 ;
        RECT 278.400 567.900 279.450 577.950 ;
        RECT 280.950 571.950 283.050 574.050 ;
        RECT 253.950 562.950 256.050 565.050 ;
        RECT 265.950 562.950 268.050 567.000 ;
        RECT 271.950 565.800 274.050 567.900 ;
        RECT 277.950 565.800 280.050 567.900 ;
        RECT 259.950 544.950 262.050 547.050 ;
        RECT 260.400 538.050 261.450 544.950 ;
        RECT 259.950 535.950 262.050 538.050 ;
        RECT 244.950 529.950 247.050 532.050 ;
        RECT 281.400 531.450 282.450 571.950 ;
        RECT 284.400 565.050 285.450 599.400 ;
        RECT 296.400 589.050 297.450 599.400 ;
        RECT 302.250 593.700 303.450 606.600 ;
        RECT 301.350 591.600 303.450 593.700 ;
        RECT 295.950 586.950 298.050 589.050 ;
        RECT 305.400 586.050 306.450 637.950 ;
        RECT 316.650 637.500 320.850 638.700 ;
        RECT 322.950 637.950 325.050 640.050 ;
        RECT 316.650 636.600 318.750 637.500 ;
        RECT 316.650 613.500 318.750 614.400 ;
        RECT 316.650 612.300 320.850 613.500 ;
        RECT 307.950 604.950 310.050 607.050 ;
        RECT 313.950 605.100 316.050 607.200 ;
        RECT 308.400 592.050 309.450 604.950 ;
        RECT 314.400 604.350 315.600 605.100 ;
        RECT 313.800 601.950 315.900 604.050 ;
        RECT 319.650 593.700 320.850 612.300 ;
        RECT 323.400 606.600 324.450 637.950 ;
        RECT 323.400 604.350 324.600 606.600 ;
        RECT 322.950 601.950 325.050 604.050 ;
        RECT 307.950 589.950 310.050 592.050 ;
        RECT 319.050 591.600 321.150 593.700 ;
        RECT 332.400 589.050 333.450 643.800 ;
        RECT 319.950 586.950 322.050 589.050 ;
        RECT 331.950 586.950 334.050 589.050 ;
        RECT 298.950 583.950 301.050 586.050 ;
        RECT 304.950 583.950 307.050 586.050 ;
        RECT 292.950 572.100 295.050 574.200 ;
        RECT 299.400 574.050 300.450 583.950 ;
        RECT 305.850 579.300 307.950 581.400 ;
        RECT 293.400 571.350 294.600 572.100 ;
        RECT 298.950 571.950 301.050 574.050 ;
        RECT 289.950 568.950 292.050 571.050 ;
        RECT 292.950 568.950 295.050 571.050 ;
        RECT 295.950 568.950 298.050 571.050 ;
        RECT 301.950 568.950 304.050 571.050 ;
        RECT 290.400 566.400 291.600 568.650 ;
        RECT 296.400 566.400 297.600 568.650 ;
        RECT 302.400 567.900 303.600 568.650 ;
        RECT 290.400 565.050 291.450 566.400 ;
        RECT 283.950 562.950 286.050 565.050 ;
        RECT 289.950 562.950 292.050 565.050 ;
        RECT 290.400 547.050 291.450 562.950 ;
        RECT 296.400 562.050 297.450 566.400 ;
        RECT 301.950 565.800 304.050 567.900 ;
        RECT 295.950 559.950 298.050 562.050 ;
        RECT 306.150 560.700 307.350 579.300 ;
        RECT 311.100 568.950 313.200 571.050 ;
        RECT 311.400 567.900 312.600 568.650 ;
        RECT 310.950 565.800 313.050 567.900 ;
        RECT 320.400 562.050 321.450 586.950 ;
        RECT 323.550 579.300 325.650 581.400 ;
        RECT 323.550 566.400 324.750 579.300 ;
        RECT 328.950 572.100 331.050 574.200 ;
        RECT 329.400 571.350 330.600 572.100 ;
        RECT 328.950 568.950 331.050 571.050 ;
        RECT 323.550 564.300 325.650 566.400 ;
        RECT 306.150 559.500 310.350 560.700 ;
        RECT 319.950 559.950 322.050 562.050 ;
        RECT 308.250 558.600 310.350 559.500 ;
        RECT 323.550 557.700 324.750 564.300 ;
        RECT 323.550 555.600 325.650 557.700 ;
        RECT 335.400 556.050 336.450 664.950 ;
        RECT 344.400 655.050 345.450 677.400 ;
        RECT 350.400 673.050 351.450 677.400 ;
        RECT 356.400 673.050 357.450 683.100 ;
        RECT 359.400 678.900 360.450 688.950 ;
        RECT 362.400 684.450 363.450 692.400 ;
        RECT 377.400 691.050 378.450 733.950 ;
        RECT 380.400 733.050 381.450 754.800 ;
        RECT 382.950 751.950 385.050 754.050 ;
        RECT 383.400 745.050 384.450 751.950 ;
        RECT 382.950 742.950 385.050 745.050 ;
        RECT 386.400 736.050 387.450 755.400 ;
        RECT 392.400 739.050 393.450 755.400 ;
        RECT 394.950 754.800 397.050 755.400 ;
        RECT 406.950 754.800 409.050 756.900 ;
        RECT 413.400 751.050 414.450 778.950 ;
        RECT 422.400 766.050 423.450 805.950 ;
        RECT 425.400 775.050 426.450 839.400 ;
        RECT 443.400 838.350 444.600 840.600 ;
        RECT 436.950 835.950 439.050 838.050 ;
        RECT 439.950 835.950 442.050 838.050 ;
        RECT 442.950 835.950 445.050 838.050 ;
        RECT 440.400 834.900 441.600 835.650 ;
        RECT 439.950 832.800 442.050 834.900 ;
        RECT 440.400 823.050 441.450 832.800 ;
        RECT 449.400 826.050 450.450 877.800 ;
        RECT 451.950 874.950 454.050 877.050 ;
        RECT 452.400 859.050 453.450 874.950 ;
        RECT 461.400 874.050 462.450 878.400 ;
        RECT 466.950 877.800 469.050 879.900 ;
        RECT 473.400 874.050 474.450 886.950 ;
        RECT 479.400 886.050 480.450 889.950 ;
        RECT 478.950 883.950 481.050 886.050 ;
        RECT 482.400 879.900 483.450 892.950 ;
        RECT 487.950 889.950 490.050 895.050 ;
        RECT 487.950 884.100 490.050 886.200 ;
        RECT 496.950 885.000 499.050 889.050 ;
        RECT 488.400 883.350 489.600 884.100 ;
        RECT 497.400 883.350 498.600 885.000 ;
        RECT 487.800 880.950 489.900 883.050 ;
        RECT 493.950 880.950 496.050 883.050 ;
        RECT 496.950 880.950 499.050 883.050 ;
        RECT 502.500 880.950 504.600 883.050 ;
        RECT 494.400 879.900 495.600 880.650 ;
        RECT 481.950 877.800 484.050 879.900 ;
        RECT 493.950 877.800 496.050 879.900 ;
        RECT 503.400 879.000 504.600 880.650 ;
        RECT 502.950 874.950 505.050 879.000 ;
        RECT 508.950 874.950 511.050 877.050 ;
        RECT 460.950 871.950 463.050 874.050 ;
        RECT 472.950 871.950 475.050 874.050 ;
        RECT 451.950 856.950 454.050 859.050 ;
        RECT 448.950 823.950 451.050 826.050 ;
        RECT 439.950 820.950 442.050 823.050 ;
        RECT 445.950 814.950 448.050 817.050 ;
        RECT 439.950 806.100 442.050 808.200 ;
        RECT 440.400 805.350 441.600 806.100 ;
        RECT 434.100 802.950 436.200 805.050 ;
        RECT 439.500 802.950 441.600 805.050 ;
        RECT 442.800 802.950 444.900 805.050 ;
        RECT 434.400 800.400 435.600 802.650 ;
        RECT 443.400 800.400 444.600 802.650 ;
        RECT 446.400 802.050 447.450 814.950 ;
        RECT 434.400 796.050 435.450 800.400 ;
        RECT 433.950 793.950 436.050 796.050 ;
        RECT 433.950 775.950 436.050 778.050 ;
        RECT 424.950 772.950 427.050 775.050 ;
        RECT 415.950 763.950 418.050 766.050 ;
        RECT 421.950 763.950 424.050 766.050 ;
        RECT 400.950 748.950 403.050 751.050 ;
        RECT 406.950 748.950 409.050 751.050 ;
        RECT 412.950 748.950 415.050 751.050 ;
        RECT 394.950 742.950 397.050 745.050 ;
        RECT 391.950 736.950 394.050 739.050 ;
        RECT 385.950 733.950 388.050 736.050 ;
        RECT 379.950 730.950 382.050 733.050 ;
        RECT 388.950 729.000 391.050 733.050 ;
        RECT 395.400 729.600 396.450 742.950 ;
        RECT 389.400 727.350 390.600 729.000 ;
        RECT 395.400 727.350 396.600 729.600 ;
        RECT 401.400 727.050 402.450 748.950 ;
        RECT 388.950 724.950 391.050 727.050 ;
        RECT 391.950 724.950 394.050 727.050 ;
        RECT 394.950 724.950 397.050 727.050 ;
        RECT 400.950 724.950 403.050 727.050 ;
        RECT 392.400 723.900 393.600 724.650 ;
        RECT 391.950 721.800 394.050 723.900 ;
        RECT 400.950 721.800 403.050 723.900 ;
        RECT 376.950 688.950 379.050 691.050 ;
        RECT 365.400 684.450 366.600 684.600 ;
        RECT 362.400 683.400 366.600 684.450 ;
        RECT 370.950 684.000 373.050 688.050 ;
        RECT 365.400 682.350 366.600 683.400 ;
        RECT 371.400 682.350 372.600 684.000 ;
        RECT 376.950 683.100 379.050 685.200 ;
        RECT 377.400 682.350 378.600 683.100 ;
        RECT 385.950 682.950 388.050 685.050 ;
        RECT 391.950 683.100 394.050 685.200 ;
        RECT 364.950 679.950 367.050 682.050 ;
        RECT 367.950 679.950 370.050 682.050 ;
        RECT 370.950 679.950 373.050 682.050 ;
        RECT 373.950 679.950 376.050 682.050 ;
        RECT 376.950 679.950 379.050 682.050 ;
        RECT 358.950 676.800 361.050 678.900 ;
        RECT 361.950 676.950 364.050 679.050 ;
        RECT 368.400 678.900 369.600 679.650 ;
        RECT 349.950 670.950 352.050 673.050 ;
        RECT 355.950 670.950 358.050 673.050 ;
        RECT 346.950 667.950 349.050 670.050 ;
        RECT 343.950 652.950 346.050 655.050 ;
        RECT 347.400 651.600 348.450 667.950 ;
        RECT 362.400 664.050 363.450 676.950 ;
        RECT 367.950 676.800 370.050 678.900 ;
        RECT 374.400 678.000 375.600 679.650 ;
        RECT 373.950 673.950 376.050 678.000 ;
        RECT 386.400 676.050 387.450 682.950 ;
        RECT 392.400 682.350 393.600 683.100 ;
        RECT 391.950 679.950 394.050 682.050 ;
        RECT 394.950 679.950 397.050 682.050 ;
        RECT 395.400 677.400 396.600 679.650 ;
        RECT 385.950 673.950 388.050 676.050 ;
        RECT 386.400 667.050 387.450 673.950 ;
        RECT 385.950 664.950 388.050 667.050 ;
        RECT 395.400 664.050 396.450 677.400 ;
        RECT 361.950 661.950 364.050 664.050 ;
        RECT 370.950 661.950 373.050 664.050 ;
        RECT 382.950 661.950 385.050 664.050 ;
        RECT 394.950 661.950 397.050 664.050 ;
        RECT 359.850 657.300 361.950 659.400 ;
        RECT 347.400 649.350 348.600 651.600 ;
        RECT 343.950 646.950 346.050 649.050 ;
        RECT 346.950 646.950 349.050 649.050 ;
        RECT 349.950 646.950 352.050 649.050 ;
        RECT 355.950 646.950 358.050 649.050 ;
        RECT 344.400 645.900 345.600 646.650 ;
        RECT 343.950 643.800 346.050 645.900 ;
        RECT 350.400 644.400 351.600 646.650 ;
        RECT 356.400 644.400 357.600 646.650 ;
        RECT 350.400 631.050 351.450 644.400 ;
        RECT 356.400 640.050 357.450 644.400 ;
        RECT 355.950 637.950 358.050 640.050 ;
        RECT 360.150 638.700 361.350 657.300 ;
        RECT 365.100 646.950 367.200 649.050 ;
        RECT 365.400 645.900 366.600 646.650 ;
        RECT 371.400 645.900 372.450 661.950 ;
        RECT 377.550 657.300 379.650 659.400 ;
        RECT 364.950 643.800 367.050 645.900 ;
        RECT 370.950 643.800 373.050 645.900 ;
        RECT 377.550 644.400 378.750 657.300 ;
        RECT 383.400 651.600 384.450 661.950 ;
        RECT 395.850 657.300 397.950 659.400 ;
        RECT 383.400 649.350 384.600 651.600 ;
        RECT 382.950 646.950 385.050 649.050 ;
        RECT 391.950 646.950 394.050 649.050 ;
        RECT 392.400 644.400 393.600 646.650 ;
        RECT 377.550 642.300 379.650 644.400 ;
        RECT 360.150 637.500 364.350 638.700 ;
        RECT 373.950 637.950 376.050 640.050 ;
        RECT 362.250 636.600 364.350 637.500 ;
        RECT 349.950 628.950 352.050 631.050 ;
        RECT 358.950 625.950 361.050 628.050 ;
        RECT 355.350 615.300 357.450 617.400 ;
        RECT 343.950 606.000 346.050 610.050 ;
        RECT 356.250 608.700 357.450 615.300 ;
        RECT 355.350 606.600 357.450 608.700 ;
        RECT 344.400 604.350 345.600 606.000 ;
        RECT 340.950 601.950 343.050 604.050 ;
        RECT 343.950 601.950 346.050 604.050 ;
        RECT 349.950 601.950 352.050 604.050 ;
        RECT 341.400 600.900 342.600 601.650 ;
        RECT 350.400 600.900 351.600 601.650 ;
        RECT 340.950 598.800 343.050 600.900 ;
        RECT 349.950 598.800 352.050 600.900 ;
        RECT 341.400 580.050 342.450 598.800 ;
        RECT 356.250 593.700 357.450 606.600 ;
        RECT 355.350 591.600 357.450 593.700 ;
        RECT 337.950 577.950 340.050 580.050 ;
        RECT 340.950 577.950 343.050 580.050 ;
        RECT 346.950 577.950 352.050 580.050 ;
        RECT 338.400 567.900 339.450 577.950 ;
        RECT 340.950 571.950 343.050 574.050 ;
        RECT 346.950 572.100 349.050 574.200 ;
        RECT 337.950 565.800 340.050 567.900 ;
        RECT 334.950 553.950 337.050 556.050 ;
        RECT 335.400 550.050 336.450 553.950 ;
        RECT 337.950 550.950 340.050 553.050 ;
        RECT 334.950 547.950 337.050 550.050 ;
        RECT 289.950 544.950 292.050 547.050 ;
        RECT 281.400 530.400 285.450 531.450 ;
        RECT 239.400 526.350 240.600 528.000 ;
        RECT 241.950 527.100 244.050 529.200 ;
        RECT 229.950 523.950 232.050 526.050 ;
        RECT 232.950 523.950 235.050 526.050 ;
        RECT 235.950 523.950 238.050 526.050 ;
        RECT 238.950 523.950 241.050 526.050 ;
        RECT 230.400 521.400 231.600 523.650 ;
        RECT 236.400 521.400 237.600 523.650 ;
        RECT 245.400 523.050 246.450 529.950 ;
        RECT 253.950 527.100 256.050 529.200 ;
        RECT 260.400 528.450 261.600 528.600 ;
        RECT 260.400 527.400 267.450 528.450 ;
        RECT 254.400 526.350 255.600 527.100 ;
        RECT 260.400 526.350 261.600 527.400 ;
        RECT 253.950 523.950 256.050 526.050 ;
        RECT 256.950 523.950 259.050 526.050 ;
        RECT 259.950 523.950 262.050 526.050 ;
        RECT 230.400 517.050 231.450 521.400 ;
        RECT 229.950 514.950 232.050 517.050 ;
        RECT 236.400 510.450 237.450 521.400 ;
        RECT 244.950 520.950 247.050 523.050 ;
        RECT 257.400 522.900 258.600 523.650 ;
        RECT 256.950 520.800 259.050 522.900 ;
        RECT 266.400 517.050 267.450 527.400 ;
        RECT 277.950 527.100 280.050 529.200 ;
        RECT 284.400 528.600 285.450 530.400 ;
        RECT 278.400 526.350 279.600 527.100 ;
        RECT 284.400 526.350 285.600 528.600 ;
        RECT 274.950 523.950 277.050 526.050 ;
        RECT 277.950 523.950 280.050 526.050 ;
        RECT 280.950 523.950 283.050 526.050 ;
        RECT 283.950 523.950 286.050 526.050 ;
        RECT 275.400 522.900 276.600 523.650 ;
        RECT 274.950 520.800 277.050 522.900 ;
        RECT 281.400 521.400 282.600 523.650 ;
        RECT 290.400 522.900 291.450 544.950 ;
        RECT 298.950 527.100 301.050 529.200 ;
        RECT 325.950 527.100 328.050 529.200 ;
        RECT 338.400 528.600 339.450 550.950 ;
        RECT 299.400 526.350 300.600 527.100 ;
        RECT 298.950 523.950 301.050 526.050 ;
        RECT 301.950 523.950 304.050 526.050 ;
        RECT 319.800 523.950 321.900 526.050 ;
        RECT 259.950 514.950 262.050 517.050 ;
        RECT 265.950 514.950 268.050 517.050 ;
        RECT 233.400 509.400 237.450 510.450 ;
        RECT 229.950 502.950 232.050 505.050 ;
        RECT 230.400 495.600 231.450 502.950 ;
        RECT 233.400 499.050 234.450 509.400 ;
        RECT 235.950 505.950 238.050 508.050 ;
        RECT 232.950 496.950 235.050 499.050 ;
        RECT 236.400 495.600 237.450 505.950 ;
        RECT 248.850 501.300 250.950 503.400 ;
        RECT 230.400 493.350 231.600 495.600 ;
        RECT 236.400 493.350 237.600 495.600 ;
        RECT 229.950 490.950 232.050 493.050 ;
        RECT 232.950 490.950 235.050 493.050 ;
        RECT 235.950 490.950 238.050 493.050 ;
        RECT 238.950 490.950 241.050 493.050 ;
        RECT 244.950 490.950 247.050 493.050 ;
        RECT 233.400 489.900 234.600 490.650 ;
        RECT 239.400 489.900 240.600 490.650 ;
        RECT 232.950 487.800 235.050 489.900 ;
        RECT 238.950 487.800 241.050 489.900 ;
        RECT 245.400 488.400 246.600 490.650 ;
        RECT 245.400 478.050 246.450 488.400 ;
        RECT 249.150 482.700 250.350 501.300 ;
        RECT 254.100 490.950 256.200 493.050 ;
        RECT 254.400 489.450 255.600 490.650 ;
        RECT 260.400 489.450 261.450 514.950 ;
        RECT 271.950 505.950 274.050 508.050 ;
        RECT 266.550 501.300 268.650 503.400 ;
        RECT 272.400 502.050 273.450 505.950 ;
        RECT 254.400 488.400 261.450 489.450 ;
        RECT 262.950 487.800 265.050 489.900 ;
        RECT 266.550 488.400 267.750 501.300 ;
        RECT 271.950 499.950 274.050 502.050 ;
        RECT 272.400 495.600 273.450 499.950 ;
        RECT 281.400 499.050 282.450 521.400 ;
        RECT 289.950 520.800 292.050 522.900 ;
        RECT 302.400 521.400 303.600 523.650 ;
        RECT 302.400 511.050 303.450 521.400 ;
        RECT 326.400 517.050 327.450 527.100 ;
        RECT 338.400 526.350 339.600 528.600 ;
        RECT 337.800 523.950 339.900 526.050 ;
        RECT 325.950 514.950 328.050 517.050 ;
        RECT 301.950 508.950 304.050 511.050 ;
        RECT 307.950 508.950 310.050 511.050 ;
        RECT 319.950 508.950 322.050 511.050 ;
        RECT 284.850 501.300 286.950 503.400 ;
        RECT 302.550 501.300 304.650 503.400 ;
        RECT 280.950 496.950 283.050 499.050 ;
        RECT 272.400 493.350 273.600 495.600 ;
        RECT 271.950 490.950 274.050 493.050 ;
        RECT 280.950 490.950 283.050 493.050 ;
        RECT 281.400 488.400 282.600 490.650 ;
        RECT 249.150 481.500 253.350 482.700 ;
        RECT 251.250 480.600 253.350 481.500 ;
        RECT 244.950 475.950 247.050 478.050 ;
        RECT 223.950 469.950 226.050 472.050 ;
        RECT 256.950 469.950 259.050 472.050 ;
        RECT 217.950 466.950 220.050 469.050 ;
        RECT 191.400 448.350 192.600 449.100 ;
        RECT 191.100 445.950 193.200 448.050 ;
        RECT 193.950 439.950 196.050 442.050 ;
        RECT 185.850 435.600 187.950 437.700 ;
        RECT 194.400 436.050 195.450 439.950 ;
        RECT 193.950 433.950 196.050 436.050 ;
        RECT 175.800 424.950 177.900 427.050 ;
        RECT 178.950 424.950 181.050 427.050 ;
        RECT 176.400 417.600 177.450 424.950 ;
        RECT 176.400 415.350 177.600 417.600 ;
        RECT 176.400 412.950 178.500 415.050 ;
        RECT 181.800 412.950 183.900 415.050 ;
        RECT 182.400 411.900 183.600 412.650 ;
        RECT 194.400 411.900 195.450 433.950 ;
        RECT 197.400 433.050 198.450 449.100 ;
        RECT 203.550 437.700 204.750 450.600 ;
        RECT 211.950 448.950 214.050 451.050 ;
        RECT 218.400 450.600 219.450 466.950 ;
        RECT 253.950 463.950 256.050 466.050 ;
        RECT 239.550 459.300 241.650 461.400 ;
        RECT 224.250 457.500 226.350 458.400 ;
        RECT 222.150 456.300 226.350 457.500 ;
        RECT 218.400 448.350 219.600 450.600 ;
        RECT 208.950 445.950 211.050 448.050 ;
        RECT 217.950 445.950 220.050 448.050 ;
        RECT 205.950 441.450 208.050 445.050 ;
        RECT 209.400 444.450 210.600 445.650 ;
        RECT 209.400 443.400 213.450 444.450 ;
        RECT 205.950 441.000 210.450 441.450 ;
        RECT 206.400 440.400 210.450 441.000 ;
        RECT 203.550 435.600 205.650 437.700 ;
        RECT 209.400 433.050 210.450 440.400 ;
        RECT 196.950 430.950 199.050 433.050 ;
        RECT 202.950 430.950 205.050 433.050 ;
        RECT 208.950 430.950 211.050 433.050 ;
        RECT 203.400 417.600 204.450 430.950 ;
        RECT 203.400 415.350 204.600 417.600 ;
        RECT 199.950 412.950 202.050 415.050 ;
        RECT 202.950 412.950 205.050 415.050 ;
        RECT 205.950 412.950 208.050 415.050 ;
        RECT 206.400 411.900 207.600 412.650 ;
        RECT 181.950 409.800 184.050 411.900 ;
        RECT 193.950 409.800 196.050 411.900 ;
        RECT 205.950 409.800 208.050 411.900 ;
        RECT 166.950 406.950 169.050 409.050 ;
        RECT 206.400 400.050 207.450 409.800 ;
        RECT 205.950 397.950 208.050 400.050 ;
        RECT 212.400 397.050 213.450 443.400 ;
        RECT 222.150 437.700 223.350 456.300 ;
        RECT 226.950 450.000 229.050 454.050 ;
        RECT 235.950 451.950 238.050 454.050 ;
        RECT 239.550 452.700 240.750 459.300 ;
        RECT 250.950 457.950 253.050 460.050 ;
        RECT 227.400 448.350 228.600 450.000 ;
        RECT 227.100 445.950 229.200 448.050 ;
        RECT 232.950 445.950 235.050 448.050 ;
        RECT 221.850 435.600 223.950 437.700 ;
        RECT 233.400 432.450 234.450 445.950 ;
        RECT 236.400 436.050 237.450 451.950 ;
        RECT 239.550 450.600 241.650 452.700 ;
        RECT 239.550 437.700 240.750 450.600 ;
        RECT 244.950 445.950 247.050 448.050 ;
        RECT 245.400 444.000 246.600 445.650 ;
        RECT 244.950 439.950 247.050 444.000 ;
        RECT 235.950 433.950 238.050 436.050 ;
        RECT 239.550 435.600 241.650 437.700 ;
        RECT 251.400 433.050 252.450 457.950 ;
        RECT 254.400 433.050 255.450 463.950 ;
        RECT 257.400 444.900 258.450 469.950 ;
        RECT 263.400 469.050 264.450 487.800 ;
        RECT 266.550 486.300 268.650 488.400 ;
        RECT 266.550 479.700 267.750 486.300 ;
        RECT 266.550 477.600 268.650 479.700 ;
        RECT 281.400 478.050 282.450 488.400 ;
        RECT 285.150 482.700 286.350 501.300 ;
        RECT 290.100 490.950 292.200 493.050 ;
        RECT 290.400 489.900 291.600 490.650 ;
        RECT 289.950 487.800 292.050 489.900 ;
        RECT 302.550 488.400 303.750 501.300 ;
        RECT 308.400 495.600 309.450 508.950 ;
        RECT 308.400 493.350 309.600 495.600 ;
        RECT 316.950 493.950 319.050 496.050 ;
        RECT 307.950 490.950 310.050 493.050 ;
        RECT 302.550 486.300 304.650 488.400 ;
        RECT 285.150 481.500 289.350 482.700 ;
        RECT 287.250 480.600 289.350 481.500 ;
        RECT 298.950 478.950 301.050 481.050 ;
        RECT 302.550 479.700 303.750 486.300 ;
        RECT 280.950 475.950 283.050 478.050 ;
        RECT 262.950 466.950 265.050 469.050 ;
        RECT 265.950 449.100 268.050 451.200 ;
        RECT 271.950 449.100 274.050 451.200 ;
        RECT 266.400 448.350 267.600 449.100 ;
        RECT 272.400 448.350 273.600 449.100 ;
        RECT 277.950 448.950 280.050 451.050 ;
        RECT 262.950 445.950 265.050 448.050 ;
        RECT 265.950 445.950 268.050 448.050 ;
        RECT 268.950 445.950 271.050 448.050 ;
        RECT 271.950 445.950 274.050 448.050 ;
        RECT 263.400 444.900 264.600 445.650 ;
        RECT 256.950 442.800 259.050 444.900 ;
        RECT 262.950 442.800 265.050 444.900 ;
        RECT 269.400 443.400 270.600 445.650 ;
        RECT 269.400 436.050 270.450 443.400 ;
        RECT 278.400 442.050 279.450 448.950 ;
        RECT 277.950 439.950 280.050 442.050 ;
        RECT 281.400 439.050 282.450 475.950 ;
        RECT 292.950 469.950 295.050 472.050 ;
        RECT 286.950 449.100 289.050 451.200 ;
        RECT 293.400 450.600 294.450 469.950 ;
        RECT 287.400 448.350 288.600 449.100 ;
        RECT 293.400 448.350 294.600 450.600 ;
        RECT 286.950 445.950 289.050 448.050 ;
        RECT 289.950 445.950 292.050 448.050 ;
        RECT 292.950 445.950 295.050 448.050 ;
        RECT 290.400 444.900 291.600 445.650 ;
        RECT 299.400 444.900 300.450 478.950 ;
        RECT 302.550 477.600 304.650 479.700 ;
        RECT 317.400 453.450 318.450 493.950 ;
        RECT 320.400 489.900 321.450 508.950 ;
        RECT 326.400 495.600 327.450 514.950 ;
        RECT 337.950 511.950 340.050 514.050 ;
        RECT 326.400 493.350 327.600 495.600 ;
        RECT 331.950 494.100 334.050 496.200 ;
        RECT 338.400 496.050 339.450 511.950 ;
        RECT 341.400 502.050 342.450 571.950 ;
        RECT 347.400 571.350 348.600 572.100 ;
        RECT 346.950 568.950 349.050 571.050 ;
        RECT 349.950 568.950 352.050 571.050 ;
        RECT 350.400 567.900 351.600 568.650 ;
        RECT 349.950 565.800 352.050 567.900 ;
        RECT 359.400 544.050 360.450 625.950 ;
        RECT 374.400 618.450 375.450 637.950 ;
        RECT 377.550 635.700 378.750 642.300 ;
        RECT 392.400 640.050 393.450 644.400 ;
        RECT 391.950 637.950 394.050 640.050 ;
        RECT 396.150 638.700 397.350 657.300 ;
        RECT 401.400 655.050 402.450 721.800 ;
        RECT 407.400 697.050 408.450 748.950 ;
        RECT 416.400 739.050 417.450 763.950 ;
        RECT 422.400 762.450 423.600 762.600 ;
        RECT 419.400 761.400 423.600 762.450 ;
        RECT 419.400 745.050 420.450 761.400 ;
        RECT 422.400 760.350 423.600 761.400 ;
        RECT 430.950 761.100 433.050 763.200 ;
        RECT 431.400 760.350 432.600 761.100 ;
        RECT 422.100 757.950 424.200 760.050 ;
        RECT 425.400 757.950 427.500 760.050 ;
        RECT 430.800 757.950 432.900 760.050 ;
        RECT 425.400 756.900 426.600 757.650 ;
        RECT 424.950 754.800 427.050 756.900 ;
        RECT 434.400 751.050 435.450 775.950 ;
        RECT 436.950 761.100 439.050 763.200 ;
        RECT 433.950 748.950 436.050 751.050 ;
        RECT 437.400 748.050 438.450 761.100 ;
        RECT 443.400 756.900 444.450 800.400 ;
        RECT 445.950 799.950 448.050 802.050 ;
        RECT 452.400 772.050 453.450 856.950 ;
        RECT 461.400 840.600 462.450 871.950 ;
        RECT 469.950 865.950 472.050 868.050 ;
        RECT 470.400 841.200 471.450 865.950 ;
        RECT 505.950 856.950 508.050 859.050 ;
        RECT 472.950 850.950 475.050 853.050 ;
        RECT 461.400 838.350 462.600 840.600 ;
        RECT 469.950 839.100 472.050 841.200 ;
        RECT 457.950 835.950 460.050 838.050 ;
        RECT 460.950 835.950 463.050 838.050 ;
        RECT 463.950 835.950 466.050 838.050 ;
        RECT 458.400 834.900 459.600 835.650 ;
        RECT 464.400 834.900 465.600 835.650 ;
        RECT 457.950 832.800 460.050 834.900 ;
        RECT 463.950 832.800 466.050 834.900 ;
        RECT 473.400 834.450 474.450 850.950 ;
        RECT 484.950 847.950 487.050 850.050 ;
        RECT 499.950 847.950 502.050 850.050 ;
        RECT 478.950 839.100 481.050 844.050 ;
        RECT 485.400 840.600 486.450 847.950 ;
        RECT 496.950 841.950 499.050 844.050 ;
        RECT 479.400 838.350 480.600 839.100 ;
        RECT 485.400 838.350 486.600 840.600 ;
        RECT 490.950 838.950 493.050 841.050 ;
        RECT 478.950 835.950 481.050 838.050 ;
        RECT 481.950 835.950 484.050 838.050 ;
        RECT 484.950 835.950 487.050 838.050 ;
        RECT 473.400 833.400 477.450 834.450 ;
        RECT 460.950 823.950 463.050 826.050 ;
        RECT 461.400 807.600 462.450 823.950 ;
        RECT 461.400 805.350 462.600 807.600 ;
        RECT 457.950 802.950 460.050 805.050 ;
        RECT 460.950 802.950 463.050 805.050 ;
        RECT 463.950 802.950 466.050 805.050 ;
        RECT 464.400 800.400 465.600 802.650 ;
        RECT 464.400 781.050 465.450 800.400 ;
        RECT 476.400 793.050 477.450 833.400 ;
        RECT 482.400 833.400 483.600 835.650 ;
        RECT 491.400 834.900 492.450 838.950 ;
        RECT 497.400 834.900 498.450 841.950 ;
        RECT 500.400 840.600 501.450 847.950 ;
        RECT 506.400 844.050 507.450 856.950 ;
        RECT 509.400 856.050 510.450 874.950 ;
        RECT 515.400 868.050 516.450 970.950 ;
        RECT 520.950 962.100 523.050 964.200 ;
        RECT 527.400 963.600 528.450 970.950 ;
        RECT 554.400 964.200 555.450 973.950 ;
        RECT 562.950 964.950 565.050 967.050 ;
        RECT 586.950 964.950 589.050 967.050 ;
        RECT 521.400 961.350 522.600 962.100 ;
        RECT 527.400 961.350 528.600 963.600 ;
        RECT 535.950 961.950 538.050 964.050 ;
        RECT 541.950 962.100 544.050 964.200 ;
        RECT 544.950 963.600 549.000 964.050 ;
        RECT 520.950 958.950 523.050 961.050 ;
        RECT 523.950 958.950 526.050 961.050 ;
        RECT 526.950 958.950 529.050 961.050 ;
        RECT 529.950 958.950 532.050 961.050 ;
        RECT 524.400 957.900 525.600 958.650 ;
        RECT 523.950 955.800 526.050 957.900 ;
        RECT 530.400 956.400 531.600 958.650 ;
        RECT 536.400 957.900 537.450 961.950 ;
        RECT 530.400 952.050 531.450 956.400 ;
        RECT 535.950 955.800 538.050 957.900 ;
        RECT 529.950 949.950 532.050 952.050 ;
        RECT 542.400 940.050 543.450 962.100 ;
        RECT 544.950 961.950 549.600 963.600 ;
        RECT 553.950 962.100 556.050 964.200 ;
        RECT 548.400 961.350 549.600 961.950 ;
        RECT 554.400 961.350 555.600 962.100 ;
        RECT 547.950 958.950 550.050 961.050 ;
        RECT 550.950 958.950 553.050 961.050 ;
        RECT 553.950 958.950 556.050 961.050 ;
        RECT 556.950 958.950 559.050 961.050 ;
        RECT 551.400 957.900 552.600 958.650 ;
        RECT 557.400 957.900 558.600 958.650 ;
        RECT 563.400 957.900 564.450 964.950 ;
        RECT 565.950 962.100 568.050 964.200 ;
        RECT 574.950 962.100 577.050 964.200 ;
        RECT 550.950 955.800 553.050 957.900 ;
        RECT 556.950 955.800 559.050 957.900 ;
        RECT 562.950 955.800 565.050 957.900 ;
        RECT 566.400 957.450 567.450 962.100 ;
        RECT 575.400 961.350 576.600 962.100 ;
        RECT 571.950 958.950 574.050 961.050 ;
        RECT 574.950 958.950 577.050 961.050 ;
        RECT 572.400 957.900 573.600 958.650 ;
        RECT 587.400 957.900 588.450 964.950 ;
        RECT 596.400 963.600 597.450 973.950 ;
        RECT 622.950 970.950 625.050 973.050 ;
        RECT 733.950 972.450 736.050 973.050 ;
        RECT 739.950 972.450 742.050 973.050 ;
        RECT 733.950 971.400 742.050 972.450 ;
        RECT 733.950 970.950 736.050 971.400 ;
        RECT 739.950 970.950 742.050 971.400 ;
        RECT 781.950 970.950 784.050 973.050 ;
        RECT 596.400 961.350 597.600 963.600 ;
        RECT 601.950 962.100 604.050 964.200 ;
        RECT 602.400 961.350 603.600 962.100 ;
        RECT 607.950 961.950 610.050 964.050 ;
        RECT 616.950 962.100 619.050 964.200 ;
        RECT 623.400 963.600 624.450 970.950 ;
        RECT 664.950 967.950 667.050 970.050 ;
        RECT 736.950 969.450 739.050 970.050 ;
        RECT 731.400 969.000 739.050 969.450 ;
        RECT 730.950 968.400 739.050 969.000 ;
        RECT 592.950 958.950 595.050 961.050 ;
        RECT 595.950 958.950 598.050 961.050 ;
        RECT 598.950 958.950 601.050 961.050 ;
        RECT 601.950 958.950 604.050 961.050 ;
        RECT 566.400 957.000 570.450 957.450 ;
        RECT 565.950 956.400 570.450 957.000 ;
        RECT 565.950 952.950 568.050 956.400 ;
        RECT 559.950 940.950 562.050 943.050 ;
        RECT 541.950 937.950 544.050 940.050 ;
        RECT 535.950 931.950 538.050 934.050 ;
        RECT 532.950 928.950 535.050 931.050 ;
        RECT 523.950 922.950 526.050 925.050 ;
        RECT 524.400 918.600 525.450 922.950 ;
        RECT 524.400 916.350 525.600 918.600 ;
        RECT 523.950 913.950 526.050 916.050 ;
        RECT 526.950 913.950 529.050 916.050 ;
        RECT 527.400 912.900 528.600 913.650 ;
        RECT 533.400 913.050 534.450 928.950 ;
        RECT 526.950 910.800 529.050 912.900 ;
        RECT 532.950 910.950 535.050 913.050 ;
        RECT 536.400 912.450 537.450 931.950 ;
        RECT 544.950 922.950 547.050 925.050 ;
        RECT 550.950 922.950 553.050 925.050 ;
        RECT 545.400 918.600 546.450 922.950 ;
        RECT 551.400 918.600 552.450 922.950 ;
        RECT 545.400 916.350 546.600 918.600 ;
        RECT 551.400 916.350 552.600 918.600 ;
        RECT 541.950 913.950 544.050 916.050 ;
        RECT 544.950 913.950 547.050 916.050 ;
        RECT 547.950 913.950 550.050 916.050 ;
        RECT 550.950 913.950 553.050 916.050 ;
        RECT 542.400 912.450 543.600 913.650 ;
        RECT 536.400 911.400 543.600 912.450 ;
        RECT 548.400 911.400 549.600 913.650 ;
        RECT 527.400 909.450 528.450 910.800 ;
        RECT 524.400 908.400 528.450 909.450 ;
        RECT 524.400 885.600 525.450 908.400 ;
        RECT 538.950 901.950 541.050 904.050 ;
        RECT 539.400 898.050 540.450 901.950 ;
        RECT 548.400 901.050 549.450 911.400 ;
        RECT 553.950 910.950 556.050 913.050 ;
        RECT 554.400 907.050 555.450 910.950 ;
        RECT 553.950 904.950 556.050 907.050 ;
        RECT 547.950 898.950 550.050 901.050 ;
        RECT 538.950 895.950 541.050 898.050 ;
        RECT 532.950 892.950 535.050 895.050 ;
        RECT 524.400 883.350 525.600 885.600 ;
        RECT 520.950 880.950 523.050 883.050 ;
        RECT 523.950 880.950 526.050 883.050 ;
        RECT 526.950 880.950 529.050 883.050 ;
        RECT 521.400 879.000 522.600 880.650 ;
        RECT 527.400 879.450 528.600 880.650 ;
        RECT 520.950 874.950 523.050 879.000 ;
        RECT 527.400 878.400 531.450 879.450 ;
        RECT 514.950 865.950 517.050 868.050 ;
        RECT 514.950 856.950 517.050 859.050 ;
        RECT 508.950 853.950 511.050 856.050 ;
        RECT 505.950 841.950 508.050 844.050 ;
        RECT 509.400 840.600 510.450 853.950 ;
        RECT 500.400 838.350 501.600 840.600 ;
        RECT 509.400 838.350 510.600 840.600 ;
        RECT 500.100 835.950 502.200 838.050 ;
        RECT 505.500 835.950 507.600 838.050 ;
        RECT 508.800 835.950 510.900 838.050 ;
        RECT 506.400 834.900 507.600 835.650 ;
        RECT 515.400 835.050 516.450 856.950 ;
        RECT 523.950 844.950 526.050 847.050 ;
        RECT 524.400 841.200 525.450 844.950 ;
        RECT 530.400 841.200 531.450 878.400 ;
        RECT 533.400 874.050 534.450 892.950 ;
        RECT 539.400 877.050 540.450 895.950 ;
        RECT 547.950 892.950 550.050 895.050 ;
        RECT 548.400 885.600 549.450 892.950 ;
        RECT 554.400 885.600 555.450 904.950 ;
        RECT 548.400 883.350 549.600 885.600 ;
        RECT 554.400 883.350 555.600 885.600 ;
        RECT 544.950 880.950 547.050 883.050 ;
        RECT 547.950 880.950 550.050 883.050 ;
        RECT 550.950 880.950 553.050 883.050 ;
        RECT 553.950 880.950 556.050 883.050 ;
        RECT 545.400 879.000 546.600 880.650 ;
        RECT 551.400 879.900 552.600 880.650 ;
        RECT 538.950 874.950 541.050 877.050 ;
        RECT 544.950 874.950 547.050 879.000 ;
        RECT 550.950 877.800 553.050 879.900 ;
        RECT 532.950 871.950 535.050 874.050 ;
        RECT 541.950 865.950 544.050 868.050 ;
        RECT 535.950 847.950 538.050 850.050 ;
        RECT 517.950 839.100 520.050 841.200 ;
        RECT 523.950 839.100 526.050 841.200 ;
        RECT 529.950 839.100 532.050 841.200 ;
        RECT 482.400 826.050 483.450 833.400 ;
        RECT 490.950 832.800 493.050 834.900 ;
        RECT 496.950 832.800 499.050 834.900 ;
        RECT 505.950 832.800 508.050 834.900 ;
        RECT 514.950 832.950 517.050 835.050 ;
        RECT 505.950 826.950 508.050 829.050 ;
        RECT 481.950 823.950 484.050 826.050 ;
        RECT 481.950 802.950 484.050 805.050 ;
        RECT 484.950 802.950 487.050 805.050 ;
        RECT 487.950 802.950 490.050 805.050 ;
        RECT 490.950 802.950 493.050 805.050 ;
        RECT 493.950 802.950 496.050 805.050 ;
        RECT 482.400 800.400 483.600 802.650 ;
        RECT 488.400 801.900 489.600 802.650 ;
        RECT 494.400 801.900 495.600 802.650 ;
        RECT 475.950 790.950 478.050 793.050 ;
        RECT 463.950 778.950 466.050 781.050 ;
        RECT 451.950 769.950 454.050 772.050 ;
        RECT 463.950 769.950 466.050 772.050 ;
        RECT 449.100 766.500 451.200 768.600 ;
        RECT 446.100 757.950 448.200 760.050 ;
        RECT 449.100 759.900 450.000 766.500 ;
        RECT 458.100 766.200 460.200 768.300 ;
        RECT 452.400 763.350 453.600 765.600 ;
        RECT 451.800 760.950 453.900 763.050 ;
        RECT 456.000 759.900 458.100 760.200 ;
        RECT 449.100 759.000 458.100 759.900 ;
        RECT 442.950 756.450 445.050 756.900 ;
        RECT 446.400 756.450 447.600 757.650 ;
        RECT 442.950 755.400 447.600 756.450 ;
        RECT 442.950 754.800 445.050 755.400 ;
        RECT 449.100 753.900 450.000 759.000 ;
        RECT 456.000 758.100 458.100 759.000 ;
        RECT 450.900 757.200 453.000 758.100 ;
        RECT 450.900 756.000 458.100 757.200 ;
        RECT 456.000 755.100 458.100 756.000 ;
        RECT 448.500 751.800 450.600 753.900 ;
        RECT 451.800 752.100 453.900 754.200 ;
        RECT 459.000 753.600 459.900 766.200 ;
        RECT 460.950 761.100 463.050 763.200 ;
        RECT 461.400 760.350 462.600 761.100 ;
        RECT 460.800 757.950 462.900 760.050 ;
        RECT 452.400 749.550 453.600 751.800 ;
        RECT 458.400 751.500 460.500 753.600 ;
        RECT 436.950 745.950 439.050 748.050 ;
        RECT 418.950 742.950 421.050 745.050 ;
        RECT 415.950 736.950 418.050 739.050 ;
        RECT 424.950 736.950 427.050 739.050 ;
        RECT 415.950 728.100 418.050 730.200 ;
        RECT 416.400 727.350 417.600 728.100 ;
        RECT 412.950 724.950 415.050 727.050 ;
        RECT 415.950 724.950 418.050 727.050 ;
        RECT 413.400 723.000 414.600 724.650 ;
        RECT 425.400 723.900 426.450 736.950 ;
        RECT 430.950 733.950 433.050 736.050 ;
        RECT 452.400 735.450 453.450 749.550 ;
        RECT 460.950 745.950 463.050 748.050 ;
        RECT 449.400 734.400 453.450 735.450 ;
        RECT 431.400 729.600 432.450 733.950 ;
        RECT 431.400 727.350 432.600 729.600 ;
        RECT 436.950 728.100 439.050 730.200 ;
        RECT 445.950 728.100 448.050 730.200 ;
        RECT 437.400 727.350 438.600 728.100 ;
        RECT 430.950 724.950 433.050 727.050 ;
        RECT 433.950 724.950 436.050 727.050 ;
        RECT 436.950 724.950 439.050 727.050 ;
        RECT 439.950 724.950 442.050 727.050 ;
        RECT 434.400 723.900 435.600 724.650 ;
        RECT 440.400 723.900 441.600 724.650 ;
        RECT 412.950 718.950 415.050 723.000 ;
        RECT 424.950 721.800 427.050 723.900 ;
        RECT 433.950 721.800 436.050 723.900 ;
        RECT 439.950 721.800 442.050 723.900 ;
        RECT 446.400 709.050 447.450 728.100 ;
        RECT 445.950 706.950 448.050 709.050 ;
        RECT 449.400 700.050 450.450 734.400 ;
        RECT 451.950 730.950 454.050 733.050 ;
        RECT 412.950 697.950 415.050 700.050 ;
        RECT 448.950 697.950 451.050 700.050 ;
        RECT 406.950 694.950 409.050 697.050 ;
        RECT 413.400 684.600 414.450 697.950 ;
        RECT 413.400 682.350 414.600 684.600 ;
        RECT 418.950 683.100 421.050 685.200 ;
        RECT 430.950 683.100 433.050 685.200 ;
        RECT 437.400 684.450 438.600 684.600 ;
        RECT 434.400 683.400 438.600 684.450 ;
        RECT 419.400 682.350 420.600 683.100 ;
        RECT 409.950 679.950 412.050 682.050 ;
        RECT 412.950 679.950 415.050 682.050 ;
        RECT 415.950 679.950 418.050 682.050 ;
        RECT 418.950 679.950 421.050 682.050 ;
        RECT 410.400 677.400 411.600 679.650 ;
        RECT 416.400 677.400 417.600 679.650 ;
        RECT 410.400 673.050 411.450 677.400 ;
        RECT 409.950 670.950 412.050 673.050 ;
        RECT 403.950 667.950 406.050 670.050 ;
        RECT 400.950 652.950 403.050 655.050 ;
        RECT 404.400 652.050 405.450 667.950 ;
        RECT 406.950 661.950 409.050 664.050 ;
        RECT 403.950 649.950 406.050 652.050 ;
        RECT 401.100 646.950 403.200 649.050 ;
        RECT 401.400 645.900 402.600 646.650 ;
        RECT 400.950 643.800 403.050 645.900 ;
        RECT 377.550 633.600 379.650 635.700 ;
        RECT 374.400 617.400 378.450 618.450 ;
        RECT 370.650 613.500 372.750 614.400 ;
        RECT 370.650 612.300 374.850 613.500 ;
        RECT 367.950 605.100 370.050 607.200 ;
        RECT 368.400 604.350 369.600 605.100 ;
        RECT 367.800 601.950 369.900 604.050 ;
        RECT 373.650 593.700 374.850 612.300 ;
        RECT 377.400 606.600 378.450 617.400 ;
        RECT 377.400 604.350 378.600 606.600 ;
        RECT 382.950 605.100 385.050 607.200 ;
        RECT 376.950 601.950 379.050 604.050 ;
        RECT 383.400 601.050 384.450 605.100 ;
        RECT 382.950 598.950 385.050 601.050 ;
        RECT 373.050 591.600 375.150 593.700 ;
        RECT 376.950 586.950 379.050 589.050 ;
        RECT 364.950 580.950 367.050 583.050 ;
        RECT 365.400 573.600 366.450 580.950 ;
        RECT 370.950 577.950 373.050 580.050 ;
        RECT 371.400 573.600 372.450 577.950 ;
        RECT 377.400 574.050 378.450 586.950 ;
        RECT 383.850 579.300 385.950 581.400 ;
        RECT 365.400 571.350 366.600 573.600 ;
        RECT 371.400 571.350 372.600 573.600 ;
        RECT 376.950 571.950 379.050 574.050 ;
        RECT 364.950 568.950 367.050 571.050 ;
        RECT 367.950 568.950 370.050 571.050 ;
        RECT 370.950 568.950 373.050 571.050 ;
        RECT 373.950 568.950 376.050 571.050 ;
        RECT 379.950 568.950 382.050 571.050 ;
        RECT 368.400 567.900 369.600 568.650 ;
        RECT 374.400 567.900 375.600 568.650 ;
        RECT 380.400 567.900 381.600 568.650 ;
        RECT 367.950 565.800 370.050 567.900 ;
        RECT 373.950 565.800 376.050 567.900 ;
        RECT 379.950 565.800 382.050 567.900 ;
        RECT 384.150 560.700 385.350 579.300 ;
        RECT 392.400 574.050 393.450 637.950 ;
        RECT 396.150 637.500 400.350 638.700 ;
        RECT 398.250 636.600 400.350 637.500 ;
        RECT 400.950 606.000 403.050 610.050 ;
        RECT 407.400 606.600 408.450 661.950 ;
        RECT 410.400 631.050 411.450 670.950 ;
        RECT 416.400 670.050 417.450 677.400 ;
        RECT 415.950 667.950 418.050 670.050 ;
        RECT 424.950 664.950 427.050 667.050 ;
        RECT 413.550 657.300 415.650 659.400 ;
        RECT 413.550 644.400 414.750 657.300 ;
        RECT 418.950 650.100 421.050 652.200 ;
        RECT 419.400 649.350 420.600 650.100 ;
        RECT 418.950 646.950 421.050 649.050 ;
        RECT 413.550 642.300 415.650 644.400 ;
        RECT 413.550 635.700 414.750 642.300 ;
        RECT 413.550 633.600 415.650 635.700 ;
        RECT 409.950 628.950 412.050 631.050 ;
        RECT 415.950 613.950 418.050 616.050 ;
        RECT 401.400 604.350 402.600 606.000 ;
        RECT 407.400 604.350 408.600 606.600 ;
        RECT 412.950 604.950 415.050 607.050 ;
        RECT 397.950 601.950 400.050 604.050 ;
        RECT 400.950 601.950 403.050 604.050 ;
        RECT 403.950 601.950 406.050 604.050 ;
        RECT 406.950 601.950 409.050 604.050 ;
        RECT 398.400 599.400 399.600 601.650 ;
        RECT 404.400 600.900 405.600 601.650 ;
        RECT 394.950 583.950 397.050 586.050 ;
        RECT 391.950 571.950 394.050 574.050 ;
        RECT 389.100 568.950 391.200 571.050 ;
        RECT 389.400 567.900 390.600 568.650 ;
        RECT 395.400 567.900 396.450 583.950 ;
        RECT 388.950 565.800 391.050 567.900 ;
        RECT 394.950 565.800 397.050 567.900 ;
        RECT 398.400 565.050 399.450 599.400 ;
        RECT 403.950 598.800 406.050 600.900 ;
        RECT 401.550 579.300 403.650 581.400 ;
        RECT 401.550 566.400 402.750 579.300 ;
        RECT 413.400 574.200 414.450 604.950 ;
        RECT 416.400 583.050 417.450 613.950 ;
        RECT 425.400 606.600 426.450 664.950 ;
        RECT 427.950 655.950 430.050 658.050 ;
        RECT 428.400 637.050 429.450 655.950 ;
        RECT 431.400 655.050 432.450 683.100 ;
        RECT 430.950 652.950 433.050 655.050 ;
        RECT 434.400 652.050 435.450 683.400 ;
        RECT 437.400 682.350 438.600 683.400 ;
        RECT 446.400 684.450 447.600 684.600 ;
        RECT 446.400 683.400 450.450 684.450 ;
        RECT 446.400 682.350 447.600 683.400 ;
        RECT 437.100 679.950 439.200 682.050 ;
        RECT 440.400 679.950 442.500 682.050 ;
        RECT 445.800 679.950 447.900 682.050 ;
        RECT 440.400 678.900 441.600 679.650 ;
        RECT 439.950 676.800 442.050 678.900 ;
        RECT 449.400 673.050 450.450 683.400 ;
        RECT 448.950 670.950 451.050 673.050 ;
        RECT 439.950 661.950 442.050 664.050 ;
        RECT 433.950 649.950 436.050 652.050 ;
        RECT 440.400 651.600 441.450 661.950 ;
        RECT 445.950 658.950 448.050 661.050 ;
        RECT 446.400 651.600 447.450 658.950 ;
        RECT 440.400 649.350 441.600 651.600 ;
        RECT 446.400 649.350 447.600 651.600 ;
        RECT 430.950 646.950 433.050 649.050 ;
        RECT 436.950 646.950 439.050 649.050 ;
        RECT 439.950 646.950 442.050 649.050 ;
        RECT 442.950 646.950 445.050 649.050 ;
        RECT 445.950 646.950 448.050 649.050 ;
        RECT 431.400 640.050 432.450 646.950 ;
        RECT 437.400 644.400 438.600 646.650 ;
        RECT 443.400 645.900 444.600 646.650 ;
        RECT 430.950 637.950 433.050 640.050 ;
        RECT 427.950 634.950 430.050 637.050 ;
        RECT 437.400 622.050 438.450 644.400 ;
        RECT 442.950 643.800 445.050 645.900 ;
        RECT 452.400 634.050 453.450 730.950 ;
        RECT 461.400 729.600 462.450 745.950 ;
        RECT 464.400 733.050 465.450 769.950 ;
        RECT 472.950 763.950 475.050 766.050 ;
        RECT 463.950 730.950 466.050 733.050 ;
        RECT 461.400 727.350 462.600 729.600 ;
        RECT 457.950 724.950 460.050 727.050 ;
        RECT 460.950 724.950 463.050 727.050 ;
        RECT 463.950 724.950 466.050 727.050 ;
        RECT 458.400 723.900 459.600 724.650 ;
        RECT 457.950 721.800 460.050 723.900 ;
        RECT 464.400 722.400 465.600 724.650 ;
        RECT 464.400 709.050 465.450 722.400 ;
        RECT 473.400 721.050 474.450 763.950 ;
        RECT 472.950 718.950 475.050 721.050 ;
        RECT 476.400 712.050 477.450 790.950 ;
        RECT 482.400 778.050 483.450 800.400 ;
        RECT 487.950 799.800 490.050 801.900 ;
        RECT 493.950 799.800 496.050 801.900 ;
        RECT 506.400 801.450 507.450 826.950 ;
        RECT 518.400 826.050 519.450 839.100 ;
        RECT 524.400 838.350 525.600 839.100 ;
        RECT 530.400 838.350 531.600 839.100 ;
        RECT 523.950 835.950 526.050 838.050 ;
        RECT 526.950 835.950 529.050 838.050 ;
        RECT 529.950 835.950 532.050 838.050 ;
        RECT 527.400 834.900 528.600 835.650 ;
        RECT 526.950 832.800 529.050 834.900 ;
        RECT 517.950 823.950 520.050 826.050 ;
        RECT 536.400 820.050 537.450 847.950 ;
        RECT 538.950 839.100 541.050 841.200 ;
        RECT 529.950 817.950 532.050 820.050 ;
        RECT 535.950 817.950 538.050 820.050 ;
        RECT 523.950 811.950 526.050 814.050 ;
        RECT 509.100 802.950 511.200 805.050 ;
        RECT 512.400 802.950 514.500 805.050 ;
        RECT 517.800 802.950 519.900 805.050 ;
        RECT 509.400 801.450 510.600 802.650 ;
        RECT 518.400 801.900 519.600 802.650 ;
        RECT 506.400 800.400 510.600 801.450 ;
        RECT 517.950 799.800 520.050 801.900 ;
        RECT 478.950 775.950 481.050 778.050 ;
        RECT 481.950 775.950 484.050 778.050 ;
        RECT 479.400 762.600 480.450 775.950 ;
        RECT 487.950 772.950 490.050 775.050 ;
        RECT 488.400 769.050 489.450 772.950 ;
        RECT 487.950 766.950 490.050 769.050 ;
        RECT 488.400 762.600 489.450 766.950 ;
        RECT 494.400 766.050 495.450 799.800 ;
        RECT 502.950 793.950 505.050 796.050 ;
        RECT 496.950 769.950 499.050 772.050 ;
        RECT 493.950 763.950 496.050 766.050 ;
        RECT 479.400 760.350 480.600 762.600 ;
        RECT 488.400 760.350 489.600 762.600 ;
        RECT 490.950 760.950 493.050 763.050 ;
        RECT 479.100 757.950 481.200 760.050 ;
        RECT 484.500 757.950 486.600 760.050 ;
        RECT 487.800 757.950 489.900 760.050 ;
        RECT 479.100 724.950 481.200 727.050 ;
        RECT 484.500 724.950 486.600 727.050 ;
        RECT 487.800 724.950 489.900 727.050 ;
        RECT 479.400 722.400 480.600 724.650 ;
        RECT 488.400 722.400 489.600 724.650 ;
        RECT 479.400 721.050 480.450 722.400 ;
        RECT 478.950 718.950 481.050 721.050 ;
        RECT 475.950 709.950 478.050 712.050 ;
        RECT 463.950 706.950 466.050 709.050 ;
        RECT 454.950 694.950 457.050 697.050 ;
        RECT 455.400 678.900 456.450 694.950 ;
        RECT 463.950 684.000 466.050 688.050 ;
        RECT 475.950 685.950 478.050 688.050 ;
        RECT 464.400 682.350 465.600 684.000 ;
        RECT 460.950 679.950 463.050 682.050 ;
        RECT 463.950 679.950 466.050 682.050 ;
        RECT 466.950 679.950 469.050 682.050 ;
        RECT 461.400 678.900 462.600 679.650 ;
        RECT 454.950 676.800 457.050 678.900 ;
        RECT 460.950 676.800 463.050 678.900 ;
        RECT 467.400 677.400 468.600 679.650 ;
        RECT 467.400 673.050 468.450 677.400 ;
        RECT 466.950 670.950 469.050 673.050 ;
        RECT 476.400 661.050 477.450 685.950 ;
        RECT 475.950 658.950 478.050 661.050 ;
        RECT 463.950 651.000 466.050 655.050 ;
        RECT 464.400 649.350 465.600 651.000 ;
        RECT 460.950 646.950 463.050 649.050 ;
        RECT 463.950 646.950 466.050 649.050 ;
        RECT 466.950 646.950 469.050 649.050 ;
        RECT 461.400 644.400 462.600 646.650 ;
        RECT 467.400 644.400 468.600 646.650 ;
        RECT 461.400 640.050 462.450 644.400 ;
        RECT 460.950 637.950 463.050 640.050 ;
        RECT 467.400 639.450 468.450 644.400 ;
        RECT 467.400 638.400 471.450 639.450 ;
        RECT 451.950 631.950 454.050 634.050 ;
        RECT 454.950 628.950 457.050 631.050 ;
        RECT 436.950 619.950 439.050 622.050 ;
        RECT 437.400 616.050 438.450 619.950 ;
        RECT 436.950 613.950 439.050 616.050 ;
        RECT 455.400 610.050 456.450 628.950 ;
        RECT 461.400 628.050 462.450 637.950 ;
        RECT 466.950 631.950 469.050 634.050 ;
        RECT 460.950 625.950 463.050 628.050 ;
        RECT 425.400 604.350 426.600 606.600 ;
        RECT 430.950 606.000 433.050 610.050 ;
        RECT 436.950 607.950 439.050 610.050 ;
        RECT 431.400 604.350 432.600 606.000 ;
        RECT 421.950 601.950 424.050 604.050 ;
        RECT 424.950 601.950 427.050 604.050 ;
        RECT 427.950 601.950 430.050 604.050 ;
        RECT 430.950 601.950 433.050 604.050 ;
        RECT 422.400 599.400 423.600 601.650 ;
        RECT 428.400 599.400 429.600 601.650 ;
        RECT 437.400 601.050 438.450 607.950 ;
        RECT 448.950 605.100 451.050 607.200 ;
        RECT 454.950 606.000 457.050 610.050 ;
        RECT 449.400 604.350 450.600 605.100 ;
        RECT 455.400 604.350 456.600 606.000 ;
        RECT 448.950 601.950 451.050 604.050 ;
        RECT 451.950 601.950 454.050 604.050 ;
        RECT 454.950 601.950 457.050 604.050 ;
        RECT 422.400 595.050 423.450 599.400 ;
        RECT 421.950 592.950 424.050 595.050 ;
        RECT 415.950 580.950 418.050 583.050 ;
        RECT 406.950 572.100 409.050 574.200 ;
        RECT 412.950 572.100 415.050 574.200 ;
        RECT 407.400 571.350 408.600 572.100 ;
        RECT 406.950 568.950 409.050 571.050 ;
        RECT 397.950 562.950 400.050 565.050 ;
        RECT 401.550 564.300 403.650 566.400 ;
        RECT 384.150 559.500 388.350 560.700 ;
        RECT 386.250 558.600 388.350 559.500 ;
        RECT 401.550 557.700 402.750 564.300 ;
        RECT 412.950 562.950 415.050 565.050 ;
        RECT 376.950 553.950 379.050 556.050 ;
        RECT 401.550 555.600 403.650 557.700 ;
        RECT 358.950 541.950 361.050 544.050 ;
        RECT 373.950 541.950 376.050 544.050 ;
        RECT 364.950 538.950 367.050 541.050 ;
        RECT 358.950 527.100 361.050 529.200 ;
        RECT 365.400 528.600 366.450 538.950 ;
        RECT 359.400 526.350 360.600 527.100 ;
        RECT 365.400 526.350 366.600 528.600 ;
        RECT 358.950 523.950 361.050 526.050 ;
        RECT 361.950 523.950 364.050 526.050 ;
        RECT 364.950 523.950 367.050 526.050 ;
        RECT 362.400 521.400 363.600 523.650 ;
        RECT 362.400 514.050 363.450 521.400 ;
        RECT 361.950 511.950 364.050 514.050 ;
        RECT 352.950 505.950 355.050 508.050 ;
        RECT 340.950 499.950 343.050 502.050 ;
        RECT 344.850 501.300 346.950 503.400 ;
        RECT 332.400 493.350 333.600 494.100 ;
        RECT 337.950 493.950 340.050 496.050 ;
        RECT 325.950 490.950 328.050 493.050 ;
        RECT 328.950 490.950 331.050 493.050 ;
        RECT 331.950 490.950 334.050 493.050 ;
        RECT 334.950 490.950 337.050 493.050 ;
        RECT 340.950 490.950 343.050 493.050 ;
        RECT 329.400 489.900 330.600 490.650 ;
        RECT 335.400 489.900 336.600 490.650 ;
        RECT 319.950 487.800 322.050 489.900 ;
        RECT 328.950 487.800 331.050 489.900 ;
        RECT 334.950 487.800 337.050 489.900 ;
        RECT 341.400 488.400 342.600 490.650 ;
        RECT 341.400 478.050 342.450 488.400 ;
        RECT 345.150 482.700 346.350 501.300 ;
        RECT 353.400 496.050 354.450 505.950 ;
        RECT 358.950 499.950 361.050 502.050 ;
        RECT 362.550 501.300 364.650 503.400 ;
        RECT 352.950 493.950 355.050 496.050 ;
        RECT 350.100 490.950 352.200 493.050 ;
        RECT 350.400 489.900 351.600 490.650 ;
        RECT 349.950 487.800 352.050 489.900 ;
        RECT 359.400 487.050 360.450 499.950 ;
        RECT 362.550 488.400 363.750 501.300 ;
        RECT 367.950 499.950 370.050 502.050 ;
        RECT 368.400 495.600 369.450 499.950 ;
        RECT 368.400 493.350 369.600 495.600 ;
        RECT 367.950 490.950 370.050 493.050 ;
        RECT 358.950 484.950 361.050 487.050 ;
        RECT 362.550 486.300 364.650 488.400 ;
        RECT 345.150 481.500 349.350 482.700 ;
        RECT 347.250 480.600 349.350 481.500 ;
        RECT 362.550 479.700 363.750 486.300 ;
        RECT 340.950 475.950 343.050 478.050 ;
        RECT 362.550 477.600 364.650 479.700 ;
        RECT 340.950 466.950 343.050 469.050 ;
        RECT 319.950 454.950 322.050 457.050 ;
        RECT 314.400 452.400 318.450 453.450 ;
        RECT 314.400 450.600 315.450 452.400 ;
        RECT 320.400 450.600 321.450 454.950 ;
        RECT 314.400 448.350 315.600 450.600 ;
        RECT 320.400 448.350 321.600 450.600 ;
        RECT 325.950 449.100 328.050 451.200 ;
        RECT 334.950 449.100 337.050 454.050 ;
        RECT 341.400 450.600 342.450 466.950 ;
        RECT 355.950 463.950 358.050 466.050 ;
        RECT 310.950 445.950 313.050 448.050 ;
        RECT 313.950 445.950 316.050 448.050 ;
        RECT 316.950 445.950 319.050 448.050 ;
        RECT 319.950 445.950 322.050 448.050 ;
        RECT 311.400 444.900 312.600 445.650 ;
        RECT 289.950 442.800 292.050 444.900 ;
        RECT 298.950 442.800 301.050 444.900 ;
        RECT 310.950 442.800 313.050 444.900 ;
        RECT 317.400 443.400 318.600 445.650 ;
        RECT 280.950 436.950 283.050 439.050 ;
        RECT 289.950 436.950 292.050 439.050 ;
        RECT 268.950 433.950 271.050 436.050 ;
        RECT 233.400 431.400 237.450 432.450 ;
        RECT 214.950 427.950 217.050 430.050 ;
        RECT 215.400 411.900 216.450 427.950 ;
        RECT 223.950 424.950 226.050 427.050 ;
        RECT 224.400 417.600 225.450 424.950 ;
        RECT 229.950 421.950 232.050 424.050 ;
        RECT 230.400 417.600 231.450 421.950 ;
        RECT 224.400 415.350 225.600 417.600 ;
        RECT 230.400 415.350 231.600 417.600 ;
        RECT 220.950 412.950 223.050 415.050 ;
        RECT 223.950 412.950 226.050 415.050 ;
        RECT 226.950 412.950 229.050 415.050 ;
        RECT 229.950 412.950 232.050 415.050 ;
        RECT 214.950 409.800 217.050 411.900 ;
        RECT 221.400 410.400 222.600 412.650 ;
        RECT 227.400 411.900 228.600 412.650 ;
        RECT 221.400 397.050 222.450 410.400 ;
        RECT 226.950 409.800 229.050 411.900 ;
        RECT 236.400 411.450 237.450 431.400 ;
        RECT 238.950 430.950 241.050 433.050 ;
        RECT 250.800 430.950 252.900 433.050 ;
        RECT 253.950 430.950 256.050 433.050 ;
        RECT 239.400 411.900 240.450 430.950 ;
        RECT 265.950 427.950 268.050 430.050 ;
        RECT 241.950 416.100 244.050 418.200 ;
        RECT 247.950 416.100 250.050 418.200 ;
        RECT 253.950 416.100 256.050 418.200 ;
        RECT 233.400 410.400 237.450 411.450 ;
        RECT 211.950 394.950 214.050 397.050 ;
        RECT 220.950 394.950 223.050 397.050 ;
        RECT 212.550 381.300 214.650 383.400 ;
        RECT 197.250 379.500 199.350 380.400 ;
        RECT 190.950 376.950 193.050 379.050 ;
        RECT 195.150 378.300 199.350 379.500 ;
        RECT 191.400 373.200 192.450 376.950 ;
        RECT 143.400 370.350 144.600 372.600 ;
        RECT 151.950 370.950 154.050 373.050 ;
        RECT 160.950 371.100 163.050 373.200 ;
        RECT 175.950 370.950 178.050 373.050 ;
        RECT 181.950 371.100 184.050 373.200 ;
        RECT 190.950 371.100 193.050 373.200 ;
        RECT 139.950 367.950 142.050 370.050 ;
        RECT 142.950 367.950 145.050 370.050 ;
        RECT 145.950 367.950 148.050 370.050 ;
        RECT 140.400 366.900 141.600 367.650 ;
        RECT 139.950 364.800 142.050 366.900 ;
        RECT 146.400 365.400 147.600 367.650 ;
        RECT 152.400 366.900 153.450 370.950 ;
        RECT 163.800 367.950 165.900 370.050 ;
        RECT 146.400 361.050 147.450 365.400 ;
        RECT 151.950 364.800 154.050 366.900 ;
        RECT 136.950 358.950 139.050 361.050 ;
        RECT 145.950 358.950 148.050 361.050 ;
        RECT 137.400 298.050 138.450 358.950 ;
        RECT 176.400 355.050 177.450 370.950 ;
        RECT 182.400 370.350 183.600 371.100 ;
        RECT 191.400 370.350 192.600 371.100 ;
        RECT 181.800 367.950 183.900 370.050 ;
        RECT 190.950 367.950 193.050 370.050 ;
        RECT 195.150 359.700 196.350 378.300 ;
        RECT 212.550 374.700 213.750 381.300 ;
        RECT 199.950 371.100 202.050 373.200 ;
        RECT 208.950 371.100 211.050 373.200 ;
        RECT 212.550 372.600 214.650 374.700 ;
        RECT 200.400 370.350 201.600 371.100 ;
        RECT 200.100 367.950 202.200 370.050 ;
        RECT 194.850 357.600 196.950 359.700 ;
        RECT 175.950 352.950 178.050 355.050 ;
        RECT 142.950 338.100 145.050 340.200 ;
        RECT 151.950 338.100 154.050 340.200 ;
        RECT 163.950 339.000 166.050 343.050 ;
        RECT 143.400 337.350 144.600 338.100 ;
        RECT 142.950 334.950 145.050 337.050 ;
        RECT 145.950 334.950 148.050 337.050 ;
        RECT 146.400 332.400 147.600 334.650 ;
        RECT 152.400 334.050 153.450 338.100 ;
        RECT 164.400 337.350 165.600 339.000 ;
        RECT 169.950 338.100 172.050 340.200 ;
        RECT 170.400 337.350 171.600 338.100 ;
        RECT 160.950 334.950 163.050 337.050 ;
        RECT 163.950 334.950 166.050 337.050 ;
        RECT 166.950 334.950 169.050 337.050 ;
        RECT 169.950 334.950 172.050 337.050 ;
        RECT 146.400 328.050 147.450 332.400 ;
        RECT 151.950 331.950 154.050 334.050 ;
        RECT 161.400 332.400 162.600 334.650 ;
        RECT 167.400 333.900 168.600 334.650 ;
        RECT 176.400 333.900 177.450 352.950 ;
        RECT 187.950 343.950 190.050 346.050 ;
        RECT 199.950 343.950 202.050 346.050 ;
        RECT 188.400 339.600 189.450 343.950 ;
        RECT 188.400 337.350 189.600 339.600 ;
        RECT 184.950 334.950 187.050 337.050 ;
        RECT 187.950 334.950 190.050 337.050 ;
        RECT 190.950 334.950 193.050 337.050 ;
        RECT 191.400 333.900 192.600 334.650 ;
        RECT 200.400 333.900 201.450 343.950 ;
        RECT 209.400 339.600 210.450 371.100 ;
        RECT 212.550 359.700 213.750 372.600 ;
        RECT 226.950 371.100 229.050 373.200 ;
        RECT 217.950 367.950 220.050 370.050 ;
        RECT 218.400 365.400 219.600 367.650 ;
        RECT 212.550 357.600 214.650 359.700 ;
        RECT 214.950 352.950 217.050 355.050 ;
        RECT 215.400 339.600 216.450 352.950 ;
        RECT 218.400 351.450 219.450 365.400 ;
        RECT 218.400 350.400 222.450 351.450 ;
        RECT 209.400 337.350 210.600 339.600 ;
        RECT 215.400 337.350 216.600 339.600 ;
        RECT 205.950 334.950 208.050 337.050 ;
        RECT 208.950 334.950 211.050 337.050 ;
        RECT 211.950 334.950 214.050 337.050 ;
        RECT 214.950 334.950 217.050 337.050 ;
        RECT 206.400 333.900 207.600 334.650 ;
        RECT 161.400 331.050 162.450 332.400 ;
        RECT 166.950 331.800 169.050 333.900 ;
        RECT 175.950 331.800 178.050 333.900 ;
        RECT 190.950 331.800 193.050 333.900 ;
        RECT 199.950 331.800 202.050 333.900 ;
        RECT 205.950 331.800 208.050 333.900 ;
        RECT 212.400 332.400 213.600 334.650 ;
        RECT 160.950 328.950 163.050 331.050 ;
        RECT 145.950 325.950 148.050 328.050 ;
        RECT 146.400 319.050 147.450 325.950 ;
        RECT 145.950 316.950 148.050 319.050 ;
        RECT 157.950 301.950 160.050 304.050 ;
        RECT 136.950 295.950 139.050 298.050 ;
        RECT 142.950 293.100 145.050 295.200 ;
        RECT 148.950 294.000 151.050 298.050 ;
        RECT 143.400 292.350 144.600 293.100 ;
        RECT 149.400 292.350 150.600 294.000 ;
        RECT 142.950 289.950 145.050 292.050 ;
        RECT 145.950 289.950 148.050 292.050 ;
        RECT 148.950 289.950 151.050 292.050 ;
        RECT 151.950 289.950 154.050 292.050 ;
        RECT 146.400 287.400 147.600 289.650 ;
        RECT 152.400 287.400 153.600 289.650 ;
        RECT 146.400 283.050 147.450 287.400 ;
        RECT 136.950 280.950 139.050 283.050 ;
        RECT 145.950 280.950 148.050 283.050 ;
        RECT 122.400 259.350 123.600 260.100 ;
        RECT 128.400 259.350 129.600 261.600 ;
        RECT 133.950 259.950 136.050 262.050 ;
        RECT 121.950 256.950 124.050 259.050 ;
        RECT 124.950 256.950 127.050 259.050 ;
        RECT 127.950 256.950 130.050 259.050 ;
        RECT 130.950 256.950 133.050 259.050 ;
        RECT 125.400 255.900 126.600 256.650 ;
        RECT 131.400 255.900 132.600 256.650 ;
        RECT 115.950 253.800 118.050 255.900 ;
        RECT 121.950 250.950 124.050 253.050 ;
        RECT 124.950 250.950 127.050 255.900 ;
        RECT 130.950 253.800 133.050 255.900 ;
        RECT 133.950 250.950 136.050 253.050 ;
        RECT 112.950 241.950 115.050 244.050 ;
        RECT 100.950 235.950 103.050 238.050 ;
        RECT 112.950 232.950 115.050 235.050 ;
        RECT 83.400 214.350 84.600 215.100 ;
        RECT 89.400 214.350 90.600 216.600 ;
        RECT 97.950 214.950 100.050 217.050 ;
        RECT 106.950 215.100 109.050 217.200 ;
        RECT 113.400 216.600 114.450 232.950 ;
        RECT 82.950 211.950 85.050 214.050 ;
        RECT 85.950 211.950 88.050 214.050 ;
        RECT 88.950 211.950 91.050 214.050 ;
        RECT 91.950 211.950 94.050 214.050 ;
        RECT 86.400 209.400 87.600 211.650 ;
        RECT 92.400 209.400 93.600 211.650 ;
        RECT 86.400 199.050 87.450 209.400 ;
        RECT 85.950 196.950 88.050 199.050 ;
        RECT 92.400 196.050 93.450 209.400 ;
        RECT 91.950 193.950 94.050 196.050 ;
        RECT 85.950 183.000 88.050 187.050 ;
        RECT 86.400 181.350 87.600 183.000 ;
        RECT 91.950 182.100 94.050 184.200 ;
        RECT 92.400 181.350 93.600 182.100 ;
        RECT 82.950 178.950 85.050 181.050 ;
        RECT 85.950 178.950 88.050 181.050 ;
        RECT 88.950 178.950 91.050 181.050 ;
        RECT 91.950 178.950 94.050 181.050 ;
        RECT 83.400 176.400 84.600 178.650 ;
        RECT 89.400 177.000 90.600 178.650 ;
        RECT 76.950 172.950 79.050 175.050 ;
        RECT 83.400 172.050 84.450 176.400 ;
        RECT 88.950 172.950 91.050 177.000 ;
        RECT 94.950 175.950 97.050 178.050 ;
        RECT 82.950 169.950 85.050 172.050 ;
        RECT 73.950 160.950 76.050 163.050 ;
        RECT 67.950 154.950 70.050 157.050 ;
        RECT 61.950 142.950 64.050 145.050 ;
        RECT 52.950 136.950 55.050 139.050 ;
        RECT 61.950 137.100 64.050 139.200 ;
        RECT 68.400 138.600 69.450 154.950 ;
        RECT 62.400 136.350 63.600 137.100 ;
        RECT 68.400 136.350 69.600 138.600 ;
        RECT 58.950 133.950 61.050 136.050 ;
        RECT 61.950 133.950 64.050 136.050 ;
        RECT 64.950 133.950 67.050 136.050 ;
        RECT 67.950 133.950 70.050 136.050 ;
        RECT 43.950 130.800 46.050 132.900 ;
        RECT 49.950 130.800 52.050 132.900 ;
        RECT 59.400 131.400 60.600 133.650 ;
        RECT 65.400 132.000 66.600 133.650 ;
        RECT 34.950 124.950 37.050 127.050 ;
        RECT 43.950 121.950 46.050 124.050 ;
        RECT 28.950 106.950 31.050 109.050 ;
        RECT 16.950 104.100 19.050 106.200 ;
        RECT 17.400 103.350 18.600 104.100 ;
        RECT 25.950 103.950 28.050 106.050 ;
        RECT 16.950 100.950 19.050 103.050 ;
        RECT 19.950 100.950 22.050 103.050 ;
        RECT 20.400 99.900 21.600 100.650 ;
        RECT 19.950 97.800 22.050 99.900 ;
        RECT 26.400 79.050 27.450 103.950 ;
        RECT 19.950 76.950 22.050 79.050 ;
        RECT 25.950 76.950 28.050 79.050 ;
        RECT 20.400 60.600 21.450 76.950 ;
        RECT 20.400 58.350 21.600 60.600 ;
        RECT 26.400 60.450 27.600 60.600 ;
        RECT 29.400 60.450 30.450 106.950 ;
        RECT 37.950 104.100 40.050 109.050 ;
        RECT 44.400 105.600 45.450 121.950 ;
        RECT 38.400 103.350 39.600 104.100 ;
        RECT 44.400 103.350 45.600 105.600 ;
        RECT 34.950 100.950 37.050 103.050 ;
        RECT 37.950 100.950 40.050 103.050 ;
        RECT 40.950 100.950 43.050 103.050 ;
        RECT 43.950 100.950 46.050 103.050 ;
        RECT 35.400 99.900 36.600 100.650 ;
        RECT 34.950 97.800 37.050 99.900 ;
        RECT 41.400 98.400 42.600 100.650 ;
        RECT 35.400 91.050 36.450 97.800 ;
        RECT 41.400 94.050 42.450 98.400 ;
        RECT 40.950 91.950 43.050 94.050 ;
        RECT 34.950 88.950 37.050 91.050 ;
        RECT 50.400 64.050 51.450 130.800 ;
        RECT 52.950 124.950 55.050 127.050 ;
        RECT 53.400 99.900 54.450 124.950 ;
        RECT 59.400 108.450 60.450 131.400 ;
        RECT 64.950 127.950 67.050 132.000 ;
        RECT 74.400 112.050 75.450 160.950 ;
        RECT 85.950 148.950 88.050 151.050 ;
        RECT 86.400 138.600 87.450 148.950 ;
        RECT 95.400 145.050 96.450 175.950 ;
        RECT 98.400 172.050 99.450 214.950 ;
        RECT 107.400 214.350 108.600 215.100 ;
        RECT 113.400 214.350 114.600 216.600 ;
        RECT 106.950 211.950 109.050 214.050 ;
        RECT 109.950 211.950 112.050 214.050 ;
        RECT 112.950 211.950 115.050 214.050 ;
        RECT 115.950 211.950 118.050 214.050 ;
        RECT 110.400 210.000 111.600 211.650 ;
        RECT 109.950 205.950 112.050 210.000 ;
        RECT 116.400 209.400 117.600 211.650 ;
        RECT 116.400 199.050 117.450 209.400 ;
        RECT 115.950 196.950 118.050 199.050 ;
        RECT 100.950 190.950 103.050 193.050 ;
        RECT 97.950 169.950 100.050 172.050 ;
        RECT 94.950 142.950 97.050 145.050 ;
        RECT 86.400 136.350 87.600 138.600 ;
        RECT 91.950 137.100 94.050 139.200 ;
        RECT 92.400 136.350 93.600 137.100 ;
        RECT 82.950 133.950 85.050 136.050 ;
        RECT 85.950 133.950 88.050 136.050 ;
        RECT 88.950 133.950 91.050 136.050 ;
        RECT 91.950 133.950 94.050 136.050 ;
        RECT 83.400 131.400 84.600 133.650 ;
        RECT 89.400 131.400 90.600 133.650 ;
        RECT 83.400 124.050 84.450 131.400 ;
        RECT 82.950 121.950 85.050 124.050 ;
        RECT 89.400 118.050 90.450 131.400 ;
        RECT 88.950 115.950 91.050 118.050 ;
        RECT 97.950 115.950 100.050 118.050 ;
        RECT 79.950 112.950 82.050 115.050 ;
        RECT 73.950 109.950 76.050 112.050 ;
        RECT 59.400 107.400 63.450 108.450 ;
        RECT 62.400 106.200 63.450 107.400 ;
        RECT 61.950 104.100 64.050 106.200 ;
        RECT 67.950 104.100 70.050 106.200 ;
        RECT 62.400 103.350 63.600 104.100 ;
        RECT 68.400 103.350 69.600 104.100 ;
        RECT 58.950 100.950 61.050 103.050 ;
        RECT 61.950 100.950 64.050 103.050 ;
        RECT 64.950 100.950 67.050 103.050 ;
        RECT 67.950 100.950 70.050 103.050 ;
        RECT 59.400 99.900 60.600 100.650 ;
        RECT 52.950 97.800 55.050 99.900 ;
        RECT 58.950 97.800 61.050 99.900 ;
        RECT 65.400 98.400 66.600 100.650 ;
        RECT 53.400 94.050 54.450 97.800 ;
        RECT 52.950 91.950 55.050 94.050 ;
        RECT 65.400 91.050 66.450 98.400 ;
        RECT 64.950 88.950 67.050 91.050 ;
        RECT 52.950 76.950 55.050 79.050 ;
        RECT 45.000 63.450 49.050 64.050 ;
        RECT 44.400 61.950 49.050 63.450 ;
        RECT 49.950 61.950 52.050 64.050 ;
        RECT 44.400 60.600 45.450 61.950 ;
        RECT 26.400 59.400 33.450 60.450 ;
        RECT 26.400 58.350 27.600 59.400 ;
        RECT 16.950 55.950 19.050 58.050 ;
        RECT 19.950 55.950 22.050 58.050 ;
        RECT 22.950 55.950 25.050 58.050 ;
        RECT 25.950 55.950 28.050 58.050 ;
        RECT 17.400 54.900 18.600 55.650 ;
        RECT 16.950 52.800 19.050 54.900 ;
        RECT 23.400 53.400 24.600 55.650 ;
        RECT 32.400 54.900 33.450 59.400 ;
        RECT 44.400 58.350 45.600 60.600 ;
        RECT 50.400 58.050 51.450 61.950 ;
        RECT 40.950 55.950 43.050 58.050 ;
        RECT 43.950 55.950 46.050 58.050 ;
        RECT 49.950 55.950 52.050 58.050 ;
        RECT 41.400 54.900 42.600 55.650 ;
        RECT 53.400 54.900 54.450 76.950 ;
        RECT 61.950 60.000 64.050 64.050 ;
        RECT 67.950 60.000 70.050 64.050 ;
        RECT 62.400 58.350 63.600 60.000 ;
        RECT 68.400 58.350 69.600 60.000 ;
        RECT 58.950 55.950 61.050 58.050 ;
        RECT 61.950 55.950 64.050 58.050 ;
        RECT 64.950 55.950 67.050 58.050 ;
        RECT 67.950 55.950 70.050 58.050 ;
        RECT 59.400 54.900 60.600 55.650 ;
        RECT 65.400 54.900 66.600 55.650 ;
        RECT 16.950 46.950 19.050 49.050 ;
        RECT 17.400 27.600 18.450 46.950 ;
        RECT 23.400 40.050 24.450 53.400 ;
        RECT 31.950 52.800 34.050 54.900 ;
        RECT 40.950 52.800 43.050 54.900 ;
        RECT 52.950 52.800 55.050 54.900 ;
        RECT 58.950 52.800 61.050 54.900 ;
        RECT 64.950 52.800 67.050 54.900 ;
        RECT 74.400 49.050 75.450 109.950 ;
        RECT 80.400 106.050 81.450 112.950 ;
        RECT 88.950 112.800 91.050 114.900 ;
        RECT 79.800 103.950 81.900 106.050 ;
        RECT 82.950 104.100 85.050 106.200 ;
        RECT 89.400 105.600 90.450 112.800 ;
        RECT 83.400 103.350 84.600 104.100 ;
        RECT 89.400 103.350 90.600 105.600 ;
        RECT 82.950 100.950 85.050 103.050 ;
        RECT 85.950 100.950 88.050 103.050 ;
        RECT 88.950 100.950 91.050 103.050 ;
        RECT 91.950 100.950 94.050 103.050 ;
        RECT 86.400 98.400 87.600 100.650 ;
        RECT 92.400 99.000 93.600 100.650 ;
        RECT 86.400 94.050 87.450 98.400 ;
        RECT 91.950 94.950 94.050 99.000 ;
        RECT 94.950 97.950 97.050 100.050 ;
        RECT 85.950 91.950 88.050 94.050 ;
        RECT 86.400 70.050 87.450 91.950 ;
        RECT 76.950 67.950 79.050 70.050 ;
        RECT 85.950 67.950 88.050 70.050 ;
        RECT 77.400 55.050 78.450 67.950 ;
        RECT 95.400 64.050 96.450 97.950 ;
        RECT 98.400 76.050 99.450 115.950 ;
        RECT 101.400 97.050 102.450 190.950 ;
        RECT 116.400 184.200 117.450 196.950 ;
        RECT 118.950 187.950 121.050 190.050 ;
        RECT 106.950 182.100 109.050 184.200 ;
        RECT 113.400 183.450 114.600 183.600 ;
        RECT 115.950 183.450 118.050 184.200 ;
        RECT 113.400 182.400 118.050 183.450 ;
        RECT 107.400 181.350 108.600 182.100 ;
        RECT 113.400 181.350 114.600 182.400 ;
        RECT 115.950 182.100 118.050 182.400 ;
        RECT 106.950 178.950 109.050 181.050 ;
        RECT 109.950 178.950 112.050 181.050 ;
        RECT 112.950 178.950 115.050 181.050 ;
        RECT 110.400 176.400 111.600 178.650 ;
        RECT 110.400 169.050 111.450 176.400 ;
        RECT 109.950 166.950 112.050 169.050 ;
        RECT 109.950 137.100 112.050 139.200 ;
        RECT 110.400 136.350 111.600 137.100 ;
        RECT 106.950 133.950 109.050 136.050 ;
        RECT 109.950 133.950 112.050 136.050 ;
        RECT 107.400 131.400 108.600 133.650 ;
        RECT 107.400 124.050 108.450 131.400 ;
        RECT 119.400 130.050 120.450 187.950 ;
        RECT 118.950 127.950 121.050 130.050 ;
        RECT 106.950 121.950 109.050 124.050 ;
        RECT 109.950 112.950 112.050 115.050 ;
        RECT 110.400 105.600 111.450 112.950 ;
        RECT 122.400 108.450 123.450 250.950 ;
        RECT 124.950 217.950 127.050 220.050 ;
        RECT 125.400 208.050 126.450 217.950 ;
        RECT 134.400 216.600 135.450 250.950 ;
        RECT 137.400 220.050 138.450 280.950 ;
        RECT 152.400 268.050 153.450 287.400 ;
        RECT 158.400 280.050 159.450 301.950 ;
        RECT 157.950 277.950 160.050 280.050 ;
        RECT 157.950 271.950 160.050 274.050 ;
        RECT 148.800 265.950 150.900 268.050 ;
        RECT 151.950 265.950 154.050 268.050 ;
        RECT 149.400 261.600 150.450 265.950 ;
        RECT 149.400 259.350 150.600 261.600 ;
        RECT 145.950 256.950 148.050 259.050 ;
        RECT 148.950 256.950 151.050 259.050 ;
        RECT 151.950 256.950 154.050 259.050 ;
        RECT 146.400 255.900 147.600 256.650 ;
        RECT 139.950 253.800 142.050 255.900 ;
        RECT 145.950 253.800 148.050 255.900 ;
        RECT 152.400 255.000 153.600 256.650 ;
        RECT 140.400 241.050 141.450 253.800 ;
        RECT 151.950 250.950 154.050 255.000 ;
        RECT 139.950 238.950 142.050 241.050 ;
        RECT 136.950 217.950 139.050 220.050 ;
        RECT 140.400 216.600 141.450 238.950 ;
        RECT 158.400 238.050 159.450 271.950 ;
        RECT 161.400 255.900 162.450 328.950 ;
        RECT 212.400 325.050 213.450 332.400 ;
        RECT 221.400 331.050 222.450 350.400 ;
        RECT 227.400 333.450 228.450 371.100 ;
        RECT 233.400 367.050 234.450 410.400 ;
        RECT 238.950 409.800 241.050 411.900 ;
        RECT 242.400 406.050 243.450 416.100 ;
        RECT 248.400 415.350 249.600 416.100 ;
        RECT 254.400 415.350 255.600 416.100 ;
        RECT 262.950 415.950 265.050 418.050 ;
        RECT 247.950 412.950 250.050 415.050 ;
        RECT 250.950 412.950 253.050 415.050 ;
        RECT 253.950 412.950 256.050 415.050 ;
        RECT 256.950 412.950 259.050 415.050 ;
        RECT 251.400 411.900 252.600 412.650 ;
        RECT 250.950 409.800 253.050 411.900 ;
        RECT 257.400 410.400 258.600 412.650 ;
        RECT 257.400 406.050 258.450 410.400 ;
        RECT 263.400 409.050 264.450 415.950 ;
        RECT 266.400 411.900 267.450 427.950 ;
        RECT 271.950 421.950 274.050 424.050 ;
        RECT 272.400 417.600 273.450 421.950 ;
        RECT 272.400 415.350 273.600 417.600 ;
        RECT 277.950 416.100 280.050 418.200 ;
        RECT 278.400 415.350 279.600 416.100 ;
        RECT 286.950 415.950 289.050 418.050 ;
        RECT 271.950 412.950 274.050 415.050 ;
        RECT 274.950 412.950 277.050 415.050 ;
        RECT 277.950 412.950 280.050 415.050 ;
        RECT 280.950 412.950 283.050 415.050 ;
        RECT 275.400 411.900 276.600 412.650 ;
        RECT 281.400 411.900 282.600 412.650 ;
        RECT 265.950 409.800 268.050 411.900 ;
        RECT 274.950 409.800 277.050 411.900 ;
        RECT 280.950 409.800 283.050 411.900 ;
        RECT 262.950 406.950 265.050 409.050 ;
        RECT 241.950 403.950 244.050 406.050 ;
        RECT 256.950 403.950 259.050 406.050 ;
        RECT 274.950 405.450 277.050 408.750 ;
        RECT 287.400 406.050 288.450 415.950 ;
        RECT 290.400 409.050 291.450 436.950 ;
        RECT 317.400 433.050 318.450 443.400 ;
        RECT 316.950 430.950 319.050 433.050 ;
        RECT 298.950 427.950 301.050 430.050 ;
        RECT 292.950 415.950 295.050 418.050 ;
        RECT 299.400 417.600 300.450 427.950 ;
        RECT 304.950 421.950 307.050 424.050 ;
        RECT 314.850 423.300 316.950 425.400 ;
        RECT 305.400 417.600 306.450 421.950 ;
        RECT 293.400 411.900 294.450 415.950 ;
        RECT 299.400 415.350 300.600 417.600 ;
        RECT 305.400 415.350 306.600 417.600 ;
        RECT 298.950 412.950 301.050 415.050 ;
        RECT 301.950 412.950 304.050 415.050 ;
        RECT 304.950 412.950 307.050 415.050 ;
        RECT 310.950 412.950 313.050 415.050 ;
        RECT 292.950 409.800 295.050 411.900 ;
        RECT 302.400 410.400 303.600 412.650 ;
        RECT 311.400 410.400 312.600 412.650 ;
        RECT 289.950 406.950 292.050 409.050 ;
        RECT 295.950 406.950 301.050 409.050 ;
        RECT 280.950 405.450 283.050 406.050 ;
        RECT 274.950 405.000 283.050 405.450 ;
        RECT 275.400 404.400 283.050 405.000 ;
        RECT 280.950 403.950 283.050 404.400 ;
        RECT 286.950 403.950 289.050 406.050 ;
        RECT 294.000 405.900 297.000 406.050 ;
        RECT 292.950 403.950 298.050 405.900 ;
        RECT 292.950 403.800 295.050 403.950 ;
        RECT 295.950 403.800 298.050 403.950 ;
        RECT 302.400 400.050 303.450 410.400 ;
        RECT 311.400 409.050 312.450 410.400 ;
        RECT 310.950 406.950 313.050 409.050 ;
        RECT 268.950 397.950 271.050 400.050 ;
        RECT 301.950 397.950 304.050 400.050 ;
        RECT 238.950 371.100 241.050 373.200 ;
        RECT 244.950 371.100 247.050 373.200 ;
        RECT 256.950 371.100 259.050 373.200 ;
        RECT 239.400 370.350 240.600 371.100 ;
        RECT 245.400 370.350 246.600 371.100 ;
        RECT 238.950 367.950 241.050 370.050 ;
        RECT 241.950 367.950 244.050 370.050 ;
        RECT 244.950 367.950 247.050 370.050 ;
        RECT 232.950 364.950 235.050 367.050 ;
        RECT 242.400 366.900 243.600 367.650 ;
        RECT 241.950 364.800 244.050 366.900 ;
        RECT 235.950 338.100 238.050 340.200 ;
        RECT 236.400 337.350 237.600 338.100 ;
        RECT 244.950 337.950 247.050 340.050 ;
        RECT 257.400 339.600 258.450 371.100 ;
        RECT 265.800 367.950 267.900 370.050 ;
        RECT 230.100 334.950 232.200 337.050 ;
        RECT 235.500 334.950 237.600 337.050 ;
        RECT 238.800 334.950 240.900 337.050 ;
        RECT 230.400 333.450 231.600 334.650 ;
        RECT 239.400 333.900 240.600 334.650 ;
        RECT 227.400 332.400 231.600 333.450 ;
        RECT 220.950 328.950 223.050 331.050 ;
        RECT 211.950 322.950 214.050 325.050 ;
        RECT 175.950 301.950 178.050 304.050 ;
        RECT 163.950 292.950 166.050 295.050 ;
        RECT 176.400 294.600 177.450 301.950 ;
        RECT 198.000 300.450 202.050 301.050 ;
        RECT 197.400 298.950 202.050 300.450 ;
        RECT 217.950 298.950 220.050 301.050 ;
        RECT 197.400 294.600 198.450 298.950 ;
        RECT 202.950 295.950 205.050 298.050 ;
        RECT 160.950 253.800 163.050 255.900 ;
        RECT 157.950 235.950 160.050 238.050 ;
        RECT 161.400 229.050 162.450 253.800 ;
        RECT 160.950 226.950 163.050 229.050 ;
        RECT 164.400 217.200 165.450 292.950 ;
        RECT 176.400 292.350 177.600 294.600 ;
        RECT 197.400 292.350 198.600 294.600 ;
        RECT 169.950 289.950 172.050 292.050 ;
        RECT 172.950 289.950 175.050 292.050 ;
        RECT 175.950 289.950 178.050 292.050 ;
        RECT 193.950 289.950 196.050 292.050 ;
        RECT 196.950 289.950 199.050 292.050 ;
        RECT 173.400 287.400 174.600 289.650 ;
        RECT 194.400 287.400 195.600 289.650 ;
        RECT 203.400 288.450 204.450 295.950 ;
        RECT 211.950 294.000 214.050 298.050 ;
        RECT 218.400 294.600 219.450 298.950 ;
        RECT 212.400 292.350 213.600 294.000 ;
        RECT 218.400 292.350 219.600 294.600 ;
        RECT 211.950 289.950 214.050 292.050 ;
        RECT 214.950 289.950 217.050 292.050 ;
        RECT 217.950 289.950 220.050 292.050 ;
        RECT 220.950 289.950 223.050 292.050 ;
        RECT 215.400 288.900 216.600 289.650 ;
        RECT 200.400 287.400 204.450 288.450 ;
        RECT 173.400 283.050 174.450 287.400 ;
        RECT 172.950 280.950 175.050 283.050 ;
        RECT 172.950 277.800 175.050 279.900 ;
        RECT 173.400 261.600 174.450 277.800 ;
        RECT 194.400 271.050 195.450 287.400 ;
        RECT 193.950 268.950 196.050 271.050 ;
        RECT 190.950 265.950 193.050 268.050 ;
        RECT 191.400 262.200 192.450 265.950 ;
        RECT 173.400 259.350 174.600 261.600 ;
        RECT 190.950 260.100 193.050 262.200 ;
        RECT 200.400 262.050 201.450 287.400 ;
        RECT 214.950 286.800 217.050 288.900 ;
        RECT 221.400 288.000 222.600 289.650 ;
        RECT 220.950 283.950 223.050 288.000 ;
        RECT 223.950 286.800 226.050 288.900 ;
        RECT 214.950 277.950 217.050 280.050 ;
        RECT 202.950 268.950 205.050 271.050 ;
        RECT 208.950 268.950 211.050 271.050 ;
        RECT 191.400 259.350 192.600 260.100 ;
        RECT 199.950 259.950 202.050 262.050 ;
        RECT 167.100 256.950 169.200 259.050 ;
        RECT 172.500 256.950 174.600 259.050 ;
        RECT 190.950 256.950 193.050 259.050 ;
        RECT 193.950 256.950 196.050 259.050 ;
        RECT 167.400 255.000 168.600 256.650 ;
        RECT 194.400 255.900 195.600 256.650 ;
        RECT 166.950 250.950 169.050 255.000 ;
        RECT 193.950 253.800 196.050 255.900 ;
        RECT 134.400 214.350 135.600 216.600 ;
        RECT 140.400 214.350 141.600 216.600 ;
        RECT 145.950 214.950 148.050 217.050 ;
        RECT 157.950 215.100 160.050 217.200 ;
        RECT 163.950 215.100 166.050 217.200 ;
        RECT 130.950 211.950 133.050 214.050 ;
        RECT 133.950 211.950 136.050 214.050 ;
        RECT 136.950 211.950 139.050 214.050 ;
        RECT 139.950 211.950 142.050 214.050 ;
        RECT 131.400 209.400 132.600 211.650 ;
        RECT 137.400 209.400 138.600 211.650 ;
        RECT 124.950 205.950 127.050 208.050 ;
        RECT 131.400 193.050 132.450 209.400 ;
        RECT 130.950 190.950 133.050 193.050 ;
        RECT 137.400 190.050 138.450 209.400 ;
        RECT 142.950 196.950 145.050 199.050 ;
        RECT 136.950 187.950 139.050 190.050 ;
        RECT 127.950 182.100 130.050 184.200 ;
        RECT 133.950 182.100 136.050 184.200 ;
        RECT 128.400 181.350 129.600 182.100 ;
        RECT 134.400 181.350 135.600 182.100 ;
        RECT 127.950 178.950 130.050 181.050 ;
        RECT 130.950 178.950 133.050 181.050 ;
        RECT 133.950 178.950 136.050 181.050 ;
        RECT 136.950 178.950 139.050 181.050 ;
        RECT 131.400 176.400 132.600 178.650 ;
        RECT 137.400 177.900 138.600 178.650 ;
        RECT 131.400 175.050 132.450 176.400 ;
        RECT 136.950 175.800 139.050 177.900 ;
        RECT 130.950 172.950 133.050 175.050 ;
        RECT 131.400 151.050 132.450 172.950 ;
        RECT 130.950 148.950 133.050 151.050 ;
        RECT 131.400 138.600 132.450 148.950 ;
        RECT 136.950 142.950 139.050 145.050 ;
        RECT 131.400 136.350 132.600 138.600 ;
        RECT 137.400 136.050 138.450 142.950 ;
        RECT 143.400 139.200 144.450 196.950 ;
        RECT 146.400 177.900 147.450 214.950 ;
        RECT 158.400 214.350 159.600 215.100 ;
        RECT 154.950 211.950 157.050 214.050 ;
        RECT 157.950 211.950 160.050 214.050 ;
        RECT 155.400 210.900 156.600 211.650 ;
        RECT 154.950 208.800 157.050 210.900 ;
        RECT 163.950 208.950 166.050 211.050 ;
        RECT 148.950 187.950 151.050 190.050 ;
        RECT 160.950 187.950 163.050 190.050 ;
        RECT 149.400 184.050 150.450 187.950 ;
        RECT 148.950 181.950 151.050 184.050 ;
        RECT 154.950 182.100 157.050 184.200 ;
        RECT 161.400 184.050 162.450 187.950 ;
        RECT 155.400 181.350 156.600 182.100 ;
        RECT 160.950 181.950 163.050 184.050 ;
        RECT 151.950 178.950 154.050 181.050 ;
        RECT 154.950 178.950 157.050 181.050 ;
        RECT 157.950 178.950 160.050 181.050 ;
        RECT 145.950 175.800 148.050 177.900 ;
        RECT 152.400 176.400 153.600 178.650 ;
        RECT 158.400 177.900 159.600 178.650 ;
        RECT 152.400 169.050 153.450 176.400 ;
        RECT 157.950 175.800 160.050 177.900 ;
        RECT 151.950 166.950 154.050 169.050 ;
        RECT 145.950 142.950 148.050 145.050 ;
        RECT 142.950 137.100 145.050 139.200 ;
        RECT 146.400 138.600 147.450 142.950 ;
        RECT 146.400 136.350 147.600 138.600 ;
        RECT 151.950 137.100 154.050 142.050 ;
        RECT 160.950 139.950 163.050 142.050 ;
        RECT 152.400 136.350 153.600 137.100 ;
        RECT 127.950 133.950 130.050 136.050 ;
        RECT 130.950 133.950 133.050 136.050 ;
        RECT 136.950 133.950 139.050 136.050 ;
        RECT 145.950 133.950 148.050 136.050 ;
        RECT 148.950 133.950 151.050 136.050 ;
        RECT 151.950 133.950 154.050 136.050 ;
        RECT 154.950 133.950 157.050 136.050 ;
        RECT 128.400 132.900 129.600 133.650 ;
        RECT 127.950 130.800 130.050 132.900 ;
        RECT 149.400 131.400 150.600 133.650 ;
        RECT 155.400 132.900 156.600 133.650 ;
        RECT 149.400 124.050 150.450 131.400 ;
        RECT 154.950 130.800 157.050 132.900 ;
        RECT 161.400 130.050 162.450 139.950 ;
        RECT 164.400 139.200 165.450 208.950 ;
        RECT 167.400 190.050 168.450 250.950 ;
        RECT 175.950 244.950 178.050 247.050 ;
        RECT 176.400 217.200 177.450 244.950 ;
        RECT 175.950 215.100 178.050 217.200 ;
        RECT 200.400 216.600 201.450 259.950 ;
        RECT 203.400 219.450 204.450 268.950 ;
        RECT 209.400 261.600 210.450 268.950 ;
        RECT 215.400 261.600 216.450 277.950 ;
        RECT 209.400 259.350 210.600 261.600 ;
        RECT 215.400 259.350 216.600 261.600 ;
        RECT 208.950 256.950 211.050 259.050 ;
        RECT 211.950 256.950 214.050 259.050 ;
        RECT 214.950 256.950 217.050 259.050 ;
        RECT 217.950 256.950 220.050 259.050 ;
        RECT 212.400 255.900 213.600 256.650 ;
        RECT 211.950 253.800 214.050 255.900 ;
        RECT 218.400 254.400 219.600 256.650 ;
        RECT 224.400 256.050 225.450 286.800 ;
        RECT 227.400 265.050 228.450 332.400 ;
        RECT 238.950 331.800 241.050 333.900 ;
        RECT 245.400 328.050 246.450 337.950 ;
        RECT 257.400 337.350 258.600 339.600 ;
        RECT 253.950 334.950 256.050 337.050 ;
        RECT 256.950 334.950 259.050 337.050 ;
        RECT 259.950 334.950 262.050 337.050 ;
        RECT 250.950 333.450 253.050 333.900 ;
        RECT 254.400 333.450 255.600 334.650 ;
        RECT 250.950 332.400 255.600 333.450 ;
        RECT 260.400 332.400 261.600 334.650 ;
        RECT 250.950 331.800 253.050 332.400 ;
        RECT 244.950 325.950 247.050 328.050 ;
        RECT 229.950 293.100 232.050 295.200 ;
        RECT 239.400 294.450 240.600 294.600 ;
        RECT 233.400 293.400 240.600 294.450 ;
        RECT 230.400 280.050 231.450 293.100 ;
        RECT 233.400 286.050 234.450 293.400 ;
        RECT 239.400 292.350 240.600 293.400 ;
        RECT 244.950 293.100 247.050 295.200 ;
        RECT 245.400 292.350 246.600 293.100 ;
        RECT 238.950 289.950 241.050 292.050 ;
        RECT 241.950 289.950 244.050 292.050 ;
        RECT 244.950 289.950 247.050 292.050 ;
        RECT 242.400 288.900 243.600 289.650 ;
        RECT 251.400 289.050 252.450 331.800 ;
        RECT 260.400 328.050 261.450 332.400 ;
        RECT 259.950 325.950 262.050 328.050 ;
        RECT 269.400 304.050 270.450 397.950 ;
        RECT 299.250 379.500 301.350 380.400 ;
        RECT 297.150 378.300 301.350 379.500 ;
        RECT 311.400 379.050 312.450 406.950 ;
        RECT 315.150 404.700 316.350 423.300 ;
        RECT 320.100 412.950 322.200 415.050 ;
        RECT 320.400 411.450 321.600 412.650 ;
        RECT 320.400 410.400 324.450 411.450 ;
        RECT 323.400 406.050 324.450 410.400 ;
        RECT 315.150 403.500 319.350 404.700 ;
        RECT 322.950 403.950 325.050 406.050 ;
        RECT 317.250 402.600 319.350 403.500 ;
        RECT 326.400 400.050 327.450 449.100 ;
        RECT 335.400 448.350 336.600 449.100 ;
        RECT 341.400 448.350 342.600 450.600 ;
        RECT 346.950 449.100 349.050 451.200 ;
        RECT 347.400 448.350 348.600 449.100 ;
        RECT 328.950 445.950 331.050 448.050 ;
        RECT 334.950 445.950 337.050 448.050 ;
        RECT 337.950 445.950 340.050 448.050 ;
        RECT 340.950 445.950 343.050 448.050 ;
        RECT 343.950 445.950 346.050 448.050 ;
        RECT 346.950 445.950 349.050 448.050 ;
        RECT 329.400 424.050 330.450 445.950 ;
        RECT 338.400 443.400 339.600 445.650 ;
        RECT 344.400 443.400 345.600 445.650 ;
        RECT 338.400 436.050 339.450 443.400 ;
        RECT 337.950 433.950 340.050 436.050 ;
        RECT 328.950 421.950 331.050 424.050 ;
        RECT 332.550 423.300 334.650 425.400 ;
        RECT 328.950 416.100 331.050 418.200 ;
        RECT 325.950 397.950 328.050 400.050 ;
        RECT 314.550 381.300 316.650 383.400 ;
        RECT 283.950 372.450 286.050 373.200 ;
        RECT 283.950 371.400 288.450 372.450 ;
        RECT 283.950 371.100 286.050 371.400 ;
        RECT 284.400 370.350 285.600 371.100 ;
        RECT 283.800 367.950 285.900 370.050 ;
        RECT 287.400 346.050 288.450 371.400 ;
        RECT 292.950 371.100 295.050 373.200 ;
        RECT 293.400 370.350 294.600 371.100 ;
        RECT 292.950 367.950 295.050 370.050 ;
        RECT 297.150 359.700 298.350 378.300 ;
        RECT 310.950 376.950 313.050 379.050 ;
        RECT 314.550 374.700 315.750 381.300 ;
        RECT 301.950 371.100 304.050 373.200 ;
        RECT 314.550 372.600 316.650 374.700 ;
        RECT 302.400 370.350 303.600 371.100 ;
        RECT 302.100 367.950 304.200 370.050 ;
        RECT 314.550 359.700 315.750 372.600 ;
        RECT 319.950 367.950 322.050 370.050 ;
        RECT 320.400 366.900 321.600 367.650 ;
        RECT 319.950 364.800 322.050 366.900 ;
        RECT 296.850 357.600 298.950 359.700 ;
        RECT 314.550 357.600 316.650 359.700 ;
        RECT 319.950 352.950 322.050 355.050 ;
        RECT 286.950 343.950 289.050 346.050 ;
        RECT 295.950 343.950 298.050 346.050 ;
        RECT 280.950 338.100 283.050 340.200 ;
        RECT 286.950 338.100 289.050 340.200 ;
        RECT 292.950 338.100 295.050 340.200 ;
        RECT 281.400 337.350 282.600 338.100 ;
        RECT 287.400 337.350 288.600 338.100 ;
        RECT 277.950 334.950 280.050 337.050 ;
        RECT 280.950 334.950 283.050 337.050 ;
        RECT 283.950 334.950 286.050 337.050 ;
        RECT 286.950 334.950 289.050 337.050 ;
        RECT 278.400 332.400 279.600 334.650 ;
        RECT 284.400 332.400 285.600 334.650 ;
        RECT 274.950 325.950 277.050 328.050 ;
        RECT 268.950 301.950 271.050 304.050 ;
        RECT 269.400 297.450 270.450 301.950 ;
        RECT 266.400 296.400 270.450 297.450 ;
        RECT 253.950 293.100 256.050 295.200 ;
        RECT 259.950 293.100 262.050 295.200 ;
        RECT 266.400 294.600 267.450 296.400 ;
        RECT 275.400 294.600 276.450 325.950 ;
        RECT 278.400 319.050 279.450 332.400 ;
        RECT 277.950 316.950 280.050 319.050 ;
        RECT 284.400 313.050 285.450 332.400 ;
        RECT 293.400 325.050 294.450 338.100 ;
        RECT 296.400 328.050 297.450 343.950 ;
        RECT 304.950 338.100 307.050 340.200 ;
        RECT 305.400 337.350 306.600 338.100 ;
        RECT 313.950 337.950 316.050 340.050 ;
        RECT 301.950 334.950 304.050 337.050 ;
        RECT 304.950 334.950 307.050 337.050 ;
        RECT 307.950 334.950 310.050 337.050 ;
        RECT 302.400 333.000 303.600 334.650 ;
        RECT 308.400 333.900 309.600 334.650 ;
        RECT 314.400 333.900 315.450 337.950 ;
        RECT 301.950 328.950 304.050 333.000 ;
        RECT 307.950 331.800 310.050 333.900 ;
        RECT 313.950 331.800 316.050 333.900 ;
        RECT 295.950 325.950 298.050 328.050 ;
        RECT 307.950 325.950 310.050 328.050 ;
        RECT 292.950 322.950 295.050 325.050 ;
        RECT 289.950 313.950 292.050 316.050 ;
        RECT 283.950 310.950 286.050 313.050 ;
        RECT 284.400 307.050 285.450 310.950 ;
        RECT 283.950 304.950 286.050 307.050 ;
        RECT 281.250 301.500 283.350 302.400 ;
        RECT 279.150 300.300 283.350 301.500 ;
        RECT 241.950 286.800 244.050 288.900 ;
        RECT 250.950 286.950 253.050 289.050 ;
        RECT 232.950 283.950 235.050 286.050 ;
        RECT 254.400 283.050 255.450 293.100 ;
        RECT 260.400 292.350 261.600 293.100 ;
        RECT 266.400 292.350 267.600 294.600 ;
        RECT 275.400 292.350 276.600 294.600 ;
        RECT 259.950 289.950 262.050 292.050 ;
        RECT 262.950 289.950 265.050 292.050 ;
        RECT 265.950 289.950 268.050 292.050 ;
        RECT 268.950 289.950 271.050 292.050 ;
        RECT 274.950 289.950 277.050 292.050 ;
        RECT 263.400 288.900 264.600 289.650 ;
        RECT 262.950 286.800 265.050 288.900 ;
        RECT 269.400 287.400 270.600 289.650 ;
        RECT 253.950 280.950 256.050 283.050 ;
        RECT 229.950 277.950 232.050 280.050 ;
        RECT 262.950 277.950 265.050 280.050 ;
        RECT 226.950 262.950 229.050 265.050 ;
        RECT 235.950 260.100 238.050 262.200 ;
        RECT 241.950 260.100 244.050 262.200 ;
        RECT 250.950 261.000 253.050 265.050 ;
        RECT 236.400 259.350 237.600 260.100 ;
        RECT 232.950 256.950 235.050 259.050 ;
        RECT 235.950 256.950 238.050 259.050 ;
        RECT 218.400 253.050 219.450 254.400 ;
        RECT 223.950 253.950 226.050 256.050 ;
        RECT 233.400 255.900 234.600 256.650 ;
        RECT 232.950 253.800 235.050 255.900 ;
        RECT 242.400 253.050 243.450 260.100 ;
        RECT 251.400 259.350 252.600 261.000 ;
        RECT 250.950 256.950 253.050 259.050 ;
        RECT 253.950 256.950 256.050 259.050 ;
        RECT 254.400 254.400 255.600 256.650 ;
        RECT 263.400 255.900 264.450 277.950 ;
        RECT 269.400 274.050 270.450 287.400 ;
        RECT 279.150 281.700 280.350 300.300 ;
        RECT 283.950 293.100 286.050 295.200 ;
        RECT 284.400 292.350 285.600 293.100 ;
        RECT 284.100 289.950 286.200 292.050 ;
        RECT 278.850 279.600 280.950 281.700 ;
        RECT 290.400 280.050 291.450 313.950 ;
        RECT 293.400 298.050 294.450 322.950 ;
        RECT 296.550 303.300 298.650 305.400 ;
        RECT 292.950 295.950 295.050 298.050 ;
        RECT 296.550 296.700 297.750 303.300 ;
        RECT 289.950 277.950 292.050 280.050 ;
        RECT 280.950 274.950 283.050 277.050 ;
        RECT 268.950 271.950 271.050 274.050 ;
        RECT 271.950 260.100 274.050 262.200 ;
        RECT 272.400 259.350 273.600 260.100 ;
        RECT 268.950 256.950 271.050 259.050 ;
        RECT 271.950 256.950 274.050 259.050 ;
        RECT 274.950 256.950 277.050 259.050 ;
        RECT 217.950 250.950 220.050 253.050 ;
        RECT 241.950 250.950 244.050 253.050 ;
        RECT 203.400 218.400 207.450 219.450 ;
        RECT 206.400 216.600 207.450 218.400 ;
        RECT 176.400 214.350 177.600 215.100 ;
        RECT 200.400 214.350 201.600 216.600 ;
        RECT 206.400 214.350 207.600 216.600 ;
        RECT 175.950 211.950 178.050 214.050 ;
        RECT 178.950 211.950 181.050 214.050 ;
        RECT 181.950 211.950 184.050 214.050 ;
        RECT 199.950 211.950 202.050 214.050 ;
        RECT 202.950 211.950 205.050 214.050 ;
        RECT 205.950 211.950 208.050 214.050 ;
        RECT 208.950 211.950 211.050 214.050 ;
        RECT 179.400 210.900 180.600 211.650 ;
        RECT 178.950 208.800 181.050 210.900 ;
        RECT 203.400 209.400 204.600 211.650 ;
        RECT 209.400 210.900 210.600 211.650 ;
        RECT 218.400 211.050 219.450 250.950 ;
        RECT 229.950 226.950 232.050 229.050 ;
        RECT 230.400 216.600 231.450 226.950 ;
        RECT 254.400 220.050 255.450 254.400 ;
        RECT 262.950 253.800 265.050 255.900 ;
        RECT 269.400 254.400 270.600 256.650 ;
        RECT 275.400 255.900 276.600 256.650 ;
        RECT 262.950 244.950 265.050 247.050 ;
        RECT 259.950 232.950 262.050 235.050 ;
        RECT 230.400 214.350 231.600 216.600 ;
        RECT 244.950 216.000 247.050 220.050 ;
        RECT 253.950 217.950 256.050 220.050 ;
        RECT 245.400 214.350 246.600 216.000 ;
        RECT 250.950 215.100 253.050 217.200 ;
        RECT 251.400 214.350 252.600 215.100 ;
        RECT 223.950 211.950 226.050 214.050 ;
        RECT 226.950 211.950 229.050 214.050 ;
        RECT 229.950 211.950 232.050 214.050 ;
        RECT 244.950 211.950 247.050 214.050 ;
        RECT 247.950 211.950 250.050 214.050 ;
        RECT 250.950 211.950 253.050 214.050 ;
        RECT 253.950 211.950 256.050 214.050 ;
        RECT 203.400 193.050 204.450 209.400 ;
        RECT 208.950 208.800 211.050 210.900 ;
        RECT 217.950 208.950 220.050 211.050 ;
        RECT 227.400 210.900 228.600 211.650 ;
        RECT 248.400 210.900 249.600 211.650 ;
        RECT 226.950 208.800 229.050 210.900 ;
        RECT 238.950 208.800 241.050 210.900 ;
        RECT 247.950 208.800 250.050 210.900 ;
        RECT 254.400 209.400 255.600 211.650 ;
        RECT 226.950 196.950 229.050 199.050 ;
        RECT 172.950 190.950 175.050 193.050 ;
        RECT 187.950 190.950 190.050 193.050 ;
        RECT 202.950 190.950 205.050 193.050 ;
        RECT 166.950 187.950 169.050 190.050 ;
        RECT 169.950 184.050 172.050 184.200 ;
        RECT 166.950 182.100 172.050 184.050 ;
        RECT 173.400 183.600 174.450 190.950 ;
        RECT 166.950 181.950 171.000 182.100 ;
        RECT 173.400 181.350 174.600 183.600 ;
        RECT 172.950 178.950 175.050 181.050 ;
        RECT 175.950 178.950 178.050 181.050 ;
        RECT 184.950 178.950 187.050 181.050 ;
        RECT 176.400 177.900 177.600 178.650 ;
        RECT 175.950 175.800 178.050 177.900 ;
        RECT 172.950 148.950 175.050 151.050 ;
        RECT 163.950 137.100 166.050 139.200 ;
        RECT 173.400 138.600 174.450 148.950 ;
        RECT 185.400 142.050 186.450 178.950 ;
        RECT 184.950 139.950 187.050 142.050 ;
        RECT 188.400 139.200 189.450 190.950 ;
        RECT 196.950 182.100 199.050 184.200 ;
        RECT 204.000 183.600 208.050 184.050 ;
        RECT 197.400 181.350 198.600 182.100 ;
        RECT 203.400 181.950 208.050 183.600 ;
        RECT 208.950 181.950 211.050 184.050 ;
        RECT 211.950 181.950 214.050 184.050 ;
        RECT 220.950 182.100 223.050 184.200 ;
        RECT 227.400 183.600 228.450 196.950 ;
        RECT 239.400 187.050 240.450 208.800 ;
        RECT 254.400 205.050 255.450 209.400 ;
        RECT 260.400 205.050 261.450 232.950 ;
        RECT 253.950 204.450 256.050 205.050 ;
        RECT 253.950 203.400 258.450 204.450 ;
        RECT 253.950 202.950 256.050 203.400 ;
        RECT 253.950 196.950 256.050 199.050 ;
        RECT 254.400 193.050 255.450 196.950 ;
        RECT 253.950 190.950 256.050 193.050 ;
        RECT 238.950 184.950 241.050 187.050 ;
        RECT 203.400 181.350 204.600 181.950 ;
        RECT 193.950 178.950 196.050 181.050 ;
        RECT 196.950 178.950 199.050 181.050 ;
        RECT 199.950 178.950 202.050 181.050 ;
        RECT 202.950 178.950 205.050 181.050 ;
        RECT 194.400 177.900 195.600 178.650 ;
        RECT 193.950 175.800 196.050 177.900 ;
        RECT 200.400 177.000 201.600 178.650 ;
        RECT 199.950 172.950 202.050 177.000 ;
        RECT 209.400 175.050 210.450 181.950 ;
        RECT 208.950 172.950 211.050 175.050 ;
        RECT 212.400 166.050 213.450 181.950 ;
        RECT 221.400 181.350 222.600 182.100 ;
        RECT 227.400 181.350 228.600 183.600 ;
        RECT 217.950 178.950 220.050 181.050 ;
        RECT 220.950 178.950 223.050 181.050 ;
        RECT 223.950 178.950 226.050 181.050 ;
        RECT 226.950 178.950 229.050 181.050 ;
        RECT 218.400 176.400 219.600 178.650 ;
        RECT 224.400 177.900 225.600 178.650 ;
        RECT 218.400 169.050 219.450 176.400 ;
        RECT 223.950 175.800 226.050 177.900 ;
        RECT 217.950 166.950 220.050 169.050 ;
        RECT 211.950 163.950 214.050 166.050 ;
        RECT 193.950 145.950 196.050 148.050 ;
        RECT 226.950 145.950 229.050 148.050 ;
        RECT 194.400 142.050 195.450 145.950 ;
        RECT 220.950 142.050 223.050 142.200 ;
        RECT 164.400 132.900 165.450 137.100 ;
        RECT 173.400 136.350 174.600 138.600 ;
        RECT 178.950 137.100 181.050 139.200 ;
        RECT 187.950 137.100 190.050 139.200 ;
        RECT 193.950 138.000 196.050 142.050 ;
        RECT 214.950 139.950 217.050 142.050 ;
        RECT 220.950 140.100 226.050 142.050 ;
        RECT 222.000 139.950 226.050 140.100 ;
        RECT 179.400 136.350 180.600 137.100 ;
        RECT 194.400 136.350 195.600 138.000 ;
        RECT 199.950 137.100 202.050 139.200 ;
        RECT 200.400 136.350 201.600 137.100 ;
        RECT 169.950 133.950 172.050 136.050 ;
        RECT 172.950 133.950 175.050 136.050 ;
        RECT 175.950 133.950 178.050 136.050 ;
        RECT 178.950 133.950 181.050 136.050 ;
        RECT 193.950 133.950 196.050 136.050 ;
        RECT 196.950 133.950 199.050 136.050 ;
        RECT 199.950 133.950 202.050 136.050 ;
        RECT 202.950 133.950 205.050 136.050 ;
        RECT 163.950 130.800 166.050 132.900 ;
        RECT 170.400 132.000 171.600 133.650 ;
        RECT 176.400 132.900 177.600 133.650 ;
        RECT 197.400 132.900 198.600 133.650 ;
        RECT 203.400 132.900 204.600 133.650 ;
        RECT 215.400 133.050 216.450 139.950 ;
        RECT 220.950 136.950 223.050 139.050 ;
        RECT 227.400 138.600 228.450 145.950 ;
        RECT 221.400 136.350 222.600 136.950 ;
        RECT 227.400 136.350 228.600 138.600 ;
        RECT 220.950 133.950 223.050 136.050 ;
        RECT 223.950 133.950 226.050 136.050 ;
        RECT 226.950 133.950 229.050 136.050 ;
        RECT 229.950 133.950 232.050 136.050 ;
        RECT 160.950 127.950 163.050 130.050 ;
        RECT 169.950 127.950 172.050 132.000 ;
        RECT 175.950 130.800 178.050 132.900 ;
        RECT 196.950 127.950 199.050 132.900 ;
        RECT 202.950 130.800 205.050 132.900 ;
        RECT 214.950 130.950 217.050 133.050 ;
        RECT 224.400 132.000 225.600 133.650 ;
        RECT 230.400 132.000 231.600 133.650 ;
        RECT 239.400 133.050 240.450 184.950 ;
        RECT 244.950 178.950 247.050 181.050 ;
        RECT 247.950 178.950 250.050 181.050 ;
        RECT 245.400 177.900 246.600 178.650 ;
        RECT 244.950 175.800 247.050 177.900 ;
        RECT 247.950 163.950 250.050 166.050 ;
        RECT 248.400 138.600 249.450 163.950 ;
        RECT 250.950 139.950 253.050 145.050 ;
        RECT 253.950 142.950 256.050 145.050 ;
        RECT 254.400 138.600 255.450 142.950 ;
        RECT 248.400 136.350 249.600 138.600 ;
        RECT 254.400 136.350 255.600 138.600 ;
        RECT 257.400 138.450 258.450 203.400 ;
        RECT 259.950 202.950 262.050 205.050 ;
        RECT 263.400 202.050 264.450 244.950 ;
        RECT 269.400 235.050 270.450 254.400 ;
        RECT 274.950 253.800 277.050 255.900 ;
        RECT 281.400 244.050 282.450 274.950 ;
        RECT 293.400 271.050 294.450 295.950 ;
        RECT 296.550 294.600 298.650 296.700 ;
        RECT 296.550 281.700 297.750 294.600 ;
        RECT 301.950 289.950 304.050 292.050 ;
        RECT 302.400 287.400 303.600 289.650 ;
        RECT 296.550 279.600 298.650 281.700 ;
        RECT 302.400 277.050 303.450 287.400 ;
        RECT 301.950 274.950 304.050 277.050 ;
        RECT 286.950 268.950 289.050 271.050 ;
        RECT 292.950 268.950 295.050 271.050 ;
        RECT 283.950 260.100 286.050 262.200 ;
        RECT 284.400 252.450 285.450 260.100 ;
        RECT 287.400 255.450 288.450 268.950 ;
        RECT 308.400 265.050 309.450 325.950 ;
        RECT 320.400 325.050 321.450 352.950 ;
        RECT 329.400 352.050 330.450 416.100 ;
        RECT 332.550 410.400 333.750 423.300 ;
        RECT 344.400 421.050 345.450 443.400 ;
        RECT 356.400 442.050 357.450 463.950 ;
        RECT 374.400 463.050 375.450 541.950 ;
        RECT 373.950 460.950 376.050 463.050 ;
        RECT 367.950 454.950 370.050 457.050 ;
        RECT 361.950 449.100 364.050 451.200 ;
        RECT 368.400 450.600 369.450 454.950 ;
        RECT 362.400 448.350 363.600 449.100 ;
        RECT 368.400 448.350 369.600 450.600 ;
        RECT 373.950 450.000 376.050 454.050 ;
        RECT 377.400 450.450 378.450 553.950 ;
        RECT 413.400 547.050 414.450 562.950 ;
        RECT 412.950 544.950 415.050 547.050 ;
        RECT 382.950 527.100 385.050 529.200 ;
        RECT 388.950 527.100 391.050 529.200 ;
        RECT 383.400 526.350 384.600 527.100 ;
        RECT 389.400 526.350 390.600 527.100 ;
        RECT 397.950 526.950 400.050 529.050 ;
        RECT 403.950 527.100 406.050 529.200 ;
        RECT 382.950 523.950 385.050 526.050 ;
        RECT 385.950 523.950 388.050 526.050 ;
        RECT 388.950 523.950 391.050 526.050 ;
        RECT 394.950 523.950 397.050 526.050 ;
        RECT 386.400 521.400 387.600 523.650 ;
        RECT 379.950 502.950 382.050 505.050 ;
        RECT 380.400 454.050 381.450 502.950 ;
        RECT 386.400 499.050 387.450 521.400 ;
        RECT 395.400 517.050 396.450 523.950 ;
        RECT 394.950 514.950 397.050 517.050 ;
        RECT 388.950 502.950 391.050 505.050 ;
        RECT 385.950 496.950 388.050 499.050 ;
        RECT 389.400 495.600 390.450 502.950 ;
        RECT 395.400 495.600 396.450 514.950 ;
        RECT 398.400 514.050 399.450 526.950 ;
        RECT 404.400 526.350 405.600 527.100 ;
        RECT 403.950 523.950 406.050 526.050 ;
        RECT 406.950 523.950 409.050 526.050 ;
        RECT 407.400 522.450 408.600 523.650 ;
        RECT 407.400 521.400 411.450 522.450 ;
        RECT 406.950 517.950 409.050 520.050 ;
        RECT 397.950 511.950 400.050 514.050 ;
        RECT 389.400 493.350 390.600 495.600 ;
        RECT 395.400 493.350 396.600 495.600 ;
        RECT 385.950 490.950 388.050 493.050 ;
        RECT 388.950 490.950 391.050 493.050 ;
        RECT 391.950 490.950 394.050 493.050 ;
        RECT 394.950 490.950 397.050 493.050 ;
        RECT 386.400 489.900 387.600 490.650 ;
        RECT 385.950 487.800 388.050 489.900 ;
        RECT 392.400 489.000 393.600 490.650 ;
        RECT 407.400 489.450 408.450 517.950 ;
        RECT 410.400 505.050 411.450 521.400 ;
        RECT 413.400 520.050 414.450 544.950 ;
        RECT 416.400 535.050 417.450 580.950 ;
        RECT 418.950 571.950 421.050 574.050 ;
        RECT 415.950 532.950 418.050 535.050 ;
        RECT 416.400 523.050 417.450 532.950 ;
        RECT 419.400 529.050 420.450 571.950 ;
        RECT 422.400 550.050 423.450 592.950 ;
        RECT 428.400 586.050 429.450 599.400 ;
        RECT 436.950 598.950 439.050 601.050 ;
        RECT 452.400 600.900 453.600 601.650 ;
        RECT 451.950 598.800 454.050 600.900 ;
        RECT 427.950 583.950 430.050 586.050 ;
        RECT 451.950 583.950 454.050 586.050 ;
        RECT 445.350 579.300 447.450 581.400 ;
        RECT 430.950 572.100 433.050 574.200 ;
        RECT 439.950 572.100 442.050 574.200 ;
        RECT 431.400 571.350 432.600 572.100 ;
        RECT 440.400 571.350 441.600 572.100 ;
        RECT 427.950 568.950 430.050 571.050 ;
        RECT 430.950 568.950 433.050 571.050 ;
        RECT 433.950 568.950 436.050 571.050 ;
        RECT 439.950 568.950 442.050 571.050 ;
        RECT 428.400 566.400 429.600 568.650 ;
        RECT 434.400 566.400 435.600 568.650 ;
        RECT 421.950 547.950 424.050 550.050 ;
        RECT 428.400 535.050 429.450 566.400 ;
        RECT 434.400 559.050 435.450 566.400 ;
        RECT 436.950 565.950 439.050 568.050 ;
        RECT 446.250 566.400 447.450 579.300 ;
        RECT 448.950 572.100 451.050 574.200 ;
        RECT 433.950 556.950 436.050 559.050 ;
        RECT 433.950 538.950 436.050 541.050 ;
        RECT 434.400 535.050 435.450 538.950 ;
        RECT 427.950 532.950 430.050 535.050 ;
        RECT 433.950 532.950 436.050 535.050 ;
        RECT 437.400 532.050 438.450 565.950 ;
        RECT 445.350 564.300 447.450 566.400 ;
        RECT 446.250 557.700 447.450 564.300 ;
        RECT 449.400 559.050 450.450 572.100 ;
        RECT 452.400 567.900 453.450 583.950 ;
        RECT 463.050 579.300 465.150 581.400 ;
        RECT 457.800 568.950 459.900 571.050 ;
        RECT 458.400 567.900 459.600 568.650 ;
        RECT 451.950 565.800 454.050 567.900 ;
        RECT 457.950 565.800 460.050 567.900 ;
        RECT 463.650 560.700 464.850 579.300 ;
        RECT 467.400 577.050 468.450 631.950 ;
        RECT 470.400 631.050 471.450 638.400 ;
        RECT 469.950 628.950 472.050 631.050 ;
        RECT 479.400 628.050 480.450 718.950 ;
        RECT 488.400 718.050 489.450 722.400 ;
        RECT 487.950 715.950 490.050 718.050 ;
        RECT 491.400 691.050 492.450 760.950 ;
        RECT 493.950 745.950 496.050 748.050 ;
        RECT 494.400 718.050 495.450 745.950 ;
        RECT 497.400 723.900 498.450 769.950 ;
        RECT 503.400 763.200 504.450 793.950 ;
        RECT 524.400 790.050 525.450 811.950 ;
        RECT 526.950 808.950 529.050 811.050 ;
        RECT 523.950 787.950 526.050 790.050 ;
        RECT 514.950 775.950 517.050 778.050 ;
        RECT 508.950 769.950 511.050 772.050 ;
        RECT 502.950 761.100 505.050 763.200 ;
        RECT 509.400 762.600 510.450 769.950 ;
        RECT 503.400 760.350 504.600 761.100 ;
        RECT 509.400 760.350 510.600 762.600 ;
        RECT 502.950 757.950 505.050 760.050 ;
        RECT 505.950 757.950 508.050 760.050 ;
        RECT 508.950 757.950 511.050 760.050 ;
        RECT 506.400 755.400 507.600 757.650 ;
        RECT 506.400 729.600 507.450 755.400 ;
        RECT 515.400 742.050 516.450 775.950 ;
        RECT 523.950 769.950 526.050 775.050 ;
        RECT 527.400 772.050 528.450 808.950 ;
        RECT 530.400 808.050 531.450 817.950 ;
        RECT 532.950 811.950 535.050 814.050 ;
        RECT 529.950 805.950 532.050 808.050 ;
        RECT 533.400 807.600 534.450 811.950 ;
        RECT 539.400 807.600 540.450 839.100 ;
        RECT 542.400 811.050 543.450 865.950 ;
        RECT 560.400 850.050 561.450 940.950 ;
        RECT 562.950 937.950 565.050 940.050 ;
        RECT 563.400 934.050 564.450 937.950 ;
        RECT 562.950 931.950 565.050 934.050 ;
        RECT 569.400 928.050 570.450 956.400 ;
        RECT 571.950 955.800 574.050 957.900 ;
        RECT 586.950 955.800 589.050 957.900 ;
        RECT 593.400 957.000 594.600 958.650 ;
        RECT 599.400 957.900 600.600 958.650 ;
        RECT 572.400 955.050 573.450 955.800 ;
        RECT 572.400 953.400 577.050 955.050 ;
        RECT 573.000 952.950 577.050 953.400 ;
        RECT 592.950 952.950 595.050 957.000 ;
        RECT 598.950 955.800 601.050 957.900 ;
        RECT 608.400 943.050 609.450 961.950 ;
        RECT 617.400 961.350 618.600 962.100 ;
        RECT 623.400 961.350 624.600 963.600 ;
        RECT 643.950 962.100 646.050 964.200 ;
        RECT 665.400 963.600 666.450 967.950 ;
        RECT 644.400 961.350 645.600 962.100 ;
        RECT 665.400 961.350 666.600 963.600 ;
        RECT 670.950 963.000 673.050 967.050 ;
        RECT 671.400 961.350 672.600 963.000 ;
        RECT 676.950 961.950 679.050 964.050 ;
        RECT 685.950 962.100 688.050 964.200 ;
        RECT 691.950 963.000 694.050 967.050 ;
        RECT 711.000 966.450 715.050 967.050 ;
        RECT 710.400 964.950 715.050 966.450 ;
        RECT 718.950 964.950 721.050 967.050 ;
        RECT 730.950 964.950 733.050 968.400 ;
        RECT 736.950 967.950 739.050 968.400 ;
        RECT 710.400 963.600 711.450 964.950 ;
        RECT 616.950 958.950 619.050 961.050 ;
        RECT 619.950 958.950 622.050 961.050 ;
        RECT 622.950 958.950 625.050 961.050 ;
        RECT 625.950 958.950 628.050 961.050 ;
        RECT 640.950 958.950 643.050 961.050 ;
        RECT 643.950 958.950 646.050 961.050 ;
        RECT 646.950 958.950 649.050 961.050 ;
        RECT 661.950 958.950 664.050 961.050 ;
        RECT 664.950 958.950 667.050 961.050 ;
        RECT 667.950 958.950 670.050 961.050 ;
        RECT 670.950 958.950 673.050 961.050 ;
        RECT 620.400 957.900 621.600 958.650 ;
        RECT 619.950 955.800 622.050 957.900 ;
        RECT 626.400 956.400 627.600 958.650 ;
        RECT 641.400 956.400 642.600 958.650 ;
        RECT 647.400 957.900 648.600 958.650 ;
        RECT 662.400 957.900 663.600 958.650 ;
        RECT 668.400 957.900 669.600 958.650 ;
        RECT 677.400 957.900 678.450 961.950 ;
        RECT 686.400 961.350 687.600 962.100 ;
        RECT 692.400 961.350 693.600 963.000 ;
        RECT 710.400 961.350 711.600 963.600 ;
        RECT 685.950 958.950 688.050 961.050 ;
        RECT 688.950 958.950 691.050 961.050 ;
        RECT 691.950 958.950 694.050 961.050 ;
        RECT 706.950 958.950 709.050 961.050 ;
        RECT 709.950 958.950 712.050 961.050 ;
        RECT 712.950 958.950 715.050 961.050 ;
        RECT 626.400 946.050 627.450 956.400 ;
        RECT 628.950 952.950 631.050 955.050 ;
        RECT 625.950 943.950 628.050 946.050 ;
        RECT 607.950 940.950 610.050 943.050 ;
        RECT 607.950 934.950 610.050 937.050 ;
        RECT 562.950 925.950 565.050 928.050 ;
        RECT 568.950 925.950 571.050 928.050 ;
        RECT 563.400 916.050 564.450 925.950 ;
        RECT 565.950 918.600 570.000 919.050 ;
        RECT 565.950 916.950 570.600 918.600 ;
        RECT 574.950 917.100 577.050 919.200 ;
        RECT 580.950 917.100 583.050 919.200 ;
        RECT 592.950 917.100 595.050 919.200 ;
        RECT 598.950 917.100 601.050 919.200 ;
        RECT 604.950 917.100 607.050 919.200 ;
        RECT 569.400 916.350 570.600 916.950 ;
        RECT 575.400 916.350 576.600 917.100 ;
        RECT 562.950 913.950 565.050 916.050 ;
        RECT 568.950 913.950 571.050 916.050 ;
        RECT 571.950 913.950 574.050 916.050 ;
        RECT 574.950 913.950 577.050 916.050 ;
        RECT 572.400 912.900 573.600 913.650 ;
        RECT 581.400 913.050 582.450 917.100 ;
        RECT 593.400 916.350 594.600 917.100 ;
        RECT 599.400 916.350 600.600 917.100 ;
        RECT 589.950 913.950 592.050 916.050 ;
        RECT 592.950 913.950 595.050 916.050 ;
        RECT 595.950 913.950 598.050 916.050 ;
        RECT 598.950 913.950 601.050 916.050 ;
        RECT 571.950 910.800 574.050 912.900 ;
        RECT 580.950 910.950 583.050 913.050 ;
        RECT 590.400 912.900 591.600 913.650 ;
        RECT 589.950 910.800 592.050 912.900 ;
        RECT 596.400 911.400 597.600 913.650 ;
        RECT 596.400 907.050 597.450 911.400 ;
        RECT 598.950 907.950 601.050 910.050 ;
        RECT 595.950 904.950 598.050 907.050 ;
        RECT 586.950 898.950 589.050 901.050 ;
        RECT 571.950 892.950 574.050 895.050 ;
        RECT 572.400 885.600 573.450 892.950 ;
        RECT 580.950 889.950 583.050 895.050 ;
        RECT 583.950 889.950 586.050 892.050 ;
        RECT 572.400 883.350 573.600 885.600 ;
        RECT 577.950 884.100 580.050 886.200 ;
        RECT 578.400 883.350 579.600 884.100 ;
        RECT 568.950 880.950 571.050 883.050 ;
        RECT 571.950 880.950 574.050 883.050 ;
        RECT 574.950 880.950 577.050 883.050 ;
        RECT 577.950 880.950 580.050 883.050 ;
        RECT 569.400 879.900 570.600 880.650 ;
        RECT 575.400 879.900 576.600 880.650 ;
        RECT 584.400 879.900 585.450 889.950 ;
        RECT 562.950 877.800 565.050 879.900 ;
        RECT 568.950 877.800 571.050 879.900 ;
        RECT 574.950 877.800 577.050 879.900 ;
        RECT 583.950 877.800 586.050 879.900 ;
        RECT 559.950 847.950 562.050 850.050 ;
        RECT 550.950 844.950 553.050 847.050 ;
        RECT 551.400 840.600 552.450 844.950 ;
        RECT 551.400 838.350 552.600 840.600 ;
        RECT 556.950 839.100 559.050 841.200 ;
        RECT 557.400 838.350 558.600 839.100 ;
        RECT 547.950 835.950 550.050 838.050 ;
        RECT 550.950 835.950 553.050 838.050 ;
        RECT 553.950 835.950 556.050 838.050 ;
        RECT 556.950 835.950 559.050 838.050 ;
        RECT 548.400 834.900 549.600 835.650 ;
        RECT 547.950 832.800 550.050 834.900 ;
        RECT 554.400 833.400 555.600 835.650 ;
        RECT 554.400 820.050 555.450 833.400 ;
        RECT 563.400 822.450 564.450 877.800 ;
        RECT 580.950 853.950 583.050 856.050 ;
        RECT 568.950 844.800 571.050 846.900 ;
        RECT 565.950 839.100 568.050 841.200 ;
        RECT 566.400 826.050 567.450 839.100 ;
        RECT 569.400 835.050 570.450 844.800 ;
        RECT 574.950 839.100 577.050 841.200 ;
        RECT 581.400 840.600 582.450 853.950 ;
        RECT 587.400 847.050 588.450 898.950 ;
        RECT 589.950 889.950 592.050 895.050 ;
        RECT 592.950 884.100 595.050 886.200 ;
        RECT 599.400 885.600 600.450 907.950 ;
        RECT 605.400 898.050 606.450 917.100 ;
        RECT 608.400 901.050 609.450 934.950 ;
        RECT 613.950 922.950 616.050 925.050 ;
        RECT 610.950 919.950 613.050 922.050 ;
        RECT 611.400 912.900 612.450 919.950 ;
        RECT 614.400 918.600 615.450 922.950 ;
        RECT 614.400 916.350 615.600 918.600 ;
        RECT 623.400 918.450 624.600 918.600 ;
        RECT 625.950 918.450 628.050 919.200 ;
        RECT 623.400 917.400 628.050 918.450 ;
        RECT 623.400 916.350 624.600 917.400 ;
        RECT 625.950 917.100 628.050 917.400 ;
        RECT 614.100 913.950 616.200 916.050 ;
        RECT 617.400 913.950 619.500 916.050 ;
        RECT 622.800 913.950 624.900 916.050 ;
        RECT 617.400 912.900 618.600 913.650 ;
        RECT 610.950 910.800 613.050 912.900 ;
        RECT 616.950 910.800 619.050 912.900 ;
        RECT 626.400 910.050 627.450 917.100 ;
        RECT 625.950 907.950 628.050 910.050 ;
        RECT 629.400 907.050 630.450 952.950 ;
        RECT 641.400 937.050 642.450 956.400 ;
        RECT 646.950 955.800 649.050 957.900 ;
        RECT 661.950 955.800 664.050 957.900 ;
        RECT 667.950 955.800 670.050 957.900 ;
        RECT 676.950 955.800 679.050 957.900 ;
        RECT 689.400 956.400 690.600 958.650 ;
        RECT 707.400 957.900 708.600 958.650 ;
        RECT 713.400 957.900 714.600 958.650 ;
        RECT 719.400 957.900 720.450 964.950 ;
        RECT 724.950 962.100 727.050 964.200 ;
        RECT 733.950 963.000 736.050 967.050 ;
        RECT 725.400 958.050 726.450 962.100 ;
        RECT 734.400 961.350 735.600 963.000 ;
        RECT 757.950 962.100 760.050 964.200 ;
        RECT 763.950 963.000 766.050 967.050 ;
        RECT 782.400 963.600 783.450 970.950 ;
        RECT 817.950 967.950 820.050 970.050 ;
        RECT 784.950 966.450 787.050 967.050 ;
        RECT 790.950 966.450 793.050 967.050 ;
        RECT 784.950 965.400 793.050 966.450 ;
        RECT 784.950 964.950 787.050 965.400 ;
        RECT 790.950 964.950 793.050 965.400 ;
        RECT 758.400 961.350 759.600 962.100 ;
        RECT 764.400 961.350 765.600 963.000 ;
        RECT 782.400 961.350 783.600 963.600 ;
        RECT 787.950 962.100 790.050 964.200 ;
        RECT 788.400 961.350 789.600 962.100 ;
        RECT 793.950 961.950 796.050 964.050 ;
        RECT 802.950 962.100 805.050 964.200 ;
        RECT 808.950 963.000 811.050 967.050 ;
        RECT 730.950 958.950 733.050 961.050 ;
        RECT 733.950 958.950 736.050 961.050 ;
        RECT 736.950 958.950 739.050 961.050 ;
        RECT 754.950 958.950 757.050 961.050 ;
        RECT 757.950 958.950 760.050 961.050 ;
        RECT 760.950 958.950 763.050 961.050 ;
        RECT 763.950 958.950 766.050 961.050 ;
        RECT 778.950 958.950 781.050 961.050 ;
        RECT 781.950 958.950 784.050 961.050 ;
        RECT 784.950 958.950 787.050 961.050 ;
        RECT 787.950 958.950 790.050 961.050 ;
        RECT 640.950 934.950 643.050 937.050 ;
        RECT 647.400 931.050 648.450 955.800 ;
        RECT 689.400 940.050 690.450 956.400 ;
        RECT 706.950 955.800 709.050 957.900 ;
        RECT 712.950 955.800 715.050 957.900 ;
        RECT 718.950 955.800 721.050 957.900 ;
        RECT 724.950 955.950 727.050 958.050 ;
        RECT 731.400 957.900 732.600 958.650 ;
        RECT 737.400 957.900 738.600 958.650 ;
        RECT 755.400 957.900 756.600 958.650 ;
        RECT 730.950 955.800 733.050 957.900 ;
        RECT 736.950 955.800 739.050 957.900 ;
        RECT 754.950 955.800 757.050 957.900 ;
        RECT 761.400 957.000 762.600 958.650 ;
        RECT 697.950 949.950 700.050 952.050 ;
        RECT 688.950 937.950 691.050 940.050 ;
        RECT 646.950 928.950 649.050 931.050 ;
        RECT 673.950 928.950 676.050 931.050 ;
        RECT 640.950 922.950 643.050 925.050 ;
        RECT 641.400 919.200 642.450 922.950 ;
        RECT 640.950 917.100 643.050 919.200 ;
        RECT 646.950 917.100 649.050 919.200 ;
        RECT 655.950 917.100 658.050 919.200 ;
        RECT 667.950 917.100 670.050 919.200 ;
        RECT 674.400 918.600 675.450 928.950 ;
        RECT 689.400 928.050 690.450 937.950 ;
        RECT 688.950 925.950 691.050 928.050 ;
        RECT 641.400 916.350 642.600 917.100 ;
        RECT 647.400 916.350 648.600 917.100 ;
        RECT 640.950 913.950 643.050 916.050 ;
        RECT 643.950 913.950 646.050 916.050 ;
        RECT 646.950 913.950 649.050 916.050 ;
        RECT 649.950 913.950 652.050 916.050 ;
        RECT 644.400 912.900 645.600 913.650 ;
        RECT 643.950 910.800 646.050 912.900 ;
        RECT 650.400 911.400 651.600 913.650 ;
        RECT 640.950 907.950 643.050 910.050 ;
        RECT 628.950 904.950 631.050 907.050 ;
        RECT 610.950 901.950 613.050 904.050 ;
        RECT 607.950 898.950 610.050 901.050 ;
        RECT 604.950 895.950 607.050 898.050 ;
        RECT 593.400 883.350 594.600 884.100 ;
        RECT 599.400 883.350 600.600 885.600 ;
        RECT 607.950 884.100 610.050 886.200 ;
        RECT 592.950 880.950 595.050 883.050 ;
        RECT 595.950 880.950 598.050 883.050 ;
        RECT 598.950 880.950 601.050 883.050 ;
        RECT 601.950 880.950 604.050 883.050 ;
        RECT 596.400 879.900 597.600 880.650 ;
        RECT 595.950 877.800 598.050 879.900 ;
        RECT 602.400 879.000 603.600 880.650 ;
        RECT 601.950 874.950 604.050 879.000 ;
        RECT 608.400 874.050 609.450 884.100 ;
        RECT 611.400 879.900 612.450 901.950 ;
        RECT 634.950 889.950 637.050 892.050 ;
        RECT 619.950 884.100 622.050 886.200 ;
        RECT 625.950 884.100 628.050 886.200 ;
        RECT 620.400 883.350 621.600 884.100 ;
        RECT 626.400 883.350 627.600 884.100 ;
        RECT 616.950 880.950 619.050 883.050 ;
        RECT 619.950 880.950 622.050 883.050 ;
        RECT 622.950 880.950 625.050 883.050 ;
        RECT 625.950 880.950 628.050 883.050 ;
        RECT 617.400 879.900 618.600 880.650 ;
        RECT 610.950 877.800 613.050 879.900 ;
        RECT 616.950 877.800 619.050 879.900 ;
        RECT 623.400 879.000 624.600 880.650 ;
        RECT 622.950 874.950 625.050 879.000 ;
        RECT 635.400 874.050 636.450 889.950 ;
        RECT 641.400 885.600 642.450 907.950 ;
        RECT 650.400 901.050 651.450 911.400 ;
        RECT 656.400 904.050 657.450 917.100 ;
        RECT 668.400 916.350 669.600 917.100 ;
        RECT 674.400 916.350 675.600 918.600 ;
        RECT 691.950 917.100 694.050 919.200 ;
        RECT 698.400 919.050 699.450 949.950 ;
        RECT 727.950 934.950 730.050 937.050 ;
        RECT 700.950 925.950 703.050 928.050 ;
        RECT 692.400 916.350 693.600 917.100 ;
        RECT 697.950 916.950 700.050 919.050 ;
        RECT 664.950 913.950 667.050 916.050 ;
        RECT 667.950 913.950 670.050 916.050 ;
        RECT 670.950 913.950 673.050 916.050 ;
        RECT 673.950 913.950 676.050 916.050 ;
        RECT 691.950 913.950 694.050 916.050 ;
        RECT 694.950 913.950 697.050 916.050 ;
        RECT 665.400 911.400 666.600 913.650 ;
        RECT 671.400 911.400 672.600 913.650 ;
        RECT 695.400 912.900 696.600 913.650 ;
        RECT 701.400 912.900 702.450 925.950 ;
        RECT 703.950 917.100 706.050 919.200 ;
        RECT 712.950 917.100 715.050 919.200 ;
        RECT 718.950 918.000 721.050 922.050 ;
        RECT 665.400 907.050 666.450 911.400 ;
        RECT 671.400 907.050 672.450 911.400 ;
        RECT 694.950 910.800 697.050 912.900 ;
        RECT 700.950 910.800 703.050 912.900 ;
        RECT 664.950 904.950 667.050 907.050 ;
        RECT 670.950 904.950 673.050 907.050 ;
        RECT 655.950 901.950 658.050 904.050 ;
        RECT 649.950 898.950 652.050 901.050 ;
        RECT 641.400 883.350 642.600 885.600 ;
        RECT 646.950 884.100 649.050 886.200 ;
        RECT 647.400 883.350 648.600 884.100 ;
        RECT 640.950 880.950 643.050 883.050 ;
        RECT 643.950 880.950 646.050 883.050 ;
        RECT 646.950 880.950 649.050 883.050 ;
        RECT 649.950 880.950 652.050 883.050 ;
        RECT 644.400 878.400 645.600 880.650 ;
        RECT 650.400 879.900 651.600 880.650 ;
        RECT 637.950 874.950 640.050 877.050 ;
        RECT 607.950 871.950 610.050 874.050 ;
        RECT 634.950 871.950 637.050 874.050 ;
        RECT 589.950 868.950 592.050 871.050 ;
        RECT 586.950 844.950 589.050 847.050 ;
        RECT 575.400 838.350 576.600 839.100 ;
        RECT 581.400 838.350 582.600 840.600 ;
        RECT 574.950 835.950 577.050 838.050 ;
        RECT 577.950 835.950 580.050 838.050 ;
        RECT 580.950 835.950 583.050 838.050 ;
        RECT 583.950 835.950 586.050 838.050 ;
        RECT 568.950 832.950 571.050 835.050 ;
        RECT 578.400 833.400 579.600 835.650 ;
        RECT 584.400 835.050 585.600 835.650 ;
        RECT 590.400 835.050 591.450 868.950 ;
        RECT 604.950 856.950 607.050 859.050 ;
        RECT 622.950 856.950 625.050 859.050 ;
        RECT 592.950 839.100 595.050 841.200 ;
        RECT 598.950 839.100 601.050 841.200 ;
        RECT 605.400 840.600 606.450 856.950 ;
        RECT 623.400 844.050 624.450 856.950 ;
        RECT 593.400 835.050 594.450 839.100 ;
        RECT 599.400 838.350 600.600 839.100 ;
        RECT 605.400 838.350 606.600 840.600 ;
        RECT 622.950 840.000 625.050 844.050 ;
        RECT 623.400 838.350 624.600 840.000 ;
        RECT 598.950 835.950 601.050 838.050 ;
        RECT 601.950 835.950 604.050 838.050 ;
        RECT 604.950 835.950 607.050 838.050 ;
        RECT 622.950 835.950 625.050 838.050 ;
        RECT 625.950 835.950 628.050 838.050 ;
        RECT 628.950 835.950 631.050 838.050 ;
        RECT 584.400 833.400 589.050 835.050 ;
        RECT 565.950 823.950 568.050 826.050 ;
        RECT 563.400 821.400 567.450 822.450 ;
        RECT 553.950 819.450 556.050 820.050 ;
        RECT 551.400 818.400 556.050 819.450 ;
        RECT 547.950 811.950 550.050 814.050 ;
        RECT 541.950 808.950 544.050 811.050 ;
        RECT 533.400 805.350 534.600 807.600 ;
        RECT 539.400 805.350 540.600 807.600 ;
        RECT 532.950 802.950 535.050 805.050 ;
        RECT 535.950 802.950 538.050 805.050 ;
        RECT 538.950 802.950 541.050 805.050 ;
        RECT 541.950 802.950 544.050 805.050 ;
        RECT 529.950 799.950 532.050 802.050 ;
        RECT 536.400 800.400 537.600 802.650 ;
        RECT 542.400 802.050 543.600 802.650 ;
        RECT 548.400 802.050 549.450 811.950 ;
        RECT 551.400 802.050 552.450 818.400 ;
        RECT 553.950 817.950 556.050 818.400 ;
        RECT 556.950 806.100 559.050 808.200 ;
        RECT 557.400 805.350 558.600 806.100 ;
        RECT 556.950 802.950 559.050 805.050 ;
        RECT 559.950 802.950 562.050 805.050 ;
        RECT 542.400 800.400 547.050 802.050 ;
        RECT 530.400 775.050 531.450 799.950 ;
        RECT 536.400 793.050 537.450 800.400 ;
        RECT 543.000 799.950 547.050 800.400 ;
        RECT 547.950 799.950 550.050 802.050 ;
        RECT 550.950 799.950 553.050 802.050 ;
        RECT 560.400 801.900 561.600 802.650 ;
        RECT 559.950 799.800 562.050 801.900 ;
        RECT 535.950 790.950 538.050 793.050 ;
        RECT 566.400 790.050 567.450 821.400 ;
        RECT 578.400 820.050 579.450 833.400 ;
        RECT 585.000 832.950 589.050 833.400 ;
        RECT 589.950 832.950 592.050 835.050 ;
        RECT 592.950 832.950 595.050 835.050 ;
        RECT 602.400 834.900 603.600 835.650 ;
        RECT 626.400 834.900 627.600 835.650 ;
        RECT 601.950 832.800 604.050 834.900 ;
        RECT 625.950 832.800 628.050 834.900 ;
        RECT 613.950 829.950 616.050 832.050 ;
        RECT 580.950 823.950 583.050 826.050 ;
        RECT 577.950 817.950 580.050 820.050 ;
        RECT 571.950 805.950 574.050 808.050 ;
        RECT 581.400 807.600 582.450 823.950 ;
        RECT 572.400 801.900 573.450 805.950 ;
        RECT 581.400 805.350 582.600 807.600 ;
        RECT 601.950 807.000 604.050 811.050 ;
        RECT 607.950 808.950 610.050 811.050 ;
        RECT 602.400 805.350 603.600 807.000 ;
        RECT 577.950 802.950 580.050 805.050 ;
        RECT 580.950 802.950 583.050 805.050 ;
        RECT 583.950 802.950 586.050 805.050 ;
        RECT 598.950 802.950 601.050 805.050 ;
        RECT 601.950 802.950 604.050 805.050 ;
        RECT 578.400 801.900 579.600 802.650 ;
        RECT 584.400 801.900 585.600 802.650 ;
        RECT 599.400 801.900 600.600 802.650 ;
        RECT 571.950 799.800 574.050 801.900 ;
        RECT 577.950 799.800 580.050 801.900 ;
        RECT 583.950 799.800 586.050 801.900 ;
        RECT 559.950 787.950 562.050 790.050 ;
        RECT 565.950 787.950 568.050 790.050 ;
        RECT 529.950 772.950 532.050 775.050 ;
        RECT 526.950 769.950 529.050 772.050 ;
        RECT 527.400 765.450 528.450 769.950 ;
        RECT 524.400 764.400 528.450 765.450 ;
        RECT 524.400 762.600 525.450 764.400 ;
        RECT 530.400 762.600 531.450 772.950 ;
        RECT 535.950 766.950 538.050 769.050 ;
        RECT 550.950 766.950 553.050 769.050 ;
        RECT 524.400 760.350 525.600 762.600 ;
        RECT 530.400 760.350 531.600 762.600 ;
        RECT 523.950 757.950 526.050 760.050 ;
        RECT 526.950 757.950 529.050 760.050 ;
        RECT 529.950 757.950 532.050 760.050 ;
        RECT 527.400 755.400 528.600 757.650 ;
        RECT 514.950 739.950 517.050 742.050 ;
        RECT 520.950 730.950 523.050 733.050 ;
        RECT 506.400 727.350 507.600 729.600 ;
        RECT 511.950 728.100 514.050 730.200 ;
        RECT 512.400 727.350 513.600 728.100 ;
        RECT 502.950 724.950 505.050 727.050 ;
        RECT 505.950 724.950 508.050 727.050 ;
        RECT 508.950 724.950 511.050 727.050 ;
        RECT 511.950 724.950 514.050 727.050 ;
        RECT 514.950 724.950 517.050 727.050 ;
        RECT 503.400 723.900 504.600 724.650 ;
        RECT 509.400 723.900 510.600 724.650 ;
        RECT 496.950 721.800 499.050 723.900 ;
        RECT 502.950 721.800 505.050 723.900 ;
        RECT 508.950 721.800 511.050 723.900 ;
        RECT 515.400 722.400 516.600 724.650 ;
        RECT 515.400 720.450 516.450 722.400 ;
        RECT 517.950 721.950 520.050 724.050 ;
        RECT 512.400 719.400 516.450 720.450 ;
        RECT 493.950 715.950 496.050 718.050 ;
        RECT 502.950 694.950 505.050 697.050 ;
        RECT 484.950 688.950 487.050 691.050 ;
        RECT 490.950 688.950 493.050 691.050 ;
        RECT 485.400 684.600 486.450 688.950 ;
        RECT 485.400 682.350 486.600 684.600 ;
        RECT 490.950 683.100 493.050 685.200 ;
        RECT 491.400 682.350 492.600 683.100 ;
        RECT 484.950 679.950 487.050 682.050 ;
        RECT 487.950 679.950 490.050 682.050 ;
        RECT 490.950 679.950 493.050 682.050 ;
        RECT 493.950 679.950 496.050 682.050 ;
        RECT 499.950 679.950 502.050 682.050 ;
        RECT 488.400 677.400 489.600 679.650 ;
        RECT 494.400 678.000 495.600 679.650 ;
        RECT 488.400 673.050 489.450 677.400 ;
        RECT 493.950 673.950 496.050 678.000 ;
        RECT 487.950 670.950 490.050 673.050 ;
        RECT 500.400 670.050 501.450 679.950 ;
        RECT 503.400 678.900 504.450 694.950 ;
        RECT 512.400 685.200 513.450 719.400 ;
        RECT 514.950 706.950 517.050 709.050 ;
        RECT 515.400 688.050 516.450 706.950 ;
        RECT 518.400 706.050 519.450 721.950 ;
        RECT 517.950 703.950 520.050 706.050 ;
        RECT 521.400 691.050 522.450 730.950 ;
        RECT 527.400 729.450 528.450 755.400 ;
        RECT 536.400 754.050 537.450 766.950 ;
        RECT 538.950 761.100 541.050 763.200 ;
        RECT 544.950 761.100 547.050 763.200 ;
        RECT 551.400 762.600 552.450 766.950 ;
        RECT 535.950 751.950 538.050 754.050 ;
        RECT 539.400 748.050 540.450 761.100 ;
        RECT 545.400 760.350 546.600 761.100 ;
        RECT 551.400 760.350 552.600 762.600 ;
        RECT 556.950 761.100 559.050 763.200 ;
        RECT 544.950 757.950 547.050 760.050 ;
        RECT 547.950 757.950 550.050 760.050 ;
        RECT 550.950 757.950 553.050 760.050 ;
        RECT 548.400 756.900 549.600 757.650 ;
        RECT 557.400 757.050 558.450 761.100 ;
        RECT 560.400 757.050 561.450 787.950 ;
        RECT 572.400 784.050 573.450 799.800 ;
        RECT 598.950 796.950 601.050 801.900 ;
        RECT 604.950 801.450 607.050 801.900 ;
        RECT 608.400 801.450 609.450 808.950 ;
        RECT 604.950 800.400 609.450 801.450 ;
        RECT 604.950 799.800 607.050 800.400 ;
        RECT 605.400 793.050 606.450 799.800 ;
        RECT 604.950 790.950 607.050 793.050 ;
        RECT 610.950 790.950 613.050 793.050 ;
        RECT 571.950 781.950 574.050 784.050 ;
        RECT 583.950 778.950 586.050 781.050 ;
        RECT 565.950 775.950 568.050 778.050 ;
        RECT 566.400 763.200 567.450 775.950 ;
        RECT 565.950 761.100 568.050 763.200 ;
        RECT 571.950 761.100 574.050 763.200 ;
        RECT 566.400 760.350 567.600 761.100 ;
        RECT 572.400 760.350 573.600 761.100 ;
        RECT 565.950 757.950 568.050 760.050 ;
        RECT 568.950 757.950 571.050 760.050 ;
        RECT 571.950 757.950 574.050 760.050 ;
        RECT 574.950 757.950 577.050 760.050 ;
        RECT 547.950 754.800 550.050 756.900 ;
        RECT 556.800 754.950 558.900 757.050 ;
        RECT 559.950 754.950 562.050 757.050 ;
        RECT 569.400 756.900 570.600 757.650 ;
        RECT 568.950 754.800 571.050 756.900 ;
        RECT 575.400 755.400 576.600 757.650 ;
        RECT 544.950 751.950 547.050 754.050 ;
        RECT 538.950 745.950 541.050 748.050 ;
        RECT 524.400 728.400 528.450 729.450 ;
        RECT 529.950 729.000 532.050 733.050 ;
        RECT 524.400 697.050 525.450 728.400 ;
        RECT 530.400 727.350 531.600 729.000 ;
        RECT 535.950 728.100 538.050 730.200 ;
        RECT 536.400 727.350 537.600 728.100 ;
        RECT 529.950 724.950 532.050 727.050 ;
        RECT 532.950 724.950 535.050 727.050 ;
        RECT 535.950 724.950 538.050 727.050 ;
        RECT 538.950 724.950 541.050 727.050 ;
        RECT 526.950 721.800 529.050 723.900 ;
        RECT 533.400 722.400 534.600 724.650 ;
        RECT 539.400 723.000 540.600 724.650 ;
        RECT 527.400 712.050 528.450 721.800 ;
        RECT 526.950 709.950 529.050 712.050 ;
        RECT 523.950 694.950 526.050 697.050 ;
        RECT 520.950 688.950 523.050 691.050 ;
        RECT 514.950 685.950 517.050 688.050 ;
        RECT 520.950 685.800 523.050 687.900 ;
        RECT 511.950 683.100 514.050 685.200 ;
        RECT 512.400 682.350 513.600 683.100 ;
        RECT 508.950 679.950 511.050 682.050 ;
        RECT 511.950 679.950 514.050 682.050 ;
        RECT 514.950 679.950 517.050 682.050 ;
        RECT 509.400 678.900 510.600 679.650 ;
        RECT 502.950 676.800 505.050 678.900 ;
        RECT 508.950 676.800 511.050 678.900 ;
        RECT 515.400 677.400 516.600 679.650 ;
        RECT 521.400 679.050 522.450 685.800 ;
        RECT 523.950 682.950 526.050 685.050 ;
        RECT 515.400 676.050 516.450 677.400 ;
        RECT 520.950 676.950 523.050 679.050 ;
        RECT 524.400 676.050 525.450 682.950 ;
        RECT 514.950 673.950 517.050 676.050 ;
        RECT 523.950 673.950 526.050 676.050 ;
        RECT 499.950 667.950 502.050 670.050 ;
        RECT 493.950 664.950 496.050 667.050 ;
        RECT 494.400 651.600 495.450 664.950 ;
        RECT 515.400 664.050 516.450 673.950 ;
        RECT 514.950 663.450 517.050 664.050 ;
        RECT 512.400 662.400 517.050 663.450 ;
        RECT 502.950 655.950 505.050 658.050 ;
        RECT 494.400 649.350 495.600 651.600 ;
        RECT 484.950 646.950 487.050 649.050 ;
        RECT 487.950 646.950 490.050 649.050 ;
        RECT 490.950 646.950 493.050 649.050 ;
        RECT 493.950 646.950 496.050 649.050 ;
        RECT 485.400 644.400 486.600 646.650 ;
        RECT 491.400 645.900 492.600 646.650 ;
        RECT 485.400 628.050 486.450 644.400 ;
        RECT 490.950 643.800 493.050 645.900 ;
        RECT 503.400 645.450 504.450 655.950 ;
        RECT 512.400 651.600 513.450 662.400 ;
        RECT 514.950 661.950 517.050 662.400 ;
        RECT 512.400 649.350 513.600 651.600 ;
        RECT 517.950 650.100 520.050 652.200 ;
        RECT 518.400 649.350 519.600 650.100 ;
        RECT 511.950 646.950 514.050 649.050 ;
        RECT 514.950 646.950 517.050 649.050 ;
        RECT 517.950 646.950 520.050 649.050 ;
        RECT 520.950 646.950 523.050 649.050 ;
        RECT 515.400 645.900 516.600 646.650 ;
        RECT 505.950 645.450 508.050 645.900 ;
        RECT 503.400 644.400 508.050 645.450 ;
        RECT 505.950 643.800 508.050 644.400 ;
        RECT 514.950 643.800 517.050 645.900 ;
        RECT 521.400 644.400 522.600 646.650 ;
        RECT 506.400 637.050 507.450 643.800 ;
        RECT 505.950 634.950 508.050 637.050 ;
        RECT 472.950 625.950 475.050 628.050 ;
        RECT 478.950 625.950 481.050 628.050 ;
        RECT 484.950 625.950 487.050 628.050 ;
        RECT 473.400 606.600 474.450 625.950 ;
        RECT 478.950 619.950 481.050 622.050 ;
        RECT 505.950 619.950 508.050 622.050 ;
        RECT 479.400 606.600 480.450 619.950 ;
        RECT 473.400 604.350 474.600 606.600 ;
        RECT 479.400 604.350 480.600 606.600 ;
        RECT 496.950 606.000 499.050 610.050 ;
        RECT 497.400 604.350 498.600 606.000 ;
        RECT 472.950 601.950 475.050 604.050 ;
        RECT 475.950 601.950 478.050 604.050 ;
        RECT 478.950 601.950 481.050 604.050 ;
        RECT 497.100 601.950 499.200 604.050 ;
        RECT 502.500 601.950 504.600 604.050 ;
        RECT 476.400 599.400 477.600 601.650 ;
        RECT 503.400 600.900 504.600 601.650 ;
        RECT 476.400 589.050 477.450 599.400 ;
        RECT 502.950 598.800 505.050 600.900 ;
        RECT 475.950 586.950 478.050 589.050 ;
        RECT 487.950 586.950 490.050 589.050 ;
        RECT 479.850 579.300 481.950 581.400 ;
        RECT 466.950 574.950 469.050 577.050 ;
        RECT 466.950 568.950 469.050 571.050 ;
        RECT 475.950 568.950 478.050 571.050 ;
        RECT 467.400 567.900 468.600 568.650 ;
        RECT 476.400 567.900 477.600 568.650 ;
        RECT 466.950 565.800 469.050 567.900 ;
        RECT 475.950 565.800 478.050 567.900 ;
        RECT 460.650 559.500 464.850 560.700 ;
        RECT 445.350 555.600 447.450 557.700 ;
        RECT 448.950 556.950 451.050 559.050 ;
        RECT 460.650 558.600 462.750 559.500 ;
        RECT 467.400 553.050 468.450 565.800 ;
        RECT 480.150 560.700 481.350 579.300 ;
        RECT 488.400 574.050 489.450 586.950 ;
        RECT 497.550 579.300 499.650 581.400 ;
        RECT 493.950 574.950 496.050 577.050 ;
        RECT 487.950 571.950 490.050 574.050 ;
        RECT 485.100 568.950 487.200 571.050 ;
        RECT 485.400 567.900 486.600 568.650 ;
        RECT 484.950 565.800 487.050 567.900 ;
        RECT 480.150 559.500 484.350 560.700 ;
        RECT 482.250 558.600 484.350 559.500 ;
        RECT 463.950 550.950 466.050 553.050 ;
        RECT 466.950 550.950 469.050 553.050 ;
        RECT 442.350 537.300 444.450 539.400 ;
        RECT 418.950 526.950 421.050 529.050 ;
        RECT 424.950 527.100 427.050 529.200 ;
        RECT 430.950 528.000 433.050 532.050 ;
        RECT 436.950 529.950 439.050 532.050 ;
        RECT 443.250 530.700 444.450 537.300 ;
        RECT 457.650 535.500 459.750 536.400 ;
        RECT 457.650 534.300 461.850 535.500 ;
        RECT 442.350 528.600 444.450 530.700 ;
        RECT 425.400 526.350 426.600 527.100 ;
        RECT 431.400 526.350 432.600 528.000 ;
        RECT 421.950 523.950 424.050 526.050 ;
        RECT 424.950 523.950 427.050 526.050 ;
        RECT 427.950 523.950 430.050 526.050 ;
        RECT 430.950 523.950 433.050 526.050 ;
        RECT 436.950 523.950 439.050 526.050 ;
        RECT 415.950 520.950 418.050 523.050 ;
        RECT 418.950 520.950 421.050 523.050 ;
        RECT 422.400 522.900 423.600 523.650 ;
        RECT 428.400 522.900 429.600 523.650 ;
        RECT 412.950 517.950 415.050 520.050 ;
        RECT 409.950 502.950 412.050 505.050 ;
        RECT 415.950 499.950 418.050 502.050 ;
        RECT 416.400 495.600 417.450 499.950 ;
        RECT 419.400 498.450 420.450 520.950 ;
        RECT 421.950 520.800 424.050 522.900 ;
        RECT 427.950 520.800 430.050 522.900 ;
        RECT 437.400 521.400 438.600 523.650 ;
        RECT 422.400 508.050 423.450 520.800 ;
        RECT 424.950 517.950 427.050 520.050 ;
        RECT 425.400 514.050 426.450 517.950 ;
        RECT 430.950 514.950 433.050 517.050 ;
        RECT 424.950 511.950 427.050 514.050 ;
        RECT 421.950 505.950 424.050 508.050 ;
        RECT 419.400 497.400 423.450 498.450 ;
        RECT 416.400 493.350 417.600 495.600 ;
        RECT 418.950 493.950 421.050 496.050 ;
        RECT 410.100 490.950 412.200 493.050 ;
        RECT 415.500 490.950 417.600 493.050 ;
        RECT 410.400 489.450 411.600 490.650 ;
        RECT 391.950 484.950 394.050 489.000 ;
        RECT 407.400 488.400 411.600 489.450 ;
        RECT 382.950 478.950 385.050 481.050 ;
        RECT 379.950 451.950 382.050 454.050 ;
        RECT 374.400 448.350 375.600 450.000 ;
        RECT 377.400 449.400 381.450 450.450 ;
        RECT 361.950 445.950 364.050 448.050 ;
        RECT 364.950 445.950 367.050 448.050 ;
        RECT 367.950 445.950 370.050 448.050 ;
        RECT 370.950 445.950 373.050 448.050 ;
        RECT 373.950 445.950 376.050 448.050 ;
        RECT 365.400 443.400 366.600 445.650 ;
        RECT 371.400 443.400 372.600 445.650 ;
        RECT 355.950 439.950 358.050 442.050 ;
        RECT 365.400 439.050 366.450 443.400 ;
        RECT 371.400 441.450 372.450 443.400 ;
        RECT 371.400 440.400 375.450 441.450 ;
        RECT 364.950 436.950 367.050 439.050 ;
        RECT 374.400 427.050 375.450 440.400 ;
        RECT 380.400 430.050 381.450 449.400 ;
        RECT 383.400 444.900 384.450 478.950 ;
        RECT 419.400 456.450 420.450 493.950 ;
        RECT 422.400 489.900 423.450 497.400 ;
        RECT 431.400 495.600 432.450 514.950 ;
        RECT 437.400 505.050 438.450 521.400 ;
        RECT 443.250 515.700 444.450 528.600 ;
        RECT 454.950 527.100 457.050 529.200 ;
        RECT 455.400 526.350 456.600 527.100 ;
        RECT 454.800 523.950 456.900 526.050 ;
        RECT 442.350 513.600 444.450 515.700 ;
        RECT 448.950 514.950 451.050 517.050 ;
        RECT 460.650 515.700 461.850 534.300 ;
        RECT 464.400 529.200 465.450 550.950 ;
        RECT 472.950 547.950 475.050 550.050 ;
        RECT 463.950 527.100 466.050 529.200 ;
        RECT 464.400 526.350 465.600 527.100 ;
        RECT 469.950 526.950 472.050 529.050 ;
        RECT 463.950 523.950 466.050 526.050 ;
        RECT 436.950 502.950 439.050 505.050 ;
        RECT 445.950 496.950 448.050 499.050 ;
        RECT 431.400 493.350 432.600 495.600 ;
        RECT 436.950 494.100 439.050 496.200 ;
        RECT 437.400 493.350 438.600 494.100 ;
        RECT 430.950 490.950 433.050 493.050 ;
        RECT 433.950 490.950 436.050 493.050 ;
        RECT 436.950 490.950 439.050 493.050 ;
        RECT 439.950 490.950 442.050 493.050 ;
        RECT 434.400 489.900 435.600 490.650 ;
        RECT 440.400 489.900 441.600 490.650 ;
        RECT 446.400 489.900 447.450 496.950 ;
        RECT 421.950 487.800 424.050 489.900 ;
        RECT 433.950 487.800 436.050 489.900 ;
        RECT 439.950 487.800 442.050 489.900 ;
        RECT 445.950 487.800 448.050 489.900 ;
        RECT 449.400 489.450 450.450 514.950 ;
        RECT 460.050 513.600 462.150 515.700 ;
        RECT 470.400 502.050 471.450 526.950 ;
        RECT 463.950 499.950 466.050 502.050 ;
        RECT 469.950 499.950 472.050 502.050 ;
        RECT 457.950 495.000 460.050 499.050 ;
        RECT 464.400 496.200 465.450 499.950 ;
        RECT 463.950 495.450 466.050 496.200 ;
        RECT 458.400 493.350 459.600 495.000 ;
        RECT 463.950 494.400 468.450 495.450 ;
        RECT 463.950 494.100 466.050 494.400 ;
        RECT 454.950 490.950 457.050 493.050 ;
        RECT 457.950 490.950 460.050 493.050 ;
        RECT 460.950 490.950 463.050 493.050 ;
        RECT 455.400 489.450 456.600 490.650 ;
        RECT 449.400 488.400 456.600 489.450 ;
        RECT 461.400 488.400 462.600 490.650 ;
        RECT 461.400 475.050 462.450 488.400 ;
        RECT 460.950 472.950 463.050 475.050 ;
        RECT 467.400 468.450 468.450 494.400 ;
        RECT 473.400 489.450 474.450 547.950 ;
        RECT 494.400 538.050 495.450 574.950 ;
        RECT 497.550 566.400 498.750 579.300 ;
        RECT 503.400 577.050 504.450 598.800 ;
        RECT 506.400 580.050 507.450 619.950 ;
        RECT 521.400 619.050 522.450 644.400 ;
        RECT 527.400 636.450 528.450 709.950 ;
        RECT 533.400 709.050 534.450 722.400 ;
        RECT 538.950 718.950 541.050 723.000 ;
        RECT 545.400 721.050 546.450 751.950 ;
        RECT 575.400 748.050 576.450 755.400 ;
        RECT 556.950 745.950 559.050 748.050 ;
        RECT 568.950 745.950 571.050 748.050 ;
        RECT 574.950 745.950 577.050 748.050 ;
        RECT 547.950 739.950 550.050 742.050 ;
        RECT 544.950 718.950 547.050 721.050 ;
        RECT 532.950 706.950 535.050 709.050 ;
        RECT 535.950 691.950 538.050 694.050 ;
        RECT 529.950 688.950 532.050 691.050 ;
        RECT 530.400 685.050 531.450 688.950 ;
        RECT 529.950 682.950 532.050 685.050 ;
        RECT 536.400 684.600 537.450 691.950 ;
        RECT 536.400 682.350 537.600 684.600 ;
        RECT 541.950 684.000 544.050 688.050 ;
        RECT 542.400 682.350 543.600 684.000 ;
        RECT 532.950 679.950 535.050 682.050 ;
        RECT 535.950 679.950 538.050 682.050 ;
        RECT 538.950 679.950 541.050 682.050 ;
        RECT 541.950 679.950 544.050 682.050 ;
        RECT 533.400 679.050 534.600 679.650 ;
        RECT 529.950 677.400 534.600 679.050 ;
        RECT 539.400 678.000 540.600 679.650 ;
        RECT 529.950 676.950 534.000 677.400 ;
        RECT 538.950 673.950 541.050 678.000 ;
        RECT 532.950 667.950 535.050 670.050 ;
        RECT 529.950 649.950 532.050 652.050 ;
        RECT 524.400 635.400 528.450 636.450 ;
        RECT 520.950 616.950 523.050 619.050 ;
        RECT 524.400 610.050 525.450 635.400 ;
        RECT 526.950 628.950 529.050 631.050 ;
        RECT 527.400 613.050 528.450 628.950 ;
        RECT 526.950 610.950 529.050 613.050 ;
        RECT 508.950 607.950 511.050 610.050 ;
        RECT 523.950 607.950 526.050 610.050 ;
        RECT 505.950 577.950 508.050 580.050 ;
        RECT 502.950 574.950 505.050 577.050 ;
        RECT 503.400 573.450 504.600 573.600 ;
        RECT 506.400 573.450 507.450 577.950 ;
        RECT 503.400 572.400 507.450 573.450 ;
        RECT 503.400 571.350 504.600 572.400 ;
        RECT 502.950 568.950 505.050 571.050 ;
        RECT 497.550 564.300 499.650 566.400 ;
        RECT 497.550 557.700 498.750 564.300 ;
        RECT 502.950 562.950 505.050 565.050 ;
        RECT 497.550 555.600 499.650 557.700 ;
        RECT 503.400 544.050 504.450 562.950 ;
        RECT 502.950 541.950 505.050 544.050 ;
        RECT 509.400 538.050 510.450 607.950 ;
        RECT 527.400 606.600 528.450 610.950 ;
        RECT 527.400 604.350 528.600 606.600 ;
        RECT 521.400 601.950 523.500 604.050 ;
        RECT 526.800 601.950 528.900 604.050 ;
        RECT 521.400 600.900 522.600 601.650 ;
        RECT 530.400 600.900 531.450 649.950 ;
        RECT 533.400 645.900 534.450 667.950 ;
        RECT 541.950 661.950 544.050 664.050 ;
        RECT 542.400 651.600 543.450 661.950 ;
        RECT 542.400 649.350 543.600 651.600 ;
        RECT 536.100 646.950 538.200 649.050 ;
        RECT 541.500 646.950 543.600 649.050 ;
        RECT 544.800 646.950 546.900 649.050 ;
        RECT 532.950 645.450 535.050 645.900 ;
        RECT 536.400 645.450 537.600 646.650 ;
        RECT 532.950 644.400 537.600 645.450 ;
        RECT 545.400 644.400 546.600 646.650 ;
        RECT 532.950 643.800 535.050 644.400 ;
        RECT 535.950 631.950 538.050 634.050 ;
        RECT 520.950 598.800 523.050 600.900 ;
        RECT 529.950 598.800 532.050 600.900 ;
        RECT 536.400 595.050 537.450 631.950 ;
        RECT 545.400 606.600 546.450 644.400 ;
        RECT 548.400 634.050 549.450 739.950 ;
        RECT 557.400 729.600 558.450 745.950 ;
        RECT 557.400 727.350 558.600 729.600 ;
        RECT 565.950 727.950 568.050 730.050 ;
        RECT 553.950 724.950 556.050 727.050 ;
        RECT 556.950 724.950 559.050 727.050 ;
        RECT 559.950 724.950 562.050 727.050 ;
        RECT 554.400 723.900 555.600 724.650 ;
        RECT 553.950 721.800 556.050 723.900 ;
        RECT 566.400 721.050 567.450 727.950 ;
        RECT 569.400 723.900 570.450 745.950 ;
        RECT 575.400 742.050 576.450 745.950 ;
        RECT 574.950 739.950 577.050 742.050 ;
        RECT 577.950 728.100 580.050 730.200 ;
        RECT 584.400 729.600 585.450 778.950 ;
        RECT 586.950 766.950 589.050 769.050 ;
        RECT 587.400 754.050 588.450 766.950 ;
        RECT 595.950 761.100 598.050 763.200 ;
        RECT 596.400 760.350 597.600 761.100 ;
        RECT 592.950 757.950 595.050 760.050 ;
        RECT 595.950 757.950 598.050 760.050 ;
        RECT 598.950 757.950 601.050 760.050 ;
        RECT 593.400 756.000 594.600 757.650 ;
        RECT 586.950 751.950 589.050 754.050 ;
        RECT 592.950 751.950 595.050 756.000 ;
        RECT 599.400 755.400 600.600 757.650 ;
        RECT 599.400 745.050 600.450 755.400 ;
        RECT 598.950 744.450 601.050 745.050 ;
        RECT 596.400 743.400 601.050 744.450 ;
        RECT 592.950 733.950 595.050 736.050 ;
        RECT 578.400 727.350 579.600 728.100 ;
        RECT 584.400 727.350 585.600 729.600 ;
        RECT 574.950 724.950 577.050 727.050 ;
        RECT 577.950 724.950 580.050 727.050 ;
        RECT 580.950 724.950 583.050 727.050 ;
        RECT 583.950 724.950 586.050 727.050 ;
        RECT 575.400 723.900 576.600 724.650 ;
        RECT 568.950 721.800 571.050 723.900 ;
        RECT 574.950 721.800 577.050 723.900 ;
        RECT 581.400 723.000 582.600 724.650 ;
        RECT 565.950 718.950 568.050 721.050 ;
        RECT 580.950 718.950 583.050 723.000 ;
        RECT 586.950 712.950 589.050 715.050 ;
        RECT 587.400 709.050 588.450 712.950 ;
        RECT 586.950 706.950 589.050 709.050 ;
        RECT 562.950 703.950 565.050 706.050 ;
        RECT 550.950 685.950 553.050 688.050 ;
        RECT 551.400 664.050 552.450 685.950 ;
        RECT 556.950 682.950 559.050 691.050 ;
        RECT 563.400 684.600 564.450 703.950 ;
        RECT 568.950 691.950 571.050 694.050 ;
        RECT 577.950 691.950 580.050 694.050 ;
        RECT 569.400 685.200 570.450 691.950 ;
        RECT 563.400 682.350 564.600 684.600 ;
        RECT 568.950 683.100 571.050 685.200 ;
        RECT 574.950 683.100 577.050 685.200 ;
        RECT 569.400 682.350 570.600 683.100 ;
        RECT 559.950 679.950 562.050 682.050 ;
        RECT 562.950 679.950 565.050 682.050 ;
        RECT 565.950 679.950 568.050 682.050 ;
        RECT 568.950 679.950 571.050 682.050 ;
        RECT 556.950 676.950 559.050 679.050 ;
        RECT 560.400 677.400 561.600 679.650 ;
        RECT 566.400 678.900 567.600 679.650 ;
        RECT 550.800 661.950 552.900 664.050 ;
        RECT 557.400 658.050 558.450 676.950 ;
        RECT 560.400 670.050 561.450 677.400 ;
        RECT 565.950 676.800 568.050 678.900 ;
        RECT 568.950 670.950 571.050 673.050 ;
        RECT 559.950 667.950 562.050 670.050 ;
        RECT 556.950 655.950 559.050 658.050 ;
        RECT 569.400 651.600 570.450 670.950 ;
        RECT 569.400 649.350 570.600 651.600 ;
        RECT 559.950 646.950 562.050 649.050 ;
        RECT 562.950 646.950 565.050 649.050 ;
        RECT 565.950 646.950 568.050 649.050 ;
        RECT 568.950 646.950 571.050 649.050 ;
        RECT 560.400 644.400 561.600 646.650 ;
        RECT 566.400 644.400 567.600 646.650 ;
        RECT 547.950 631.950 550.050 634.050 ;
        RECT 560.400 631.050 561.450 644.400 ;
        RECT 566.400 637.050 567.450 644.400 ;
        RECT 565.950 634.950 568.050 637.050 ;
        RECT 553.950 628.950 556.050 631.050 ;
        RECT 559.950 628.950 562.050 631.050 ;
        RECT 547.950 610.950 553.050 613.050 ;
        RECT 545.400 604.350 546.600 606.600 ;
        RECT 550.950 606.000 553.050 609.900 ;
        RECT 554.400 607.050 555.450 628.950 ;
        RECT 556.950 619.950 559.050 622.050 ;
        RECT 562.950 619.950 565.050 622.050 ;
        RECT 557.400 613.050 558.450 619.950 ;
        RECT 559.950 613.950 562.050 616.050 ;
        RECT 556.950 610.950 559.050 613.050 ;
        RECT 556.950 607.800 559.050 609.900 ;
        RECT 551.400 604.350 552.600 606.000 ;
        RECT 553.950 604.950 556.050 607.050 ;
        RECT 541.950 601.950 544.050 604.050 ;
        RECT 544.950 601.950 547.050 604.050 ;
        RECT 547.950 601.950 550.050 604.050 ;
        RECT 550.950 601.950 553.050 604.050 ;
        RECT 542.400 600.900 543.600 601.650 ;
        RECT 541.950 598.800 544.050 600.900 ;
        RECT 548.400 599.400 549.600 601.650 ;
        RECT 529.950 592.950 532.050 595.050 ;
        RECT 535.950 592.950 538.050 595.050 ;
        RECT 511.950 577.950 514.050 580.050 ;
        RECT 493.950 535.950 496.050 538.050 ;
        RECT 499.950 535.950 502.050 538.050 ;
        RECT 508.950 535.950 511.050 538.050 ;
        RECT 484.950 532.950 487.050 535.050 ;
        RECT 485.400 528.600 486.450 532.950 ;
        RECT 485.400 526.350 486.600 528.600 ;
        RECT 490.950 527.100 493.050 529.200 ;
        RECT 496.950 527.100 499.050 529.200 ;
        RECT 491.400 526.350 492.600 527.100 ;
        RECT 481.950 523.950 484.050 526.050 ;
        RECT 484.950 523.950 487.050 526.050 ;
        RECT 487.950 523.950 490.050 526.050 ;
        RECT 490.950 523.950 493.050 526.050 ;
        RECT 482.400 522.900 483.600 523.650 ;
        RECT 481.950 520.800 484.050 522.900 ;
        RECT 488.400 521.400 489.600 523.650 ;
        RECT 482.400 519.450 483.450 520.800 ;
        RECT 482.400 518.400 486.450 519.450 ;
        RECT 481.950 514.950 484.050 517.050 ;
        RECT 482.400 495.600 483.450 514.950 ;
        RECT 482.400 493.350 483.600 495.600 ;
        RECT 476.100 490.950 478.200 493.050 ;
        RECT 481.500 490.950 483.600 493.050 ;
        RECT 476.400 489.450 477.600 490.650 ;
        RECT 473.400 488.400 477.600 489.450 ;
        RECT 464.400 467.400 468.450 468.450 ;
        RECT 416.400 455.400 420.450 456.450 ;
        RECT 391.950 450.000 394.050 454.050 ;
        RECT 392.400 448.350 393.600 450.000 ;
        RECT 397.950 449.100 400.050 451.200 ;
        RECT 403.950 449.100 406.050 451.200 ;
        RECT 416.400 450.600 417.450 455.400 ;
        RECT 433.950 454.950 436.050 457.050 ;
        RECT 451.950 454.950 454.050 457.050 ;
        RECT 398.400 448.350 399.600 449.100 ;
        RECT 388.950 445.950 391.050 448.050 ;
        RECT 391.950 445.950 394.050 448.050 ;
        RECT 394.950 445.950 397.050 448.050 ;
        RECT 397.950 445.950 400.050 448.050 ;
        RECT 389.400 444.900 390.600 445.650 ;
        RECT 382.950 442.800 385.050 444.900 ;
        RECT 388.950 442.800 391.050 444.900 ;
        RECT 395.400 444.000 396.600 445.650 ;
        RECT 394.950 439.950 397.050 444.000 ;
        RECT 400.950 439.950 403.050 442.050 ;
        RECT 385.950 433.950 388.050 436.050 ;
        RECT 379.950 427.950 382.050 430.050 ;
        RECT 350.850 423.300 352.950 425.400 ;
        RECT 368.550 423.300 370.650 425.400 ;
        RECT 373.950 424.950 376.050 427.050 ;
        RECT 343.950 418.950 346.050 421.050 ;
        RECT 337.950 416.100 340.050 418.200 ;
        RECT 338.400 415.350 339.600 416.100 ;
        RECT 337.950 412.950 340.050 415.050 ;
        RECT 346.950 412.950 349.050 415.050 ;
        RECT 347.400 411.000 348.600 412.650 ;
        RECT 332.550 408.300 334.650 410.400 ;
        RECT 332.550 401.700 333.750 408.300 ;
        RECT 346.950 406.950 349.050 411.000 ;
        RECT 351.150 404.700 352.350 423.300 ;
        RECT 356.100 412.950 358.200 415.050 ;
        RECT 356.400 410.400 357.600 412.650 ;
        RECT 368.550 410.400 369.750 423.300 ;
        RECT 373.950 417.000 376.050 421.050 ;
        RECT 374.400 415.350 375.600 417.000 ;
        RECT 373.950 412.950 376.050 415.050 ;
        RECT 356.400 408.450 357.450 410.400 ;
        RECT 356.400 407.400 360.450 408.450 ;
        RECT 351.150 403.500 355.350 404.700 ;
        RECT 332.550 399.600 334.650 401.700 ;
        RECT 340.950 400.950 343.050 403.050 ;
        RECT 353.250 402.600 355.350 403.500 ;
        RECT 341.400 397.050 342.450 400.950 ;
        RECT 340.950 394.950 343.050 397.050 ;
        RECT 334.950 370.950 337.050 373.050 ;
        RECT 340.950 371.100 343.050 373.200 ;
        RECT 346.950 371.100 349.050 373.200 ;
        RECT 352.800 371.100 354.900 373.200 ;
        RECT 355.950 371.100 358.050 373.200 ;
        RECT 359.400 373.050 360.450 407.400 ;
        RECT 368.550 408.300 370.650 410.400 ;
        RECT 368.550 401.700 369.750 408.300 ;
        RECT 379.950 406.950 382.050 409.050 ;
        RECT 368.550 399.600 370.650 401.700 ;
        RECT 367.950 385.950 370.050 388.050 ;
        RECT 335.400 358.050 336.450 370.950 ;
        RECT 341.400 370.350 342.600 371.100 ;
        RECT 347.400 370.350 348.600 371.100 ;
        RECT 340.950 367.950 343.050 370.050 ;
        RECT 343.950 367.950 346.050 370.050 ;
        RECT 346.950 367.950 349.050 370.050 ;
        RECT 344.400 366.000 345.600 367.650 ;
        RECT 343.950 361.950 346.050 366.000 ;
        RECT 349.950 361.950 352.050 367.050 ;
        RECT 334.950 355.950 337.050 358.050 ;
        RECT 328.950 349.950 331.050 352.050 ;
        RECT 325.950 343.950 328.050 346.050 ;
        RECT 344.850 345.300 346.950 347.400 ;
        RECT 326.400 339.600 327.450 343.950 ;
        RECT 326.400 337.350 327.600 339.600 ;
        RECT 331.950 338.100 334.050 340.200 ;
        RECT 332.400 337.350 333.600 338.100 ;
        RECT 325.950 334.950 328.050 337.050 ;
        RECT 328.950 334.950 331.050 337.050 ;
        RECT 331.950 334.950 334.050 337.050 ;
        RECT 334.950 334.950 337.050 337.050 ;
        RECT 340.950 334.950 343.050 337.050 ;
        RECT 329.400 333.900 330.600 334.650 ;
        RECT 328.950 331.800 331.050 333.900 ;
        RECT 335.400 332.400 336.600 334.650 ;
        RECT 341.400 332.400 342.600 334.650 ;
        RECT 335.400 325.050 336.450 332.400 ;
        RECT 341.400 328.050 342.450 332.400 ;
        RECT 340.950 325.950 343.050 328.050 ;
        RECT 345.150 326.700 346.350 345.300 ;
        RECT 353.400 340.050 354.450 371.100 ;
        RECT 356.400 367.050 357.450 371.100 ;
        RECT 358.950 370.950 361.050 373.050 ;
        RECT 361.950 372.000 364.050 376.050 ;
        RECT 368.400 372.600 369.450 385.950 ;
        RECT 362.400 370.350 363.600 372.000 ;
        RECT 368.400 370.350 369.600 372.600 ;
        RECT 361.950 367.950 364.050 370.050 ;
        RECT 364.950 367.950 367.050 370.050 ;
        RECT 367.950 367.950 370.050 370.050 ;
        RECT 370.950 367.950 373.050 370.050 ;
        RECT 355.950 364.950 358.050 367.050 ;
        RECT 358.950 361.950 361.050 367.050 ;
        RECT 365.400 366.000 366.600 367.650 ;
        RECT 371.400 366.900 372.600 367.650 ;
        RECT 364.950 361.950 367.050 366.000 ;
        RECT 370.950 364.800 373.050 366.900 ;
        RECT 355.950 349.950 358.050 352.050 ;
        RECT 352.950 337.950 355.050 340.050 ;
        RECT 350.100 334.950 352.200 337.050 ;
        RECT 350.400 333.900 351.600 334.650 ;
        RECT 349.800 331.800 351.900 333.900 ;
        RECT 352.950 331.950 355.050 334.050 ;
        RECT 345.150 325.500 349.350 326.700 ;
        RECT 319.950 322.950 322.050 325.050 ;
        RECT 334.950 322.950 337.050 325.050 ;
        RECT 347.250 324.600 349.350 325.500 ;
        RECT 346.950 313.950 349.050 316.050 ;
        RECT 334.950 307.950 337.050 310.050 ;
        RECT 343.950 307.950 346.050 310.050 ;
        RECT 313.950 293.100 316.050 295.200 ;
        RECT 322.950 293.100 325.050 295.200 ;
        RECT 330.000 294.600 334.050 295.050 ;
        RECT 314.400 288.450 315.450 293.100 ;
        RECT 323.400 292.350 324.600 293.100 ;
        RECT 329.400 292.950 334.050 294.600 ;
        RECT 329.400 292.350 330.600 292.950 ;
        RECT 335.400 292.050 336.450 307.950 ;
        RECT 337.950 292.950 340.050 295.050 ;
        RECT 344.400 294.600 345.450 307.950 ;
        RECT 347.400 298.050 348.450 313.950 ;
        RECT 346.950 295.950 349.050 298.050 ;
        RECT 319.950 289.950 322.050 292.050 ;
        RECT 322.950 289.950 325.050 292.050 ;
        RECT 325.950 289.950 328.050 292.050 ;
        RECT 328.950 289.950 331.050 292.050 ;
        RECT 334.950 289.950 337.050 292.050 ;
        RECT 320.400 288.900 321.600 289.650 ;
        RECT 314.400 287.400 318.450 288.450 ;
        RECT 317.400 271.050 318.450 287.400 ;
        RECT 319.950 286.800 322.050 288.900 ;
        RECT 326.400 287.400 327.600 289.650 ;
        RECT 326.400 283.050 327.450 287.400 ;
        RECT 325.950 280.950 328.050 283.050 ;
        RECT 335.400 280.050 336.450 289.950 ;
        RECT 338.400 289.050 339.450 292.950 ;
        RECT 344.400 292.350 345.600 294.600 ;
        RECT 349.950 294.450 352.050 295.200 ;
        RECT 353.400 294.450 354.450 331.950 ;
        RECT 356.400 298.050 357.450 349.950 ;
        RECT 358.950 343.950 361.050 346.050 ;
        RECT 362.550 345.300 364.650 347.400 ;
        RECT 371.400 345.450 372.450 364.800 ;
        RECT 380.400 346.050 381.450 406.950 ;
        RECT 386.400 373.200 387.450 433.950 ;
        RECT 394.950 417.000 397.050 421.050 ;
        RECT 395.400 415.350 396.600 417.000 ;
        RECT 391.950 412.950 394.050 415.050 ;
        RECT 394.950 412.950 397.050 415.050 ;
        RECT 392.400 410.400 393.600 412.650 ;
        RECT 392.400 388.050 393.450 410.400 ;
        RECT 391.950 385.950 394.050 388.050 ;
        RECT 385.950 371.100 388.050 373.200 ;
        RECT 391.950 371.100 394.050 373.200 ;
        RECT 397.950 371.100 400.050 373.200 ;
        RECT 386.400 370.350 387.600 371.100 ;
        RECT 392.400 370.350 393.600 371.100 ;
        RECT 385.950 367.950 388.050 370.050 ;
        RECT 388.950 367.950 391.050 370.050 ;
        RECT 391.950 367.950 394.050 370.050 ;
        RECT 389.400 366.000 390.600 367.650 ;
        RECT 388.950 361.950 391.050 366.000 ;
        RECT 398.400 364.050 399.450 371.100 ;
        RECT 397.950 361.950 400.050 364.050 ;
        RECT 388.950 352.950 391.050 355.050 ;
        RECT 359.400 310.050 360.450 343.950 ;
        RECT 362.550 332.400 363.750 345.300 ;
        RECT 371.400 344.400 375.450 345.450 ;
        RECT 367.950 338.100 370.050 340.200 ;
        RECT 368.400 337.350 369.600 338.100 ;
        RECT 367.950 334.950 370.050 337.050 ;
        RECT 362.550 330.300 364.650 332.400 ;
        RECT 362.550 323.700 363.750 330.300 ;
        RECT 374.400 325.050 375.450 344.400 ;
        RECT 379.950 343.950 382.050 346.050 ;
        RECT 389.400 339.600 390.450 352.950 ;
        RECT 389.400 337.350 390.600 339.600 ;
        RECT 385.950 334.950 388.050 337.050 ;
        RECT 388.950 334.950 391.050 337.050 ;
        RECT 391.950 334.950 394.050 337.050 ;
        RECT 386.400 333.900 387.600 334.650 ;
        RECT 385.950 331.800 388.050 333.900 ;
        RECT 392.400 333.000 393.600 334.650 ;
        RECT 386.400 328.050 387.450 331.800 ;
        RECT 391.950 328.950 394.050 333.000 ;
        RECT 382.800 325.950 384.900 328.050 ;
        RECT 385.950 325.950 388.050 328.050 ;
        RECT 362.550 321.600 364.650 323.700 ;
        RECT 373.950 322.950 376.050 325.050 ;
        RECT 367.950 319.950 370.050 322.050 ;
        RECT 368.400 313.050 369.450 319.950 ;
        RECT 374.400 319.050 375.450 322.950 ;
        RECT 373.950 316.950 376.050 319.050 ;
        RECT 367.950 310.950 370.050 313.050 ;
        RECT 358.950 307.950 361.050 310.050 ;
        RECT 361.350 303.300 363.450 305.400 ;
        RECT 355.950 295.950 358.050 298.050 ;
        RECT 362.250 296.700 363.450 303.300 ;
        RECT 361.350 294.600 363.450 296.700 ;
        RECT 349.950 293.400 354.450 294.450 ;
        RECT 349.950 293.100 352.050 293.400 ;
        RECT 350.400 292.350 351.600 293.100 ;
        RECT 343.950 289.950 346.050 292.050 ;
        RECT 346.950 289.950 349.050 292.050 ;
        RECT 349.950 289.950 352.050 292.050 ;
        RECT 355.950 289.950 358.050 292.050 ;
        RECT 337.950 286.950 340.050 289.050 ;
        RECT 347.400 288.900 348.600 289.650 ;
        RECT 356.400 288.900 357.600 289.650 ;
        RECT 346.950 286.800 349.050 288.900 ;
        RECT 355.950 286.800 358.050 288.900 ;
        RECT 362.250 281.700 363.450 294.600 ;
        RECT 364.950 293.100 367.050 295.200 ;
        RECT 365.400 283.050 366.450 293.100 ;
        RECT 334.950 277.950 337.050 280.050 ;
        RECT 346.950 277.950 349.050 280.050 ;
        RECT 361.350 279.600 363.450 281.700 ;
        RECT 364.950 280.950 367.050 283.050 ;
        RECT 322.950 274.950 325.050 277.050 ;
        RECT 311.850 267.300 313.950 269.400 ;
        RECT 316.950 268.950 319.050 271.050 ;
        RECT 307.950 262.950 310.050 265.050 ;
        RECT 292.950 260.100 295.050 262.200 ;
        RECT 298.950 260.100 301.050 262.200 ;
        RECT 293.400 259.350 294.600 260.100 ;
        RECT 299.400 259.350 300.600 260.100 ;
        RECT 292.950 256.950 295.050 259.050 ;
        RECT 295.950 256.950 298.050 259.050 ;
        RECT 298.950 256.950 301.050 259.050 ;
        RECT 301.950 256.950 304.050 259.050 ;
        RECT 307.950 256.950 310.050 259.050 ;
        RECT 296.400 255.900 297.600 256.650 ;
        RECT 287.400 254.400 291.450 255.450 ;
        RECT 284.400 251.400 288.450 252.450 ;
        RECT 280.950 241.950 283.050 244.050 ;
        RECT 281.400 238.050 282.450 241.950 ;
        RECT 280.950 235.950 283.050 238.050 ;
        RECT 268.950 232.950 271.050 235.050 ;
        RECT 265.950 220.950 268.050 223.050 ;
        RECT 262.950 199.950 265.050 202.050 ;
        RECT 266.400 183.600 267.450 220.950 ;
        RECT 274.950 216.000 277.050 220.050 ;
        RECT 275.400 214.350 276.600 216.000 ;
        RECT 280.950 215.100 283.050 217.200 ;
        RECT 281.400 214.350 282.600 215.100 ;
        RECT 271.950 211.950 274.050 214.050 ;
        RECT 274.950 211.950 277.050 214.050 ;
        RECT 277.950 211.950 280.050 214.050 ;
        RECT 280.950 211.950 283.050 214.050 ;
        RECT 272.400 210.900 273.600 211.650 ;
        RECT 271.950 208.800 274.050 210.900 ;
        RECT 278.400 209.400 279.600 211.650 ;
        RECT 287.400 211.050 288.450 251.400 ;
        RECT 290.400 226.050 291.450 254.400 ;
        RECT 295.950 253.800 298.050 255.900 ;
        RECT 302.400 254.400 303.600 256.650 ;
        RECT 308.400 255.000 309.600 256.650 ;
        RECT 302.400 250.050 303.450 254.400 ;
        RECT 307.950 250.950 310.050 255.000 ;
        RECT 301.950 247.950 304.050 250.050 ;
        RECT 301.950 232.950 304.050 235.050 ;
        RECT 289.950 223.950 292.050 226.050 ;
        RECT 274.950 193.950 277.050 196.050 ;
        RECT 266.400 181.350 267.600 183.600 ;
        RECT 262.950 178.950 265.050 181.050 ;
        RECT 265.950 178.950 268.050 181.050 ;
        RECT 268.950 178.950 271.050 181.050 ;
        RECT 263.400 176.400 264.600 178.650 ;
        RECT 269.400 176.400 270.600 178.650 ;
        RECT 263.400 166.050 264.450 176.400 ;
        RECT 262.950 163.950 265.050 166.050 ;
        RECT 257.400 137.400 261.450 138.450 ;
        RECT 244.950 133.950 247.050 136.050 ;
        RECT 247.950 133.950 250.050 136.050 ;
        RECT 250.950 133.950 253.050 136.050 ;
        RECT 253.950 133.950 256.050 136.050 ;
        RECT 223.950 127.950 226.050 132.000 ;
        RECT 229.950 127.950 232.050 132.000 ;
        RECT 238.950 130.950 241.050 133.050 ;
        RECT 245.400 132.900 246.600 133.650 ;
        RECT 244.950 130.800 247.050 132.900 ;
        RECT 251.400 132.000 252.600 133.650 ;
        RECT 127.950 121.950 130.050 124.050 ;
        RECT 148.950 121.950 151.050 124.050 ;
        RECT 122.400 107.400 126.450 108.450 ;
        RECT 110.400 103.350 111.600 105.600 ;
        RECT 115.950 104.100 118.050 106.200 ;
        RECT 116.400 103.350 117.600 104.100 ;
        RECT 121.950 103.950 124.050 106.050 ;
        RECT 106.950 100.950 109.050 103.050 ;
        RECT 109.950 100.950 112.050 103.050 ;
        RECT 112.950 100.950 115.050 103.050 ;
        RECT 115.950 100.950 118.050 103.050 ;
        RECT 107.400 99.450 108.600 100.650 ;
        RECT 113.400 99.900 114.600 100.650 ;
        RECT 104.400 98.400 108.600 99.450 ;
        RECT 100.950 94.950 103.050 97.050 ;
        RECT 97.950 73.950 100.050 76.050 ;
        RECT 97.950 64.950 100.050 67.050 ;
        RECT 94.950 61.950 97.050 64.050 ;
        RECT 88.950 59.100 91.050 61.200 ;
        RECT 89.400 58.350 90.600 59.100 ;
        RECT 85.950 55.950 88.050 58.050 ;
        RECT 88.950 55.950 91.050 58.050 ;
        RECT 76.800 52.950 78.900 55.050 ;
        RECT 79.950 52.950 82.050 55.050 ;
        RECT 86.400 54.900 87.600 55.650 ;
        RECT 46.950 46.950 49.050 49.050 ;
        RECT 73.950 46.950 76.050 49.050 ;
        RECT 22.950 37.950 25.050 40.050 ;
        RECT 31.950 34.950 34.050 37.050 ;
        RECT 32.400 27.600 33.450 34.950 ;
        RECT 17.400 25.350 18.600 27.600 ;
        RECT 32.400 25.350 33.600 27.600 ;
        RECT 13.950 22.950 16.050 25.050 ;
        RECT 16.950 22.950 19.050 25.050 ;
        RECT 31.950 22.950 34.050 25.050 ;
        RECT 34.950 22.950 37.050 25.050 ;
        RECT 14.400 20.400 15.600 22.650 ;
        RECT 35.400 20.400 36.600 22.650 ;
        RECT 47.400 21.900 48.450 46.950 ;
        RECT 80.400 31.050 81.450 52.950 ;
        RECT 85.950 52.800 88.050 54.900 ;
        RECT 98.400 37.050 99.450 64.950 ;
        RECT 101.400 54.900 102.450 94.950 ;
        RECT 104.400 94.050 105.450 98.400 ;
        RECT 112.950 94.950 115.050 99.900 ;
        RECT 122.400 94.050 123.450 103.950 ;
        RECT 125.400 99.900 126.450 107.400 ;
        RECT 128.400 103.050 129.450 121.950 ;
        RECT 232.950 115.950 235.050 118.050 ;
        RECT 139.950 112.950 142.050 115.050 ;
        RECT 133.950 109.950 136.050 112.050 ;
        RECT 134.400 105.600 135.450 109.950 ;
        RECT 140.400 105.600 141.450 112.950 ;
        RECT 134.400 103.350 135.600 105.600 ;
        RECT 140.400 103.350 141.600 105.600 ;
        RECT 154.950 104.100 157.050 106.200 ;
        RECT 160.950 104.100 163.050 106.200 ;
        RECT 169.950 104.100 172.050 106.200 ;
        RECT 178.950 104.100 181.050 106.200 ;
        RECT 184.950 105.000 187.050 109.050 ;
        RECT 202.950 106.950 208.050 109.050 ;
        RECT 211.950 106.950 217.050 109.050 ;
        RECT 223.950 106.950 226.050 109.050 ;
        RECT 127.950 100.950 130.050 103.050 ;
        RECT 133.950 100.950 136.050 103.050 ;
        RECT 136.950 100.950 139.050 103.050 ;
        RECT 139.950 100.950 142.050 103.050 ;
        RECT 142.950 100.950 145.050 103.050 ;
        RECT 124.950 97.800 127.050 99.900 ;
        RECT 137.400 99.000 138.600 100.650 ;
        RECT 143.400 99.900 144.600 100.650 ;
        RECT 103.950 91.950 106.050 94.050 ;
        RECT 121.950 91.950 124.050 94.050 ;
        RECT 122.400 70.050 123.450 91.950 ;
        RECT 121.950 67.950 124.050 70.050 ;
        RECT 125.400 67.050 126.450 97.800 ;
        RECT 136.950 94.950 139.050 99.000 ;
        RECT 142.950 97.800 145.050 99.900 ;
        RECT 145.950 70.950 148.050 73.050 ;
        RECT 136.950 67.950 139.050 70.050 ;
        RECT 106.950 64.950 109.050 67.050 ;
        RECT 124.950 64.950 127.050 67.050 ;
        RECT 107.400 60.600 108.450 64.950 ;
        RECT 107.400 58.350 108.600 60.600 ;
        RECT 112.950 59.100 115.050 61.200 ;
        RECT 113.400 58.350 114.600 59.100 ;
        RECT 121.950 58.950 124.050 61.050 ;
        RECT 130.950 60.000 133.050 64.050 ;
        RECT 137.400 60.600 138.450 67.950 ;
        RECT 106.950 55.950 109.050 58.050 ;
        RECT 109.950 55.950 112.050 58.050 ;
        RECT 112.950 55.950 115.050 58.050 ;
        RECT 115.950 55.950 118.050 58.050 ;
        RECT 100.950 52.800 103.050 54.900 ;
        RECT 110.400 53.400 111.600 55.650 ;
        RECT 116.400 53.400 117.600 55.650 ;
        RECT 110.400 49.050 111.450 53.400 ;
        RECT 109.950 46.950 112.050 49.050 ;
        RECT 116.400 43.050 117.450 53.400 ;
        RECT 115.950 40.950 118.050 43.050 ;
        RECT 85.950 31.950 88.050 34.050 ;
        RECT 94.950 31.950 97.050 37.050 ;
        RECT 97.800 34.950 99.900 37.050 ;
        RECT 55.950 26.100 58.050 28.200 ;
        RECT 61.950 27.000 64.050 31.050 ;
        RECT 79.950 28.950 82.050 31.050 ;
        RECT 56.400 25.350 57.600 26.100 ;
        RECT 62.400 25.350 63.600 27.000 ;
        RECT 73.950 25.950 76.050 28.050 ;
        RECT 80.400 27.600 81.450 28.950 ;
        RECT 86.400 27.600 87.450 31.950 ;
        RECT 52.950 22.950 55.050 25.050 ;
        RECT 55.950 22.950 58.050 25.050 ;
        RECT 58.950 22.950 61.050 25.050 ;
        RECT 61.950 22.950 64.050 25.050 ;
        RECT 53.400 21.900 54.600 22.650 ;
        RECT 14.400 13.050 15.450 20.400 ;
        RECT 35.400 16.050 36.450 20.400 ;
        RECT 46.950 19.800 49.050 21.900 ;
        RECT 52.950 19.800 55.050 21.900 ;
        RECT 59.400 20.400 60.600 22.650 ;
        RECT 59.400 19.050 60.450 20.400 ;
        RECT 74.400 19.050 75.450 25.950 ;
        RECT 80.400 25.350 81.600 27.600 ;
        RECT 86.400 25.350 87.600 27.600 ;
        RECT 94.950 26.100 97.050 28.200 ;
        RECT 79.950 22.950 82.050 25.050 ;
        RECT 82.950 22.950 85.050 25.050 ;
        RECT 85.950 22.950 88.050 25.050 ;
        RECT 88.950 22.950 91.050 25.050 ;
        RECT 83.400 21.000 84.600 22.650 ;
        RECT 34.950 13.950 37.050 16.050 ;
        RECT 58.950 13.950 61.050 19.050 ;
        RECT 73.950 16.950 76.050 19.050 ;
        RECT 82.950 16.950 85.050 21.000 ;
        RECT 89.400 20.400 90.600 22.650 ;
        RECT 89.400 13.050 90.450 20.400 ;
        RECT 91.950 13.950 94.050 19.050 ;
        RECT 95.400 13.050 96.450 26.100 ;
        RECT 98.400 21.900 99.450 34.950 ;
        RECT 100.950 31.950 103.050 37.050 ;
        RECT 106.950 26.100 109.050 28.200 ;
        RECT 112.950 26.100 115.050 28.200 ;
        RECT 107.400 25.350 108.600 26.100 ;
        RECT 113.400 25.350 114.600 26.100 ;
        RECT 103.950 22.950 106.050 25.050 ;
        RECT 106.950 22.950 109.050 25.050 ;
        RECT 109.950 22.950 112.050 25.050 ;
        RECT 112.950 22.950 115.050 25.050 ;
        RECT 104.400 21.900 105.600 22.650 ;
        RECT 110.400 21.900 111.600 22.650 ;
        RECT 122.400 21.900 123.450 58.950 ;
        RECT 131.400 58.350 132.600 60.000 ;
        RECT 137.400 58.350 138.600 60.600 ;
        RECT 130.950 55.950 133.050 58.050 ;
        RECT 133.950 55.950 136.050 58.050 ;
        RECT 136.950 55.950 139.050 58.050 ;
        RECT 139.950 55.950 142.050 58.050 ;
        RECT 134.400 53.400 135.600 55.650 ;
        RECT 140.400 54.450 141.600 55.650 ;
        RECT 146.400 54.450 147.450 70.950 ;
        RECT 155.400 64.050 156.450 104.100 ;
        RECT 161.400 103.350 162.600 104.100 ;
        RECT 160.950 100.950 163.050 103.050 ;
        RECT 163.950 100.950 166.050 103.050 ;
        RECT 164.400 99.900 165.600 100.650 ;
        RECT 163.950 97.800 166.050 99.900 ;
        RECT 170.400 94.050 171.450 104.100 ;
        RECT 179.400 103.350 180.600 104.100 ;
        RECT 185.400 103.350 186.600 105.000 ;
        RECT 199.950 104.100 202.050 106.200 ;
        RECT 208.950 104.100 211.050 106.200 ;
        RECT 215.400 105.450 216.600 105.600 ;
        RECT 215.400 104.400 222.450 105.450 ;
        RECT 178.950 100.950 181.050 103.050 ;
        RECT 181.950 100.950 184.050 103.050 ;
        RECT 184.950 100.950 187.050 103.050 ;
        RECT 187.950 100.950 190.050 103.050 ;
        RECT 182.400 99.900 183.600 100.650 ;
        RECT 188.400 99.900 189.600 100.650 ;
        RECT 181.950 97.800 184.050 99.900 ;
        RECT 187.950 97.800 190.050 99.900 ;
        RECT 182.400 94.050 183.450 97.800 ;
        RECT 169.950 91.950 172.050 94.050 ;
        RECT 181.950 91.950 184.050 94.050 ;
        RECT 193.950 88.950 196.050 91.050 ;
        RECT 184.950 73.950 187.050 76.050 ;
        RECT 157.950 70.950 160.050 73.050 ;
        RECT 178.950 70.950 181.050 73.050 ;
        RECT 154.950 61.950 157.050 64.050 ;
        RECT 158.400 60.600 159.450 70.950 ;
        RECT 166.950 67.950 169.050 70.050 ;
        RECT 158.400 58.350 159.600 60.600 ;
        RECT 157.950 55.950 160.050 58.050 ;
        RECT 160.950 55.950 163.050 58.050 ;
        RECT 140.400 53.400 147.450 54.450 ;
        RECT 161.400 54.450 162.600 55.650 ;
        RECT 167.400 54.450 168.450 67.950 ;
        RECT 172.950 61.950 175.050 64.050 ;
        RECT 173.400 54.900 174.450 61.950 ;
        RECT 179.400 60.600 180.450 70.950 ;
        RECT 185.400 60.600 186.450 73.950 ;
        RECT 179.400 58.350 180.600 60.600 ;
        RECT 185.400 58.350 186.600 60.600 ;
        RECT 178.950 55.950 181.050 58.050 ;
        RECT 181.950 55.950 184.050 58.050 ;
        RECT 184.950 55.950 187.050 58.050 ;
        RECT 187.950 55.950 190.050 58.050 ;
        RECT 182.400 54.900 183.600 55.650 ;
        RECT 188.400 54.900 189.600 55.650 ;
        RECT 194.400 55.050 195.450 88.950 ;
        RECT 200.400 76.050 201.450 104.100 ;
        RECT 209.400 103.350 210.600 104.100 ;
        RECT 215.400 103.350 216.600 104.400 ;
        RECT 205.950 100.950 208.050 103.050 ;
        RECT 208.950 100.950 211.050 103.050 ;
        RECT 211.950 100.950 214.050 103.050 ;
        RECT 214.950 100.950 217.050 103.050 ;
        RECT 206.400 99.900 207.600 100.650 ;
        RECT 205.950 97.800 208.050 99.900 ;
        RECT 212.400 98.400 213.600 100.650 ;
        RECT 199.950 73.950 202.050 76.050 ;
        RECT 206.400 70.050 207.450 97.800 ;
        RECT 212.400 94.050 213.450 98.400 ;
        RECT 211.950 91.950 214.050 94.050 ;
        RECT 208.950 73.950 211.050 76.050 ;
        RECT 202.950 67.950 205.050 70.050 ;
        RECT 205.950 67.950 208.050 70.050 ;
        RECT 196.950 61.950 199.050 64.050 ;
        RECT 161.400 53.400 168.450 54.450 ;
        RECT 134.400 49.050 135.450 53.400 ;
        RECT 172.950 52.800 175.050 54.900 ;
        RECT 181.950 52.800 184.050 54.900 ;
        RECT 187.950 52.800 190.050 54.900 ;
        RECT 193.800 52.950 195.900 55.050 ;
        RECT 197.400 54.900 198.450 61.950 ;
        RECT 203.400 60.600 204.450 67.950 ;
        RECT 209.400 60.600 210.450 73.950 ;
        RECT 221.400 73.050 222.450 104.400 ;
        RECT 224.400 99.900 225.450 106.950 ;
        RECT 233.400 105.600 234.450 115.950 ;
        RECT 233.400 103.350 234.600 105.600 ;
        RECT 229.950 100.950 232.050 103.050 ;
        RECT 232.950 100.950 235.050 103.050 ;
        RECT 235.950 100.950 238.050 103.050 ;
        RECT 223.950 97.800 226.050 99.900 ;
        RECT 230.400 98.400 231.600 100.650 ;
        RECT 236.400 99.900 237.600 100.650 ;
        RECT 230.400 94.050 231.450 98.400 ;
        RECT 235.950 97.800 238.050 99.900 ;
        RECT 230.400 91.950 235.050 94.050 ;
        RECT 230.400 91.050 231.450 91.950 ;
        RECT 229.950 88.950 232.050 91.050 ;
        RECT 245.400 88.050 246.450 130.800 ;
        RECT 250.950 127.950 253.050 132.000 ;
        RECT 260.400 112.050 261.450 137.400 ;
        RECT 262.950 137.100 265.050 139.200 ;
        RECT 269.400 139.050 270.450 176.400 ;
        RECT 275.400 166.050 276.450 193.950 ;
        RECT 278.400 187.050 279.450 209.400 ;
        RECT 286.950 208.950 289.050 211.050 ;
        RECT 290.400 208.050 291.450 223.950 ;
        RECT 295.950 220.950 298.050 223.050 ;
        RECT 296.400 216.600 297.450 220.950 ;
        RECT 302.400 216.600 303.450 232.950 ;
        RECT 296.400 214.350 297.600 216.600 ;
        RECT 302.400 214.350 303.600 216.600 ;
        RECT 308.400 216.450 309.450 250.950 ;
        RECT 312.150 248.700 313.350 267.300 ;
        RECT 317.100 256.950 319.200 259.050 ;
        RECT 317.400 255.900 318.600 256.650 ;
        RECT 316.950 253.800 319.050 255.900 ;
        RECT 323.400 250.050 324.450 274.950 ;
        RECT 343.950 271.950 346.050 274.050 ;
        RECT 329.550 267.300 331.650 269.400 ;
        RECT 340.950 268.950 343.050 271.050 ;
        RECT 325.950 262.950 328.050 265.050 ;
        RECT 326.400 253.050 327.450 262.950 ;
        RECT 329.550 254.400 330.750 267.300 ;
        RECT 334.950 260.100 337.050 262.200 ;
        RECT 335.400 259.350 336.600 260.100 ;
        RECT 334.950 256.950 337.050 259.050 ;
        RECT 325.950 250.950 328.050 253.050 ;
        RECT 329.550 252.300 331.650 254.400 ;
        RECT 312.150 247.500 316.350 248.700 ;
        RECT 322.950 247.950 325.050 250.050 ;
        RECT 314.250 246.600 316.350 247.500 ;
        RECT 329.550 245.700 330.750 252.300 ;
        RECT 329.550 243.600 331.650 245.700 ;
        RECT 341.400 241.050 342.450 268.950 ;
        RECT 344.400 247.050 345.450 271.950 ;
        RECT 347.400 255.900 348.450 277.950 ;
        RECT 358.950 274.950 361.050 277.050 ;
        RECT 349.950 260.100 352.050 262.200 ;
        RECT 359.400 261.600 360.450 274.950 ;
        RECT 368.400 271.050 369.450 310.950 ;
        RECT 376.650 301.500 378.750 302.400 ;
        RECT 376.650 300.300 380.850 301.500 ;
        RECT 373.950 293.100 376.050 295.200 ;
        RECT 374.400 292.350 375.600 293.100 ;
        RECT 373.800 289.950 375.900 292.050 ;
        RECT 370.950 286.950 373.050 289.050 ;
        RECT 371.400 277.050 372.450 286.950 ;
        RECT 379.650 281.700 380.850 300.300 ;
        RECT 383.400 295.200 384.450 325.950 ;
        RECT 401.400 325.050 402.450 439.950 ;
        RECT 404.400 418.050 405.450 449.100 ;
        RECT 416.400 448.350 417.600 450.600 ;
        RECT 421.950 450.000 424.050 454.050 ;
        RECT 422.400 448.350 423.600 450.000 ;
        RECT 430.950 449.100 433.050 451.200 ;
        RECT 412.950 445.950 415.050 448.050 ;
        RECT 415.950 445.950 418.050 448.050 ;
        RECT 418.950 445.950 421.050 448.050 ;
        RECT 421.950 445.950 424.050 448.050 ;
        RECT 413.400 444.900 414.600 445.650 ;
        RECT 419.400 444.900 420.600 445.650 ;
        RECT 412.950 442.800 415.050 444.900 ;
        RECT 418.950 442.800 421.050 444.900 ;
        RECT 424.950 442.800 427.050 444.900 ;
        RECT 421.950 436.950 424.050 439.050 ;
        RECT 418.950 421.950 421.050 424.050 ;
        RECT 403.950 415.950 406.050 418.050 ;
        RECT 412.800 412.950 414.900 415.050 ;
        RECT 419.400 411.900 420.450 421.950 ;
        RECT 418.950 409.800 421.050 411.900 ;
        RECT 406.950 371.100 409.050 373.200 ;
        RECT 412.950 371.100 415.050 373.200 ;
        RECT 407.400 370.350 408.600 371.100 ;
        RECT 413.400 370.350 414.600 371.100 ;
        RECT 406.950 367.950 409.050 370.050 ;
        RECT 409.950 367.950 412.050 370.050 ;
        RECT 412.950 367.950 415.050 370.050 ;
        RECT 415.950 367.950 418.050 370.050 ;
        RECT 403.950 364.950 406.050 367.050 ;
        RECT 410.400 365.400 411.600 367.650 ;
        RECT 416.400 365.400 417.600 367.650 ;
        RECT 404.400 358.050 405.450 364.950 ;
        RECT 403.950 355.950 406.050 358.050 ;
        RECT 404.400 331.050 405.450 355.950 ;
        RECT 410.400 355.050 411.450 365.400 ;
        RECT 412.950 361.950 415.050 364.050 ;
        RECT 409.950 352.950 412.050 355.050 ;
        RECT 413.400 339.600 414.450 361.950 ;
        RECT 416.400 358.050 417.450 365.400 ;
        RECT 418.950 364.950 421.050 367.050 ;
        RECT 415.950 355.950 418.050 358.050 ;
        RECT 419.400 348.450 420.450 364.950 ;
        RECT 422.400 351.450 423.450 436.950 ;
        RECT 425.400 366.450 426.450 442.800 ;
        RECT 431.400 424.050 432.450 449.100 ;
        RECT 430.950 421.950 433.050 424.050 ;
        RECT 430.800 412.950 432.900 415.050 ;
        RECT 431.400 410.400 432.600 412.650 ;
        RECT 431.400 391.050 432.450 410.400 ;
        RECT 434.400 400.050 435.450 454.950 ;
        RECT 442.950 453.450 447.000 454.050 ;
        RECT 442.950 451.950 447.450 453.450 ;
        RECT 439.950 449.100 442.050 451.200 ;
        RECT 446.400 450.600 447.450 451.950 ;
        RECT 452.400 450.600 453.450 454.950 ;
        RECT 440.400 448.350 441.600 449.100 ;
        RECT 446.400 448.350 447.600 450.600 ;
        RECT 452.400 448.350 453.600 450.600 ;
        RECT 439.950 445.950 442.050 448.050 ;
        RECT 442.950 445.950 445.050 448.050 ;
        RECT 445.950 445.950 448.050 448.050 ;
        RECT 448.950 445.950 451.050 448.050 ;
        RECT 451.950 445.950 454.050 448.050 ;
        RECT 443.400 443.400 444.600 445.650 ;
        RECT 449.400 444.000 450.600 445.650 ;
        RECT 443.400 436.050 444.450 443.400 ;
        RECT 448.950 439.950 451.050 444.000 ;
        RECT 442.950 433.950 445.050 436.050 ;
        RECT 445.950 430.950 448.050 433.050 ;
        RECT 446.400 427.050 447.450 430.950 ;
        RECT 445.950 424.950 448.050 427.050 ;
        RECT 464.400 424.050 465.450 467.400 ;
        RECT 469.950 463.950 472.050 466.050 ;
        RECT 470.400 450.600 471.450 463.950 ;
        RECT 481.950 451.950 484.050 454.050 ;
        RECT 470.400 448.350 471.600 450.600 ;
        RECT 475.950 449.100 478.050 451.200 ;
        RECT 476.400 448.350 477.600 449.100 ;
        RECT 469.950 445.950 472.050 448.050 ;
        RECT 472.950 445.950 475.050 448.050 ;
        RECT 475.950 445.950 478.050 448.050 ;
        RECT 473.400 444.900 474.600 445.650 ;
        RECT 482.400 445.050 483.450 451.950 ;
        RECT 485.400 451.200 486.450 518.400 ;
        RECT 488.400 511.050 489.450 521.400 ;
        RECT 497.400 520.050 498.450 527.100 ;
        RECT 496.950 517.950 499.050 520.050 ;
        RECT 500.400 517.050 501.450 535.950 ;
        RECT 505.950 527.100 508.050 529.200 ;
        RECT 512.400 528.600 513.450 577.950 ;
        RECT 514.950 571.950 517.050 574.050 ;
        RECT 520.950 572.100 523.050 574.200 ;
        RECT 515.400 546.450 516.450 571.950 ;
        RECT 521.400 571.350 522.600 572.100 ;
        RECT 520.950 568.950 523.050 571.050 ;
        RECT 523.950 568.950 526.050 571.050 ;
        RECT 524.400 566.400 525.600 568.650 ;
        RECT 530.400 568.050 531.450 592.950 ;
        RECT 548.400 589.050 549.450 599.400 ;
        RECT 553.950 598.950 556.050 601.050 ;
        RECT 554.400 594.450 555.450 598.950 ;
        RECT 557.400 598.050 558.450 607.800 ;
        RECT 556.950 595.950 559.050 598.050 ;
        RECT 554.400 593.400 558.450 594.450 ;
        RECT 547.950 586.950 550.050 589.050 ;
        RECT 541.950 583.950 544.050 586.050 ;
        RECT 542.400 580.050 543.450 583.950 ;
        RECT 547.950 580.950 550.050 583.050 ;
        RECT 541.950 577.950 544.050 580.050 ;
        RECT 541.950 572.100 544.050 574.200 ;
        RECT 548.400 573.600 549.450 580.950 ;
        RECT 542.400 571.350 543.600 572.100 ;
        RECT 548.400 571.350 549.600 573.600 ;
        RECT 553.950 572.100 556.050 574.200 ;
        RECT 538.950 568.950 541.050 571.050 ;
        RECT 541.950 568.950 544.050 571.050 ;
        RECT 544.950 568.950 547.050 571.050 ;
        RECT 547.950 568.950 550.050 571.050 ;
        RECT 524.400 565.050 525.450 566.400 ;
        RECT 529.950 565.950 532.050 568.050 ;
        RECT 539.400 567.450 540.600 568.650 ;
        RECT 545.400 567.900 546.600 568.650 ;
        RECT 536.400 566.400 540.600 567.450 ;
        RECT 524.400 563.400 529.050 565.050 ;
        RECT 525.000 562.950 529.050 563.400 ;
        RECT 523.950 559.950 526.050 562.050 ;
        RECT 515.400 545.400 519.450 546.450 ;
        RECT 514.950 541.950 517.050 544.050 ;
        RECT 515.400 537.450 516.450 541.950 ;
        RECT 518.400 541.050 519.450 545.400 ;
        RECT 517.950 538.950 520.050 541.050 ;
        RECT 515.400 536.400 519.450 537.450 ;
        RECT 506.400 526.350 507.600 527.100 ;
        RECT 512.400 526.350 513.600 528.600 ;
        RECT 505.950 523.950 508.050 526.050 ;
        RECT 508.950 523.950 511.050 526.050 ;
        RECT 511.950 523.950 514.050 526.050 ;
        RECT 509.400 521.400 510.600 523.650 ;
        RECT 509.400 520.050 510.450 521.400 ;
        RECT 514.950 520.950 517.050 523.050 ;
        RECT 505.950 518.400 510.450 520.050 ;
        RECT 505.950 517.950 510.000 518.400 ;
        RECT 499.950 516.450 502.050 517.050 ;
        RECT 497.400 515.400 502.050 516.450 ;
        RECT 487.950 508.950 490.050 511.050 ;
        RECT 497.400 484.050 498.450 515.400 ;
        RECT 499.950 514.950 502.050 515.400 ;
        RECT 508.950 514.950 511.050 517.050 ;
        RECT 499.950 494.100 502.050 496.200 ;
        RECT 500.400 493.350 501.600 494.100 ;
        RECT 500.400 490.950 502.500 493.050 ;
        RECT 505.800 490.950 507.900 493.050 ;
        RECT 506.400 489.900 507.600 490.650 ;
        RECT 505.950 487.800 508.050 489.900 ;
        RECT 496.950 481.950 499.050 484.050 ;
        RECT 505.950 481.950 508.050 484.050 ;
        RECT 484.950 449.100 487.050 451.200 ;
        RECT 490.950 450.000 493.050 454.050 ;
        RECT 496.950 450.000 499.050 454.050 ;
        RECT 472.950 442.800 475.050 444.900 ;
        RECT 481.950 442.950 484.050 445.050 ;
        RECT 466.950 439.950 469.050 442.050 ;
        RECT 463.950 421.950 466.050 424.050 ;
        RECT 442.950 418.950 445.050 421.050 ;
        RECT 433.950 397.950 436.050 400.050 ;
        RECT 430.950 388.950 433.050 391.050 ;
        RECT 430.950 371.100 433.050 373.200 ;
        RECT 436.950 372.000 439.050 376.050 ;
        RECT 443.400 373.050 444.450 418.950 ;
        RECT 451.950 417.000 454.050 421.050 ;
        RECT 452.400 415.350 453.600 417.000 ;
        RECT 457.950 416.100 460.050 418.200 ;
        RECT 458.400 415.350 459.600 416.100 ;
        RECT 448.950 412.950 451.050 415.050 ;
        RECT 451.950 412.950 454.050 415.050 ;
        RECT 454.950 412.950 457.050 415.050 ;
        RECT 457.950 412.950 460.050 415.050 ;
        RECT 460.950 412.950 463.050 415.050 ;
        RECT 449.400 411.900 450.600 412.650 ;
        RECT 455.400 411.900 456.600 412.650 ;
        RECT 448.950 409.800 451.050 411.900 ;
        RECT 454.950 409.800 457.050 411.900 ;
        RECT 461.400 410.400 462.600 412.650 ;
        RECT 461.400 400.050 462.450 410.400 ;
        RECT 445.950 397.950 448.050 400.050 ;
        RECT 460.950 397.950 463.050 400.050 ;
        RECT 431.400 370.350 432.600 371.100 ;
        RECT 437.400 370.350 438.600 372.000 ;
        RECT 442.950 370.950 445.050 373.050 ;
        RECT 430.950 367.950 433.050 370.050 ;
        RECT 433.950 367.950 436.050 370.050 ;
        RECT 436.950 367.950 439.050 370.050 ;
        RECT 439.950 367.950 442.050 370.050 ;
        RECT 425.400 365.400 429.450 366.450 ;
        RECT 422.400 350.400 426.450 351.450 ;
        RECT 419.400 347.400 423.450 348.450 ;
        RECT 413.400 337.350 414.600 339.600 ;
        RECT 409.950 334.950 412.050 337.050 ;
        RECT 412.950 334.950 415.050 337.050 ;
        RECT 415.950 334.950 418.050 337.050 ;
        RECT 410.400 332.400 411.600 334.650 ;
        RECT 416.400 333.900 417.600 334.650 ;
        RECT 403.950 328.950 406.050 331.050 ;
        RECT 410.400 328.050 411.450 332.400 ;
        RECT 415.950 331.800 418.050 333.900 ;
        RECT 409.950 325.950 412.050 328.050 ;
        RECT 416.400 325.050 417.450 331.800 ;
        RECT 422.400 325.050 423.450 347.400 ;
        RECT 400.950 322.950 403.050 325.050 ;
        RECT 406.950 322.950 409.050 325.050 ;
        RECT 398.250 301.500 400.350 302.400 ;
        RECT 396.150 300.300 400.350 301.500 ;
        RECT 382.950 293.100 385.050 295.200 ;
        RECT 391.950 293.100 394.050 295.200 ;
        RECT 383.400 292.350 384.600 293.100 ;
        RECT 392.400 292.350 393.600 293.100 ;
        RECT 382.950 289.950 385.050 292.050 ;
        RECT 391.950 289.950 394.050 292.050 ;
        RECT 379.050 279.600 381.150 281.700 ;
        RECT 382.950 280.950 385.050 283.050 ;
        RECT 396.150 281.700 397.350 300.300 ;
        RECT 400.950 293.100 403.050 295.200 ;
        RECT 401.400 292.350 402.600 293.100 ;
        RECT 401.100 289.950 403.200 292.050 ;
        RECT 370.950 274.950 373.050 277.050 ;
        RECT 367.950 268.950 370.050 271.050 ;
        RECT 346.950 253.800 349.050 255.900 ;
        RECT 343.950 244.950 346.050 247.050 ;
        RECT 328.950 238.950 331.050 241.050 ;
        RECT 340.950 238.950 343.050 241.050 ;
        RECT 317.250 223.500 319.350 224.400 ;
        RECT 315.150 222.300 319.350 223.500 ;
        RECT 310.950 216.450 313.050 220.050 ;
        RECT 308.400 216.000 313.050 216.450 ;
        RECT 308.400 215.400 312.600 216.000 ;
        RECT 311.400 214.350 312.600 215.400 ;
        RECT 295.950 211.950 298.050 214.050 ;
        RECT 298.950 211.950 301.050 214.050 ;
        RECT 301.950 211.950 304.050 214.050 ;
        RECT 304.950 211.950 307.050 214.050 ;
        RECT 310.950 211.950 313.050 214.050 ;
        RECT 299.400 210.900 300.600 211.650 ;
        RECT 298.950 208.800 301.050 210.900 ;
        RECT 305.400 210.000 306.600 211.650 ;
        RECT 289.950 205.950 292.050 208.050 ;
        RECT 304.950 205.950 307.050 210.000 ;
        RECT 310.950 205.950 313.050 208.050 ;
        RECT 311.400 198.450 312.450 205.950 ;
        RECT 315.150 203.700 316.350 222.300 ;
        RECT 319.950 215.100 322.050 217.200 ;
        RECT 320.400 214.350 321.600 215.100 ;
        RECT 320.100 211.950 322.200 214.050 ;
        RECT 329.400 211.050 330.450 238.950 ;
        RECT 347.400 229.050 348.450 253.800 ;
        RECT 350.400 253.050 351.450 260.100 ;
        RECT 359.400 259.350 360.600 261.600 ;
        RECT 373.950 259.950 376.050 262.050 ;
        RECT 383.400 261.600 384.450 280.950 ;
        RECT 391.950 277.950 394.050 280.050 ;
        RECT 395.850 279.600 397.950 281.700 ;
        RECT 392.400 271.050 393.450 277.950 ;
        RECT 394.950 271.950 397.050 274.050 ;
        RECT 391.950 268.950 394.050 271.050 ;
        RECT 391.950 262.950 394.050 265.050 ;
        RECT 355.950 256.950 358.050 259.050 ;
        RECT 358.950 256.950 361.050 259.050 ;
        RECT 361.950 256.950 364.050 259.050 ;
        RECT 356.400 255.000 357.600 256.650 ;
        RECT 362.400 255.900 363.600 256.650 ;
        RECT 374.400 255.900 375.450 259.950 ;
        RECT 383.400 259.350 384.600 261.600 ;
        RECT 379.950 256.950 382.050 259.050 ;
        RECT 382.950 256.950 385.050 259.050 ;
        RECT 385.950 256.950 388.050 259.050 ;
        RECT 380.400 255.900 381.600 256.650 ;
        RECT 386.400 255.900 387.600 256.650 ;
        RECT 392.400 255.900 393.450 262.950 ;
        RECT 349.950 250.950 352.050 253.050 ;
        RECT 355.950 250.950 358.050 255.000 ;
        RECT 361.950 253.800 364.050 255.900 ;
        RECT 373.950 253.800 376.050 255.900 ;
        RECT 379.950 253.800 382.050 255.900 ;
        RECT 385.950 253.800 388.050 255.900 ;
        RECT 391.950 253.800 394.050 255.900 ;
        RECT 395.400 250.050 396.450 271.950 ;
        RECT 407.400 265.050 408.450 322.950 ;
        RECT 409.950 322.800 412.050 324.900 ;
        RECT 415.950 322.950 418.050 325.050 ;
        RECT 421.950 322.950 424.050 325.050 ;
        RECT 410.400 276.450 411.450 322.800 ;
        RECT 413.550 303.300 415.650 305.400 ;
        RECT 413.550 296.700 414.750 303.300 ;
        RECT 413.550 294.600 415.650 296.700 ;
        RECT 413.550 281.700 414.750 294.600 ;
        RECT 418.950 289.950 421.050 292.050 ;
        RECT 419.400 288.000 420.600 289.650 ;
        RECT 418.950 283.950 421.050 288.000 ;
        RECT 425.400 286.050 426.450 350.400 ;
        RECT 424.950 283.950 427.050 286.050 ;
        RECT 413.550 279.600 415.650 281.700 ;
        RECT 421.950 277.950 424.050 280.050 ;
        RECT 410.400 275.400 414.450 276.450 ;
        RECT 406.950 262.950 409.050 265.050 ;
        RECT 403.950 260.100 406.050 262.200 ;
        RECT 404.400 259.350 405.600 260.100 ;
        RECT 400.950 256.950 403.050 259.050 ;
        RECT 403.950 256.950 406.050 259.050 ;
        RECT 406.950 256.950 409.050 259.050 ;
        RECT 407.400 254.400 408.600 256.650 ;
        RECT 413.400 255.450 414.450 275.400 ;
        RECT 422.400 262.050 423.450 277.950 ;
        RECT 428.400 274.050 429.450 365.400 ;
        RECT 434.400 365.400 435.600 367.650 ;
        RECT 440.400 365.400 441.600 367.650 ;
        RECT 434.400 355.050 435.450 365.400 ;
        RECT 433.950 352.950 436.050 355.050 ;
        RECT 430.950 338.100 433.050 340.200 ;
        RECT 431.400 337.350 432.600 338.100 ;
        RECT 431.400 334.950 433.500 337.050 ;
        RECT 436.800 334.950 438.900 337.050 ;
        RECT 437.400 333.900 438.600 334.650 ;
        RECT 436.950 333.450 439.050 333.900 ;
        RECT 440.400 333.450 441.450 365.400 ;
        RECT 446.400 333.900 447.450 397.950 ;
        RECT 467.400 397.050 468.450 439.950 ;
        RECT 485.400 439.050 486.450 449.100 ;
        RECT 491.400 448.350 492.600 450.000 ;
        RECT 497.400 448.350 498.600 450.000 ;
        RECT 490.950 445.950 493.050 448.050 ;
        RECT 493.950 445.950 496.050 448.050 ;
        RECT 496.950 445.950 499.050 448.050 ;
        RECT 499.950 445.950 502.050 448.050 ;
        RECT 494.400 444.900 495.600 445.650 ;
        RECT 493.950 442.800 496.050 444.900 ;
        RECT 500.400 443.400 501.600 445.650 ;
        RECT 500.400 441.450 501.450 443.400 ;
        RECT 494.400 440.400 501.450 441.450 ;
        RECT 494.400 439.050 495.450 440.400 ;
        RECT 484.950 436.950 487.050 439.050 ;
        RECT 493.950 436.950 496.050 439.050 ;
        RECT 487.950 427.950 490.050 430.050 ;
        RECT 469.950 421.950 472.050 424.050 ;
        RECT 466.950 394.950 469.050 397.050 ;
        RECT 470.400 388.050 471.450 421.950 ;
        RECT 472.950 416.100 475.050 418.200 ;
        RECT 481.950 416.100 484.050 418.200 ;
        RECT 473.400 406.050 474.450 416.100 ;
        RECT 482.400 415.350 483.600 416.100 ;
        RECT 476.100 412.950 478.200 415.050 ;
        RECT 481.500 412.950 483.600 415.050 ;
        RECT 476.400 411.900 477.600 412.650 ;
        RECT 475.950 409.800 478.050 411.900 ;
        RECT 472.950 403.950 475.050 406.050 ;
        RECT 481.950 400.950 484.050 403.050 ;
        RECT 475.950 394.950 478.050 397.050 ;
        RECT 448.950 385.950 451.050 388.050 ;
        RECT 469.950 385.950 472.050 388.050 ;
        RECT 449.400 340.200 450.450 385.950 ;
        RECT 469.350 381.300 471.450 383.400 ;
        RECT 451.950 375.450 456.000 376.050 ;
        RECT 451.950 373.950 456.450 375.450 ;
        RECT 470.250 374.700 471.450 381.300 ;
        RECT 472.950 379.950 475.050 382.050 ;
        RECT 455.400 372.600 456.450 373.950 ;
        RECT 469.350 372.600 471.450 374.700 ;
        RECT 455.400 370.350 456.600 372.600 ;
        RECT 454.950 367.950 457.050 370.050 ;
        RECT 457.950 367.950 460.050 370.050 ;
        RECT 463.950 367.950 466.050 370.050 ;
        RECT 458.400 366.900 459.600 367.650 ;
        RECT 464.400 366.900 465.600 367.650 ;
        RECT 457.950 364.800 460.050 366.900 ;
        RECT 463.950 364.800 466.050 366.900 ;
        RECT 454.950 358.950 457.050 361.050 ;
        RECT 470.250 359.700 471.450 372.600 ;
        RECT 473.400 361.050 474.450 379.950 ;
        RECT 448.950 338.100 451.050 340.200 ;
        RECT 455.400 339.600 456.450 358.950 ;
        RECT 469.350 357.600 471.450 359.700 ;
        RECT 472.950 358.950 475.050 361.050 ;
        RECT 472.950 352.950 475.050 355.050 ;
        RECT 473.400 348.450 474.450 352.950 ;
        RECT 476.400 352.050 477.450 394.950 ;
        RECT 482.400 388.050 483.450 400.950 ;
        RECT 488.400 400.050 489.450 427.950 ;
        RECT 494.400 412.050 495.450 436.950 ;
        RECT 496.950 421.950 499.050 424.050 ;
        RECT 497.400 417.600 498.450 421.950 ;
        RECT 506.400 418.200 507.450 481.950 ;
        RECT 509.400 472.050 510.450 514.950 ;
        RECT 511.950 502.950 514.050 505.050 ;
        RECT 512.400 496.200 513.450 502.950 ;
        RECT 511.950 494.100 514.050 496.200 ;
        RECT 512.400 490.050 513.450 494.100 ;
        RECT 511.950 487.950 514.050 490.050 ;
        RECT 511.950 478.950 514.050 481.050 ;
        RECT 508.950 469.950 511.050 472.050 ;
        RECT 497.400 415.350 498.600 417.600 ;
        RECT 505.950 416.100 508.050 418.200 ;
        RECT 497.400 412.950 499.500 415.050 ;
        RECT 502.800 412.950 504.900 415.050 ;
        RECT 493.950 409.950 496.050 412.050 ;
        RECT 503.400 411.900 504.600 412.650 ;
        RECT 502.950 409.800 505.050 411.900 ;
        RECT 509.400 409.050 510.450 469.950 ;
        RECT 512.400 463.050 513.450 478.950 ;
        RECT 511.950 460.950 514.050 463.050 ;
        RECT 515.400 460.050 516.450 520.950 ;
        RECT 518.400 469.050 519.450 536.400 ;
        RECT 520.950 535.950 523.050 538.050 ;
        RECT 521.400 517.050 522.450 535.950 ;
        RECT 524.400 529.050 525.450 559.950 ;
        RECT 532.950 553.950 535.050 556.050 ;
        RECT 533.400 550.050 534.450 553.950 ;
        RECT 532.950 547.950 535.050 550.050 ;
        RECT 536.400 544.050 537.450 566.400 ;
        RECT 538.950 562.950 541.050 565.050 ;
        RECT 544.950 562.950 547.050 567.900 ;
        RECT 550.950 562.950 553.050 568.050 ;
        RECT 539.400 559.050 540.450 562.950 ;
        RECT 538.950 556.950 541.050 559.050 ;
        RECT 554.400 556.050 555.450 572.100 ;
        RECT 557.400 558.450 558.450 593.400 ;
        RECT 560.400 592.050 561.450 613.950 ;
        RECT 563.400 600.450 564.450 619.950 ;
        RECT 575.400 616.050 576.450 683.100 ;
        RECT 578.400 667.050 579.450 691.950 ;
        RECT 587.400 685.200 588.450 706.950 ;
        RECT 593.400 694.050 594.450 733.950 ;
        RECT 596.400 723.900 597.450 743.400 ;
        RECT 598.950 742.950 601.050 743.400 ;
        RECT 605.400 736.050 606.450 790.950 ;
        RECT 611.400 784.050 612.450 790.950 ;
        RECT 610.950 781.950 613.050 784.050 ;
        RECT 614.400 765.450 615.450 829.950 ;
        RECT 625.950 826.950 628.050 829.050 ;
        RECT 626.400 813.450 627.450 826.950 ;
        RECT 619.500 809.400 621.600 811.500 ;
        RECT 626.400 811.200 627.600 813.450 ;
        RECT 617.100 802.950 619.200 805.050 ;
        RECT 617.400 801.900 618.600 802.650 ;
        RECT 616.950 799.800 619.050 801.900 ;
        RECT 620.100 796.800 621.000 809.400 ;
        RECT 626.100 808.800 628.200 810.900 ;
        RECT 629.400 809.100 631.500 811.200 ;
        RECT 621.900 807.000 624.000 807.900 ;
        RECT 621.900 805.800 629.100 807.000 ;
        RECT 627.000 804.900 629.100 805.800 ;
        RECT 621.900 804.000 624.000 804.900 ;
        RECT 630.000 804.000 630.900 809.100 ;
        RECT 631.950 806.100 634.050 808.200 ;
        RECT 632.400 805.350 633.600 806.100 ;
        RECT 621.900 803.100 630.900 804.000 ;
        RECT 621.900 802.800 624.000 803.100 ;
        RECT 626.100 799.950 628.200 802.050 ;
        RECT 626.400 797.400 627.600 799.650 ;
        RECT 619.800 794.700 621.900 796.800 ;
        RECT 630.000 796.500 630.900 803.100 ;
        RECT 631.800 802.950 633.900 805.050 ;
        RECT 634.950 796.950 637.050 799.050 ;
        RECT 628.800 794.400 630.900 796.500 ;
        RECT 628.950 787.950 631.050 790.050 ;
        RECT 619.950 781.950 622.050 784.050 ;
        RECT 620.400 778.050 621.450 781.950 ;
        RECT 619.950 775.950 622.050 778.050 ;
        RECT 622.950 772.950 625.050 775.050 ;
        RECT 623.400 769.050 624.450 772.950 ;
        RECT 622.950 766.950 625.050 769.050 ;
        RECT 611.400 764.400 615.450 765.450 ;
        RECT 607.950 754.950 610.050 757.050 ;
        RECT 608.400 742.050 609.450 754.950 ;
        RECT 607.950 739.950 610.050 742.050 ;
        RECT 611.400 736.050 612.450 764.400 ;
        RECT 613.950 761.100 616.050 763.200 ;
        RECT 623.400 762.600 624.450 766.950 ;
        RECT 614.400 760.350 615.600 761.100 ;
        RECT 623.400 760.350 624.600 762.600 ;
        RECT 614.100 757.950 616.200 760.050 ;
        RECT 617.400 757.950 619.500 760.050 ;
        RECT 622.800 757.950 624.900 760.050 ;
        RECT 617.400 755.400 618.600 757.650 ;
        RECT 617.400 745.050 618.450 755.400 ;
        RECT 629.400 754.050 630.450 787.950 ;
        RECT 631.950 769.950 634.050 772.050 ;
        RECT 628.950 751.950 631.050 754.050 ;
        RECT 616.950 742.950 619.050 745.050 ;
        RECT 604.950 733.950 607.050 736.050 ;
        RECT 610.950 733.950 613.050 736.050 ;
        RECT 616.950 733.950 619.050 736.050 ;
        RECT 604.950 728.100 607.050 730.200 ;
        RECT 610.950 728.100 613.050 730.200 ;
        RECT 605.400 727.350 606.600 728.100 ;
        RECT 611.400 727.350 612.600 728.100 ;
        RECT 601.950 724.950 604.050 727.050 ;
        RECT 604.950 724.950 607.050 727.050 ;
        RECT 607.950 724.950 610.050 727.050 ;
        RECT 610.950 724.950 613.050 727.050 ;
        RECT 602.400 723.900 603.600 724.650 ;
        RECT 595.950 721.800 598.050 723.900 ;
        RECT 601.950 721.800 604.050 723.900 ;
        RECT 608.400 722.400 609.600 724.650 ;
        RECT 604.950 706.950 607.050 709.050 ;
        RECT 592.950 691.950 595.050 694.050 ;
        RECT 586.950 683.100 589.050 685.200 ;
        RECT 592.950 683.100 595.050 685.200 ;
        RECT 601.950 683.100 604.050 685.200 ;
        RECT 587.400 682.350 588.600 683.100 ;
        RECT 593.400 682.350 594.600 683.100 ;
        RECT 583.950 679.950 586.050 682.050 ;
        RECT 586.950 679.950 589.050 682.050 ;
        RECT 589.950 679.950 592.050 682.050 ;
        RECT 592.950 679.950 595.050 682.050 ;
        RECT 595.950 679.950 598.050 682.050 ;
        RECT 580.950 676.950 583.050 679.050 ;
        RECT 584.400 677.400 585.600 679.650 ;
        RECT 590.400 678.900 591.600 679.650 ;
        RECT 577.950 664.950 580.050 667.050 ;
        RECT 581.400 631.050 582.450 676.950 ;
        RECT 584.400 658.050 585.450 677.400 ;
        RECT 589.950 676.800 592.050 678.900 ;
        RECT 596.400 678.450 597.600 679.650 ;
        RECT 596.400 677.400 600.450 678.450 ;
        RECT 599.400 664.050 600.450 677.400 ;
        RECT 598.950 661.950 601.050 664.050 ;
        RECT 583.950 655.950 586.050 658.050 ;
        RECT 599.400 652.200 600.450 661.950 ;
        RECT 589.950 650.100 592.050 652.200 ;
        RECT 598.950 650.100 601.050 652.200 ;
        RECT 590.400 649.350 591.600 650.100 ;
        RECT 586.950 646.950 589.050 649.050 ;
        RECT 589.950 646.950 592.050 649.050 ;
        RECT 587.400 644.400 588.600 646.650 ;
        RECT 587.400 634.050 588.450 644.400 ;
        RECT 592.950 643.800 595.050 645.900 ;
        RECT 586.950 631.950 589.050 634.050 ;
        RECT 580.950 628.950 583.050 631.050 ;
        RECT 583.950 616.950 586.050 619.050 ;
        RECT 574.950 613.950 577.050 616.050 ;
        RECT 568.950 610.950 571.050 613.050 ;
        RECT 569.400 607.200 570.450 610.950 ;
        RECT 574.950 610.800 577.050 612.900 ;
        RECT 568.950 605.100 571.050 607.200 ;
        RECT 575.400 606.600 576.450 610.800 ;
        RECT 580.950 607.950 583.050 610.050 ;
        RECT 569.400 604.350 570.600 605.100 ;
        RECT 575.400 604.350 576.600 606.600 ;
        RECT 568.950 601.950 571.050 604.050 ;
        RECT 571.950 601.950 574.050 604.050 ;
        RECT 574.950 601.950 577.050 604.050 ;
        RECT 563.400 599.400 567.450 600.450 ;
        RECT 572.400 600.000 573.600 601.650 ;
        RECT 559.950 589.950 562.050 592.050 ;
        RECT 566.400 573.600 567.450 599.400 ;
        RECT 571.950 595.950 574.050 600.000 ;
        RECT 581.400 597.450 582.450 607.950 ;
        RECT 584.400 601.050 585.450 616.950 ;
        RECT 586.950 610.950 589.050 616.050 ;
        RECT 593.400 613.050 594.450 643.800 ;
        RECT 599.400 616.050 600.450 650.100 ;
        RECT 598.950 613.950 601.050 616.050 ;
        RECT 592.950 610.950 595.050 613.050 ;
        RECT 587.400 607.050 588.450 610.950 ;
        RECT 586.950 604.950 589.050 607.050 ;
        RECT 589.950 606.000 592.050 610.050 ;
        RECT 590.400 604.350 591.600 606.000 ;
        RECT 595.950 605.100 598.050 607.200 ;
        RECT 596.400 604.350 597.600 605.100 ;
        RECT 589.950 601.950 592.050 604.050 ;
        RECT 592.950 601.950 595.050 604.050 ;
        RECT 595.950 601.950 598.050 604.050 ;
        RECT 583.950 598.950 586.050 601.050 ;
        RECT 593.400 600.900 594.600 601.650 ;
        RECT 592.950 598.800 595.050 600.900 ;
        RECT 578.400 596.400 582.450 597.450 ;
        RECT 574.950 589.950 577.050 592.050 ;
        RECT 566.400 571.350 567.600 573.600 ;
        RECT 562.950 568.950 565.050 571.050 ;
        RECT 565.950 568.950 568.050 571.050 ;
        RECT 568.950 568.950 571.050 571.050 ;
        RECT 563.400 567.000 564.600 568.650 ;
        RECT 569.400 567.900 570.600 568.650 ;
        RECT 562.950 562.950 565.050 567.000 ;
        RECT 568.950 565.800 571.050 567.900 ;
        RECT 571.950 565.950 574.050 568.050 ;
        RECT 559.950 558.450 562.050 559.050 ;
        RECT 557.400 557.400 562.050 558.450 ;
        RECT 559.950 556.950 562.050 557.400 ;
        RECT 553.950 553.950 556.050 556.050 ;
        RECT 560.400 544.050 561.450 556.950 ;
        RECT 562.950 550.950 565.050 553.050 ;
        RECT 535.950 541.950 538.050 544.050 ;
        RECT 559.950 541.950 562.050 544.050 ;
        RECT 563.400 541.050 564.450 550.950 ;
        RECT 541.350 537.300 543.450 539.400 ;
        RECT 562.950 538.950 565.050 541.050 ;
        RECT 526.950 532.950 529.050 535.050 ;
        RECT 523.950 526.950 526.050 529.050 ;
        RECT 527.400 528.600 528.450 532.950 ;
        RECT 542.250 530.700 543.450 537.300 ;
        RECT 556.650 535.500 558.750 536.400 ;
        RECT 556.650 534.300 560.850 535.500 ;
        RECT 541.350 528.600 543.450 530.700 ;
        RECT 527.400 526.350 528.600 528.600 ;
        RECT 526.950 523.950 529.050 526.050 ;
        RECT 529.950 523.950 532.050 526.050 ;
        RECT 535.950 523.950 538.050 526.050 ;
        RECT 530.400 522.450 531.600 523.650 ;
        RECT 536.400 522.450 537.600 523.650 ;
        RECT 530.400 521.400 537.600 522.450 ;
        RECT 520.950 514.950 523.050 517.050 ;
        RECT 542.250 515.700 543.450 528.600 ;
        RECT 547.950 526.950 550.050 529.050 ;
        RECT 553.950 527.100 556.050 529.200 ;
        RECT 535.950 511.950 538.050 514.050 ;
        RECT 541.350 513.600 543.450 515.700 ;
        RECT 529.950 494.100 532.050 496.200 ;
        RECT 530.400 493.350 531.600 494.100 ;
        RECT 523.800 490.950 525.900 493.050 ;
        RECT 529.800 490.950 531.900 493.050 ;
        RECT 524.400 488.400 525.600 490.650 ;
        RECT 524.400 484.050 525.450 488.400 ;
        RECT 523.950 481.950 526.050 484.050 ;
        RECT 517.950 466.950 520.050 469.050 ;
        RECT 514.950 457.950 517.050 460.050 ;
        RECT 520.950 457.950 523.050 460.050 ;
        RECT 529.350 459.300 531.450 461.400 ;
        RECT 511.950 453.450 516.000 454.050 ;
        RECT 511.950 451.950 516.450 453.450 ;
        RECT 515.400 450.600 516.450 451.950 ;
        RECT 521.400 451.050 522.450 457.950 ;
        RECT 530.250 452.700 531.450 459.300 ;
        RECT 515.400 448.350 516.600 450.600 ;
        RECT 520.950 448.950 523.050 451.050 ;
        RECT 529.350 450.600 531.450 452.700 ;
        RECT 514.950 445.950 517.050 448.050 ;
        RECT 517.950 445.950 520.050 448.050 ;
        RECT 523.950 445.950 526.050 448.050 ;
        RECT 511.950 442.950 514.050 445.050 ;
        RECT 518.400 444.900 519.600 445.650 ;
        RECT 524.400 444.900 525.600 445.650 ;
        RECT 508.950 406.950 511.050 409.050 ;
        RECT 487.950 397.950 490.050 400.050 ;
        RECT 512.400 394.050 513.450 442.950 ;
        RECT 517.950 442.800 520.050 444.900 ;
        RECT 523.950 442.800 526.050 444.900 ;
        RECT 518.400 436.050 519.450 442.800 ;
        RECT 530.250 437.700 531.450 450.600 ;
        RECT 536.400 439.050 537.450 511.950 ;
        RECT 548.400 511.050 549.450 526.950 ;
        RECT 554.400 526.350 555.600 527.100 ;
        RECT 553.800 523.950 555.900 526.050 ;
        RECT 559.650 515.700 560.850 534.300 ;
        RECT 568.950 532.950 571.050 535.050 ;
        RECT 563.400 528.450 564.600 528.600 ;
        RECT 569.400 528.450 570.450 532.950 ;
        RECT 563.400 527.400 570.450 528.450 ;
        RECT 563.400 526.350 564.600 527.400 ;
        RECT 562.950 523.950 565.050 526.050 ;
        RECT 569.400 522.450 570.450 527.400 ;
        RECT 566.400 521.400 570.450 522.450 ;
        RECT 559.050 513.600 561.150 515.700 ;
        RECT 566.400 511.050 567.450 521.400 ;
        RECT 572.400 517.050 573.450 565.950 ;
        RECT 575.400 550.050 576.450 589.950 ;
        RECT 578.400 565.050 579.450 596.400 ;
        RECT 583.950 595.800 586.050 597.900 ;
        RECT 580.950 592.950 583.050 595.050 ;
        RECT 577.950 562.950 580.050 565.050 ;
        RECT 581.400 562.050 582.450 592.950 ;
        RECT 584.400 574.050 585.450 595.800 ;
        RECT 602.400 595.050 603.450 683.100 ;
        RECT 605.400 679.050 606.450 706.950 ;
        RECT 608.400 685.050 609.450 722.400 ;
        RECT 610.950 691.950 613.050 694.050 ;
        RECT 607.950 682.950 610.050 685.050 ;
        RECT 611.400 684.600 612.450 691.950 ;
        RECT 617.400 688.200 618.450 733.950 ;
        RECT 619.950 728.100 622.050 730.200 ;
        RECT 625.950 728.100 628.050 730.200 ;
        RECT 632.400 729.600 633.450 769.950 ;
        RECT 635.400 733.050 636.450 796.950 ;
        RECT 638.400 790.050 639.450 874.950 ;
        RECT 644.400 874.050 645.450 878.400 ;
        RECT 649.950 877.800 652.050 879.900 ;
        RECT 643.950 871.950 646.050 874.050 ;
        RECT 656.400 871.050 657.450 901.950 ;
        RECT 704.400 901.050 705.450 917.100 ;
        RECT 713.400 916.350 714.600 917.100 ;
        RECT 719.400 916.350 720.600 918.000 ;
        RECT 709.950 913.950 712.050 916.050 ;
        RECT 712.950 913.950 715.050 916.050 ;
        RECT 715.950 913.950 718.050 916.050 ;
        RECT 718.950 913.950 721.050 916.050 ;
        RECT 710.400 912.900 711.600 913.650 ;
        RECT 709.950 910.800 712.050 912.900 ;
        RECT 716.400 911.400 717.600 913.650 ;
        RECT 716.400 907.050 717.450 911.400 ;
        RECT 728.400 907.050 729.450 934.950 ;
        RECT 731.400 922.050 732.450 955.800 ;
        RECT 733.950 931.950 736.050 934.050 ;
        RECT 734.400 922.050 735.450 931.950 ;
        RECT 737.400 925.050 738.450 955.800 ;
        RECT 751.950 952.950 754.050 955.050 ;
        RECT 760.950 952.950 763.050 957.000 ;
        RECT 779.400 956.400 780.600 958.650 ;
        RECT 785.400 957.900 786.600 958.650 ;
        RECT 794.400 957.900 795.450 961.950 ;
        RECT 803.400 961.350 804.600 962.100 ;
        RECT 809.400 961.350 810.600 963.000 ;
        RECT 802.950 958.950 805.050 961.050 ;
        RECT 805.950 958.950 808.050 961.050 ;
        RECT 808.950 958.950 811.050 961.050 ;
        RECT 811.950 958.950 814.050 961.050 ;
        RECT 742.950 943.950 745.050 946.050 ;
        RECT 736.950 922.950 739.050 925.050 ;
        RECT 730.950 919.950 733.050 922.050 ;
        RECT 733.950 919.950 736.050 922.050 ;
        RECT 736.950 917.100 739.050 919.200 ;
        RECT 743.400 918.600 744.450 943.950 ;
        RECT 748.950 925.950 751.050 928.050 ;
        RECT 737.400 916.350 738.600 917.100 ;
        RECT 743.400 916.350 744.600 918.600 ;
        RECT 733.950 913.950 736.050 916.050 ;
        RECT 736.950 913.950 739.050 916.050 ;
        RECT 739.950 913.950 742.050 916.050 ;
        RECT 742.950 913.950 745.050 916.050 ;
        RECT 734.400 912.900 735.600 913.650 ;
        RECT 733.950 910.800 736.050 912.900 ;
        RECT 740.400 911.400 741.600 913.650 ;
        RECT 740.400 907.050 741.450 911.400 ;
        RECT 742.950 907.950 745.050 910.050 ;
        RECT 715.950 904.950 718.050 907.050 ;
        RECT 727.950 904.950 730.050 907.050 ;
        RECT 739.950 904.950 742.050 907.050 ;
        RECT 703.950 898.950 706.050 901.050 ;
        RECT 664.950 895.950 667.050 898.050 ;
        RECT 665.400 892.050 666.450 895.950 ;
        RECT 727.950 892.950 730.050 895.050 ;
        RECT 664.950 889.950 667.050 892.050 ;
        RECT 712.950 889.950 715.050 892.050 ;
        RECT 665.400 885.600 666.450 889.950 ;
        RECT 665.400 883.350 666.600 885.600 ;
        RECT 700.950 884.100 703.050 886.200 ;
        RECT 713.400 885.600 714.450 889.950 ;
        RECT 664.950 880.950 667.050 883.050 ;
        RECT 667.950 880.950 670.050 883.050 ;
        RECT 683.100 880.950 685.200 883.050 ;
        RECT 686.400 880.950 688.500 883.050 ;
        RECT 691.800 880.950 693.900 883.050 ;
        RECT 668.400 879.900 669.600 880.650 ;
        RECT 667.950 877.800 670.050 879.900 ;
        RECT 683.400 878.400 684.600 880.650 ;
        RECT 692.400 878.400 693.600 880.650 ;
        RECT 679.950 874.950 682.050 877.050 ;
        RECT 655.950 868.950 658.050 871.050 ;
        RECT 640.950 847.950 643.050 850.050 ;
        RECT 641.400 835.050 642.450 847.950 ;
        RECT 649.950 839.100 652.050 841.200 ;
        RECT 664.950 839.100 667.050 841.200 ;
        RECT 670.950 839.100 673.050 841.200 ;
        RECT 676.950 839.100 679.050 841.200 ;
        RECT 650.400 838.350 651.600 839.100 ;
        RECT 665.400 838.350 666.600 839.100 ;
        RECT 671.400 838.350 672.600 839.100 ;
        RECT 646.950 835.950 649.050 838.050 ;
        RECT 649.950 835.950 652.050 838.050 ;
        RECT 664.950 835.950 667.050 838.050 ;
        RECT 667.950 835.950 670.050 838.050 ;
        RECT 670.950 835.950 673.050 838.050 ;
        RECT 640.950 832.950 643.050 835.050 ;
        RECT 647.400 833.400 648.600 835.650 ;
        RECT 668.400 833.400 669.600 835.650 ;
        RECT 647.400 829.050 648.450 833.400 ;
        RECT 640.950 826.950 643.050 829.050 ;
        RECT 646.950 826.950 649.050 829.050 ;
        RECT 664.950 826.950 667.050 829.050 ;
        RECT 641.400 801.900 642.450 826.950 ;
        RECT 655.950 823.950 658.050 826.050 ;
        RECT 656.400 820.050 657.450 823.950 ;
        RECT 655.950 817.950 658.050 820.050 ;
        RECT 649.950 806.100 652.050 808.200 ;
        RECT 656.400 807.600 657.450 817.950 ;
        RECT 650.400 805.350 651.600 806.100 ;
        RECT 656.400 805.350 657.600 807.600 ;
        RECT 661.950 806.100 664.050 808.200 ;
        RECT 646.950 802.950 649.050 805.050 ;
        RECT 649.950 802.950 652.050 805.050 ;
        RECT 652.950 802.950 655.050 805.050 ;
        RECT 655.950 802.950 658.050 805.050 ;
        RECT 647.400 801.900 648.600 802.650 ;
        RECT 653.400 801.900 654.600 802.650 ;
        RECT 640.950 799.800 643.050 801.900 ;
        RECT 646.950 799.800 649.050 801.900 ;
        RECT 652.950 799.800 655.050 801.900 ;
        RECT 637.950 787.950 640.050 790.050 ;
        RECT 649.950 781.950 652.050 784.050 ;
        RECT 650.400 769.050 651.450 781.950 ;
        RECT 653.400 781.050 654.450 799.800 ;
        RECT 662.400 790.050 663.450 806.100 ;
        RECT 661.950 787.950 664.050 790.050 ;
        RECT 652.950 778.950 655.050 781.050 ;
        RECT 649.950 766.950 652.050 769.050 ;
        RECT 643.950 761.100 646.050 763.200 ;
        RECT 649.950 761.100 652.050 763.200 ;
        RECT 644.400 760.350 645.600 761.100 ;
        RECT 650.400 760.350 651.600 761.100 ;
        RECT 640.950 757.950 643.050 760.050 ;
        RECT 643.950 757.950 646.050 760.050 ;
        RECT 646.950 757.950 649.050 760.050 ;
        RECT 649.950 757.950 652.050 760.050 ;
        RECT 641.400 756.000 642.600 757.650 ;
        RECT 647.400 756.900 648.600 757.650 ;
        RECT 640.950 751.950 643.050 756.000 ;
        RECT 646.950 754.800 649.050 756.900 ;
        RECT 662.400 756.450 663.450 787.950 ;
        RECT 665.400 778.050 666.450 826.950 ;
        RECT 668.400 820.050 669.450 833.400 ;
        RECT 673.950 832.950 676.050 835.050 ;
        RECT 667.950 817.950 670.050 820.050 ;
        RECT 674.400 807.600 675.450 832.950 ;
        RECT 677.400 829.050 678.450 839.100 ;
        RECT 680.400 829.050 681.450 874.950 ;
        RECT 683.400 865.050 684.450 878.400 ;
        RECT 682.950 862.950 685.050 865.050 ;
        RECT 683.400 847.050 684.450 862.950 ;
        RECT 692.400 859.050 693.450 878.400 ;
        RECT 685.950 856.950 688.050 859.050 ;
        RECT 691.950 856.950 694.050 859.050 ;
        RECT 682.950 844.950 685.050 847.050 ;
        RECT 686.400 840.450 687.450 856.950 ;
        RECT 694.950 847.950 697.050 850.050 ;
        RECT 695.400 844.200 696.450 847.950 ;
        RECT 701.400 847.050 702.450 884.100 ;
        RECT 713.400 883.350 714.600 885.600 ;
        RECT 718.950 884.100 721.050 886.200 ;
        RECT 719.400 883.350 720.600 884.100 ;
        RECT 709.950 880.950 712.050 883.050 ;
        RECT 712.950 880.950 715.050 883.050 ;
        RECT 715.950 880.950 718.050 883.050 ;
        RECT 718.950 880.950 721.050 883.050 ;
        RECT 710.400 879.000 711.600 880.650 ;
        RECT 709.950 874.950 712.050 879.000 ;
        RECT 716.400 878.400 717.600 880.650 ;
        RECT 710.400 871.050 711.450 874.950 ;
        RECT 709.950 868.950 712.050 871.050 ;
        RECT 709.950 853.950 712.050 856.050 ;
        RECT 700.950 844.950 703.050 847.050 ;
        RECT 694.950 842.100 697.050 844.200 ;
        RECT 683.400 839.400 687.450 840.450 ;
        RECT 676.800 826.950 678.900 829.050 ;
        RECT 679.950 826.950 682.050 829.050 ;
        RECT 674.400 805.350 675.600 807.600 ;
        RECT 670.950 802.950 673.050 805.050 ;
        RECT 673.950 802.950 676.050 805.050 ;
        RECT 676.950 802.950 679.050 805.050 ;
        RECT 671.400 801.900 672.600 802.650 ;
        RECT 670.950 799.800 673.050 801.900 ;
        RECT 677.400 800.400 678.600 802.650 ;
        RECT 677.400 790.050 678.450 800.400 ;
        RECT 676.950 787.950 679.050 790.050 ;
        RECT 683.400 787.050 684.450 839.400 ;
        RECT 688.950 839.100 691.050 841.200 ;
        RECT 689.400 838.350 690.600 839.100 ;
        RECT 694.950 838.950 697.050 841.050 ;
        RECT 695.400 838.350 696.600 838.950 ;
        RECT 688.950 835.950 691.050 838.050 ;
        RECT 691.950 835.950 694.050 838.050 ;
        RECT 694.950 835.950 697.050 838.050 ;
        RECT 692.400 833.400 693.600 835.650 ;
        RECT 688.950 829.950 691.050 832.050 ;
        RECT 689.400 817.050 690.450 829.950 ;
        RECT 692.400 829.050 693.450 833.400 ;
        RECT 691.950 826.950 694.050 829.050 ;
        RECT 701.400 823.050 702.450 844.950 ;
        RECT 703.950 841.950 706.050 844.050 ;
        RECT 704.400 832.050 705.450 841.950 ;
        RECT 710.400 840.600 711.450 853.950 ;
        RECT 716.400 853.050 717.450 878.400 ;
        RECT 721.950 853.950 724.050 856.050 ;
        RECT 715.950 850.950 718.050 853.050 ;
        RECT 710.400 838.350 711.600 840.600 ;
        RECT 715.950 839.100 718.050 841.200 ;
        RECT 716.400 838.350 717.600 839.100 ;
        RECT 709.950 835.950 712.050 838.050 ;
        RECT 712.950 835.950 715.050 838.050 ;
        RECT 715.950 835.950 718.050 838.050 ;
        RECT 713.400 833.400 714.600 835.650 ;
        RECT 703.950 829.950 706.050 832.050 ;
        RECT 703.950 823.950 706.050 826.050 ;
        RECT 694.950 820.950 697.050 823.050 ;
        RECT 700.950 820.950 703.050 823.050 ;
        RECT 688.950 814.950 691.050 817.050 ;
        RECT 695.400 807.600 696.450 820.950 ;
        RECT 695.400 805.350 696.600 807.600 ;
        RECT 691.950 802.950 694.050 805.050 ;
        RECT 694.950 802.950 697.050 805.050 ;
        RECT 697.950 802.950 700.050 805.050 ;
        RECT 698.400 800.400 699.600 802.650 ;
        RECT 698.400 790.050 699.450 800.400 ;
        RECT 700.950 796.950 703.050 799.050 ;
        RECT 701.400 793.050 702.450 796.950 ;
        RECT 700.950 790.950 703.050 793.050 ;
        RECT 704.400 790.050 705.450 823.950 ;
        RECT 706.950 820.950 709.050 823.050 ;
        RECT 707.400 796.050 708.450 820.950 ;
        RECT 713.400 817.050 714.450 833.400 ;
        RECT 722.400 823.050 723.450 853.950 ;
        RECT 728.400 841.200 729.450 892.950 ;
        RECT 733.950 884.100 736.050 886.200 ;
        RECT 734.400 883.350 735.600 884.100 ;
        RECT 733.950 880.950 736.050 883.050 ;
        RECT 736.950 880.950 739.050 883.050 ;
        RECT 737.400 879.000 738.600 880.650 ;
        RECT 736.950 874.950 739.050 879.000 ;
        RECT 743.400 853.050 744.450 907.950 ;
        RECT 749.400 907.050 750.450 925.950 ;
        RECT 748.950 904.950 751.050 907.050 ;
        RECT 752.400 904.050 753.450 952.950 ;
        RECT 779.400 952.050 780.450 956.400 ;
        RECT 784.950 955.800 787.050 957.900 ;
        RECT 793.950 955.800 796.050 957.900 ;
        RECT 806.400 956.400 807.600 958.650 ;
        RECT 812.400 957.000 813.600 958.650 ;
        RECT 769.950 949.950 772.050 952.050 ;
        RECT 778.950 949.950 781.050 952.050 ;
        RECT 757.950 917.100 760.050 919.200 ;
        RECT 758.400 916.350 759.600 917.100 ;
        RECT 766.950 916.950 769.050 919.050 ;
        RECT 757.950 913.950 760.050 916.050 ;
        RECT 760.950 913.950 763.050 916.050 ;
        RECT 761.400 912.000 762.600 913.650 ;
        RECT 760.950 907.950 763.050 912.000 ;
        RECT 751.950 901.950 754.050 904.050 ;
        RECT 767.400 889.050 768.450 916.950 ;
        RECT 770.400 912.900 771.450 949.950 ;
        RECT 806.400 946.050 807.450 956.400 ;
        RECT 811.950 952.950 814.050 957.000 ;
        RECT 818.400 955.050 819.450 967.950 ;
        RECT 823.950 966.750 826.050 967.200 ;
        RECT 829.950 966.750 832.050 967.200 ;
        RECT 823.950 965.700 832.050 966.750 ;
        RECT 823.950 965.100 826.050 965.700 ;
        RECT 829.950 965.100 832.050 965.700 ;
        RECT 820.950 961.950 823.050 964.050 ;
        RECT 829.950 961.950 832.050 964.050 ;
        RECT 817.950 952.950 820.050 955.050 ;
        RECT 805.950 943.950 808.050 946.050 ;
        RECT 775.950 940.950 778.050 943.050 ;
        RECT 776.400 937.050 777.450 940.950 ;
        RECT 778.950 937.950 781.050 940.050 ;
        RECT 775.950 934.950 778.050 937.050 ;
        RECT 776.400 918.600 777.450 934.950 ;
        RECT 779.400 928.050 780.450 937.950 ;
        RECT 781.950 928.950 784.050 931.050 ;
        RECT 805.950 928.950 808.050 931.050 ;
        RECT 778.950 925.950 781.050 928.050 ;
        RECT 782.400 925.050 783.450 928.950 ;
        RECT 781.950 922.950 784.050 925.050 ;
        RECT 782.400 918.600 783.450 922.950 ;
        RECT 806.400 918.600 807.450 928.950 ;
        RECT 821.400 925.050 822.450 961.950 ;
        RECT 830.400 961.350 831.600 961.950 ;
        RECT 826.950 958.950 829.050 961.050 ;
        RECT 829.950 958.950 832.050 961.050 ;
        RECT 827.400 957.900 828.600 958.650 ;
        RECT 826.950 955.800 829.050 957.900 ;
        RECT 836.400 931.050 837.450 973.950 ;
        RECT 856.950 970.950 859.050 973.050 ;
        RECT 844.950 966.450 847.050 967.050 ;
        RECT 853.950 966.450 856.050 967.050 ;
        RECT 844.950 965.400 856.050 966.450 ;
        RECT 844.950 964.950 847.050 965.400 ;
        RECT 853.950 964.950 856.050 965.400 ;
        RECT 850.950 962.100 853.050 964.200 ;
        RECT 857.400 963.600 858.450 970.950 ;
        RECT 883.950 967.950 886.050 973.050 ;
        RECT 886.950 967.950 889.050 970.050 ;
        RECT 889.950 967.950 895.050 970.050 ;
        RECT 868.950 966.450 871.050 967.050 ;
        RECT 868.950 965.400 879.450 966.450 ;
        RECT 868.950 964.950 871.050 965.400 ;
        RECT 878.400 964.200 879.450 965.400 ;
        RECT 851.400 961.350 852.600 962.100 ;
        RECT 857.400 961.350 858.600 963.600 ;
        RECT 871.950 962.100 874.050 964.200 ;
        RECT 877.950 962.100 880.050 964.200 ;
        RECT 872.400 961.350 873.600 962.100 ;
        RECT 878.400 961.350 879.600 962.100 ;
        RECT 847.950 958.950 850.050 961.050 ;
        RECT 850.950 958.950 853.050 961.050 ;
        RECT 853.950 958.950 856.050 961.050 ;
        RECT 856.950 958.950 859.050 961.050 ;
        RECT 871.950 958.950 874.050 961.050 ;
        RECT 874.950 958.950 877.050 961.050 ;
        RECT 877.950 958.950 880.050 961.050 ;
        RECT 880.950 958.950 883.050 961.050 ;
        RECT 844.950 952.950 847.050 958.050 ;
        RECT 848.400 957.000 849.600 958.650 ;
        RECT 854.400 957.900 855.600 958.650 ;
        RECT 847.950 952.950 850.050 957.000 ;
        RECT 853.950 955.800 856.050 957.900 ;
        RECT 862.950 955.800 865.050 957.900 ;
        RECT 875.400 957.000 876.600 958.650 ;
        RECT 881.400 957.900 882.600 958.650 ;
        RECT 887.400 958.050 888.450 967.950 ;
        RECT 910.950 964.950 913.050 967.050 ;
        RECT 898.950 962.100 901.050 964.200 ;
        RECT 904.950 962.100 907.050 964.200 ;
        RECT 899.400 961.350 900.600 962.100 ;
        RECT 905.400 961.350 906.600 962.100 ;
        RECT 895.950 958.950 898.050 961.050 ;
        RECT 898.950 958.950 901.050 961.050 ;
        RECT 901.950 958.950 904.050 961.050 ;
        RECT 904.950 958.950 907.050 961.050 ;
        RECT 853.950 954.450 856.050 954.750 ;
        RECT 859.950 954.450 862.050 955.050 ;
        RECT 853.950 953.400 862.050 954.450 ;
        RECT 853.950 952.650 856.050 953.400 ;
        RECT 859.950 952.950 862.050 953.400 ;
        RECT 863.400 943.050 864.450 955.800 ;
        RECT 865.950 952.950 871.050 955.050 ;
        RECT 874.950 952.950 877.050 957.000 ;
        RECT 880.950 955.800 883.050 957.900 ;
        RECT 886.950 955.950 889.050 958.050 ;
        RECT 896.400 957.900 897.600 958.650 ;
        RECT 895.950 955.800 898.050 957.900 ;
        RECT 902.400 956.400 903.600 958.650 ;
        RECT 875.400 946.050 876.450 952.950 ;
        RECT 886.950 952.800 889.050 954.900 ;
        RECT 874.950 943.950 877.050 946.050 ;
        RECT 862.950 940.950 865.050 943.050 ;
        RECT 835.950 928.950 838.050 931.050 ;
        RECT 865.950 925.950 868.050 928.050 ;
        RECT 820.950 922.950 823.050 925.050 ;
        RECT 850.950 922.950 853.050 925.050 ;
        RECT 776.400 916.350 777.600 918.600 ;
        RECT 782.400 916.350 783.600 918.600 ;
        RECT 806.400 916.350 807.600 918.600 ;
        RECT 811.950 917.100 814.050 919.200 ;
        RECT 817.950 917.100 820.050 919.200 ;
        RECT 812.400 916.350 813.600 917.100 ;
        RECT 775.950 913.950 778.050 916.050 ;
        RECT 778.950 913.950 781.050 916.050 ;
        RECT 781.950 913.950 784.050 916.050 ;
        RECT 784.950 913.950 787.050 916.050 ;
        RECT 802.950 913.950 805.050 916.050 ;
        RECT 805.950 913.950 808.050 916.050 ;
        RECT 808.950 913.950 811.050 916.050 ;
        RECT 811.950 913.950 814.050 916.050 ;
        RECT 779.400 912.900 780.600 913.650 ;
        RECT 785.400 912.900 786.600 913.650 ;
        RECT 803.400 912.900 804.600 913.650 ;
        RECT 769.950 910.800 772.050 912.900 ;
        RECT 778.950 910.800 781.050 912.900 ;
        RECT 784.950 910.800 787.050 912.900 ;
        RECT 802.950 910.800 805.050 912.900 ;
        RECT 809.400 911.400 810.600 913.650 ;
        RECT 772.950 898.950 775.050 901.050 ;
        RECT 757.950 885.000 760.050 889.050 ;
        RECT 766.950 886.950 769.050 889.050 ;
        RECT 764.400 885.450 765.600 885.600 ;
        RECT 758.400 883.350 759.600 885.000 ;
        RECT 764.400 884.400 771.450 885.450 ;
        RECT 764.400 883.350 765.600 884.400 ;
        RECT 754.950 880.950 757.050 883.050 ;
        RECT 757.950 880.950 760.050 883.050 ;
        RECT 760.950 880.950 763.050 883.050 ;
        RECT 763.950 880.950 766.050 883.050 ;
        RECT 755.400 879.900 756.600 880.650 ;
        RECT 754.950 877.800 757.050 879.900 ;
        RECT 761.400 878.400 762.600 880.650 ;
        RECT 761.400 871.050 762.450 878.400 ;
        RECT 760.950 868.950 763.050 871.050 ;
        RECT 770.400 868.050 771.450 884.400 ;
        RECT 769.950 865.950 772.050 868.050 ;
        RECT 773.400 856.050 774.450 898.950 ;
        RECT 809.400 895.050 810.450 911.400 ;
        RECT 808.950 892.950 811.050 895.050 ;
        RECT 781.950 885.000 784.050 889.050 ;
        RECT 782.400 883.350 783.600 885.000 ;
        RECT 787.950 884.100 790.050 886.200 ;
        RECT 788.400 883.350 789.600 884.100 ;
        RECT 796.950 883.950 799.050 886.050 ;
        RECT 805.950 884.100 808.050 886.200 ;
        RECT 811.950 884.100 814.050 886.200 ;
        RECT 778.950 880.950 781.050 883.050 ;
        RECT 781.950 880.950 784.050 883.050 ;
        RECT 784.950 880.950 787.050 883.050 ;
        RECT 787.950 880.950 790.050 883.050 ;
        RECT 779.400 878.400 780.600 880.650 ;
        RECT 785.400 879.900 786.600 880.650 ;
        RECT 779.400 871.050 780.450 878.400 ;
        RECT 784.950 877.800 787.050 879.900 ;
        RECT 778.950 868.950 781.050 871.050 ;
        RECT 772.950 853.950 775.050 856.050 ;
        RECT 742.950 850.950 745.050 853.050 ;
        RECT 727.950 839.100 730.050 841.200 ;
        RECT 733.950 839.100 736.050 841.200 ;
        RECT 734.400 838.350 735.600 839.100 ;
        RECT 730.950 835.950 733.050 838.050 ;
        RECT 733.950 835.950 736.050 838.050 ;
        RECT 736.950 835.950 739.050 838.050 ;
        RECT 731.400 833.400 732.600 835.650 ;
        RECT 737.400 834.000 738.600 835.650 ;
        RECT 721.950 820.950 724.050 823.050 ;
        RECT 712.950 814.950 715.050 817.050 ;
        RECT 712.950 802.950 715.050 805.050 ;
        RECT 715.950 802.950 718.050 805.050 ;
        RECT 718.950 802.950 721.050 805.050 ;
        RECT 721.950 802.950 724.050 805.050 ;
        RECT 724.950 802.950 727.050 805.050 ;
        RECT 713.400 801.000 714.600 802.650 ;
        RECT 712.950 796.950 715.050 801.000 ;
        RECT 719.400 800.400 720.600 802.650 ;
        RECT 725.400 800.400 726.600 802.650 ;
        RECT 719.400 799.050 720.450 800.400 ;
        RECT 719.400 797.400 724.050 799.050 ;
        RECT 720.000 796.950 724.050 797.400 ;
        RECT 706.950 793.950 709.050 796.050 ;
        RECT 706.950 790.800 709.050 792.900 ;
        RECT 691.950 787.950 694.050 790.050 ;
        RECT 697.950 787.950 700.050 790.050 ;
        RECT 703.950 787.950 706.050 790.050 ;
        RECT 682.950 784.950 685.050 787.050 ;
        RECT 664.950 775.950 667.050 778.050 ;
        RECT 688.950 775.950 691.050 778.050 ;
        RECT 670.950 766.950 673.050 769.050 ;
        RECT 671.400 762.600 672.450 766.950 ;
        RECT 682.950 763.950 685.050 766.050 ;
        RECT 671.400 760.350 672.600 762.600 ;
        RECT 676.950 761.100 679.050 763.200 ;
        RECT 677.400 760.350 678.600 761.100 ;
        RECT 667.950 757.950 670.050 760.050 ;
        RECT 670.950 757.950 673.050 760.050 ;
        RECT 673.950 757.950 676.050 760.050 ;
        RECT 676.950 757.950 679.050 760.050 ;
        RECT 668.400 756.450 669.600 757.650 ;
        RECT 674.400 756.900 675.600 757.650 ;
        RECT 662.400 755.400 669.600 756.450 ;
        RECT 673.950 754.800 676.050 756.900 ;
        RECT 634.950 730.950 637.050 733.050 ;
        RECT 620.400 711.450 621.450 728.100 ;
        RECT 626.400 727.350 627.600 728.100 ;
        RECT 632.400 727.350 633.600 729.600 ;
        RECT 625.950 724.950 628.050 727.050 ;
        RECT 628.950 724.950 631.050 727.050 ;
        RECT 631.950 724.950 634.050 727.050 ;
        RECT 634.950 724.950 637.050 727.050 ;
        RECT 629.400 722.400 630.600 724.650 ;
        RECT 635.400 723.900 636.600 724.650 ;
        RECT 625.950 715.950 628.050 718.050 ;
        RECT 620.400 710.400 624.450 711.450 ;
        RECT 616.950 686.100 619.050 688.200 ;
        RECT 611.400 682.350 612.600 684.600 ;
        RECT 616.950 682.950 619.050 685.050 ;
        RECT 617.400 682.350 618.600 682.950 ;
        RECT 610.950 679.950 613.050 682.050 ;
        RECT 613.950 679.950 616.050 682.050 ;
        RECT 616.950 679.950 619.050 682.050 ;
        RECT 604.950 676.950 607.050 679.050 ;
        RECT 614.400 678.000 615.600 679.650 ;
        RECT 613.950 673.950 616.050 678.000 ;
        RECT 623.400 664.050 624.450 710.400 ;
        RECT 626.400 676.050 627.450 715.950 ;
        RECT 629.400 715.050 630.450 722.400 ;
        RECT 634.950 721.800 637.050 723.900 ;
        RECT 643.950 721.800 646.050 723.900 ;
        RECT 637.950 715.950 640.050 718.050 ;
        RECT 628.950 712.950 631.050 715.050 ;
        RECT 638.400 709.050 639.450 715.950 ;
        RECT 644.400 712.050 645.450 721.800 ;
        RECT 647.400 718.050 648.450 754.800 ;
        RECT 679.950 753.450 682.050 757.050 ;
        RECT 677.400 753.000 682.050 753.450 ;
        RECT 676.950 752.400 681.450 753.000 ;
        RECT 667.950 748.950 670.050 751.050 ;
        RECT 676.950 748.950 679.050 752.400 ;
        RECT 655.950 739.950 658.050 742.050 ;
        RECT 656.400 730.200 657.450 739.950 ;
        RECT 655.950 728.100 658.050 730.200 ;
        RECT 656.400 727.350 657.600 728.100 ;
        RECT 652.950 724.950 655.050 727.050 ;
        RECT 655.950 724.950 658.050 727.050 ;
        RECT 658.950 724.950 661.050 727.050 ;
        RECT 659.400 723.900 660.600 724.650 ;
        RECT 658.950 721.800 661.050 723.900 ;
        RECT 668.400 718.050 669.450 748.950 ;
        RECT 683.400 742.050 684.450 763.950 ;
        RECT 689.400 753.450 690.450 775.950 ;
        RECT 692.400 763.050 693.450 787.950 ;
        RECT 697.950 766.050 700.050 766.200 ;
        RECT 697.950 764.100 703.050 766.050 ;
        RECT 699.000 763.950 703.050 764.100 ;
        RECT 691.950 760.950 694.050 763.050 ;
        RECT 697.950 760.950 700.050 763.050 ;
        RECT 703.950 761.100 706.050 763.200 ;
        RECT 698.400 760.350 699.600 760.950 ;
        RECT 694.950 757.950 697.050 760.050 ;
        RECT 697.950 757.950 700.050 760.050 ;
        RECT 695.400 756.000 696.600 757.650 ;
        RECT 689.400 752.400 693.450 753.450 ;
        RECT 682.950 739.950 685.050 742.050 ;
        RECT 670.950 730.950 673.050 733.050 ;
        RECT 646.950 715.950 649.050 718.050 ;
        RECT 658.950 715.950 661.050 718.050 ;
        RECT 667.950 715.950 670.050 718.050 ;
        RECT 643.950 709.950 646.050 712.050 ;
        RECT 637.950 706.950 640.050 709.050 ;
        RECT 655.950 688.950 658.050 691.050 ;
        RECT 637.950 683.100 640.050 685.200 ;
        RECT 638.400 682.350 639.600 683.100 ;
        RECT 643.950 682.950 646.050 685.050 ;
        RECT 656.400 684.600 657.450 688.950 ;
        RECT 659.400 688.050 660.450 715.950 ;
        RECT 671.400 715.050 672.450 730.950 ;
        RECT 688.950 727.950 691.050 730.050 ;
        RECT 674.100 724.950 676.200 727.050 ;
        RECT 679.500 724.950 681.600 727.050 ;
        RECT 682.800 724.950 684.900 727.050 ;
        RECT 674.400 723.900 675.600 724.650 ;
        RECT 673.950 721.800 676.050 723.900 ;
        RECT 683.400 722.400 684.600 724.650 ;
        RECT 670.950 712.950 673.050 715.050 ;
        RECT 667.950 703.950 670.050 706.050 ;
        RECT 658.950 685.950 661.050 688.050 ;
        RECT 664.950 685.950 667.050 688.050 ;
        RECT 634.950 679.950 637.050 682.050 ;
        RECT 637.950 679.950 640.050 682.050 ;
        RECT 635.400 677.400 636.600 679.650 ;
        RECT 625.950 673.950 628.050 676.050 ;
        RECT 635.400 673.050 636.450 677.400 ;
        RECT 634.950 670.950 637.050 673.050 ;
        RECT 622.950 661.950 625.050 664.050 ;
        RECT 628.950 661.950 631.050 664.050 ;
        RECT 625.950 658.950 628.050 661.050 ;
        RECT 616.950 655.950 619.050 658.050 ;
        RECT 617.400 655.200 618.600 655.950 ;
        RECT 604.950 649.950 607.050 652.050 ;
        RECT 612.900 651.900 615.000 653.700 ;
        RECT 616.800 652.800 618.900 654.900 ;
        RECT 620.100 654.300 622.200 656.400 ;
        RECT 611.400 650.700 620.100 651.900 ;
        RECT 605.400 645.450 606.450 649.950 ;
        RECT 608.100 646.950 610.200 649.050 ;
        RECT 608.400 645.900 609.600 646.650 ;
        RECT 607.950 645.450 610.050 645.900 ;
        RECT 605.400 644.400 610.050 645.450 ;
        RECT 607.950 643.800 610.050 644.400 ;
        RECT 611.400 641.700 612.300 650.700 ;
        RECT 618.000 649.800 620.100 650.700 ;
        RECT 621.000 648.900 621.900 654.300 ;
        RECT 622.950 650.100 625.050 652.200 ;
        RECT 623.400 649.350 624.600 650.100 ;
        RECT 615.000 647.700 621.900 648.900 ;
        RECT 615.000 645.300 615.900 647.700 ;
        RECT 613.800 643.200 615.900 645.300 ;
        RECT 616.800 643.950 618.900 646.050 ;
        RECT 610.500 639.600 612.600 641.700 ;
        RECT 617.400 641.400 618.600 643.650 ;
        RECT 620.700 640.500 621.900 647.700 ;
        RECT 622.800 646.950 624.900 649.050 ;
        RECT 620.100 638.400 622.200 640.500 ;
        RECT 626.400 637.050 627.450 658.950 ;
        RECT 629.400 652.200 630.450 661.950 ;
        RECT 640.950 658.950 643.050 661.050 ;
        RECT 631.950 655.950 634.050 658.050 ;
        RECT 628.950 650.100 631.050 652.200 ;
        RECT 604.950 634.950 607.050 637.050 ;
        RECT 625.950 634.950 628.050 637.050 ;
        RECT 601.950 592.950 604.050 595.050 ;
        RECT 589.950 586.950 592.050 589.050 ;
        RECT 590.400 574.200 591.450 586.950 ;
        RECT 605.400 586.050 606.450 634.950 ;
        RECT 610.950 631.950 613.050 634.050 ;
        RECT 611.400 616.050 612.450 631.950 ;
        RECT 625.950 628.950 628.050 631.050 ;
        RECT 619.950 616.950 622.050 619.050 ;
        RECT 610.950 613.950 613.050 616.050 ;
        RECT 613.950 606.000 616.050 610.050 ;
        RECT 620.400 606.600 621.450 616.950 ;
        RECT 614.400 604.350 615.600 606.000 ;
        RECT 620.400 604.350 621.600 606.600 ;
        RECT 610.950 601.950 613.050 604.050 ;
        RECT 613.950 601.950 616.050 604.050 ;
        RECT 616.950 601.950 619.050 604.050 ;
        RECT 619.950 601.950 622.050 604.050 ;
        RECT 611.400 600.900 612.600 601.650 ;
        RECT 610.950 598.800 613.050 600.900 ;
        RECT 617.400 599.400 618.600 601.650 ;
        RECT 604.950 583.950 607.050 586.050 ;
        RECT 610.950 583.950 613.050 586.050 ;
        RECT 617.400 585.450 618.450 599.400 ;
        RECT 626.400 598.050 627.450 628.950 ;
        RECT 632.400 610.050 633.450 655.950 ;
        RECT 641.400 651.600 642.450 658.950 ;
        RECT 644.400 655.050 645.450 682.950 ;
        RECT 656.400 682.350 657.600 684.600 ;
        RECT 652.950 679.950 655.050 682.050 ;
        RECT 655.950 679.950 658.050 682.050 ;
        RECT 658.950 679.950 661.050 682.050 ;
        RECT 653.400 677.400 654.600 679.650 ;
        RECT 659.400 679.050 660.600 679.650 ;
        RECT 659.400 677.400 664.050 679.050 ;
        RECT 653.400 664.050 654.450 677.400 ;
        RECT 660.000 676.950 664.050 677.400 ;
        RECT 665.400 667.050 666.450 685.950 ;
        RECT 668.400 679.050 669.450 703.950 ;
        RECT 667.950 676.800 670.050 679.050 ;
        RECT 664.950 664.950 667.050 667.050 ;
        RECT 652.950 661.950 655.050 664.050 ;
        RECT 653.400 658.050 654.450 661.950 ;
        RECT 652.950 655.950 655.050 658.050 ;
        RECT 671.400 655.050 672.450 712.950 ;
        RECT 683.400 712.050 684.450 722.400 ;
        RECT 689.400 712.050 690.450 727.950 ;
        RECT 682.950 709.950 685.050 712.050 ;
        RECT 688.950 709.950 691.050 712.050 ;
        RECT 692.400 700.050 693.450 752.400 ;
        RECT 694.950 751.950 697.050 756.000 ;
        RECT 704.400 733.050 705.450 761.100 ;
        RECT 700.950 729.000 703.050 733.050 ;
        RECT 703.950 730.950 706.050 733.050 ;
        RECT 707.400 730.050 708.450 790.800 ;
        RECT 713.400 769.050 714.450 796.950 ;
        RECT 715.950 793.950 718.050 796.050 ;
        RECT 716.400 772.050 717.450 793.950 ;
        RECT 725.400 787.050 726.450 800.400 ;
        RECT 724.950 784.950 727.050 787.050 ;
        RECT 715.950 769.950 718.050 772.050 ;
        RECT 712.950 766.950 715.050 769.050 ;
        RECT 712.950 761.100 715.050 763.200 ;
        RECT 718.950 761.100 721.050 766.050 ;
        RECT 713.400 760.350 714.600 761.100 ;
        RECT 719.400 760.350 720.600 761.100 ;
        RECT 712.950 757.950 715.050 760.050 ;
        RECT 715.950 757.950 718.050 760.050 ;
        RECT 718.950 757.950 721.050 760.050 ;
        RECT 721.950 757.950 724.050 760.050 ;
        RECT 722.400 756.900 723.600 757.650 ;
        RECT 721.950 754.800 724.050 756.900 ;
        RECT 731.400 754.050 732.450 833.400 ;
        RECT 736.950 829.950 739.050 834.000 ;
        RECT 743.400 826.050 744.450 850.950 ;
        RECT 775.950 847.950 778.050 850.050 ;
        RECT 760.950 844.950 763.050 847.050 ;
        RECT 766.950 844.950 769.050 847.050 ;
        RECT 754.950 839.100 757.050 841.200 ;
        RECT 761.400 840.600 762.450 844.950 ;
        RECT 755.400 838.350 756.600 839.100 ;
        RECT 761.400 838.350 762.600 840.600 ;
        RECT 751.950 835.950 754.050 838.050 ;
        RECT 754.950 835.950 757.050 838.050 ;
        RECT 757.950 835.950 760.050 838.050 ;
        RECT 760.950 835.950 763.050 838.050 ;
        RECT 752.400 834.900 753.600 835.650 ;
        RECT 758.400 834.900 759.600 835.650 ;
        RECT 751.950 832.800 754.050 834.900 ;
        RECT 757.950 832.800 760.050 834.900 ;
        RECT 752.400 826.050 753.450 832.800 ;
        RECT 767.400 829.050 768.450 844.950 ;
        RECT 772.950 838.950 775.050 841.050 ;
        RECT 773.400 832.050 774.450 838.950 ;
        RECT 776.400 835.050 777.450 847.950 ;
        RECT 797.400 847.050 798.450 883.950 ;
        RECT 806.400 883.350 807.600 884.100 ;
        RECT 812.400 883.350 813.600 884.100 ;
        RECT 802.950 880.950 805.050 883.050 ;
        RECT 805.950 880.950 808.050 883.050 ;
        RECT 808.950 880.950 811.050 883.050 ;
        RECT 811.950 880.950 814.050 883.050 ;
        RECT 803.400 878.400 804.600 880.650 ;
        RECT 809.400 879.000 810.600 880.650 ;
        RECT 799.950 874.950 802.050 877.050 ;
        RECT 796.950 844.950 799.050 847.050 ;
        RECT 787.950 839.100 790.050 841.200 ;
        RECT 796.950 839.100 799.050 841.200 ;
        RECT 788.400 838.350 789.600 839.100 ;
        RECT 797.400 838.350 798.600 839.100 ;
        RECT 781.800 835.950 783.900 838.050 ;
        RECT 787.950 835.950 790.050 838.050 ;
        RECT 790.950 835.950 793.050 838.050 ;
        RECT 796.500 835.950 798.600 838.050 ;
        RECT 775.950 832.950 778.050 835.050 ;
        RECT 782.400 833.400 783.600 835.650 ;
        RECT 791.400 834.000 792.600 835.650 ;
        RECT 772.950 829.950 775.050 832.050 ;
        RECT 782.400 829.050 783.450 833.400 ;
        RECT 790.950 829.950 793.050 834.000 ;
        RECT 766.950 826.950 769.050 829.050 ;
        RECT 781.950 826.950 784.050 829.050 ;
        RECT 733.950 823.950 736.050 826.050 ;
        RECT 742.950 823.950 745.050 826.050 ;
        RECT 751.950 823.950 754.050 826.050 ;
        RECT 734.400 799.050 735.450 823.950 ;
        RECT 781.950 823.800 784.050 825.900 ;
        RECT 742.950 814.950 745.050 817.050 ;
        RECT 743.400 808.200 744.450 814.950 ;
        RECT 742.950 806.100 745.050 808.200 ;
        RECT 763.950 806.100 766.050 808.200 ;
        RECT 769.950 806.100 772.050 808.200 ;
        RECT 778.950 806.100 781.050 808.200 ;
        RECT 743.400 805.350 744.600 806.100 ;
        RECT 764.400 805.350 765.600 806.100 ;
        RECT 770.400 805.350 771.600 806.100 ;
        RECT 739.950 802.950 742.050 805.050 ;
        RECT 742.950 802.950 745.050 805.050 ;
        RECT 745.950 802.950 748.050 805.050 ;
        RECT 754.950 802.950 757.050 805.050 ;
        RECT 760.950 802.950 763.050 805.050 ;
        RECT 763.950 802.950 766.050 805.050 ;
        RECT 766.950 802.950 769.050 805.050 ;
        RECT 769.950 802.950 772.050 805.050 ;
        RECT 772.950 802.950 775.050 805.050 ;
        RECT 740.400 800.400 741.600 802.650 ;
        RECT 733.950 796.950 736.050 799.050 ;
        RECT 740.400 787.050 741.450 800.400 ;
        RECT 739.950 784.950 742.050 787.050 ;
        RECT 755.400 775.050 756.450 802.950 ;
        RECT 761.400 800.400 762.600 802.650 ;
        RECT 767.400 801.900 768.600 802.650 ;
        RECT 757.950 793.950 760.050 796.050 ;
        RECT 758.400 787.050 759.450 793.950 ;
        RECT 761.400 793.050 762.450 800.400 ;
        RECT 766.950 799.800 769.050 801.900 ;
        RECT 773.400 800.400 774.600 802.650 ;
        RECT 779.400 802.050 780.450 806.100 ;
        RECT 782.400 805.050 783.450 823.800 ;
        RECT 787.950 814.950 790.050 817.050 ;
        RECT 788.400 807.600 789.450 814.950 ;
        RECT 788.400 805.350 789.600 807.600 ;
        RECT 781.950 802.950 784.050 805.050 ;
        RECT 787.950 802.950 790.050 805.050 ;
        RECT 790.950 802.950 793.050 805.050 ;
        RECT 763.950 796.950 766.050 799.050 ;
        RECT 760.950 790.950 763.050 793.050 ;
        RECT 757.950 784.950 760.050 787.050 ;
        RECT 754.950 772.950 757.050 775.050 ;
        RECT 736.950 766.950 739.050 769.050 ;
        RECT 748.950 766.950 751.050 769.050 ;
        RECT 733.950 760.950 736.050 766.050 ;
        RECT 733.950 754.950 736.050 757.050 ;
        RECT 730.950 751.950 733.050 754.050 ;
        RECT 724.950 745.950 727.050 748.050 ;
        RECT 725.400 742.050 726.450 745.950 ;
        RECT 734.400 745.050 735.450 754.950 ;
        RECT 733.950 742.950 736.050 745.050 ;
        RECT 709.950 739.950 712.050 742.050 ;
        RECT 724.950 739.950 727.050 742.050 ;
        RECT 710.400 733.050 711.450 739.950 ;
        RECT 730.950 736.950 733.050 739.050 ;
        RECT 709.950 730.950 712.050 733.050 ;
        RECT 715.950 730.950 718.050 733.050 ;
        RECT 701.400 727.350 702.600 729.000 ;
        RECT 706.950 727.950 709.050 730.050 ;
        RECT 697.950 724.950 700.050 727.050 ;
        RECT 700.950 724.950 703.050 727.050 ;
        RECT 703.950 724.950 706.050 727.050 ;
        RECT 704.400 723.450 705.600 724.650 ;
        RECT 706.950 723.450 709.050 724.050 ;
        RECT 704.400 722.400 709.050 723.450 ;
        RECT 706.950 721.950 709.050 722.400 ;
        RECT 673.950 697.950 676.050 700.050 ;
        RECT 691.950 697.950 694.050 700.050 ;
        RECT 697.950 697.950 700.050 700.050 ;
        RECT 643.950 652.950 646.050 655.050 ;
        RECT 670.950 652.950 673.050 655.050 ;
        RECT 641.400 649.350 642.600 651.600 ;
        RECT 646.950 650.100 649.050 652.200 ;
        RECT 647.400 649.350 648.600 650.100 ;
        RECT 658.950 649.950 661.050 652.050 ;
        RECT 637.950 646.950 640.050 649.050 ;
        RECT 640.950 646.950 643.050 649.050 ;
        RECT 643.950 646.950 646.050 649.050 ;
        RECT 646.950 646.950 649.050 649.050 ;
        RECT 638.400 644.400 639.600 646.650 ;
        RECT 644.400 645.000 645.600 646.650 ;
        RECT 638.400 618.450 639.450 644.400 ;
        RECT 640.950 640.950 643.050 643.050 ;
        RECT 643.950 640.950 646.050 645.000 ;
        RECT 659.400 643.050 660.450 649.950 ;
        RECT 662.100 646.950 664.200 649.050 ;
        RECT 667.500 646.950 669.600 649.050 ;
        RECT 670.800 646.950 672.900 649.050 ;
        RECT 662.400 644.400 663.600 646.650 ;
        RECT 671.400 645.450 672.600 646.650 ;
        RECT 674.400 645.450 675.450 697.950 ;
        RECT 680.100 688.500 682.200 690.600 ;
        RECT 677.100 679.950 679.200 682.050 ;
        RECT 680.100 681.900 681.000 688.500 ;
        RECT 689.100 688.200 691.200 690.300 ;
        RECT 683.400 685.350 684.600 687.600 ;
        RECT 682.800 682.950 684.900 685.050 ;
        RECT 687.000 681.900 689.100 682.200 ;
        RECT 680.100 681.000 689.100 681.900 ;
        RECT 677.400 678.900 678.600 679.650 ;
        RECT 676.950 676.800 679.050 678.900 ;
        RECT 680.100 675.900 681.000 681.000 ;
        RECT 687.000 680.100 689.100 681.000 ;
        RECT 681.900 679.200 684.000 680.100 ;
        RECT 681.900 678.000 689.100 679.200 ;
        RECT 687.000 677.100 689.100 678.000 ;
        RECT 679.500 673.800 681.600 675.900 ;
        RECT 682.800 674.100 684.900 676.200 ;
        RECT 690.000 675.600 690.900 688.200 ;
        RECT 698.400 685.200 699.450 697.950 ;
        RECT 703.950 691.800 706.050 693.900 ;
        RECT 704.400 688.050 705.450 691.800 ;
        RECT 703.950 685.950 706.050 688.050 ;
        RECT 691.950 683.100 694.050 685.200 ;
        RECT 697.950 683.100 700.050 685.200 ;
        RECT 707.400 684.450 708.450 721.950 ;
        RECT 710.400 721.050 711.450 730.950 ;
        RECT 712.950 727.950 715.050 730.050 ;
        RECT 709.950 718.950 712.050 721.050 ;
        RECT 713.400 715.050 714.450 727.950 ;
        RECT 716.400 724.050 717.450 730.950 ;
        RECT 731.400 729.600 732.450 736.950 ;
        RECT 731.400 727.350 732.600 729.600 ;
        RECT 721.950 724.950 724.050 727.050 ;
        RECT 724.950 724.950 727.050 727.050 ;
        RECT 727.950 724.950 730.050 727.050 ;
        RECT 730.950 724.950 733.050 727.050 ;
        RECT 715.950 721.950 718.050 724.050 ;
        RECT 722.400 723.900 723.600 724.650 ;
        RECT 721.950 721.800 724.050 723.900 ;
        RECT 728.400 723.000 729.600 724.650 ;
        RECT 727.950 718.950 730.050 723.000 ;
        RECT 709.800 712.950 711.900 715.050 ;
        RECT 712.950 712.950 715.050 715.050 ;
        RECT 721.950 712.950 724.050 715.050 ;
        RECT 710.400 687.450 711.450 712.950 ;
        RECT 710.400 686.400 714.450 687.450 ;
        RECT 704.400 683.400 708.450 684.450 ;
        RECT 713.400 684.600 714.450 686.400 ;
        RECT 692.400 682.350 693.600 683.100 ;
        RECT 691.800 679.950 693.900 682.050 ;
        RECT 683.400 671.550 684.600 673.800 ;
        RECT 689.400 673.500 691.500 675.600 ;
        RECT 676.950 664.950 679.050 667.050 ;
        RECT 671.400 644.400 675.450 645.450 ;
        RECT 658.950 640.950 661.050 643.050 ;
        RECT 635.400 617.400 639.450 618.450 ;
        RECT 635.400 610.050 636.450 617.400 ;
        RECT 631.950 607.950 634.050 610.050 ;
        RECT 634.950 607.950 637.050 610.050 ;
        RECT 641.400 607.200 642.450 640.950 ;
        RECT 662.400 634.050 663.450 644.400 ;
        RECT 661.950 631.950 664.050 634.050 ;
        RECT 661.950 610.950 664.050 613.050 ;
        RECT 635.400 606.450 636.600 606.600 ;
        RECT 629.400 605.400 636.600 606.450 ;
        RECT 625.950 595.950 628.050 598.050 ;
        RECT 614.400 584.400 618.450 585.450 ;
        RECT 602.850 579.300 604.950 581.400 ;
        RECT 583.950 571.950 586.050 574.050 ;
        RECT 589.950 572.100 592.050 574.200 ;
        RECT 590.400 571.350 591.600 572.100 ;
        RECT 586.950 568.950 589.050 571.050 ;
        RECT 589.950 568.950 592.050 571.050 ;
        RECT 592.950 568.950 595.050 571.050 ;
        RECT 598.950 568.950 601.050 571.050 ;
        RECT 587.400 566.400 588.600 568.650 ;
        RECT 593.400 566.400 594.600 568.650 ;
        RECT 599.400 566.400 600.600 568.650 ;
        RECT 580.950 559.950 583.050 562.050 ;
        RECT 587.400 556.050 588.450 566.400 ;
        RECT 589.950 559.950 592.050 562.050 ;
        RECT 586.950 553.950 589.050 556.050 ;
        RECT 574.950 547.950 577.050 550.050 ;
        RECT 580.950 523.950 583.050 526.050 ;
        RECT 583.950 523.950 586.050 526.050 ;
        RECT 584.400 522.900 585.600 523.650 ;
        RECT 590.400 523.050 591.450 559.950 ;
        RECT 593.400 559.050 594.450 566.400 ;
        RECT 592.950 556.950 595.050 559.050 ;
        RECT 592.950 553.800 595.050 555.900 ;
        RECT 583.950 520.800 586.050 522.900 ;
        RECT 589.950 520.950 592.050 523.050 ;
        RECT 571.950 514.950 574.050 517.050 ;
        RECT 547.950 508.950 550.050 511.050 ;
        RECT 559.950 508.950 562.050 511.050 ;
        RECT 565.950 508.950 568.050 511.050 ;
        RECT 560.400 502.050 561.450 508.950 ;
        RECT 568.950 505.950 571.050 508.050 ;
        RECT 544.950 499.950 547.050 502.050 ;
        RECT 559.950 499.950 562.050 502.050 ;
        RECT 565.350 501.300 567.450 503.400 ;
        RECT 545.400 463.050 546.450 499.950 ;
        RECT 553.950 494.100 556.050 496.200 ;
        RECT 559.950 494.100 562.050 496.200 ;
        RECT 554.400 493.350 555.600 494.100 ;
        RECT 560.400 493.350 561.600 494.100 ;
        RECT 550.950 490.950 553.050 493.050 ;
        RECT 553.950 490.950 556.050 493.050 ;
        RECT 559.950 490.950 562.050 493.050 ;
        RECT 551.400 488.400 552.600 490.650 ;
        RECT 566.250 488.400 567.450 501.300 ;
        RECT 551.400 475.050 552.450 488.400 ;
        RECT 565.350 486.300 567.450 488.400 ;
        RECT 566.250 479.700 567.450 486.300 ;
        RECT 565.350 477.600 567.450 479.700 ;
        RECT 550.950 472.950 553.050 475.050 ;
        RECT 544.950 460.950 547.050 463.050 ;
        RECT 550.950 460.950 553.050 463.050 ;
        RECT 544.650 457.500 546.750 458.400 ;
        RECT 544.650 456.300 548.850 457.500 ;
        RECT 541.950 450.000 544.050 454.050 ;
        RECT 542.400 448.350 543.600 450.000 ;
        RECT 541.800 445.950 543.900 448.050 ;
        RECT 517.950 433.950 520.050 436.050 ;
        RECT 529.350 435.600 531.450 437.700 ;
        RECT 535.950 436.950 538.050 439.050 ;
        RECT 547.650 437.700 548.850 456.300 ;
        RECT 551.400 450.600 552.450 460.950 ;
        RECT 565.350 459.300 567.450 461.400 ;
        RECT 566.250 452.700 567.450 459.300 ;
        RECT 565.350 450.600 567.450 452.700 ;
        RECT 551.400 448.350 552.600 450.600 ;
        RECT 550.950 445.950 553.050 448.050 ;
        RECT 559.950 445.950 562.050 448.050 ;
        RECT 553.950 442.950 556.050 445.050 ;
        RECT 560.400 443.400 561.600 445.650 ;
        RECT 547.050 435.600 549.150 437.700 ;
        RECT 550.950 436.950 553.050 439.050 ;
        RECT 526.950 424.950 529.050 427.050 ;
        RECT 517.950 416.100 520.050 418.200 ;
        RECT 518.400 415.350 519.600 416.100 ;
        RECT 518.400 412.950 520.500 415.050 ;
        RECT 523.800 412.950 525.900 415.050 ;
        RECT 524.400 410.400 525.600 412.650 ;
        RECT 517.950 406.950 520.050 409.050 ;
        RECT 511.950 391.950 514.050 394.050 ;
        RECT 490.950 388.950 493.050 391.050 ;
        RECT 481.950 385.950 484.050 388.050 ;
        RECT 484.650 379.500 486.750 380.400 ;
        RECT 484.650 378.300 488.850 379.500 ;
        RECT 481.950 372.000 484.050 376.050 ;
        RECT 482.400 370.350 483.600 372.000 ;
        RECT 481.800 367.950 483.900 370.050 ;
        RECT 481.950 361.950 484.050 364.050 ;
        RECT 475.950 349.950 478.050 352.050 ;
        RECT 482.400 348.450 483.450 361.950 ;
        RECT 487.650 359.700 488.850 378.300 ;
        RECT 491.400 373.200 492.450 388.950 ;
        RECT 511.950 387.450 516.000 388.050 ;
        RECT 511.950 387.000 516.450 387.450 ;
        RECT 511.950 385.950 517.050 387.000 ;
        RECT 514.950 382.950 517.050 385.950 ;
        RECT 506.250 379.500 508.350 380.400 ;
        RECT 511.950 379.950 514.050 382.050 ;
        RECT 504.150 378.300 508.350 379.500 ;
        RECT 490.950 371.100 493.050 373.200 ;
        RECT 499.950 371.100 502.050 373.200 ;
        RECT 491.400 370.350 492.600 371.100 ;
        RECT 500.400 370.350 501.600 371.100 ;
        RECT 490.950 367.950 493.050 370.050 ;
        RECT 499.950 367.950 502.050 370.050 ;
        RECT 504.150 359.700 505.350 378.300 ;
        RECT 512.400 375.450 513.450 379.950 ;
        RECT 509.400 374.400 513.450 375.450 ;
        RECT 509.400 372.600 510.450 374.400 ;
        RECT 509.400 370.350 510.600 372.600 ;
        RECT 514.950 370.950 517.050 373.050 ;
        RECT 509.100 367.950 511.200 370.050 ;
        RECT 511.950 364.950 514.050 367.050 ;
        RECT 487.050 357.600 489.150 359.700 ;
        RECT 503.850 357.600 505.950 359.700 ;
        RECT 512.400 352.050 513.450 364.950 ;
        RECT 493.950 349.950 496.050 352.050 ;
        RECT 502.950 349.950 505.050 352.050 ;
        RECT 511.950 349.950 514.050 352.050 ;
        RECT 473.400 347.400 483.450 348.450 ;
        RECT 460.950 343.950 463.050 346.050 ;
        RECT 461.400 339.600 462.450 343.950 ;
        RECT 455.400 337.350 456.600 339.600 ;
        RECT 461.400 337.350 462.600 339.600 ;
        RECT 475.950 339.000 478.050 343.050 ;
        RECT 476.400 337.350 477.600 339.000 ;
        RECT 451.950 334.950 454.050 337.050 ;
        RECT 454.950 334.950 457.050 337.050 ;
        RECT 457.950 334.950 460.050 337.050 ;
        RECT 460.950 334.950 463.050 337.050 ;
        RECT 476.400 334.950 478.500 337.050 ;
        RECT 481.800 334.950 483.900 337.050 ;
        RECT 436.950 332.400 441.450 333.450 ;
        RECT 436.950 331.800 439.050 332.400 ;
        RECT 440.400 301.050 441.450 332.400 ;
        RECT 445.950 331.800 448.050 333.900 ;
        RECT 452.400 332.400 453.600 334.650 ;
        RECT 458.400 333.900 459.600 334.650 ;
        RECT 482.400 333.900 483.600 334.650 ;
        RECT 448.950 319.950 451.050 322.050 ;
        RECT 449.400 316.050 450.450 319.950 ;
        RECT 448.950 313.950 451.050 316.050 ;
        RECT 452.400 307.050 453.450 332.400 ;
        RECT 457.950 331.800 460.050 333.900 ;
        RECT 481.950 331.800 484.050 333.900 ;
        RECT 451.950 304.950 454.050 307.050 ;
        RECT 439.950 298.950 442.050 301.050 ;
        RECT 451.950 298.950 454.050 301.050 ;
        RECT 458.400 300.450 459.450 331.800 ;
        RECT 466.950 316.950 469.050 319.050 ;
        RECT 467.400 313.050 468.450 316.950 ;
        RECT 469.950 313.950 472.050 316.050 ;
        RECT 466.950 310.950 469.050 313.050 ;
        RECT 455.400 299.400 459.450 300.450 ;
        RECT 430.950 293.100 433.050 295.200 ;
        RECT 436.950 293.100 439.050 295.200 ;
        RECT 442.950 293.100 445.050 295.200 ;
        RECT 431.400 283.050 432.450 293.100 ;
        RECT 437.400 292.350 438.600 293.100 ;
        RECT 443.400 292.350 444.600 293.100 ;
        RECT 436.950 289.950 439.050 292.050 ;
        RECT 439.950 289.950 442.050 292.050 ;
        RECT 442.950 289.950 445.050 292.050 ;
        RECT 445.950 289.950 448.050 292.050 ;
        RECT 440.400 288.900 441.600 289.650 ;
        RECT 439.950 286.800 442.050 288.900 ;
        RECT 446.400 287.400 447.600 289.650 ;
        RECT 446.400 283.050 447.450 287.400 ;
        RECT 452.400 283.050 453.450 298.950 ;
        RECT 430.950 280.950 433.050 283.050 ;
        RECT 445.950 280.950 448.050 283.050 ;
        RECT 451.950 280.950 454.050 283.050 ;
        RECT 433.950 277.950 436.050 280.050 ;
        RECT 427.950 271.950 430.050 274.050 ;
        RECT 427.950 265.950 430.050 268.050 ;
        RECT 418.950 259.950 421.050 262.050 ;
        RECT 421.950 259.950 424.050 262.050 ;
        RECT 428.400 261.600 429.450 265.950 ;
        RECT 434.400 262.200 435.450 277.950 ;
        RECT 442.950 268.950 445.050 271.050 ;
        RECT 439.950 265.950 442.050 268.050 ;
        RECT 415.950 256.950 418.050 259.050 ;
        RECT 410.400 254.400 414.450 255.450 ;
        RECT 376.950 247.950 379.050 250.050 ;
        RECT 394.950 247.950 397.050 250.050 ;
        RECT 349.950 235.950 352.050 238.050 ;
        RECT 332.550 225.300 334.650 227.400 ;
        RECT 343.800 226.950 345.900 229.050 ;
        RECT 346.950 226.950 349.050 229.050 ;
        RECT 332.550 218.700 333.750 225.300 ;
        RECT 332.550 216.600 334.650 218.700 ;
        RECT 322.950 208.950 325.050 211.050 ;
        RECT 328.950 208.950 331.050 211.050 ;
        RECT 314.850 201.600 316.950 203.700 ;
        RECT 311.400 197.400 315.450 198.450 ;
        RECT 301.950 193.950 304.050 196.050 ;
        RECT 310.950 193.950 313.050 196.050 ;
        RECT 280.950 187.950 283.050 190.050 ;
        RECT 277.950 184.950 280.050 187.050 ;
        RECT 281.400 177.900 282.450 187.950 ;
        RECT 289.950 182.100 292.050 184.200 ;
        RECT 290.400 181.350 291.600 182.100 ;
        RECT 298.950 181.950 301.050 184.050 ;
        RECT 286.950 178.950 289.050 181.050 ;
        RECT 289.950 178.950 292.050 181.050 ;
        RECT 292.950 178.950 295.050 181.050 ;
        RECT 287.400 177.900 288.600 178.650 ;
        RECT 280.950 175.800 283.050 177.900 ;
        RECT 286.950 175.800 289.050 177.900 ;
        RECT 299.400 175.050 300.450 181.950 ;
        RECT 302.400 177.900 303.450 193.950 ;
        RECT 307.950 187.950 310.050 190.050 ;
        RECT 308.400 184.200 309.450 187.950 ;
        RECT 311.400 187.050 312.450 193.950 ;
        RECT 310.950 184.950 313.050 187.050 ;
        RECT 307.950 182.100 310.050 184.200 ;
        RECT 314.400 183.600 315.450 197.400 ;
        RECT 308.400 181.350 309.600 182.100 ;
        RECT 314.400 181.350 315.600 183.600 ;
        RECT 307.950 178.950 310.050 181.050 ;
        RECT 310.950 178.950 313.050 181.050 ;
        RECT 313.950 178.950 316.050 181.050 ;
        RECT 316.950 178.950 319.050 181.050 ;
        RECT 311.400 177.900 312.600 178.650 ;
        RECT 301.950 175.800 304.050 177.900 ;
        RECT 310.950 175.800 313.050 177.900 ;
        RECT 317.400 176.400 318.600 178.650 ;
        RECT 323.400 178.050 324.450 208.950 ;
        RECT 332.550 203.700 333.750 216.600 ;
        RECT 337.950 211.950 340.050 214.050 ;
        RECT 338.400 209.400 339.600 211.650 ;
        RECT 344.400 210.900 345.450 226.950 ;
        RECT 343.950 210.450 346.050 210.900 ;
        RECT 343.950 209.400 348.450 210.450 ;
        RECT 332.550 201.600 334.650 203.700 ;
        RECT 338.400 202.050 339.450 209.400 ;
        RECT 343.950 208.800 346.050 209.400 ;
        RECT 337.950 201.450 340.050 202.050 ;
        RECT 337.950 200.400 342.450 201.450 ;
        RECT 337.950 199.950 340.050 200.400 ;
        RECT 334.950 190.950 337.050 193.050 ;
        RECT 335.400 183.600 336.450 190.950 ;
        RECT 341.400 184.050 342.450 200.400 ;
        RECT 343.950 190.950 346.050 193.050 ;
        RECT 335.400 181.350 336.600 183.600 ;
        RECT 340.950 181.950 343.050 184.050 ;
        RECT 331.950 178.950 334.050 181.050 ;
        RECT 334.950 178.950 337.050 181.050 ;
        RECT 337.950 178.950 340.050 181.050 ;
        RECT 298.950 172.950 301.050 175.050 ;
        RECT 310.950 174.450 313.050 174.750 ;
        RECT 317.400 174.450 318.450 176.400 ;
        RECT 322.950 175.950 325.050 178.050 ;
        RECT 328.950 175.950 331.050 178.050 ;
        RECT 332.400 177.900 333.600 178.650 ;
        RECT 338.400 177.900 339.600 178.650 ;
        RECT 310.950 173.400 318.450 174.450 ;
        RECT 310.950 172.650 313.050 173.400 ;
        RECT 274.950 163.950 277.050 166.050 ;
        RECT 271.950 144.450 276.000 145.050 ;
        RECT 271.950 142.950 276.450 144.450 ;
        RECT 295.950 142.950 298.050 145.050 ;
        RECT 275.400 141.450 276.450 142.950 ;
        RECT 275.400 140.400 279.450 141.450 ;
        RECT 263.400 130.050 264.450 137.100 ;
        RECT 268.950 136.950 271.050 139.050 ;
        RECT 271.950 137.100 274.050 139.200 ;
        RECT 278.400 138.600 279.450 140.400 ;
        RECT 296.400 138.600 297.450 142.950 ;
        RECT 272.400 136.350 273.600 137.100 ;
        RECT 278.400 136.350 279.600 138.600 ;
        RECT 296.400 136.350 297.600 138.600 ;
        RECT 307.950 137.100 310.050 139.200 ;
        RECT 313.950 137.100 316.050 139.200 ;
        RECT 319.950 137.100 322.050 139.200 ;
        RECT 271.950 133.950 274.050 136.050 ;
        RECT 274.950 133.950 277.050 136.050 ;
        RECT 277.950 133.950 280.050 136.050 ;
        RECT 280.950 133.950 283.050 136.050 ;
        RECT 295.950 133.950 298.050 136.050 ;
        RECT 298.950 133.950 301.050 136.050 ;
        RECT 275.400 131.400 276.600 133.650 ;
        RECT 281.400 132.900 282.600 133.650 ;
        RECT 299.400 132.900 300.600 133.650 ;
        RECT 262.950 127.950 265.050 130.050 ;
        RECT 259.950 109.950 262.050 112.050 ;
        RECT 247.950 104.100 250.050 106.200 ;
        RECT 256.950 104.100 259.050 106.200 ;
        RECT 263.400 105.600 264.450 127.950 ;
        RECT 275.400 106.200 276.450 131.400 ;
        RECT 280.950 130.800 283.050 132.900 ;
        RECT 298.950 130.800 301.050 132.900 ;
        RECT 299.400 118.050 300.450 130.800 ;
        RECT 286.950 115.950 289.050 118.050 ;
        RECT 298.950 115.950 301.050 118.050 ;
        RECT 248.400 94.050 249.450 104.100 ;
        RECT 257.400 103.350 258.600 104.100 ;
        RECT 263.400 103.350 264.600 105.600 ;
        RECT 274.950 104.100 277.050 106.200 ;
        RECT 280.950 104.100 283.050 106.200 ;
        RECT 287.400 105.600 288.450 115.950 ;
        RECT 292.950 109.950 295.050 112.050 ;
        RECT 281.400 103.350 282.600 104.100 ;
        RECT 287.400 103.350 288.600 105.600 ;
        RECT 253.950 100.950 256.050 103.050 ;
        RECT 256.950 100.950 259.050 103.050 ;
        RECT 259.950 100.950 262.050 103.050 ;
        RECT 262.950 100.950 265.050 103.050 ;
        RECT 265.950 100.950 268.050 103.050 ;
        RECT 280.950 100.950 283.050 103.050 ;
        RECT 283.950 100.950 286.050 103.050 ;
        RECT 286.950 100.950 289.050 103.050 ;
        RECT 254.400 99.900 255.600 100.650 ;
        RECT 260.400 99.900 261.600 100.650 ;
        RECT 253.950 97.800 256.050 99.900 ;
        RECT 259.950 97.800 262.050 99.900 ;
        RECT 266.400 98.400 267.600 100.650 ;
        RECT 284.400 99.000 285.600 100.650 ;
        RECT 247.950 91.950 250.050 94.050 ;
        RECT 266.400 88.050 267.450 98.400 ;
        RECT 283.950 94.950 286.050 99.000 ;
        RECT 293.400 97.050 294.450 109.950 ;
        RECT 295.950 104.100 298.050 106.200 ;
        RECT 301.950 104.100 304.050 106.200 ;
        RECT 308.400 105.600 309.450 137.100 ;
        RECT 314.400 136.350 315.600 137.100 ;
        RECT 320.400 136.350 321.600 137.100 ;
        RECT 313.950 133.950 316.050 136.050 ;
        RECT 316.950 133.950 319.050 136.050 ;
        RECT 319.950 133.950 322.050 136.050 ;
        RECT 317.400 132.900 318.600 133.650 ;
        RECT 329.400 133.050 330.450 175.950 ;
        RECT 331.950 175.800 334.050 177.900 ;
        RECT 337.950 175.800 340.050 177.900 ;
        RECT 338.400 154.050 339.450 175.800 ;
        RECT 344.400 175.050 345.450 190.950 ;
        RECT 343.950 172.950 346.050 175.050 ;
        RECT 337.950 151.950 340.050 154.050 ;
        RECT 347.400 139.200 348.450 209.400 ;
        RECT 350.400 187.050 351.450 235.950 ;
        RECT 361.950 220.950 364.050 223.050 ;
        RECT 362.400 216.600 363.450 220.950 ;
        RECT 362.400 214.350 363.600 216.600 ;
        RECT 358.950 211.950 361.050 214.050 ;
        RECT 361.950 211.950 364.050 214.050 ;
        RECT 359.400 210.900 360.600 211.650 ;
        RECT 377.400 211.050 378.450 247.950 ;
        RECT 407.400 247.050 408.450 254.400 ;
        RECT 406.950 244.950 409.050 247.050 ;
        RECT 406.950 226.950 409.050 229.050 ;
        RECT 398.250 223.500 400.350 224.400 ;
        RECT 396.150 222.300 400.350 223.500 ;
        RECT 391.950 216.000 394.050 220.050 ;
        RECT 392.400 214.350 393.600 216.000 ;
        RECT 380.100 211.950 382.200 214.050 ;
        RECT 385.500 211.950 387.600 214.050 ;
        RECT 391.950 211.950 394.050 214.050 ;
        RECT 358.950 208.800 361.050 210.900 ;
        RECT 376.950 208.950 379.050 211.050 ;
        RECT 386.400 210.900 387.600 211.650 ;
        RECT 385.950 208.800 388.050 210.900 ;
        RECT 373.950 205.950 376.050 208.050 ;
        RECT 361.950 187.950 364.050 190.050 ;
        RECT 367.950 187.950 370.050 190.050 ;
        RECT 349.950 184.950 352.050 187.050 ;
        RECT 355.950 182.100 358.050 184.200 ;
        RECT 362.400 183.600 363.450 187.950 ;
        RECT 356.400 181.350 357.600 182.100 ;
        RECT 362.400 181.350 363.600 183.600 ;
        RECT 352.950 178.950 355.050 181.050 ;
        RECT 355.950 178.950 358.050 181.050 ;
        RECT 358.950 178.950 361.050 181.050 ;
        RECT 361.950 178.950 364.050 181.050 ;
        RECT 349.950 175.950 352.050 178.050 ;
        RECT 353.400 177.000 354.600 178.650 ;
        RECT 359.400 177.900 360.600 178.650 ;
        RECT 368.400 177.900 369.450 187.950 ;
        RECT 374.400 178.050 375.450 205.950 ;
        RECT 396.150 203.700 397.350 222.300 ;
        RECT 400.950 215.100 403.050 217.200 ;
        RECT 401.400 214.350 402.600 215.100 ;
        RECT 401.100 211.950 403.200 214.050 ;
        RECT 403.950 208.950 406.050 211.050 ;
        RECT 395.850 201.600 397.950 203.700 ;
        RECT 382.950 182.100 385.050 184.200 ;
        RECT 383.400 181.350 384.600 182.100 ;
        RECT 391.950 181.950 394.050 184.050 ;
        RECT 404.400 183.600 405.450 208.950 ;
        RECT 407.400 186.450 408.450 226.950 ;
        RECT 410.400 199.050 411.450 254.400 ;
        RECT 416.400 241.050 417.450 256.950 ;
        RECT 419.400 255.900 420.450 259.950 ;
        RECT 428.400 259.350 429.600 261.600 ;
        RECT 433.950 260.100 436.050 262.200 ;
        RECT 434.400 259.350 435.600 260.100 ;
        RECT 424.950 256.950 427.050 259.050 ;
        RECT 427.950 256.950 430.050 259.050 ;
        RECT 430.950 256.950 433.050 259.050 ;
        RECT 433.950 256.950 436.050 259.050 ;
        RECT 418.950 253.800 421.050 255.900 ;
        RECT 421.950 253.950 424.050 256.050 ;
        RECT 425.400 255.900 426.600 256.650 ;
        RECT 422.400 250.050 423.450 253.950 ;
        RECT 424.950 253.800 427.050 255.900 ;
        RECT 431.400 254.400 432.600 256.650 ;
        RECT 418.800 247.950 420.900 250.050 ;
        RECT 421.950 247.950 424.050 250.050 ;
        RECT 427.950 247.950 430.050 250.050 ;
        RECT 415.950 238.950 418.050 241.050 ;
        RECT 419.400 229.050 420.450 247.950 ;
        RECT 424.950 238.950 427.050 241.050 ;
        RECT 413.550 225.300 415.650 227.400 ;
        RECT 418.950 226.950 421.050 229.050 ;
        RECT 413.550 218.700 414.750 225.300 ;
        RECT 413.550 216.600 415.650 218.700 ;
        RECT 413.550 203.700 414.750 216.600 ;
        RECT 418.950 211.950 421.050 214.050 ;
        RECT 419.400 210.000 420.600 211.650 ;
        RECT 418.950 205.950 421.050 210.000 ;
        RECT 413.550 201.600 415.650 203.700 ;
        RECT 409.950 196.950 412.050 199.050 ;
        RECT 415.950 196.950 418.050 199.050 ;
        RECT 407.400 185.400 411.450 186.450 ;
        RECT 410.400 184.200 411.450 185.400 ;
        RECT 379.950 178.950 382.050 181.050 ;
        RECT 382.950 178.950 385.050 181.050 ;
        RECT 385.950 178.950 388.050 181.050 ;
        RECT 337.950 137.100 340.050 139.200 ;
        RECT 346.950 137.100 349.050 139.200 ;
        RECT 338.400 136.350 339.600 137.100 ;
        RECT 337.950 133.950 340.050 136.050 ;
        RECT 340.950 133.950 343.050 136.050 ;
        RECT 316.950 130.800 319.050 132.900 ;
        RECT 328.950 130.950 331.050 133.050 ;
        RECT 341.400 131.400 342.600 133.650 ;
        RECT 341.400 121.050 342.450 131.400 ;
        RECT 340.950 118.950 343.050 121.050 ;
        RECT 341.400 112.050 342.450 118.950 ;
        RECT 340.950 109.950 343.050 112.050 ;
        RECT 346.950 109.950 349.050 112.050 ;
        RECT 316.950 106.950 319.050 109.050 ;
        RECT 296.400 100.050 297.450 104.100 ;
        RECT 302.400 103.350 303.600 104.100 ;
        RECT 308.400 103.350 309.600 105.600 ;
        RECT 301.950 100.950 304.050 103.050 ;
        RECT 304.950 100.950 307.050 103.050 ;
        RECT 307.950 100.950 310.050 103.050 ;
        RECT 310.950 100.950 313.050 103.050 ;
        RECT 295.950 97.950 298.050 100.050 ;
        RECT 305.400 99.900 306.600 100.650 ;
        RECT 304.950 97.800 307.050 99.900 ;
        RECT 311.400 99.000 312.600 100.650 ;
        RECT 317.400 100.050 318.450 106.950 ;
        RECT 328.950 104.100 331.050 106.200 ;
        RECT 337.950 105.000 340.050 109.050 ;
        RECT 329.400 103.350 330.600 104.100 ;
        RECT 338.400 103.350 339.600 105.000 ;
        RECT 328.800 100.950 330.900 103.050 ;
        RECT 334.950 100.950 337.050 103.050 ;
        RECT 337.950 100.950 340.050 103.050 ;
        RECT 343.500 100.950 345.600 103.050 ;
        RECT 292.950 94.950 295.050 97.050 ;
        RECT 303.000 96.750 306.000 97.050 ;
        RECT 301.950 94.950 307.050 96.750 ;
        RECT 310.950 94.950 313.050 99.000 ;
        RECT 316.950 97.950 319.050 100.050 ;
        RECT 335.400 99.000 336.600 100.650 ;
        RECT 344.400 99.450 345.600 100.650 ;
        RECT 347.400 99.450 348.450 109.950 ;
        RECT 334.950 94.950 337.050 99.000 ;
        RECT 344.400 98.400 348.450 99.450 ;
        RECT 301.950 94.650 304.050 94.950 ;
        RECT 304.950 94.650 307.050 94.950 ;
        RECT 244.950 85.950 247.050 88.050 ;
        RECT 265.950 85.950 268.050 88.050 ;
        RECT 232.950 73.950 235.050 76.050 ;
        RECT 220.950 70.950 223.050 73.050 ;
        RECT 203.400 58.350 204.600 60.600 ;
        RECT 209.400 58.350 210.600 60.600 ;
        RECT 226.950 60.000 229.050 64.050 ;
        RECT 233.400 60.600 234.450 73.950 ;
        RECT 259.950 70.950 262.050 73.050 ;
        RECT 268.950 70.950 271.050 73.050 ;
        RECT 247.950 64.950 250.050 67.050 ;
        RECT 227.400 58.350 228.600 60.000 ;
        RECT 233.400 58.350 234.600 60.600 ;
        RECT 238.950 59.100 241.050 61.200 ;
        RECT 244.950 59.100 247.050 61.200 ;
        RECT 239.400 58.350 240.600 59.100 ;
        RECT 202.950 55.950 205.050 58.050 ;
        RECT 205.950 55.950 208.050 58.050 ;
        RECT 208.950 55.950 211.050 58.050 ;
        RECT 211.950 55.950 214.050 58.050 ;
        RECT 226.950 55.950 229.050 58.050 ;
        RECT 229.950 55.950 232.050 58.050 ;
        RECT 232.950 55.950 235.050 58.050 ;
        RECT 235.950 55.950 238.050 58.050 ;
        RECT 238.950 55.950 241.050 58.050 ;
        RECT 206.400 54.900 207.600 55.650 ;
        RECT 212.400 54.900 213.600 55.650 ;
        RECT 230.400 54.900 231.600 55.650 ;
        RECT 196.950 52.800 199.050 54.900 ;
        RECT 205.950 52.800 208.050 54.900 ;
        RECT 211.950 52.800 214.050 54.900 ;
        RECT 229.950 52.800 232.050 54.900 ;
        RECT 236.400 53.400 237.600 55.650 ;
        RECT 133.950 46.950 136.050 49.050 ;
        RECT 236.400 43.050 237.450 53.400 ;
        RECT 245.400 43.050 246.450 59.100 ;
        RECT 248.400 49.050 249.450 64.950 ;
        RECT 253.950 59.100 256.050 61.200 ;
        RECT 260.400 60.600 261.450 70.950 ;
        RECT 254.400 58.350 255.600 59.100 ;
        RECT 260.400 58.350 261.600 60.600 ;
        RECT 253.950 55.950 256.050 58.050 ;
        RECT 256.950 55.950 259.050 58.050 ;
        RECT 259.950 55.950 262.050 58.050 ;
        RECT 262.950 55.950 265.050 58.050 ;
        RECT 257.400 54.900 258.600 55.650 ;
        RECT 263.400 54.900 264.600 55.650 ;
        RECT 269.400 55.050 270.450 70.950 ;
        RECT 304.950 64.950 307.050 67.050 ;
        RECT 337.950 64.950 340.050 67.050 ;
        RECT 271.950 59.100 274.050 61.200 ;
        RECT 280.950 59.100 283.050 61.200 ;
        RECT 286.950 59.100 289.050 61.200 ;
        RECT 305.400 60.600 306.450 64.950 ;
        RECT 256.950 52.800 259.050 54.900 ;
        RECT 262.950 52.800 265.050 54.900 ;
        RECT 268.950 52.950 271.050 55.050 ;
        RECT 247.950 46.950 250.050 49.050 ;
        RECT 187.950 40.950 190.050 43.050 ;
        RECT 208.950 40.950 211.050 43.050 ;
        RECT 235.950 40.950 238.050 43.050 ;
        RECT 244.950 40.950 247.050 43.050 ;
        RECT 145.950 37.950 148.050 40.050 ;
        RECT 175.950 37.950 178.050 40.050 ;
        RECT 136.950 34.950 139.050 37.050 ;
        RECT 130.950 26.100 133.050 28.200 ;
        RECT 137.400 27.600 138.450 34.950 ;
        RECT 131.400 25.350 132.600 26.100 ;
        RECT 137.400 25.350 138.600 27.600 ;
        RECT 127.950 22.950 130.050 25.050 ;
        RECT 130.950 22.950 133.050 25.050 ;
        RECT 133.950 22.950 136.050 25.050 ;
        RECT 136.950 22.950 139.050 25.050 ;
        RECT 97.950 19.800 100.050 21.900 ;
        RECT 103.950 19.800 106.050 21.900 ;
        RECT 109.950 19.800 112.050 21.900 ;
        RECT 121.950 19.800 124.050 21.900 ;
        RECT 128.400 21.000 129.600 22.650 ;
        RECT 127.950 16.950 130.050 21.000 ;
        RECT 134.400 20.400 135.600 22.650 ;
        RECT 146.400 21.900 147.450 37.950 ;
        RECT 154.950 26.100 157.050 28.200 ;
        RECT 160.950 26.100 163.050 28.200 ;
        RECT 176.400 27.600 177.450 37.950 ;
        RECT 155.400 25.350 156.600 26.100 ;
        RECT 161.400 25.350 162.600 26.100 ;
        RECT 176.400 25.350 177.600 27.600 ;
        RECT 151.950 22.950 154.050 25.050 ;
        RECT 154.950 22.950 157.050 25.050 ;
        RECT 157.950 22.950 160.050 25.050 ;
        RECT 160.950 22.950 163.050 25.050 ;
        RECT 175.950 22.950 178.050 25.050 ;
        RECT 178.950 22.950 181.050 25.050 ;
        RECT 134.400 16.050 135.450 20.400 ;
        RECT 145.950 19.800 148.050 21.900 ;
        RECT 152.400 20.400 153.600 22.650 ;
        RECT 158.400 21.900 159.600 22.650 ;
        RECT 152.400 16.050 153.450 20.400 ;
        RECT 157.950 19.800 160.050 21.900 ;
        RECT 179.400 21.000 180.600 22.650 ;
        RECT 188.400 21.900 189.450 40.950 ;
        RECT 196.950 31.950 199.050 34.050 ;
        RECT 197.400 27.600 198.450 31.950 ;
        RECT 197.400 25.350 198.600 27.600 ;
        RECT 202.950 26.100 205.050 28.200 ;
        RECT 203.400 25.350 204.600 26.100 ;
        RECT 209.400 25.050 210.450 40.950 ;
        RECT 257.400 34.050 258.450 52.800 ;
        RECT 262.950 46.950 265.050 49.050 ;
        RECT 220.950 31.950 223.050 34.050 ;
        RECT 250.950 31.950 253.050 34.050 ;
        RECT 256.950 31.950 259.050 34.050 ;
        RECT 211.950 25.950 214.050 28.050 ;
        RECT 221.400 27.600 222.450 31.950 ;
        RECT 193.950 22.950 196.050 25.050 ;
        RECT 196.950 22.950 199.050 25.050 ;
        RECT 199.950 22.950 202.050 25.050 ;
        RECT 202.950 22.950 205.050 25.050 ;
        RECT 208.950 22.950 211.050 25.050 ;
        RECT 194.400 21.900 195.600 22.650 ;
        RECT 178.950 16.950 181.050 21.000 ;
        RECT 187.950 19.800 190.050 21.900 ;
        RECT 193.950 19.800 196.050 21.900 ;
        RECT 200.400 21.000 201.600 22.650 ;
        RECT 212.400 21.900 213.450 25.950 ;
        RECT 221.400 25.350 222.600 27.600 ;
        RECT 226.950 27.000 229.050 31.050 ;
        RECT 227.400 25.350 228.600 27.000 ;
        RECT 244.950 26.100 247.050 28.200 ;
        RECT 251.400 27.600 252.450 31.950 ;
        RECT 259.950 28.950 262.050 31.050 ;
        RECT 245.400 25.350 246.600 26.100 ;
        RECT 251.400 25.350 252.600 27.600 ;
        RECT 217.950 22.950 220.050 25.050 ;
        RECT 220.950 22.950 223.050 25.050 ;
        RECT 223.950 22.950 226.050 25.050 ;
        RECT 226.950 22.950 229.050 25.050 ;
        RECT 244.950 22.950 247.050 25.050 ;
        RECT 247.950 22.950 250.050 25.050 ;
        RECT 250.950 22.950 253.050 25.050 ;
        RECT 253.950 22.950 256.050 25.050 ;
        RECT 218.400 22.050 219.600 22.650 ;
        RECT 199.950 16.950 202.050 21.000 ;
        RECT 211.950 19.800 214.050 21.900 ;
        RECT 214.950 20.400 219.600 22.050 ;
        RECT 224.400 21.000 225.600 22.650 ;
        RECT 248.400 21.900 249.600 22.650 ;
        RECT 254.400 22.050 255.600 22.650 ;
        RECT 214.950 19.950 219.000 20.400 ;
        RECT 205.950 16.950 211.050 19.050 ;
        RECT 223.950 16.950 226.050 21.000 ;
        RECT 247.950 19.800 250.050 21.900 ;
        RECT 254.400 20.400 259.050 22.050 ;
        RECT 260.400 21.900 261.450 28.950 ;
        RECT 263.400 22.050 264.450 46.950 ;
        RECT 268.950 40.950 271.050 43.050 ;
        RECT 269.400 27.600 270.450 40.950 ;
        RECT 272.400 31.050 273.450 59.100 ;
        RECT 281.400 58.350 282.600 59.100 ;
        RECT 287.400 58.350 288.600 59.100 ;
        RECT 305.400 58.350 306.600 60.600 ;
        RECT 310.950 59.100 313.050 61.200 ;
        RECT 322.950 59.100 325.050 61.200 ;
        RECT 331.950 59.100 334.050 61.200 ;
        RECT 338.400 60.600 339.450 64.950 ;
        RECT 311.400 58.350 312.600 59.100 ;
        RECT 280.950 55.950 283.050 58.050 ;
        RECT 283.950 55.950 286.050 58.050 ;
        RECT 286.950 55.950 289.050 58.050 ;
        RECT 289.950 55.950 292.050 58.050 ;
        RECT 295.950 55.950 298.050 58.050 ;
        RECT 304.950 55.950 307.050 58.050 ;
        RECT 307.950 55.950 310.050 58.050 ;
        RECT 310.950 55.950 313.050 58.050 ;
        RECT 313.950 55.950 316.050 58.050 ;
        RECT 284.400 53.400 285.600 55.650 ;
        RECT 290.400 54.900 291.600 55.650 ;
        RECT 274.950 37.950 277.050 40.050 ;
        RECT 271.950 28.950 274.050 31.050 ;
        RECT 275.400 27.600 276.450 37.950 ;
        RECT 284.400 37.050 285.450 53.400 ;
        RECT 289.950 52.800 292.050 54.900 ;
        RECT 296.400 49.050 297.450 55.950 ;
        RECT 308.400 54.900 309.600 55.650 ;
        RECT 307.950 52.800 310.050 54.900 ;
        RECT 314.400 53.400 315.600 55.650 ;
        RECT 295.950 46.950 298.050 49.050 ;
        RECT 314.400 46.050 315.450 53.400 ;
        RECT 313.950 43.950 316.050 46.050 ;
        RECT 310.950 37.950 313.050 40.050 ;
        RECT 283.950 34.950 286.050 37.050 ;
        RECT 301.950 34.950 304.050 37.050 ;
        RECT 269.400 25.350 270.600 27.600 ;
        RECT 275.400 25.350 276.600 27.600 ;
        RECT 268.950 22.950 271.050 25.050 ;
        RECT 271.950 22.950 274.050 25.050 ;
        RECT 274.950 22.950 277.050 25.050 ;
        RECT 277.950 22.950 280.050 25.050 ;
        RECT 255.000 19.950 259.050 20.400 ;
        RECT 259.950 19.800 262.050 21.900 ;
        RECT 262.950 19.950 265.050 22.050 ;
        RECT 272.400 21.900 273.600 22.650 ;
        RECT 278.400 21.900 279.600 22.650 ;
        RECT 284.400 21.900 285.450 34.950 ;
        RECT 286.950 25.950 289.050 28.050 ;
        RECT 295.950 26.100 298.050 28.200 ;
        RECT 302.400 27.600 303.450 34.950 ;
        RECT 311.400 28.050 312.450 37.950 ;
        RECT 271.950 19.800 274.050 21.900 ;
        RECT 277.950 19.800 280.050 21.900 ;
        RECT 283.950 19.800 286.050 21.900 ;
        RECT 106.950 13.950 112.050 16.050 ;
        RECT 133.950 13.950 136.050 16.050 ;
        RECT 151.950 13.950 154.050 16.050 ;
        RECT 248.400 13.050 249.450 19.800 ;
        RECT 287.400 16.050 288.450 25.950 ;
        RECT 296.400 25.350 297.600 26.100 ;
        RECT 302.400 25.350 303.600 27.600 ;
        RECT 310.950 25.950 313.050 28.050 ;
        RECT 316.950 26.100 319.050 28.200 ;
        RECT 323.400 27.600 324.450 59.100 ;
        RECT 332.400 58.350 333.600 59.100 ;
        RECT 338.400 58.350 339.600 60.600 ;
        RECT 331.950 55.950 334.050 58.050 ;
        RECT 334.950 55.950 337.050 58.050 ;
        RECT 337.950 55.950 340.050 58.050 ;
        RECT 340.950 55.950 343.050 58.050 ;
        RECT 335.400 54.900 336.600 55.650 ;
        RECT 341.400 54.900 342.600 55.650 ;
        RECT 334.950 52.800 337.050 54.900 ;
        RECT 340.950 52.800 343.050 54.900 ;
        RECT 331.950 34.950 334.050 37.050 ;
        RECT 317.400 25.350 318.600 26.100 ;
        RECT 323.400 25.350 324.600 27.600 ;
        RECT 292.950 22.950 295.050 25.050 ;
        RECT 295.950 22.950 298.050 25.050 ;
        RECT 298.950 22.950 301.050 25.050 ;
        RECT 301.950 22.950 304.050 25.050 ;
        RECT 316.950 22.950 319.050 25.050 ;
        RECT 319.950 22.950 322.050 25.050 ;
        RECT 322.950 22.950 325.050 25.050 ;
        RECT 325.950 22.950 328.050 25.050 ;
        RECT 293.400 21.900 294.600 22.650 ;
        RECT 299.400 21.900 300.600 22.650 ;
        RECT 292.950 19.800 295.050 21.900 ;
        RECT 298.950 19.800 301.050 21.900 ;
        RECT 320.400 21.000 321.600 22.650 ;
        RECT 326.400 21.450 327.600 22.650 ;
        RECT 332.400 21.450 333.450 34.950 ;
        RECT 350.400 34.050 351.450 175.950 ;
        RECT 352.950 172.950 355.050 177.000 ;
        RECT 358.950 175.800 361.050 177.900 ;
        RECT 367.950 175.800 370.050 177.900 ;
        RECT 373.950 175.950 376.050 178.050 ;
        RECT 380.400 177.900 381.600 178.650 ;
        RECT 386.400 177.900 387.600 178.650 ;
        RECT 379.950 175.800 382.050 177.900 ;
        RECT 385.950 175.800 388.050 177.900 ;
        RECT 392.400 175.050 393.450 181.950 ;
        RECT 404.400 181.350 405.600 183.600 ;
        RECT 409.950 182.100 412.050 184.200 ;
        RECT 410.400 181.350 411.600 182.100 ;
        RECT 400.950 178.950 403.050 181.050 ;
        RECT 403.950 178.950 406.050 181.050 ;
        RECT 406.950 178.950 409.050 181.050 ;
        RECT 409.950 178.950 412.050 181.050 ;
        RECT 401.400 177.000 402.600 178.650 ;
        RECT 391.950 172.950 394.050 175.050 ;
        RECT 400.950 172.950 403.050 177.000 ;
        RECT 407.400 176.400 408.600 178.650 ;
        RECT 403.950 172.950 406.050 175.050 ;
        RECT 382.950 160.950 385.050 163.050 ;
        RECT 383.400 154.050 384.450 160.950 ;
        RECT 382.950 151.950 385.050 154.050 ;
        RECT 358.950 137.100 361.050 139.200 ;
        RECT 359.400 136.350 360.600 137.100 ;
        RECT 370.950 136.950 373.050 139.050 ;
        RECT 383.400 138.600 384.450 151.950 ;
        RECT 358.950 133.950 361.050 136.050 ;
        RECT 361.950 133.950 364.050 136.050 ;
        RECT 364.950 133.950 367.050 136.050 ;
        RECT 362.400 131.400 363.600 133.650 ;
        RECT 362.400 118.050 363.450 131.400 ;
        RECT 361.950 115.950 364.050 118.050 ;
        RECT 371.400 112.050 372.450 136.950 ;
        RECT 383.400 136.350 384.600 138.600 ;
        RECT 388.950 137.100 391.050 139.200 ;
        RECT 394.950 138.000 397.050 142.050 ;
        RECT 389.400 136.350 390.600 137.100 ;
        RECT 395.400 136.350 396.600 138.000 ;
        RECT 382.950 133.950 385.050 136.050 ;
        RECT 385.950 133.950 388.050 136.050 ;
        RECT 388.950 133.950 391.050 136.050 ;
        RECT 391.950 133.950 394.050 136.050 ;
        RECT 394.950 133.950 397.050 136.050 ;
        RECT 404.400 133.050 405.450 172.950 ;
        RECT 397.950 130.950 400.050 133.050 ;
        RECT 403.950 130.950 406.050 133.050 ;
        RECT 379.950 118.950 382.050 121.050 ;
        RECT 388.950 118.950 391.050 121.050 ;
        RECT 380.400 112.050 381.450 118.950 ;
        RECT 382.950 115.950 385.050 118.050 ;
        RECT 361.950 109.950 364.050 112.050 ;
        RECT 370.950 109.950 373.050 112.050 ;
        RECT 379.950 109.950 382.050 112.050 ;
        RECT 362.400 105.600 363.450 109.950 ;
        RECT 362.400 103.350 363.600 105.600 ;
        RECT 367.950 105.000 370.050 109.050 ;
        RECT 376.950 106.950 379.050 109.050 ;
        RECT 368.400 103.350 369.600 105.000 ;
        RECT 361.950 100.950 364.050 103.050 ;
        RECT 364.950 100.950 367.050 103.050 ;
        RECT 367.950 100.950 370.050 103.050 ;
        RECT 365.400 98.400 366.600 100.650 ;
        RECT 358.950 79.950 361.050 82.050 ;
        RECT 355.950 70.950 358.050 73.050 ;
        RECT 352.950 64.950 355.050 67.050 ;
        RECT 353.400 55.050 354.450 64.950 ;
        RECT 356.400 61.200 357.450 70.950 ;
        RECT 355.950 59.100 358.050 61.200 ;
        RECT 359.400 60.600 360.450 79.950 ;
        RECT 365.400 70.050 366.450 98.400 ;
        RECT 377.400 82.050 378.450 106.950 ;
        RECT 383.400 105.600 384.450 115.950 ;
        RECT 389.400 105.600 390.450 118.950 ;
        RECT 383.400 103.350 384.600 105.600 ;
        RECT 389.400 103.350 390.600 105.600 ;
        RECT 382.950 100.950 385.050 103.050 ;
        RECT 385.950 100.950 388.050 103.050 ;
        RECT 388.950 100.950 391.050 103.050 ;
        RECT 386.400 98.400 387.600 100.650 ;
        RECT 398.400 99.450 399.450 130.950 ;
        RECT 407.400 118.050 408.450 176.400 ;
        RECT 416.400 175.050 417.450 196.950 ;
        RECT 425.400 190.050 426.450 238.950 ;
        RECT 428.400 199.050 429.450 247.950 ;
        RECT 431.400 247.050 432.450 254.400 ;
        RECT 433.950 250.950 436.050 253.050 ;
        RECT 430.950 244.950 433.050 247.050 ;
        RECT 430.950 215.100 433.050 217.200 ;
        RECT 431.400 208.050 432.450 215.100 ;
        RECT 434.400 211.050 435.450 250.950 ;
        RECT 440.400 250.050 441.450 265.950 ;
        RECT 443.400 253.050 444.450 268.950 ;
        RECT 455.400 265.050 456.450 299.400 ;
        RECT 460.950 293.100 463.050 295.200 ;
        RECT 461.400 292.350 462.600 293.100 ;
        RECT 460.950 289.950 463.050 292.050 ;
        RECT 463.950 289.950 466.050 292.050 ;
        RECT 464.400 288.000 465.600 289.650 ;
        RECT 463.950 283.950 466.050 288.000 ;
        RECT 466.950 286.950 469.050 289.050 ;
        RECT 470.400 288.900 471.450 313.950 ;
        RECT 472.950 304.950 475.050 307.050 ;
        RECT 467.400 274.050 468.450 286.950 ;
        RECT 469.950 286.800 472.050 288.900 ;
        RECT 466.950 271.950 469.050 274.050 ;
        RECT 464.850 267.300 466.950 269.400 ;
        RECT 454.950 262.950 457.050 265.050 ;
        RECT 451.950 260.100 454.050 262.200 ;
        RECT 452.400 259.350 453.600 260.100 ;
        RECT 448.950 256.950 451.050 259.050 ;
        RECT 451.950 256.950 454.050 259.050 ;
        RECT 454.950 256.950 457.050 259.050 ;
        RECT 460.950 256.950 463.050 259.050 ;
        RECT 449.400 254.400 450.600 256.650 ;
        RECT 461.400 255.900 462.600 256.650 ;
        RECT 442.950 250.950 445.050 253.050 ;
        RECT 439.950 247.950 442.050 250.050 ;
        RECT 449.400 247.050 450.450 254.400 ;
        RECT 460.950 253.800 463.050 255.900 ;
        RECT 465.150 248.700 466.350 267.300 ;
        RECT 473.400 262.050 474.450 304.950 ;
        RECT 484.950 301.950 487.050 304.050 ;
        RECT 475.950 294.600 480.000 295.050 ;
        RECT 485.400 294.600 486.450 301.950 ;
        RECT 475.950 292.950 480.600 294.600 ;
        RECT 479.400 292.350 480.600 292.950 ;
        RECT 485.400 292.350 486.600 294.600 ;
        RECT 478.950 289.950 481.050 292.050 ;
        RECT 481.950 289.950 484.050 292.050 ;
        RECT 484.950 289.950 487.050 292.050 ;
        RECT 487.950 289.950 490.050 292.050 ;
        RECT 482.400 288.900 483.600 289.650 ;
        RECT 488.400 288.900 489.600 289.650 ;
        RECT 494.400 289.050 495.450 349.950 ;
        RECT 503.400 339.600 504.450 349.950 ;
        RECT 503.400 337.350 504.600 339.600 ;
        RECT 499.950 334.950 502.050 337.050 ;
        RECT 502.950 334.950 505.050 337.050 ;
        RECT 505.950 334.950 508.050 337.050 ;
        RECT 500.400 333.900 501.600 334.650 ;
        RECT 499.950 331.800 502.050 333.900 ;
        RECT 506.400 332.400 507.600 334.650 ;
        RECT 496.950 325.950 499.050 328.050 ;
        RECT 481.950 286.800 484.050 288.900 ;
        RECT 487.950 286.800 490.050 288.900 ;
        RECT 493.950 286.950 496.050 289.050 ;
        RECT 488.400 271.050 489.450 286.800 ;
        RECT 478.950 268.950 481.050 271.050 ;
        RECT 475.950 262.950 478.050 265.050 ;
        RECT 472.950 259.950 475.050 262.050 ;
        RECT 470.100 256.950 472.200 259.050 ;
        RECT 470.400 255.000 471.600 256.650 ;
        RECT 469.950 253.050 472.050 255.000 ;
        RECT 469.800 252.000 472.050 253.050 ;
        RECT 469.800 250.950 471.900 252.000 ;
        RECT 472.950 250.950 475.050 253.050 ;
        RECT 465.150 247.500 469.350 248.700 ;
        RECT 448.950 244.950 451.050 247.050 ;
        RECT 467.250 246.600 469.350 247.500 ;
        RECT 473.400 244.050 474.450 250.950 ;
        RECT 476.400 247.050 477.450 262.950 ;
        RECT 479.400 253.050 480.450 268.950 ;
        RECT 482.550 267.300 484.650 269.400 ;
        RECT 487.950 268.950 490.050 271.050 ;
        RECT 482.550 254.400 483.750 267.300 ;
        RECT 487.950 260.100 490.050 262.200 ;
        RECT 488.400 259.350 489.600 260.100 ;
        RECT 487.950 256.950 490.050 259.050 ;
        RECT 478.950 250.950 481.050 253.050 ;
        RECT 482.550 252.300 484.650 254.400 ;
        RECT 490.950 253.950 493.050 256.050 ;
        RECT 497.400 255.900 498.450 325.950 ;
        RECT 500.400 295.050 501.450 331.800 ;
        RECT 502.950 301.950 505.050 304.050 ;
        RECT 499.950 292.950 502.050 295.050 ;
        RECT 503.400 294.600 504.450 301.950 ;
        RECT 506.400 298.050 507.450 332.400 ;
        RECT 515.400 328.050 516.450 370.950 ;
        RECT 518.400 361.050 519.450 406.950 ;
        RECT 524.400 387.450 525.450 410.400 ;
        RECT 527.400 391.050 528.450 424.950 ;
        RECT 541.950 417.000 544.050 421.050 ;
        RECT 542.400 415.350 543.600 417.000 ;
        RECT 547.950 416.100 550.050 418.200 ;
        RECT 551.400 418.050 552.450 436.950 ;
        RECT 554.400 418.200 555.450 442.950 ;
        RECT 560.400 439.050 561.450 443.400 ;
        RECT 559.950 436.950 562.050 439.050 ;
        RECT 566.250 437.700 567.450 450.600 ;
        RECT 569.400 445.050 570.450 505.950 ;
        RECT 583.050 501.300 585.150 503.400 ;
        RECT 577.800 490.950 579.900 493.050 ;
        RECT 578.400 489.900 579.600 490.650 ;
        RECT 577.950 487.800 580.050 489.900 ;
        RECT 583.650 482.700 584.850 501.300 ;
        RECT 590.400 495.450 591.450 520.950 ;
        RECT 593.400 514.050 594.450 553.800 ;
        RECT 599.400 535.050 600.450 566.400 ;
        RECT 603.150 560.700 604.350 579.300 ;
        RECT 611.400 574.050 612.450 583.950 ;
        RECT 614.400 580.050 615.450 584.400 ;
        RECT 616.950 580.950 619.050 583.050 ;
        RECT 613.950 577.950 616.050 580.050 ;
        RECT 613.950 574.800 616.050 576.900 ;
        RECT 610.950 571.950 613.050 574.050 ;
        RECT 608.100 568.950 610.200 571.050 ;
        RECT 608.400 567.900 609.600 568.650 ;
        RECT 607.950 565.800 610.050 567.900 ;
        RECT 603.150 559.500 607.350 560.700 ;
        RECT 605.250 558.600 607.350 559.500 ;
        RECT 614.400 559.050 615.450 574.800 ;
        RECT 617.400 562.050 618.450 580.950 ;
        RECT 620.550 579.300 622.650 581.400 ;
        RECT 620.550 566.400 621.750 579.300 ;
        RECT 626.400 573.450 627.600 573.600 ;
        RECT 629.400 573.450 630.450 605.400 ;
        RECT 635.400 604.350 636.600 605.400 ;
        RECT 640.950 605.100 643.050 607.200 ;
        RECT 649.950 605.100 652.050 607.200 ;
        RECT 655.950 605.100 658.050 607.200 ;
        RECT 662.400 606.600 663.450 610.950 ;
        RECT 641.400 604.350 642.600 605.100 ;
        RECT 634.950 601.950 637.050 604.050 ;
        RECT 637.950 601.950 640.050 604.050 ;
        RECT 640.950 601.950 643.050 604.050 ;
        RECT 631.950 595.950 634.050 601.050 ;
        RECT 638.400 600.900 639.600 601.650 ;
        RECT 637.950 598.800 640.050 600.900 ;
        RECT 634.950 595.950 637.050 598.050 ;
        RECT 626.400 572.400 633.450 573.450 ;
        RECT 626.400 571.350 627.600 572.400 ;
        RECT 625.950 568.950 628.050 571.050 ;
        RECT 620.550 564.300 622.650 566.400 ;
        RECT 616.950 559.950 619.050 562.050 ;
        RECT 613.950 556.950 616.050 559.050 ;
        RECT 620.550 557.700 621.750 564.300 ;
        RECT 620.550 555.600 622.650 557.700 ;
        RECT 632.400 541.050 633.450 572.400 ;
        RECT 604.950 538.950 607.050 541.050 ;
        RECT 631.950 538.950 634.050 541.050 ;
        RECT 598.950 532.950 601.050 535.050 ;
        RECT 598.950 528.000 601.050 531.900 ;
        RECT 605.400 528.600 606.450 538.950 ;
        RECT 613.950 532.950 616.050 535.050 ;
        RECT 610.950 529.950 613.050 532.050 ;
        RECT 599.400 526.350 600.600 528.000 ;
        RECT 605.400 526.350 606.600 528.600 ;
        RECT 598.950 523.950 601.050 526.050 ;
        RECT 601.950 523.950 604.050 526.050 ;
        RECT 604.950 523.950 607.050 526.050 ;
        RECT 602.400 521.400 603.600 523.650 ;
        RECT 592.950 511.950 595.050 514.050 ;
        RECT 602.400 504.450 603.450 521.400 ;
        RECT 611.400 508.050 612.450 529.950 ;
        RECT 614.400 523.050 615.450 532.950 ;
        RECT 625.950 527.100 628.050 529.200 ;
        RECT 631.950 527.100 634.050 529.200 ;
        RECT 626.400 526.350 627.600 527.100 ;
        RECT 619.950 523.950 622.050 526.050 ;
        RECT 622.950 523.950 625.050 526.050 ;
        RECT 625.950 523.950 628.050 526.050 ;
        RECT 613.950 520.950 616.050 523.050 ;
        RECT 623.400 522.900 624.600 523.650 ;
        RECT 632.400 523.050 633.450 527.100 ;
        RECT 622.950 520.800 625.050 522.900 ;
        RECT 631.950 520.950 634.050 523.050 ;
        RECT 625.950 517.950 628.050 520.050 ;
        RECT 622.950 511.950 625.050 514.050 ;
        RECT 610.950 505.950 613.050 508.050 ;
        RECT 616.950 505.950 619.050 508.050 ;
        RECT 599.400 503.400 603.450 504.450 ;
        RECT 590.400 494.400 594.450 495.450 ;
        RECT 586.950 490.950 589.050 493.050 ;
        RECT 580.650 481.500 584.850 482.700 ;
        RECT 587.400 488.400 588.600 490.650 ;
        RECT 580.650 480.600 582.750 481.500 ;
        RECT 587.400 463.050 588.450 488.400 ;
        RECT 586.950 460.950 589.050 463.050 ;
        RECT 580.650 457.500 582.750 458.400 ;
        RECT 580.650 456.300 584.850 457.500 ;
        RECT 571.950 448.950 574.050 451.050 ;
        RECT 577.950 449.100 580.050 451.200 ;
        RECT 568.950 442.950 571.050 445.050 ;
        RECT 560.400 433.050 561.450 436.950 ;
        RECT 565.350 435.600 567.450 437.700 ;
        RECT 559.950 430.950 562.050 433.050 ;
        RECT 572.400 424.050 573.450 448.950 ;
        RECT 578.400 448.350 579.600 449.100 ;
        RECT 577.800 445.950 579.900 448.050 ;
        RECT 583.650 437.700 584.850 456.300 ;
        RECT 587.400 450.600 588.450 460.950 ;
        RECT 587.400 448.350 588.600 450.600 ;
        RECT 586.950 445.950 589.050 448.050 ;
        RECT 583.050 435.600 585.150 437.700 ;
        RECT 586.950 436.950 589.050 439.050 ;
        RECT 580.950 430.950 583.050 433.050 ;
        RECT 571.950 421.950 574.050 424.050 ;
        RECT 577.350 423.300 579.450 425.400 ;
        RECT 548.400 415.350 549.600 416.100 ;
        RECT 550.950 415.950 553.050 418.050 ;
        RECT 553.950 416.100 556.050 418.200 ;
        RECT 538.950 412.950 541.050 415.050 ;
        RECT 541.950 412.950 544.050 415.050 ;
        RECT 544.950 412.950 547.050 415.050 ;
        RECT 547.950 412.950 550.050 415.050 ;
        RECT 539.400 411.000 540.600 412.650 ;
        RECT 529.950 406.950 532.050 409.050 ;
        RECT 535.950 406.950 538.050 409.050 ;
        RECT 538.950 406.950 541.050 411.000 ;
        RECT 545.400 410.400 546.600 412.650 ;
        RECT 554.400 412.050 555.450 416.100 ;
        RECT 556.950 415.950 559.050 421.050 ;
        RECT 565.950 416.100 568.050 418.200 ;
        RECT 571.950 416.100 574.050 418.200 ;
        RECT 566.400 415.350 567.600 416.100 ;
        RECT 572.400 415.350 573.600 416.100 ;
        RECT 556.950 412.800 559.050 414.900 ;
        RECT 562.950 412.950 565.050 415.050 ;
        RECT 565.950 412.950 568.050 415.050 ;
        RECT 571.950 412.950 574.050 415.050 ;
        RECT 526.950 388.950 529.050 391.050 ;
        RECT 524.400 386.400 528.450 387.450 ;
        RECT 521.550 381.300 523.650 383.400 ;
        RECT 521.550 374.700 522.750 381.300 ;
        RECT 527.400 376.050 528.450 386.400 ;
        RECT 521.550 372.600 523.650 374.700 ;
        RECT 526.950 373.950 529.050 376.050 ;
        RECT 530.400 373.050 531.450 406.950 ;
        RECT 517.950 358.950 520.050 361.050 ;
        RECT 521.550 359.700 522.750 372.600 ;
        RECT 529.950 370.950 532.050 373.050 ;
        RECT 526.950 367.950 529.050 370.050 ;
        RECT 527.400 365.400 528.600 367.650 ;
        RECT 521.550 357.600 523.650 359.700 ;
        RECT 527.400 355.050 528.450 365.400 ;
        RECT 526.950 352.950 529.050 355.050 ;
        RECT 523.950 339.000 526.050 343.050 ;
        RECT 529.950 340.950 532.050 343.050 ;
        RECT 524.400 337.350 525.600 339.000 ;
        RECT 520.950 334.950 523.050 337.050 ;
        RECT 523.950 334.950 526.050 337.050 ;
        RECT 521.400 332.400 522.600 334.650 ;
        RECT 530.400 334.050 531.450 340.950 ;
        RECT 514.950 325.950 517.050 328.050 ;
        RECT 508.950 316.950 511.050 319.050 ;
        RECT 509.400 301.050 510.450 316.950 ;
        RECT 521.400 313.050 522.450 332.400 ;
        RECT 529.950 331.950 532.050 334.050 ;
        RECT 526.950 313.950 529.050 316.050 ;
        RECT 520.950 310.950 523.050 313.050 ;
        RECT 517.350 303.300 519.450 305.400 ;
        RECT 520.950 304.800 523.050 306.900 ;
        RECT 508.950 298.950 511.050 301.050 ;
        RECT 505.950 295.950 508.050 298.050 ;
        RECT 518.250 296.700 519.450 303.300 ;
        RECT 517.350 294.600 519.450 296.700 ;
        RECT 503.400 292.350 504.600 294.600 ;
        RECT 502.950 289.950 505.050 292.050 ;
        RECT 505.950 289.950 508.050 292.050 ;
        RECT 511.950 289.950 514.050 292.050 ;
        RECT 506.400 288.900 507.600 289.650 ;
        RECT 512.400 288.900 513.600 289.650 ;
        RECT 505.950 286.800 508.050 288.900 ;
        RECT 511.950 286.800 514.050 288.900 ;
        RECT 508.950 283.950 511.050 286.050 ;
        RECT 509.400 280.050 510.450 283.950 ;
        RECT 518.250 281.700 519.450 294.600 ;
        RECT 508.950 277.950 511.050 280.050 ;
        RECT 517.350 279.600 519.450 281.700 ;
        RECT 502.950 271.950 505.050 274.050 ;
        RECT 499.950 265.950 502.050 268.050 ;
        RECT 500.400 262.200 501.450 265.950 ;
        RECT 499.950 260.100 502.050 262.200 ;
        RECT 475.800 244.950 477.900 247.050 ;
        RECT 478.950 244.950 481.050 247.050 ;
        RECT 482.550 245.700 483.750 252.300 ;
        RECT 445.950 241.950 448.050 244.050 ;
        RECT 472.950 241.950 475.050 244.050 ;
        RECT 439.950 215.100 442.050 217.200 ;
        RECT 446.400 216.600 447.450 241.950 ;
        RECT 448.950 238.950 451.050 241.050 ;
        RECT 449.400 223.050 450.450 238.950 ;
        RECT 460.950 232.950 463.050 235.050 ;
        RECT 457.350 225.300 459.450 227.400 ;
        RECT 448.950 220.950 451.050 223.050 ;
        RECT 458.250 218.700 459.450 225.300 ;
        RECT 457.350 216.600 459.450 218.700 ;
        RECT 440.400 214.350 441.600 215.100 ;
        RECT 446.400 214.350 447.600 216.600 ;
        RECT 439.950 211.950 442.050 214.050 ;
        RECT 442.950 211.950 445.050 214.050 ;
        RECT 445.950 211.950 448.050 214.050 ;
        RECT 451.950 211.950 454.050 214.050 ;
        RECT 433.950 208.950 436.050 211.050 ;
        RECT 443.400 210.900 444.600 211.650 ;
        RECT 442.950 208.800 445.050 210.900 ;
        RECT 452.400 209.400 453.600 211.650 ;
        RECT 430.950 205.950 433.050 208.050 ;
        RECT 452.400 199.050 453.450 209.400 ;
        RECT 458.250 203.700 459.450 216.600 ;
        RECT 457.350 201.600 459.450 203.700 ;
        RECT 461.400 199.050 462.450 232.950 ;
        RECT 479.400 229.050 480.450 244.950 ;
        RECT 482.550 243.600 484.650 245.700 ;
        RECT 478.950 226.950 481.050 229.050 ;
        RECT 472.650 223.500 474.750 224.400 ;
        RECT 472.650 222.300 476.850 223.500 ;
        RECT 469.950 215.100 472.050 217.200 ;
        RECT 470.400 214.350 471.600 215.100 ;
        RECT 469.800 211.950 471.900 214.050 ;
        RECT 466.950 208.950 469.050 211.050 ;
        RECT 427.950 196.950 430.050 199.050 ;
        RECT 451.950 196.950 454.050 199.050 ;
        RECT 460.950 196.950 463.050 199.050 ;
        RECT 467.400 196.050 468.450 208.950 ;
        RECT 475.650 203.700 476.850 222.300 ;
        RECT 487.950 219.450 490.050 223.050 ;
        RECT 485.400 218.400 490.050 219.450 ;
        RECT 478.950 215.100 481.050 217.200 ;
        RECT 479.400 214.350 480.600 215.100 ;
        RECT 478.950 211.950 481.050 214.050 ;
        RECT 485.400 205.050 486.450 218.400 ;
        RECT 487.950 217.950 490.050 218.400 ;
        RECT 491.400 217.200 492.450 253.950 ;
        RECT 496.950 253.800 499.050 255.900 ;
        RECT 500.400 253.050 501.450 260.100 ;
        RECT 499.950 250.950 502.050 253.050 ;
        RECT 503.400 250.050 504.450 271.950 ;
        RECT 521.400 271.050 522.450 304.800 ;
        RECT 523.950 295.950 526.050 298.050 ;
        RECT 527.400 297.450 528.450 313.950 ;
        RECT 530.400 307.050 531.450 331.950 ;
        RECT 536.400 316.050 537.450 406.950 ;
        RECT 545.400 403.050 546.450 410.400 ;
        RECT 550.950 406.950 553.050 412.050 ;
        RECT 553.950 409.950 556.050 412.050 ;
        RECT 557.400 406.050 558.450 412.800 ;
        RECT 559.950 406.950 562.050 412.050 ;
        RECT 563.400 410.400 564.600 412.650 ;
        RECT 578.250 410.400 579.450 423.300 ;
        RECT 556.950 403.950 559.050 406.050 ;
        RECT 563.400 403.050 564.450 410.400 ;
        RECT 577.350 408.300 579.450 410.400 ;
        RECT 544.950 400.950 547.050 403.050 ;
        RECT 562.950 400.950 565.050 403.050 ;
        RECT 578.250 401.700 579.450 408.300 ;
        RECT 541.950 397.950 544.050 400.050 ;
        RECT 577.350 399.600 579.450 401.700 ;
        RECT 538.950 391.950 541.050 394.050 ;
        RECT 539.400 355.050 540.450 391.950 ;
        RECT 542.400 370.050 543.450 397.950 ;
        RECT 556.950 388.950 559.050 391.050 ;
        RECT 550.950 376.950 553.050 379.050 ;
        RECT 551.400 372.600 552.450 376.950 ;
        RECT 553.950 373.950 556.050 376.050 ;
        RECT 551.400 370.350 552.600 372.600 ;
        RECT 541.950 367.950 544.050 370.050 ;
        RECT 545.400 367.950 547.500 370.050 ;
        RECT 550.800 367.950 552.900 370.050 ;
        RECT 538.950 352.950 541.050 355.050 ;
        RECT 542.400 349.050 543.450 367.950 ;
        RECT 550.950 361.950 553.050 364.050 ;
        RECT 541.950 346.950 544.050 349.050 ;
        RECT 539.400 334.950 541.500 337.050 ;
        RECT 544.800 334.950 546.900 337.050 ;
        RECT 545.400 333.900 546.600 334.650 ;
        RECT 544.950 331.800 547.050 333.900 ;
        RECT 538.950 325.950 541.050 328.050 ;
        RECT 535.950 313.950 538.050 316.050 ;
        RECT 529.950 304.950 532.050 307.050 ;
        RECT 532.650 301.500 534.750 302.400 ;
        RECT 532.650 300.300 536.850 301.500 ;
        RECT 527.400 296.400 531.450 297.450 ;
        RECT 524.400 274.050 525.450 295.950 ;
        RECT 530.400 294.600 531.450 296.400 ;
        RECT 530.400 292.350 531.600 294.600 ;
        RECT 529.800 289.950 531.900 292.050 ;
        RECT 535.650 281.700 536.850 300.300 ;
        RECT 539.400 294.600 540.450 325.950 ;
        RECT 551.400 318.450 552.450 361.950 ;
        RECT 554.400 358.050 555.450 373.950 ;
        RECT 557.400 373.200 558.450 388.950 ;
        RECT 556.950 371.100 559.050 373.200 ;
        RECT 571.950 371.100 574.050 373.200 ;
        RECT 553.950 355.950 556.050 358.050 ;
        RECT 553.950 349.950 556.050 352.050 ;
        RECT 554.400 322.050 555.450 349.950 ;
        RECT 553.950 319.950 556.050 322.050 ;
        RECT 551.400 317.400 555.450 318.450 ;
        RECT 550.950 313.950 553.050 316.050 ;
        RECT 544.950 307.950 547.050 310.050 ;
        RECT 539.400 292.350 540.600 294.600 ;
        RECT 538.950 289.950 541.050 292.050 ;
        RECT 545.400 286.050 546.450 307.950 ;
        RECT 551.400 292.050 552.450 313.950 ;
        RECT 550.950 289.950 553.050 292.050 ;
        RECT 544.950 283.950 547.050 286.050 ;
        RECT 535.050 279.600 537.150 281.700 ;
        RECT 554.400 280.050 555.450 317.400 ;
        RECT 557.400 310.050 558.450 371.100 ;
        RECT 572.400 370.350 573.600 371.100 ;
        RECT 562.950 367.950 565.050 370.050 ;
        RECT 568.950 367.950 571.050 370.050 ;
        RECT 571.950 367.950 574.050 370.050 ;
        RECT 563.400 339.600 564.450 367.950 ;
        RECT 569.400 366.000 570.600 367.650 ;
        RECT 568.950 361.950 571.050 366.000 ;
        RECT 581.400 364.050 582.450 430.950 ;
        RECT 583.950 427.950 586.050 430.050 ;
        RECT 580.950 361.950 583.050 364.050 ;
        RECT 584.400 361.050 585.450 427.950 ;
        RECT 587.400 418.050 588.450 436.950 ;
        RECT 593.400 430.050 594.450 494.400 ;
        RECT 599.400 489.900 600.450 503.400 ;
        RECT 601.950 499.950 604.050 502.050 ;
        RECT 598.950 487.800 601.050 489.900 ;
        RECT 595.950 466.950 598.050 469.050 ;
        RECT 596.400 457.050 597.450 466.950 ;
        RECT 598.950 460.950 601.050 463.050 ;
        RECT 595.950 454.950 598.050 457.050 ;
        RECT 595.950 451.800 598.050 453.900 ;
        RECT 596.400 436.050 597.450 451.800 ;
        RECT 595.950 433.950 598.050 436.050 ;
        RECT 592.950 427.950 595.050 430.050 ;
        RECT 595.050 423.300 597.150 425.400 ;
        RECT 586.950 415.950 589.050 418.050 ;
        RECT 589.800 412.950 591.900 415.050 ;
        RECT 590.400 411.900 591.600 412.650 ;
        RECT 589.950 409.800 592.050 411.900 ;
        RECT 595.650 404.700 596.850 423.300 ;
        RECT 599.400 421.050 600.450 460.950 ;
        RECT 602.400 454.050 603.450 499.950 ;
        RECT 610.950 494.100 613.050 496.200 ;
        RECT 617.400 495.600 618.450 505.950 ;
        RECT 611.400 493.350 612.600 494.100 ;
        RECT 617.400 493.350 618.600 495.600 ;
        RECT 607.950 490.950 610.050 493.050 ;
        RECT 610.950 490.950 613.050 493.050 ;
        RECT 613.950 490.950 616.050 493.050 ;
        RECT 616.950 490.950 619.050 493.050 ;
        RECT 608.400 489.900 609.600 490.650 ;
        RECT 607.950 487.800 610.050 489.900 ;
        RECT 614.400 488.400 615.600 490.650 ;
        RECT 604.950 478.950 607.050 481.050 ;
        RECT 605.400 469.050 606.450 478.950 ;
        RECT 614.400 475.050 615.450 488.400 ;
        RECT 616.950 475.950 619.050 478.050 ;
        RECT 613.950 472.950 616.050 475.050 ;
        RECT 617.400 469.050 618.450 475.950 ;
        RECT 604.950 466.950 607.050 469.050 ;
        RECT 616.950 466.950 619.050 469.050 ;
        RECT 601.950 451.950 604.050 454.050 ;
        RECT 607.950 450.000 610.050 454.050 ;
        RECT 613.950 450.000 616.050 454.050 ;
        RECT 608.400 448.350 609.600 450.000 ;
        RECT 614.400 448.350 615.600 450.000 ;
        RECT 604.950 445.950 607.050 448.050 ;
        RECT 607.950 445.950 610.050 448.050 ;
        RECT 610.950 445.950 613.050 448.050 ;
        RECT 613.950 445.950 616.050 448.050 ;
        RECT 605.400 443.400 606.600 445.650 ;
        RECT 611.400 444.900 612.600 445.650 ;
        RECT 605.400 427.050 606.450 443.400 ;
        RECT 610.950 442.800 613.050 444.900 ;
        RECT 616.950 439.950 619.050 445.050 ;
        RECT 623.400 439.050 624.450 511.950 ;
        RECT 626.400 466.050 627.450 517.950 ;
        RECT 635.400 504.450 636.450 595.950 ;
        RECT 637.950 592.950 640.050 595.050 ;
        RECT 638.400 514.050 639.450 592.950 ;
        RECT 640.950 586.950 643.050 589.050 ;
        RECT 641.400 574.050 642.450 586.950 ;
        RECT 650.400 580.050 651.450 605.100 ;
        RECT 656.400 604.350 657.600 605.100 ;
        RECT 662.400 604.350 663.600 606.600 ;
        RECT 655.950 601.950 658.050 604.050 ;
        RECT 658.950 601.950 661.050 604.050 ;
        RECT 661.950 601.950 664.050 604.050 ;
        RECT 664.950 601.950 667.050 604.050 ;
        RECT 659.400 600.900 660.600 601.650 ;
        RECT 665.400 600.900 666.600 601.650 ;
        RECT 658.950 598.800 661.050 600.900 ;
        RECT 664.950 598.800 667.050 600.900 ;
        RECT 659.400 595.050 660.450 598.800 ;
        RECT 658.950 592.950 661.050 595.050 ;
        RECT 661.950 589.950 664.050 592.050 ;
        RECT 649.950 577.950 652.050 580.050 ;
        RECT 640.950 571.950 643.050 574.050 ;
        RECT 646.950 572.100 649.050 574.200 ;
        RECT 647.400 571.350 648.600 572.100 ;
        RECT 643.950 568.950 646.050 571.050 ;
        RECT 646.950 568.950 649.050 571.050 ;
        RECT 649.950 568.950 652.050 571.050 ;
        RECT 644.400 567.900 645.600 568.650 ;
        RECT 643.950 565.800 646.050 567.900 ;
        RECT 650.400 566.400 651.600 568.650 ;
        RECT 650.400 564.450 651.450 566.400 ;
        RECT 647.400 563.400 651.450 564.450 ;
        RECT 647.400 553.050 648.450 563.400 ;
        RECT 646.950 550.950 649.050 553.050 ;
        RECT 643.950 527.100 646.050 529.200 ;
        RECT 649.950 527.100 652.050 529.200 ;
        RECT 644.400 526.350 645.600 527.100 ;
        RECT 650.400 526.350 651.600 527.100 ;
        RECT 643.950 523.950 646.050 526.050 ;
        RECT 646.950 523.950 649.050 526.050 ;
        RECT 649.950 523.950 652.050 526.050 ;
        RECT 652.950 523.950 655.050 526.050 ;
        RECT 640.950 520.950 643.050 523.050 ;
        RECT 647.400 522.000 648.600 523.650 ;
        RECT 637.950 511.950 640.050 514.050 ;
        RECT 632.400 504.000 636.450 504.450 ;
        RECT 631.950 503.400 636.450 504.000 ;
        RECT 631.950 499.950 634.050 503.400 ;
        RECT 631.950 490.950 634.050 493.050 ;
        RECT 634.950 490.950 637.050 493.050 ;
        RECT 632.400 488.400 633.600 490.650 ;
        RECT 632.400 478.050 633.450 488.400 ;
        RECT 637.950 487.950 640.050 490.050 ;
        RECT 631.950 475.950 634.050 478.050 ;
        RECT 631.950 469.950 634.050 472.050 ;
        RECT 625.950 463.950 628.050 466.050 ;
        RECT 626.400 445.050 627.450 463.950 ;
        RECT 632.400 463.050 633.450 469.950 ;
        RECT 631.950 460.950 634.050 463.050 ;
        RECT 632.400 450.600 633.450 460.950 ;
        RECT 638.400 454.050 639.450 487.950 ;
        RECT 641.400 469.050 642.450 520.950 ;
        RECT 643.950 517.950 646.050 520.050 ;
        RECT 646.950 517.950 649.050 522.000 ;
        RECT 653.400 521.400 654.600 523.650 ;
        RECT 662.400 523.050 663.450 589.950 ;
        RECT 671.400 589.050 672.450 644.400 ;
        RECT 673.950 613.950 676.050 616.050 ;
        RECT 674.400 601.050 675.450 613.950 ;
        RECT 677.400 607.050 678.450 664.950 ;
        RECT 683.400 652.050 684.450 671.550 ;
        RECT 691.950 667.950 694.050 670.050 ;
        RECT 682.950 649.950 685.050 652.050 ;
        RECT 685.950 651.000 688.050 655.050 ;
        RECT 692.400 651.600 693.450 667.950 ;
        RECT 686.400 649.350 687.600 651.000 ;
        RECT 692.400 649.350 693.600 651.600 ;
        RECT 685.950 646.950 688.050 649.050 ;
        RECT 688.950 646.950 691.050 649.050 ;
        RECT 691.950 646.950 694.050 649.050 ;
        RECT 689.400 644.400 690.600 646.650 ;
        RECT 679.950 637.950 682.050 640.050 ;
        RECT 680.400 634.050 681.450 637.950 ;
        RECT 689.400 634.050 690.450 644.400 ;
        RECT 679.950 631.950 682.050 634.050 ;
        RECT 688.950 631.950 691.050 634.050 ;
        RECT 704.400 619.050 705.450 683.400 ;
        RECT 713.400 682.350 714.600 684.600 ;
        RECT 718.950 683.100 721.050 685.200 ;
        RECT 722.400 685.050 723.450 712.950 ;
        RECT 727.950 709.950 730.050 712.050 ;
        RECT 724.950 697.950 727.050 700.050 ;
        RECT 719.400 682.350 720.600 683.100 ;
        RECT 721.950 682.950 724.050 685.050 ;
        RECT 709.950 679.950 712.050 682.050 ;
        RECT 712.950 679.950 715.050 682.050 ;
        RECT 715.950 679.950 718.050 682.050 ;
        RECT 718.950 679.950 721.050 682.050 ;
        RECT 710.400 677.400 711.600 679.650 ;
        RECT 716.400 678.900 717.600 679.650 ;
        RECT 710.400 670.050 711.450 677.400 ;
        RECT 715.950 676.800 718.050 678.900 ;
        RECT 721.950 676.950 724.050 679.050 ;
        RECT 709.950 667.950 712.050 670.050 ;
        RECT 712.950 650.100 715.050 652.200 ;
        RECT 713.400 649.350 714.600 650.100 ;
        RECT 709.950 646.950 712.050 649.050 ;
        RECT 712.950 646.950 715.050 649.050 ;
        RECT 715.950 646.950 718.050 649.050 ;
        RECT 716.400 644.400 717.600 646.650 ;
        RECT 716.400 640.050 717.450 644.400 ;
        RECT 715.950 637.950 718.050 640.050 ;
        RECT 703.950 616.950 706.050 619.050 ;
        RECT 712.950 616.950 715.050 619.050 ;
        RECT 685.950 610.950 688.050 613.050 ;
        RECT 686.400 607.200 687.450 610.950 ;
        RECT 676.950 604.950 679.050 607.050 ;
        RECT 679.950 605.100 682.050 607.200 ;
        RECT 685.950 605.100 688.050 607.200 ;
        RECT 694.950 605.100 697.050 607.200 ;
        RECT 713.400 606.600 714.450 616.950 ;
        RECT 722.400 609.450 723.450 676.950 ;
        RECT 725.400 673.050 726.450 697.950 ;
        RECT 724.950 670.950 727.050 673.050 ;
        RECT 724.950 651.450 727.050 652.050 ;
        RECT 728.400 651.450 729.450 709.950 ;
        RECT 737.400 700.050 738.450 766.950 ;
        RECT 739.950 762.000 742.050 766.050 ;
        RECT 749.400 762.600 750.450 766.950 ;
        RECT 740.400 760.350 741.600 762.000 ;
        RECT 749.400 760.350 750.600 762.600 ;
        RECT 740.100 757.950 742.200 760.050 ;
        RECT 745.500 757.950 747.600 760.050 ;
        RECT 748.800 757.950 750.900 760.050 ;
        RECT 746.400 755.400 747.600 757.650 ;
        RECT 739.950 751.950 742.050 754.050 ;
        RECT 740.400 712.050 741.450 751.950 ;
        RECT 746.400 748.050 747.450 755.400 ;
        RECT 748.950 748.950 751.050 751.050 ;
        RECT 745.950 745.950 748.050 748.050 ;
        RECT 749.400 729.600 750.450 748.950 ;
        RECT 755.400 730.050 756.450 772.950 ;
        RECT 757.950 763.950 760.050 766.050 ;
        RECT 758.400 739.050 759.450 763.950 ;
        RECT 764.400 763.200 765.450 796.950 ;
        RECT 773.400 787.050 774.450 800.400 ;
        RECT 778.950 799.950 781.050 802.050 ;
        RECT 791.400 801.900 792.600 802.650 ;
        RECT 800.400 802.050 801.450 874.950 ;
        RECT 803.400 868.050 804.450 878.400 ;
        RECT 808.950 874.950 811.050 879.000 ;
        RECT 814.950 877.950 817.050 880.050 ;
        RECT 802.950 865.950 805.050 868.050 ;
        RECT 815.400 850.050 816.450 877.950 ;
        RECT 818.400 859.050 819.450 917.100 ;
        RECT 821.400 913.050 822.450 922.950 ;
        RECT 830.400 918.450 831.600 918.600 ;
        RECT 824.400 917.400 831.600 918.450 ;
        RECT 820.950 910.950 823.050 913.050 ;
        RECT 824.400 886.050 825.450 917.400 ;
        RECT 830.400 916.350 831.600 917.400 ;
        RECT 835.950 917.100 838.050 919.200 ;
        RECT 841.950 917.100 844.050 919.200 ;
        RECT 851.400 918.600 852.450 922.950 ;
        RECT 862.950 919.950 865.050 922.050 ;
        RECT 836.400 916.350 837.600 917.100 ;
        RECT 829.950 913.950 832.050 916.050 ;
        RECT 832.950 913.950 835.050 916.050 ;
        RECT 835.950 913.950 838.050 916.050 ;
        RECT 833.400 912.900 834.600 913.650 ;
        RECT 832.950 910.800 835.050 912.900 ;
        RECT 842.400 912.450 843.450 917.100 ;
        RECT 851.400 916.350 852.600 918.600 ;
        RECT 856.950 917.100 859.050 919.200 ;
        RECT 857.400 916.350 858.600 917.100 ;
        RECT 850.950 913.950 853.050 916.050 ;
        RECT 853.950 913.950 856.050 916.050 ;
        RECT 856.950 913.950 859.050 916.050 ;
        RECT 839.400 911.400 843.450 912.450 ;
        RECT 854.400 912.000 855.600 913.650 ;
        RECT 839.400 907.050 840.450 911.400 ;
        RECT 847.950 907.950 850.050 910.050 ;
        RECT 853.950 907.950 856.050 912.000 ;
        RECT 863.400 910.050 864.450 919.950 ;
        RECT 862.950 907.950 865.050 910.050 ;
        RECT 838.950 904.950 841.050 907.050 ;
        RECT 823.950 883.950 826.050 886.050 ;
        RECT 832.950 884.100 835.050 886.200 ;
        RECT 839.400 885.600 840.450 904.950 ;
        RECT 833.400 883.350 834.600 884.100 ;
        RECT 839.400 883.350 840.600 885.600 ;
        RECT 829.950 880.950 832.050 883.050 ;
        RECT 832.950 880.950 835.050 883.050 ;
        RECT 835.950 880.950 838.050 883.050 ;
        RECT 838.950 880.950 841.050 883.050 ;
        RECT 830.400 878.400 831.600 880.650 ;
        RECT 836.400 878.400 837.600 880.650 ;
        RECT 817.950 856.950 820.050 859.050 ;
        RECT 814.950 847.950 817.050 850.050 ;
        RECT 805.950 844.950 808.050 847.050 ;
        RECT 806.400 834.900 807.450 844.950 ;
        RECT 808.950 838.950 811.050 841.050 ;
        RECT 817.950 839.100 820.050 841.200 ;
        RECT 823.950 839.100 826.050 841.200 ;
        RECT 805.950 832.800 808.050 834.900 ;
        RECT 809.400 814.050 810.450 838.950 ;
        RECT 818.400 838.350 819.600 839.100 ;
        RECT 824.400 838.350 825.600 839.100 ;
        RECT 814.950 835.950 817.050 838.050 ;
        RECT 817.950 835.950 820.050 838.050 ;
        RECT 820.950 835.950 823.050 838.050 ;
        RECT 823.950 835.950 826.050 838.050 ;
        RECT 815.400 834.900 816.600 835.650 ;
        RECT 821.400 834.900 822.600 835.650 ;
        RECT 814.950 832.800 817.050 834.900 ;
        RECT 820.950 832.800 823.050 834.900 ;
        RECT 808.950 811.950 811.050 814.050 ;
        RECT 808.950 806.100 811.050 808.200 ;
        RECT 815.400 807.600 816.450 832.800 ;
        RECT 830.400 829.050 831.450 878.400 ;
        RECT 836.400 876.450 837.450 878.400 ;
        RECT 848.400 877.050 849.450 907.950 ;
        RECT 866.400 906.450 867.450 925.950 ;
        RECT 868.950 922.950 871.050 925.050 ;
        RECT 869.400 919.050 870.450 922.950 ;
        RECT 868.950 916.950 871.050 919.050 ;
        RECT 874.950 918.000 877.050 922.050 ;
        RECT 880.950 918.000 883.050 922.050 ;
        RECT 875.400 916.350 876.600 918.000 ;
        RECT 881.400 916.350 882.600 918.000 ;
        RECT 871.950 913.950 874.050 916.050 ;
        RECT 874.950 913.950 877.050 916.050 ;
        RECT 877.950 913.950 880.050 916.050 ;
        RECT 880.950 913.950 883.050 916.050 ;
        RECT 872.400 911.400 873.600 913.650 ;
        RECT 878.400 912.900 879.600 913.650 ;
        RECT 887.400 913.050 888.450 952.800 ;
        RECT 902.400 952.050 903.450 956.400 ;
        RECT 889.950 949.950 892.050 952.050 ;
        RECT 901.950 949.950 904.050 952.050 ;
        RECT 890.400 937.050 891.450 949.950 ;
        RECT 911.400 943.050 912.450 964.950 ;
        RECT 920.400 963.600 921.450 973.950 ;
        RECT 991.950 970.950 994.050 973.050 ;
        RECT 1003.950 970.950 1006.050 973.050 ;
        RECT 973.950 967.950 976.050 970.050 ;
        RECT 920.400 961.350 921.600 963.600 ;
        RECT 925.950 963.000 928.050 967.050 ;
        RECT 926.400 961.350 927.600 963.000 ;
        RECT 934.950 961.950 937.050 964.050 ;
        RECT 943.950 962.100 946.050 967.050 ;
        RECT 949.950 962.100 952.050 964.200 ;
        RECT 955.950 962.100 958.050 964.200 ;
        RECT 919.950 958.950 922.050 961.050 ;
        RECT 922.950 958.950 925.050 961.050 ;
        RECT 925.950 958.950 928.050 961.050 ;
        RECT 928.950 958.950 931.050 961.050 ;
        RECT 923.400 957.000 924.600 958.650 ;
        RECT 929.400 957.900 930.600 958.650 ;
        RECT 935.400 957.900 936.450 961.950 ;
        RECT 950.400 961.350 951.600 962.100 ;
        RECT 956.400 961.350 957.600 962.100 ;
        RECT 961.800 961.950 963.900 964.050 ;
        RECT 964.950 961.950 967.050 964.050 ;
        RECT 974.400 963.600 975.450 967.950 ;
        RECT 946.950 958.950 949.050 961.050 ;
        RECT 949.950 958.950 952.050 961.050 ;
        RECT 952.950 958.950 955.050 961.050 ;
        RECT 955.950 958.950 958.050 961.050 ;
        RECT 922.950 952.950 925.050 957.000 ;
        RECT 928.950 955.800 931.050 957.900 ;
        RECT 934.950 952.950 937.050 957.900 ;
        RECT 947.400 957.000 948.600 958.650 ;
        RECT 953.400 957.000 954.600 958.650 ;
        RECT 962.400 957.900 963.450 961.950 ;
        RECT 946.950 952.950 949.050 957.000 ;
        RECT 952.950 952.950 955.050 957.000 ;
        RECT 961.950 955.800 964.050 957.900 ;
        RECT 910.950 940.950 913.050 943.050 ;
        RECT 916.950 940.950 919.050 943.050 ;
        RECT 889.950 934.950 892.050 937.050 ;
        RECT 890.400 913.050 891.450 934.950 ;
        RECT 898.950 925.950 901.050 928.050 ;
        RECT 913.950 925.950 916.050 928.050 ;
        RECT 899.400 918.600 900.450 925.950 ;
        RECT 899.400 916.350 900.600 918.600 ;
        RECT 904.950 918.000 907.050 922.050 ;
        RECT 910.950 919.950 913.050 922.050 ;
        RECT 905.400 916.350 906.600 918.000 ;
        RECT 895.950 913.950 898.050 916.050 ;
        RECT 898.950 913.950 901.050 916.050 ;
        RECT 901.950 913.950 904.050 916.050 ;
        RECT 904.950 913.950 907.050 916.050 ;
        RECT 866.400 905.400 870.450 906.450 ;
        RECT 862.950 898.950 865.050 901.050 ;
        RECT 856.950 889.950 859.050 892.050 ;
        RECT 857.400 885.600 858.450 889.950 ;
        RECT 863.400 886.200 864.450 898.950 ;
        RECT 857.400 883.350 858.600 885.600 ;
        RECT 862.950 884.100 865.050 886.200 ;
        RECT 863.400 883.350 864.600 884.100 ;
        RECT 853.950 880.950 856.050 883.050 ;
        RECT 856.950 880.950 859.050 883.050 ;
        RECT 859.950 880.950 862.050 883.050 ;
        RECT 862.950 880.950 865.050 883.050 ;
        RECT 854.400 879.000 855.600 880.650 ;
        RECT 860.400 879.000 861.600 880.650 ;
        RECT 869.400 880.050 870.450 905.400 ;
        RECT 872.400 901.050 873.450 911.400 ;
        RECT 877.950 910.800 880.050 912.900 ;
        RECT 886.800 910.950 888.900 913.050 ;
        RECT 889.950 910.950 892.050 913.050 ;
        RECT 896.400 912.900 897.600 913.650 ;
        RECT 902.400 912.900 903.600 913.650 ;
        RECT 895.950 910.800 898.050 912.900 ;
        RECT 901.950 910.800 904.050 912.900 ;
        RECT 871.950 898.950 874.050 901.050 ;
        RECT 892.950 895.950 895.050 898.050 ;
        RECT 889.950 889.950 892.050 892.050 ;
        RECT 871.950 884.100 874.050 886.200 ;
        RECT 877.950 884.100 880.050 886.200 ;
        RECT 883.950 884.100 886.050 886.200 ;
        RECT 865.800 879.000 867.900 880.050 ;
        RECT 833.400 875.400 837.450 876.450 ;
        RECT 833.400 835.050 834.450 875.400 ;
        RECT 847.950 874.950 850.050 877.050 ;
        RECT 853.950 876.450 856.050 879.000 ;
        RECT 853.950 875.400 858.450 876.450 ;
        RECT 853.950 874.950 856.050 875.400 ;
        RECT 841.950 865.950 844.050 868.050 ;
        RECT 835.950 839.100 838.050 841.200 ;
        RECT 842.400 840.600 843.450 865.950 ;
        RECT 853.950 853.950 856.050 856.050 ;
        RECT 847.950 847.950 850.050 850.050 ;
        RECT 848.400 840.600 849.450 847.950 ;
        RECT 854.400 841.050 855.450 853.950 ;
        RECT 832.950 832.950 835.050 835.050 ;
        RECT 832.950 829.800 835.050 831.900 ;
        RECT 823.950 826.950 826.050 829.050 ;
        RECT 829.950 826.950 832.050 829.050 ;
        RECT 820.950 811.950 823.050 814.050 ;
        RECT 809.400 805.350 810.600 806.100 ;
        RECT 815.400 805.350 816.600 807.600 ;
        RECT 805.950 802.950 808.050 805.050 ;
        RECT 808.950 802.950 811.050 805.050 ;
        RECT 811.950 802.950 814.050 805.050 ;
        RECT 814.950 802.950 817.050 805.050 ;
        RECT 790.950 799.800 793.050 801.900 ;
        RECT 799.950 799.950 802.050 802.050 ;
        RECT 806.400 801.900 807.600 802.650 ;
        RECT 812.400 801.900 813.600 802.650 ;
        RECT 821.400 801.900 822.450 811.950 ;
        RECT 805.950 799.800 808.050 801.900 ;
        RECT 811.950 799.800 814.050 801.900 ;
        RECT 820.950 799.800 823.050 801.900 ;
        RECT 772.950 784.950 775.050 787.050 ;
        RECT 791.400 769.050 792.450 799.800 ;
        RECT 787.800 768.000 789.900 769.050 ;
        RECT 787.800 766.950 790.050 768.000 ;
        RECT 790.950 766.950 793.050 769.050 ;
        RECT 763.950 761.100 766.050 763.200 ;
        RECT 769.950 762.000 772.050 766.050 ;
        RECT 781.950 763.950 784.050 766.050 ;
        RECT 787.950 765.450 790.050 766.950 ;
        RECT 787.950 765.000 792.450 765.450 ;
        RECT 788.400 764.400 792.450 765.000 ;
        RECT 764.400 760.350 765.600 761.100 ;
        RECT 770.400 760.350 771.600 762.000 ;
        RECT 763.950 757.950 766.050 760.050 ;
        RECT 766.950 757.950 769.050 760.050 ;
        RECT 769.950 757.950 772.050 760.050 ;
        RECT 772.950 757.950 775.050 760.050 ;
        RECT 767.400 755.400 768.600 757.650 ;
        RECT 773.400 756.900 774.600 757.650 ;
        RECT 782.400 757.050 783.450 763.950 ;
        RECT 791.400 762.600 792.450 764.400 ;
        RECT 791.400 760.350 792.600 762.600 ;
        RECT 796.950 761.100 799.050 763.200 ;
        RECT 802.950 761.100 805.050 763.200 ;
        RECT 797.400 760.350 798.600 761.100 ;
        RECT 787.950 757.950 790.050 760.050 ;
        RECT 790.950 757.950 793.050 760.050 ;
        RECT 793.950 757.950 796.050 760.050 ;
        RECT 796.950 757.950 799.050 760.050 ;
        RECT 767.400 745.050 768.450 755.400 ;
        RECT 772.950 754.800 775.050 756.900 ;
        RECT 781.950 754.950 784.050 757.050 ;
        RECT 788.400 756.900 789.600 757.650 ;
        RECT 794.400 756.900 795.600 757.650 ;
        RECT 787.950 754.800 790.050 756.900 ;
        RECT 793.950 754.800 796.050 756.900 ;
        RECT 799.950 751.950 802.050 757.050 ;
        RECT 803.400 751.050 804.450 761.100 ;
        RECT 806.400 757.050 807.450 799.800 ;
        RECT 824.400 796.050 825.450 826.950 ;
        RECT 833.400 807.600 834.450 829.800 ;
        RECT 836.400 826.050 837.450 839.100 ;
        RECT 842.400 838.350 843.600 840.600 ;
        RECT 848.400 838.350 849.600 840.600 ;
        RECT 853.950 838.950 856.050 841.050 ;
        RECT 841.950 835.950 844.050 838.050 ;
        RECT 844.950 835.950 847.050 838.050 ;
        RECT 847.950 835.950 850.050 838.050 ;
        RECT 850.950 835.950 853.050 838.050 ;
        RECT 838.950 832.950 841.050 835.050 ;
        RECT 845.400 833.400 846.600 835.650 ;
        RECT 851.400 834.000 852.600 835.650 ;
        RECT 835.950 823.950 838.050 826.050 ;
        RECT 839.400 807.600 840.450 832.950 ;
        RECT 845.400 826.050 846.450 833.400 ;
        RECT 850.950 829.950 853.050 834.000 ;
        RECT 844.950 823.950 847.050 826.050 ;
        RECT 844.950 817.950 847.050 820.050 ;
        RECT 833.400 805.350 834.600 807.600 ;
        RECT 839.400 805.350 840.600 807.600 ;
        RECT 829.950 802.950 832.050 805.050 ;
        RECT 832.950 802.950 835.050 805.050 ;
        RECT 835.950 802.950 838.050 805.050 ;
        RECT 838.950 802.950 841.050 805.050 ;
        RECT 830.400 800.400 831.600 802.650 ;
        RECT 836.400 801.900 837.600 802.650 ;
        RECT 845.400 801.900 846.450 817.950 ;
        RECT 850.950 811.950 853.050 814.050 ;
        RECT 847.950 808.950 850.050 811.050 ;
        RECT 830.400 798.450 831.450 800.400 ;
        RECT 835.950 799.800 838.050 801.900 ;
        RECT 844.950 799.800 847.050 801.900 ;
        RECT 830.400 797.400 834.450 798.450 ;
        RECT 823.950 793.950 826.050 796.050 ;
        RECT 829.950 793.950 832.050 796.050 ;
        RECT 808.950 784.950 811.050 787.050 ;
        RECT 805.950 754.950 808.050 757.050 ;
        RECT 809.400 756.900 810.450 784.950 ;
        RECT 814.950 766.950 817.050 769.050 ;
        RECT 815.400 762.600 816.450 766.950 ;
        RECT 815.400 760.350 816.600 762.600 ;
        RECT 820.950 761.100 823.050 763.200 ;
        RECT 821.400 760.350 822.600 761.100 ;
        RECT 814.950 757.950 817.050 760.050 ;
        RECT 817.950 757.950 820.050 760.050 ;
        RECT 820.950 757.950 823.050 760.050 ;
        RECT 823.950 757.950 826.050 760.050 ;
        RECT 818.400 756.900 819.600 757.650 ;
        RECT 824.400 756.900 825.600 757.650 ;
        RECT 808.950 754.800 811.050 756.900 ;
        RECT 817.950 754.800 820.050 756.900 ;
        RECT 823.950 754.800 826.050 756.900 ;
        RECT 802.950 748.950 805.050 751.050 ;
        RECT 805.950 745.950 808.050 748.050 ;
        RECT 766.950 742.950 769.050 745.050 ;
        RECT 757.950 736.950 760.050 739.050 ;
        RECT 772.950 736.950 775.050 739.050 ;
        RECT 749.400 727.350 750.600 729.600 ;
        RECT 754.950 727.950 757.050 730.050 ;
        RECT 763.950 727.950 766.050 730.050 ;
        RECT 773.400 729.600 774.450 736.950 ;
        RECT 781.950 733.950 784.050 736.050 ;
        RECT 787.950 733.950 793.050 736.050 ;
        RECT 782.400 730.050 783.450 733.950 ;
        RECT 745.950 724.950 748.050 727.050 ;
        RECT 748.950 724.950 751.050 727.050 ;
        RECT 751.950 724.950 754.050 727.050 ;
        RECT 746.400 723.900 747.600 724.650 ;
        RECT 745.950 721.800 748.050 723.900 ;
        RECT 752.400 722.400 753.600 724.650 ;
        RECT 752.400 715.050 753.450 722.400 ;
        RECT 764.400 718.050 765.450 727.950 ;
        RECT 773.400 727.350 774.600 729.600 ;
        RECT 781.800 727.950 783.900 730.050 ;
        RECT 784.950 728.100 787.050 730.200 ;
        RECT 790.950 728.100 793.050 730.200 ;
        RECT 796.950 728.100 799.050 730.200 ;
        RECT 802.950 728.100 805.050 730.200 ;
        RECT 769.950 724.950 772.050 727.050 ;
        RECT 772.950 724.950 775.050 727.050 ;
        RECT 775.950 724.950 778.050 727.050 ;
        RECT 770.400 722.400 771.600 724.650 ;
        RECT 776.400 723.900 777.600 724.650 ;
        RECT 770.400 718.050 771.450 722.400 ;
        RECT 775.950 721.800 778.050 723.900 ;
        RECT 763.950 715.950 766.050 718.050 ;
        RECT 769.950 715.950 772.050 718.050 ;
        RECT 751.950 712.950 754.050 715.050 ;
        RECT 739.950 709.950 742.050 712.050 ;
        RECT 770.400 700.050 771.450 715.950 ;
        RECT 772.950 706.950 775.050 709.050 ;
        RECT 730.950 697.950 733.050 700.050 ;
        RECT 736.950 697.950 739.050 700.050 ;
        RECT 751.950 697.950 754.050 700.050 ;
        RECT 769.950 697.950 772.050 700.050 ;
        RECT 731.400 655.050 732.450 697.950 ;
        RECT 736.950 691.950 739.050 694.050 ;
        RECT 737.400 684.600 738.450 691.950 ;
        RECT 737.400 682.350 738.600 684.600 ;
        RECT 742.950 683.100 745.050 685.200 ;
        RECT 743.400 682.350 744.600 683.100 ;
        RECT 736.950 679.950 739.050 682.050 ;
        RECT 739.950 679.950 742.050 682.050 ;
        RECT 742.950 679.950 745.050 682.050 ;
        RECT 745.950 679.950 748.050 682.050 ;
        RECT 740.400 677.400 741.600 679.650 ;
        RECT 746.400 677.400 747.600 679.650 ;
        RECT 740.400 661.050 741.450 677.400 ;
        RECT 746.400 673.050 747.450 677.400 ;
        RECT 748.950 676.950 751.050 679.050 ;
        RECT 745.950 670.950 748.050 673.050 ;
        RECT 733.950 658.950 736.050 661.050 ;
        RECT 739.950 658.950 742.050 661.050 ;
        RECT 745.950 658.950 748.050 661.050 ;
        RECT 730.950 652.950 733.050 655.050 ;
        RECT 724.950 650.400 729.450 651.450 ;
        RECT 734.400 651.600 735.450 658.950 ;
        RECT 742.950 652.950 745.050 655.050 ;
        RECT 724.950 649.950 727.050 650.400 ;
        RECT 719.400 608.400 723.450 609.450 ;
        RECT 680.400 604.350 681.600 605.100 ;
        RECT 686.400 604.350 687.600 605.100 ;
        RECT 679.950 601.950 682.050 604.050 ;
        RECT 682.950 601.950 685.050 604.050 ;
        RECT 685.950 601.950 688.050 604.050 ;
        RECT 688.950 601.950 691.050 604.050 ;
        RECT 673.950 598.950 676.050 601.050 ;
        RECT 683.400 600.900 684.600 601.650 ;
        RECT 682.950 598.800 685.050 600.900 ;
        RECT 689.400 599.400 690.600 601.650 ;
        RECT 679.950 595.950 682.050 598.050 ;
        RECT 685.950 595.950 688.050 598.050 ;
        RECT 670.950 586.950 673.050 589.050 ;
        RECT 670.950 580.950 673.050 583.050 ;
        RECT 671.400 574.200 672.450 580.950 ;
        RECT 670.950 572.100 673.050 574.200 ;
        RECT 676.950 572.100 679.050 574.200 ;
        RECT 680.400 574.050 681.450 595.950 ;
        RECT 682.950 586.950 685.050 589.050 ;
        RECT 671.400 571.350 672.600 572.100 ;
        RECT 677.400 571.350 678.600 572.100 ;
        RECT 679.950 571.950 682.050 574.050 ;
        RECT 667.950 568.950 670.050 571.050 ;
        RECT 670.950 568.950 673.050 571.050 ;
        RECT 673.950 568.950 676.050 571.050 ;
        RECT 676.950 568.950 679.050 571.050 ;
        RECT 668.400 566.400 669.600 568.650 ;
        RECT 674.400 566.400 675.600 568.650 ;
        RECT 668.400 562.050 669.450 566.400 ;
        RECT 667.950 559.950 670.050 562.050 ;
        RECT 674.400 556.050 675.450 566.400 ;
        RECT 679.950 559.950 682.050 565.050 ;
        RECT 673.950 553.950 676.050 556.050 ;
        RECT 683.400 538.050 684.450 586.950 ;
        RECT 686.400 550.050 687.450 595.950 ;
        RECT 689.400 589.050 690.450 599.400 ;
        RECT 695.400 598.050 696.450 605.100 ;
        RECT 713.400 604.350 714.600 606.600 ;
        RECT 706.950 601.950 709.050 604.050 ;
        RECT 709.950 601.950 712.050 604.050 ;
        RECT 712.950 601.950 715.050 604.050 ;
        RECT 710.400 599.400 711.600 601.650 ;
        RECT 694.950 595.950 697.050 598.050 ;
        RECT 688.950 586.950 691.050 589.050 ;
        RECT 694.950 580.950 697.050 583.050 ;
        RECT 695.400 573.600 696.450 580.950 ;
        RECT 710.400 580.050 711.450 599.400 ;
        RECT 712.950 595.950 715.050 598.050 ;
        RECT 709.950 577.950 712.050 580.050 ;
        RECT 695.400 571.350 696.600 573.600 ;
        RECT 700.950 572.100 703.050 574.200 ;
        RECT 701.400 571.350 702.600 572.100 ;
        RECT 691.950 568.950 694.050 571.050 ;
        RECT 694.950 568.950 697.050 571.050 ;
        RECT 697.950 568.950 700.050 571.050 ;
        RECT 700.950 568.950 703.050 571.050 ;
        RECT 688.950 565.950 691.050 568.050 ;
        RECT 692.400 567.000 693.600 568.650 ;
        RECT 698.400 567.000 699.600 568.650 ;
        RECT 685.950 547.950 688.050 550.050 ;
        RECT 685.950 538.950 688.050 541.050 ;
        RECT 682.950 535.950 685.050 538.050 ;
        RECT 673.950 527.100 676.050 529.200 ;
        RECT 680.400 528.450 681.600 528.600 ;
        RECT 683.400 528.450 684.450 535.950 ;
        RECT 686.400 529.200 687.450 538.950 ;
        RECT 680.400 527.400 684.450 528.450 ;
        RECT 674.400 526.350 675.600 527.100 ;
        RECT 680.400 526.350 681.600 527.400 ;
        RECT 685.950 527.100 688.050 529.200 ;
        RECT 670.950 523.950 673.050 526.050 ;
        RECT 673.950 523.950 676.050 526.050 ;
        RECT 676.950 523.950 679.050 526.050 ;
        RECT 679.950 523.950 682.050 526.050 ;
        RECT 644.400 508.050 645.450 517.950 ;
        RECT 653.400 511.050 654.450 521.400 ;
        RECT 655.950 520.950 658.050 523.050 ;
        RECT 661.950 520.950 664.050 523.050 ;
        RECT 667.950 522.450 670.050 523.050 ;
        RECT 671.400 522.450 672.600 523.650 ;
        RECT 677.400 522.900 678.600 523.650 ;
        RECT 667.950 521.400 672.600 522.450 ;
        RECT 667.950 520.950 670.050 521.400 ;
        RECT 652.950 508.950 655.050 511.050 ;
        RECT 643.950 505.950 646.050 508.050 ;
        RECT 656.400 502.050 657.450 520.950 ;
        RECT 643.950 499.950 646.050 502.050 ;
        RECT 655.950 499.950 658.050 502.050 ;
        RECT 664.950 499.950 667.050 502.050 ;
        RECT 644.400 490.050 645.450 499.950 ;
        RECT 665.400 496.200 666.450 499.950 ;
        RECT 649.950 494.100 652.050 496.200 ;
        RECT 655.950 494.100 658.050 496.200 ;
        RECT 664.800 494.100 666.900 496.200 ;
        RECT 668.400 496.050 669.450 520.950 ;
        RECT 676.950 520.800 679.050 522.900 ;
        RECT 686.400 522.450 687.450 527.100 ;
        RECT 683.400 521.400 687.450 522.450 ;
        RECT 679.950 499.950 682.050 502.050 ;
        RECT 670.950 496.950 679.050 499.050 ;
        RECT 650.400 493.350 651.600 494.100 ;
        RECT 656.400 493.350 657.600 494.100 ;
        RECT 649.950 490.950 652.050 493.050 ;
        RECT 652.950 490.950 655.050 493.050 ;
        RECT 655.950 490.950 658.050 493.050 ;
        RECT 643.950 487.950 646.050 490.050 ;
        RECT 653.400 489.900 654.600 490.650 ;
        RECT 652.950 487.800 655.050 489.900 ;
        RECT 649.950 475.950 652.050 478.050 ;
        RECT 646.950 469.950 649.050 472.050 ;
        RECT 640.950 466.950 643.050 469.050 ;
        RECT 647.400 457.050 648.450 469.950 ;
        RECT 646.950 454.950 649.050 457.050 ;
        RECT 637.950 451.950 640.050 454.050 ;
        RECT 638.400 450.600 639.450 451.950 ;
        RECT 632.400 448.350 633.600 450.600 ;
        RECT 638.400 448.350 639.600 450.600 ;
        RECT 631.950 445.950 634.050 448.050 ;
        RECT 634.950 445.950 637.050 448.050 ;
        RECT 637.950 445.950 640.050 448.050 ;
        RECT 640.950 445.950 643.050 448.050 ;
        RECT 625.950 442.950 628.050 445.050 ;
        RECT 641.400 443.400 642.600 445.650 ;
        RECT 610.950 436.950 613.050 439.050 ;
        RECT 622.950 436.950 625.050 439.050 ;
        RECT 604.950 424.950 607.050 427.050 ;
        RECT 598.950 418.950 601.050 421.050 ;
        RECT 604.950 418.950 607.050 421.050 ;
        RECT 598.950 412.950 601.050 415.050 ;
        RECT 599.400 411.900 600.600 412.650 ;
        RECT 605.400 411.900 606.450 418.950 ;
        RECT 598.950 409.800 601.050 411.900 ;
        RECT 604.950 409.800 607.050 411.900 ;
        RECT 592.650 403.500 596.850 404.700 ;
        RECT 592.650 402.600 594.750 403.500 ;
        RECT 607.950 385.800 610.050 387.900 ;
        RECT 595.950 382.950 598.050 385.050 ;
        RECT 587.400 367.950 589.500 370.050 ;
        RECT 592.500 367.950 594.600 370.050 ;
        RECT 593.400 366.000 594.600 367.650 ;
        RECT 596.400 367.050 597.450 382.950 ;
        RECT 601.950 373.950 604.050 376.050 ;
        RECT 592.950 361.950 595.050 366.000 ;
        RECT 595.950 364.950 598.050 367.050 ;
        RECT 583.950 358.950 586.050 361.050 ;
        RECT 592.950 358.800 595.050 360.900 ;
        RECT 581.850 345.300 583.950 347.400 ;
        RECT 563.400 337.350 564.600 339.600 ;
        RECT 568.950 338.100 571.050 340.200 ;
        RECT 569.400 337.350 570.600 338.100 ;
        RECT 562.950 334.950 565.050 337.050 ;
        RECT 565.950 334.950 568.050 337.050 ;
        RECT 568.950 334.950 571.050 337.050 ;
        RECT 571.950 334.950 574.050 337.050 ;
        RECT 577.950 334.950 580.050 337.050 ;
        RECT 566.400 332.400 567.600 334.650 ;
        RECT 572.400 333.900 573.600 334.650 ;
        RECT 562.950 322.950 565.050 325.050 ;
        RECT 563.400 316.050 564.450 322.950 ;
        RECT 562.950 313.950 565.050 316.050 ;
        RECT 556.950 307.950 559.050 310.050 ;
        RECT 563.400 294.600 564.450 313.950 ;
        RECT 566.400 313.050 567.450 332.400 ;
        RECT 571.950 331.800 574.050 333.900 ;
        RECT 578.400 332.400 579.600 334.650 ;
        RECT 578.400 328.050 579.450 332.400 ;
        RECT 577.950 325.950 580.050 328.050 ;
        RECT 582.150 326.700 583.350 345.300 ;
        RECT 587.100 334.950 589.200 337.050 ;
        RECT 587.400 333.900 588.600 334.650 ;
        RECT 586.950 331.800 589.050 333.900 ;
        RECT 565.950 310.950 568.050 313.050 ;
        RECT 574.350 303.300 576.450 305.400 ;
        RECT 578.400 304.050 579.450 325.950 ;
        RECT 582.150 325.500 586.350 326.700 ;
        RECT 584.250 324.600 586.350 325.500 ;
        RECT 593.400 325.050 594.450 358.800 ;
        RECT 596.400 343.050 597.450 364.950 ;
        RECT 602.400 358.050 603.450 373.950 ;
        RECT 608.400 372.600 609.450 385.800 ;
        RECT 611.400 379.050 612.450 436.950 ;
        RECT 641.400 436.050 642.450 443.400 ;
        RECT 640.950 433.950 643.050 436.050 ;
        RECT 613.950 427.950 616.050 430.050 ;
        RECT 640.950 427.950 643.050 430.050 ;
        RECT 614.400 424.050 615.450 427.950 ;
        RECT 613.950 421.950 616.050 424.050 ;
        RECT 619.950 416.100 622.050 418.200 ;
        RECT 620.400 415.350 621.600 416.100 ;
        RECT 631.950 415.950 634.050 418.050 ;
        RECT 641.400 417.600 642.450 427.950 ;
        RECT 616.950 412.950 619.050 415.050 ;
        RECT 619.950 412.950 622.050 415.050 ;
        RECT 622.950 412.950 625.050 415.050 ;
        RECT 617.400 411.000 618.600 412.650 ;
        RECT 616.950 406.950 619.050 411.000 ;
        RECT 623.400 410.400 624.600 412.650 ;
        RECT 632.400 411.900 633.450 415.950 ;
        RECT 641.400 415.350 642.600 417.600 ;
        RECT 646.950 416.100 649.050 418.200 ;
        RECT 650.400 418.050 651.450 475.950 ;
        RECT 661.950 460.950 664.050 463.050 ;
        RECT 662.400 450.600 663.450 460.950 ;
        RECT 665.400 451.050 666.450 494.100 ;
        RECT 667.950 493.950 670.050 496.050 ;
        RECT 674.400 495.600 675.450 496.950 ;
        RECT 680.400 496.200 681.450 499.950 ;
        RECT 674.400 493.350 675.600 495.600 ;
        RECT 679.950 494.100 682.050 496.200 ;
        RECT 670.950 490.950 673.050 493.050 ;
        RECT 673.950 490.950 676.050 493.050 ;
        RECT 676.950 490.950 679.050 493.050 ;
        RECT 667.950 487.950 670.050 490.050 ;
        RECT 671.400 488.400 672.600 490.650 ;
        RECT 662.400 448.350 663.600 450.600 ;
        RECT 664.950 448.950 667.050 451.050 ;
        RECT 655.950 445.950 658.050 448.050 ;
        RECT 658.950 445.950 661.050 448.050 ;
        RECT 661.950 445.950 664.050 448.050 ;
        RECT 659.400 444.900 660.600 445.650 ;
        RECT 668.400 445.050 669.450 487.950 ;
        RECT 671.400 472.050 672.450 488.400 ;
        RECT 683.400 478.050 684.450 521.400 ;
        RECT 689.400 487.050 690.450 565.950 ;
        RECT 691.950 562.950 694.050 567.000 ;
        RECT 697.950 562.950 700.050 567.000 ;
        RECT 710.400 565.050 711.450 577.950 ;
        RECT 713.400 574.050 714.450 595.950 ;
        RECT 719.400 586.050 720.450 608.400 ;
        RECT 721.950 605.100 724.050 607.200 ;
        RECT 725.400 606.450 726.450 649.950 ;
        RECT 734.400 649.350 735.600 651.600 ;
        RECT 730.950 646.950 733.050 649.050 ;
        RECT 733.950 646.950 736.050 649.050 ;
        RECT 736.950 646.950 739.050 649.050 ;
        RECT 731.400 645.000 732.600 646.650 ;
        RECT 737.400 645.000 738.600 646.650 ;
        RECT 730.950 640.950 733.050 645.000 ;
        RECT 736.950 640.950 739.050 645.000 ;
        RECT 743.400 640.050 744.450 652.950 ;
        RECT 746.400 643.050 747.450 658.950 ;
        RECT 749.400 643.050 750.450 676.950 ;
        RECT 752.400 652.050 753.450 697.950 ;
        RECT 769.950 685.950 772.050 688.050 ;
        RECT 760.950 683.100 763.050 685.200 ;
        RECT 761.400 682.350 762.600 683.100 ;
        RECT 760.950 679.950 763.050 682.050 ;
        RECT 763.950 679.950 766.050 682.050 ;
        RECT 764.400 678.900 765.600 679.650 ;
        RECT 763.950 676.800 766.050 678.900 ;
        RECT 766.950 676.950 769.050 679.050 ;
        RECT 770.400 678.900 771.450 685.950 ;
        RECT 773.400 679.050 774.450 706.950 ;
        RECT 776.400 682.050 777.450 721.800 ;
        RECT 782.400 697.050 783.450 727.950 ;
        RECT 785.400 718.050 786.450 728.100 ;
        RECT 791.400 727.350 792.600 728.100 ;
        RECT 797.400 727.350 798.600 728.100 ;
        RECT 790.950 724.950 793.050 727.050 ;
        RECT 793.950 724.950 796.050 727.050 ;
        RECT 796.950 724.950 799.050 727.050 ;
        RECT 794.400 722.400 795.600 724.650 ;
        RECT 803.400 724.050 804.450 728.100 ;
        RECT 784.950 715.950 787.050 718.050 ;
        RECT 794.400 715.050 795.450 722.400 ;
        RECT 802.950 721.950 805.050 724.050 ;
        RECT 793.950 712.950 796.050 715.050 ;
        RECT 806.400 709.050 807.450 745.950 ;
        RECT 814.950 733.950 817.050 736.050 ;
        RECT 815.400 729.600 816.450 733.950 ;
        RECT 826.950 730.950 829.050 733.050 ;
        RECT 815.400 727.350 816.600 729.600 ;
        RECT 820.950 728.100 823.050 730.200 ;
        RECT 821.400 727.350 822.600 728.100 ;
        RECT 814.950 724.950 817.050 727.050 ;
        RECT 817.950 724.950 820.050 727.050 ;
        RECT 820.950 724.950 823.050 727.050 ;
        RECT 818.400 723.900 819.600 724.650 ;
        RECT 817.950 721.800 820.050 723.900 ;
        RECT 823.950 721.950 826.050 724.050 ;
        RECT 805.950 706.950 808.050 709.050 ;
        RECT 781.950 694.950 784.050 697.050 ;
        RECT 796.950 694.950 799.050 697.050 ;
        RECT 781.950 691.800 784.050 693.900 ;
        RECT 782.400 688.200 783.450 691.800 ;
        RECT 781.950 686.100 784.050 688.200 ;
        RECT 781.950 682.950 784.050 685.050 ;
        RECT 787.950 684.000 790.050 688.050 ;
        RECT 782.400 682.350 783.600 682.950 ;
        RECT 788.400 682.350 789.600 684.000 ;
        RECT 793.950 682.950 796.050 688.050 ;
        RECT 775.950 679.950 778.050 682.050 ;
        RECT 781.950 679.950 784.050 682.050 ;
        RECT 784.950 679.950 787.050 682.050 ;
        RECT 787.950 679.950 790.050 682.050 ;
        RECT 790.950 679.950 793.050 682.050 ;
        RECT 763.950 664.950 766.050 667.050 ;
        RECT 751.950 649.950 754.050 652.050 ;
        RECT 757.950 651.000 760.050 655.050 ;
        RECT 764.400 651.600 765.450 664.950 ;
        RECT 767.400 652.050 768.450 676.950 ;
        RECT 769.950 676.800 772.050 678.900 ;
        RECT 772.950 676.950 775.050 679.050 ;
        RECT 776.400 655.050 777.450 679.950 ;
        RECT 778.950 676.950 781.050 679.050 ;
        RECT 785.400 678.000 786.600 679.650 ;
        RECT 779.400 667.050 780.450 676.950 ;
        RECT 784.950 673.950 787.050 678.000 ;
        RECT 791.400 677.400 792.600 679.650 ;
        RECT 791.400 670.050 792.450 677.400 ;
        RECT 790.950 667.950 793.050 670.050 ;
        RECT 778.950 664.950 781.050 667.050 ;
        RECT 769.950 652.950 772.050 655.050 ;
        RECT 775.950 652.950 778.050 655.050 ;
        RECT 758.400 649.350 759.600 651.000 ;
        RECT 764.400 649.350 765.600 651.600 ;
        RECT 766.950 649.950 769.050 652.050 ;
        RECT 754.950 646.950 757.050 649.050 ;
        RECT 757.950 646.950 760.050 649.050 ;
        RECT 760.950 646.950 763.050 649.050 ;
        RECT 763.950 646.950 766.050 649.050 ;
        RECT 755.400 644.400 756.600 646.650 ;
        RECT 761.400 645.900 762.600 646.650 ;
        RECT 745.950 640.950 748.050 643.050 ;
        RECT 748.950 640.950 751.050 643.050 ;
        RECT 742.950 637.950 745.050 640.050 ;
        RECT 733.950 631.950 736.050 634.050 ;
        RECT 734.400 628.050 735.450 631.950 ;
        RECT 733.950 625.950 736.050 628.050 ;
        RECT 743.400 607.200 744.450 637.950 ;
        RECT 755.400 616.050 756.450 644.400 ;
        RECT 760.950 643.800 763.050 645.900 ;
        RECT 761.400 628.050 762.450 643.800 ;
        RECT 760.950 625.950 763.050 628.050 ;
        RECT 754.950 613.950 757.050 616.050 ;
        RECT 760.950 613.950 763.050 616.050 ;
        RECT 745.950 607.950 748.050 610.050 ;
        RECT 728.400 606.450 729.600 606.600 ;
        RECT 725.400 605.400 729.600 606.450 ;
        RECT 722.400 598.050 723.450 605.100 ;
        RECT 728.400 604.350 729.600 605.400 ;
        RECT 733.950 605.100 736.050 607.200 ;
        RECT 742.950 605.100 745.050 607.200 ;
        RECT 734.400 604.350 735.600 605.100 ;
        RECT 727.950 601.950 730.050 604.050 ;
        RECT 730.950 601.950 733.050 604.050 ;
        RECT 733.950 601.950 736.050 604.050 ;
        RECT 736.950 601.950 739.050 604.050 ;
        RECT 731.400 600.000 732.600 601.650 ;
        RECT 721.950 595.950 724.050 598.050 ;
        RECT 730.950 597.450 733.050 600.000 ;
        RECT 728.400 596.400 733.050 597.450 ;
        RECT 718.950 583.950 721.050 586.050 ;
        RECT 724.950 583.950 727.050 586.050 ;
        RECT 718.950 580.800 721.050 582.900 ;
        RECT 712.950 571.950 715.050 574.050 ;
        RECT 719.400 573.600 720.450 580.800 ;
        RECT 725.400 574.050 726.450 583.950 ;
        RECT 719.400 571.350 720.600 573.600 ;
        RECT 724.950 571.950 727.050 574.050 ;
        RECT 715.950 568.950 718.050 571.050 ;
        RECT 718.950 568.950 721.050 571.050 ;
        RECT 721.950 568.950 724.050 571.050 ;
        RECT 712.950 565.950 715.050 568.050 ;
        RECT 716.400 567.000 717.600 568.650 ;
        RECT 703.950 562.950 706.050 565.050 ;
        RECT 709.950 562.950 712.050 565.050 ;
        RECT 692.400 556.050 693.450 562.950 ;
        RECT 691.950 553.950 694.050 556.050 ;
        RECT 704.400 538.050 705.450 562.950 ;
        RECT 713.400 541.050 714.450 565.950 ;
        RECT 715.950 562.950 718.050 567.000 ;
        RECT 722.400 566.400 723.600 568.650 ;
        RECT 722.400 564.450 723.450 566.400 ;
        RECT 724.950 565.950 727.050 568.050 ;
        RECT 719.400 563.400 723.450 564.450 ;
        RECT 712.950 538.950 715.050 541.050 ;
        RECT 703.950 535.950 706.050 538.050 ;
        RECT 691.950 529.950 694.050 532.050 ;
        RECT 692.400 505.050 693.450 529.950 ;
        RECT 697.950 528.000 700.050 532.050 ;
        RECT 703.950 528.000 706.050 532.050 ;
        RECT 712.950 529.950 715.050 532.050 ;
        RECT 698.400 526.350 699.600 528.000 ;
        RECT 704.400 526.350 705.600 528.000 ;
        RECT 697.950 523.950 700.050 526.050 ;
        RECT 700.950 523.950 703.050 526.050 ;
        RECT 703.950 523.950 706.050 526.050 ;
        RECT 706.950 523.950 709.050 526.050 ;
        RECT 701.400 522.900 702.600 523.650 ;
        RECT 700.950 517.950 703.050 522.900 ;
        RECT 707.400 521.400 708.600 523.650 ;
        RECT 707.400 514.050 708.450 521.400 ;
        RECT 713.400 520.050 714.450 529.950 ;
        RECT 719.400 529.050 720.450 563.400 ;
        RECT 725.400 541.050 726.450 565.950 ;
        RECT 728.400 559.050 729.450 596.400 ;
        RECT 730.950 595.950 733.050 596.400 ;
        RECT 737.400 599.400 738.600 601.650 ;
        RECT 737.400 592.050 738.450 599.400 ;
        RECT 739.950 595.950 742.050 598.050 ;
        RECT 736.950 589.950 739.050 592.050 ;
        RECT 730.950 583.950 733.050 586.050 ;
        RECT 727.950 556.950 730.050 559.050 ;
        RECT 731.400 544.050 732.450 583.950 ;
        RECT 740.400 579.450 741.450 595.950 ;
        RECT 743.400 586.050 744.450 605.100 ;
        RECT 746.400 589.050 747.450 607.950 ;
        RECT 754.950 606.000 757.050 610.050 ;
        RECT 761.400 606.600 762.450 613.950 ;
        RECT 755.400 604.350 756.600 606.000 ;
        RECT 761.400 604.350 762.600 606.600 ;
        RECT 751.950 601.950 754.050 604.050 ;
        RECT 754.950 601.950 757.050 604.050 ;
        RECT 757.950 601.950 760.050 604.050 ;
        RECT 760.950 601.950 763.050 604.050 ;
        RECT 752.400 600.450 753.600 601.650 ;
        RECT 758.400 600.900 759.600 601.650 ;
        RECT 770.400 601.050 771.450 652.950 ;
        RECT 778.950 650.100 781.050 652.200 ;
        RECT 784.950 650.100 787.050 655.050 ;
        RECT 793.950 650.100 796.050 652.200 ;
        RECT 779.400 649.350 780.600 650.100 ;
        RECT 785.400 649.350 786.600 650.100 ;
        RECT 778.950 646.950 781.050 649.050 ;
        RECT 781.950 646.950 784.050 649.050 ;
        RECT 784.950 646.950 787.050 649.050 ;
        RECT 787.950 646.950 790.050 649.050 ;
        RECT 782.400 645.000 783.600 646.650 ;
        RECT 788.400 645.900 789.600 646.650 ;
        RECT 781.950 640.950 784.050 645.000 ;
        RECT 787.950 643.800 790.050 645.900 ;
        RECT 788.400 616.050 789.450 643.800 ;
        RECT 794.400 640.050 795.450 650.100 ;
        RECT 797.400 646.050 798.450 694.950 ;
        RECT 799.950 683.100 802.050 685.200 ;
        RECT 805.950 683.100 808.050 685.200 ;
        RECT 811.950 684.000 814.050 688.050 ;
        RECT 820.950 685.950 823.050 688.050 ;
        RECT 800.400 676.050 801.450 683.100 ;
        RECT 806.400 682.350 807.600 683.100 ;
        RECT 812.400 682.350 813.600 684.000 ;
        RECT 805.950 679.950 808.050 682.050 ;
        RECT 808.950 679.950 811.050 682.050 ;
        RECT 811.950 679.950 814.050 682.050 ;
        RECT 814.950 679.950 817.050 682.050 ;
        RECT 809.400 678.000 810.600 679.650 ;
        RECT 799.950 673.950 802.050 676.050 ;
        RECT 808.950 673.950 811.050 678.000 ;
        RECT 815.400 677.400 816.600 679.650 ;
        RECT 815.400 664.050 816.450 677.400 ;
        RECT 821.400 676.050 822.450 685.950 ;
        RECT 824.400 676.050 825.450 721.950 ;
        RECT 827.400 688.050 828.450 730.950 ;
        RECT 830.400 688.050 831.450 793.950 ;
        RECT 833.400 730.050 834.450 797.400 ;
        RECT 848.400 781.050 849.450 808.950 ;
        RECT 847.950 778.950 850.050 781.050 ;
        RECT 851.400 772.050 852.450 811.950 ;
        RECT 857.400 811.050 858.450 875.400 ;
        RECT 859.950 874.950 862.050 879.000 ;
        RECT 865.800 877.950 868.050 879.000 ;
        RECT 868.950 877.950 871.050 880.050 ;
        RECT 865.950 876.450 868.050 877.950 ;
        RECT 863.400 876.000 868.050 876.450 ;
        RECT 863.400 875.400 867.450 876.000 ;
        RECT 859.950 841.950 862.050 844.050 ;
        RECT 860.400 826.050 861.450 841.950 ;
        RECT 863.400 841.050 864.450 875.400 ;
        RECT 872.400 847.050 873.450 884.100 ;
        RECT 878.400 883.350 879.600 884.100 ;
        RECT 884.400 883.350 885.600 884.100 ;
        RECT 877.950 880.950 880.050 883.050 ;
        RECT 880.950 880.950 883.050 883.050 ;
        RECT 883.950 880.950 886.050 883.050 ;
        RECT 881.400 879.900 882.600 880.650 ;
        RECT 880.950 877.800 883.050 879.900 ;
        RECT 890.400 868.050 891.450 889.950 ;
        RECT 889.950 865.950 892.050 868.050 ;
        RECT 893.400 865.050 894.450 895.950 ;
        RECT 902.400 885.600 903.450 910.800 ;
        RECT 911.400 886.200 912.450 919.950 ;
        RECT 914.400 904.050 915.450 925.950 ;
        RECT 913.950 901.950 916.050 904.050 ;
        RECT 902.400 883.350 903.600 885.600 ;
        RECT 910.950 884.100 913.050 886.200 ;
        RECT 917.400 885.450 918.450 940.950 ;
        RECT 943.950 931.950 946.050 934.050 ;
        RECT 922.950 921.750 925.050 922.200 ;
        RECT 933.000 921.750 937.050 922.050 ;
        RECT 922.950 920.700 937.050 921.750 ;
        RECT 922.950 920.100 925.050 920.700 ;
        RECT 932.400 919.950 937.050 920.700 ;
        RECT 922.950 916.950 925.050 919.050 ;
        RECT 932.400 918.600 933.450 919.950 ;
        RECT 923.400 916.350 924.600 916.950 ;
        RECT 932.400 916.350 933.600 918.600 ;
        RECT 937.950 916.950 940.050 919.050 ;
        RECT 923.100 913.950 925.200 916.050 ;
        RECT 928.500 913.950 930.600 916.050 ;
        RECT 931.800 913.950 933.900 916.050 ;
        RECT 929.400 911.400 930.600 913.650 ;
        RECT 929.400 907.050 930.450 911.400 ;
        RECT 934.950 910.950 937.050 913.050 ;
        RECT 922.950 904.950 925.050 907.050 ;
        RECT 928.950 904.950 931.050 907.050 ;
        RECT 914.400 884.400 918.450 885.450 ;
        RECT 923.400 885.600 924.450 904.950 ;
        RECT 898.950 880.950 901.050 883.050 ;
        RECT 901.950 880.950 904.050 883.050 ;
        RECT 904.950 880.950 907.050 883.050 ;
        RECT 899.400 878.400 900.600 880.650 ;
        RECT 905.400 879.900 906.600 880.650 ;
        RECT 880.950 862.950 883.050 865.050 ;
        RECT 892.950 862.950 895.050 865.050 ;
        RECT 871.950 844.950 874.050 847.050 ;
        RECT 862.950 838.950 865.050 841.050 ;
        RECT 868.950 840.000 871.050 844.050 ;
        RECT 869.400 838.350 870.600 840.000 ;
        RECT 874.950 839.100 877.050 841.200 ;
        RECT 875.400 838.350 876.600 839.100 ;
        RECT 865.950 835.950 868.050 838.050 ;
        RECT 868.950 835.950 871.050 838.050 ;
        RECT 871.950 835.950 874.050 838.050 ;
        RECT 874.950 835.950 877.050 838.050 ;
        RECT 866.400 834.900 867.600 835.650 ;
        RECT 872.400 834.900 873.600 835.650 ;
        RECT 865.950 832.800 868.050 834.900 ;
        RECT 871.950 832.800 874.050 834.900 ;
        RECT 877.950 832.950 880.050 835.050 ;
        RECT 872.400 831.450 873.450 832.800 ;
        RECT 869.400 830.400 873.450 831.450 ;
        RECT 859.950 823.950 862.050 826.050 ;
        RECT 859.950 811.950 862.050 814.050 ;
        RECT 856.950 808.950 859.050 811.050 ;
        RECT 860.400 807.600 861.450 811.950 ;
        RECT 869.400 808.200 870.450 830.400 ;
        RECT 874.950 829.950 877.050 832.050 ;
        RECT 871.950 823.950 874.050 826.050 ;
        RECT 860.400 805.350 861.600 807.600 ;
        RECT 868.950 806.100 871.050 808.200 ;
        RECT 856.950 802.950 859.050 805.050 ;
        RECT 859.950 802.950 862.050 805.050 ;
        RECT 862.950 802.950 865.050 805.050 ;
        RECT 857.400 801.450 858.600 802.650 ;
        RECT 863.400 801.900 864.600 802.650 ;
        RECT 854.400 800.400 858.600 801.450 ;
        RECT 854.400 796.050 855.450 800.400 ;
        RECT 862.950 799.800 865.050 801.900 ;
        RECT 869.400 796.050 870.450 806.100 ;
        RECT 853.950 793.950 856.050 796.050 ;
        RECT 868.950 793.950 871.050 796.050 ;
        RECT 854.400 790.050 855.450 793.950 ;
        RECT 853.950 787.950 856.050 790.050 ;
        RECT 850.950 769.950 853.050 772.050 ;
        RECT 838.950 762.000 841.050 766.050 ;
        RECT 839.400 760.350 840.600 762.000 ;
        RECT 844.950 761.100 847.050 766.050 ;
        RECT 853.950 763.950 856.050 766.050 ;
        RECT 856.950 763.950 862.050 766.050 ;
        RECT 845.400 760.350 846.600 761.100 ;
        RECT 838.950 757.950 841.050 760.050 ;
        RECT 841.950 757.950 844.050 760.050 ;
        RECT 844.950 757.950 847.050 760.050 ;
        RECT 842.400 755.400 843.600 757.650 ;
        RECT 854.400 756.900 855.450 763.950 ;
        RECT 860.400 762.450 861.600 762.600 ;
        RECT 857.400 761.400 861.600 762.450 ;
        RECT 868.950 762.000 871.050 766.050 ;
        RECT 842.400 733.200 843.450 755.400 ;
        RECT 853.950 754.800 856.050 756.900 ;
        RECT 857.400 739.050 858.450 761.400 ;
        RECT 860.400 760.350 861.600 761.400 ;
        RECT 869.400 760.350 870.600 762.000 ;
        RECT 860.100 757.950 862.200 760.050 ;
        RECT 863.400 757.950 865.500 760.050 ;
        RECT 868.800 757.950 870.900 760.050 ;
        RECT 863.400 756.900 864.600 757.650 ;
        RECT 862.950 754.800 865.050 756.900 ;
        RECT 872.400 753.450 873.450 823.950 ;
        RECT 875.400 808.050 876.450 829.950 ;
        RECT 878.400 814.050 879.450 832.950 ;
        RECT 881.400 832.050 882.450 862.950 ;
        RECT 899.400 847.050 900.450 878.400 ;
        RECT 904.950 877.800 907.050 879.900 ;
        RECT 905.400 876.450 906.450 877.800 ;
        RECT 902.400 875.400 906.450 876.450 ;
        RECT 886.950 844.950 889.050 847.050 ;
        RECT 898.950 844.950 901.050 847.050 ;
        RECT 883.950 839.100 886.050 841.200 ;
        RECT 887.400 841.050 888.450 844.950 ;
        RECT 880.950 829.950 883.050 832.050 ;
        RECT 884.400 820.050 885.450 839.100 ;
        RECT 886.950 838.950 889.050 841.050 ;
        RECT 889.950 839.100 892.050 841.200 ;
        RECT 895.950 840.000 898.050 844.050 ;
        RECT 902.400 841.050 903.450 875.400 ;
        RECT 904.950 868.950 907.050 871.050 ;
        RECT 890.400 838.350 891.600 839.100 ;
        RECT 896.400 838.350 897.600 840.000 ;
        RECT 901.950 838.950 904.050 841.050 ;
        RECT 889.950 835.950 892.050 838.050 ;
        RECT 892.950 835.950 895.050 838.050 ;
        RECT 895.950 835.950 898.050 838.050 ;
        RECT 898.950 835.950 901.050 838.050 ;
        RECT 893.400 834.900 894.600 835.650 ;
        RECT 899.400 834.900 900.600 835.650 ;
        RECT 892.950 832.800 895.050 834.900 ;
        RECT 898.950 832.800 901.050 834.900 ;
        RECT 901.950 832.950 904.050 835.050 ;
        RECT 895.950 823.950 898.050 826.050 ;
        RECT 883.950 817.950 886.050 820.050 ;
        RECT 892.950 817.950 895.050 820.050 ;
        RECT 877.950 811.950 880.050 814.050 ;
        RECT 874.950 805.950 877.050 808.050 ;
        RECT 880.950 806.100 883.050 808.200 ;
        RECT 886.950 806.100 889.050 808.200 ;
        RECT 881.400 805.350 882.600 806.100 ;
        RECT 887.400 805.350 888.600 806.100 ;
        RECT 877.950 802.950 880.050 805.050 ;
        RECT 880.950 802.950 883.050 805.050 ;
        RECT 883.950 802.950 886.050 805.050 ;
        RECT 886.950 802.950 889.050 805.050 ;
        RECT 874.950 799.950 877.050 802.050 ;
        RECT 878.400 801.900 879.600 802.650 ;
        RECT 884.400 801.900 885.600 802.650 ;
        RECT 893.400 802.050 894.450 817.950 ;
        RECT 869.400 752.400 873.450 753.450 ;
        RECT 850.950 736.950 853.050 739.050 ;
        RECT 856.950 736.950 859.050 739.050 ;
        RECT 841.950 731.100 844.050 733.200 ;
        RECT 832.950 727.950 835.050 730.050 ;
        RECT 835.950 728.100 838.050 730.200 ;
        RECT 836.400 727.350 837.600 728.100 ;
        RECT 841.950 727.950 844.050 730.050 ;
        RECT 842.400 727.350 843.600 727.950 ;
        RECT 835.950 724.950 838.050 727.050 ;
        RECT 838.950 724.950 841.050 727.050 ;
        RECT 841.950 724.950 844.050 727.050 ;
        RECT 844.950 724.950 847.050 727.050 ;
        RECT 839.400 723.000 840.600 724.650 ;
        RECT 845.400 724.050 846.600 724.650 ;
        RECT 832.950 718.950 835.050 721.050 ;
        RECT 838.950 718.950 841.050 723.000 ;
        RECT 845.400 722.400 850.050 724.050 ;
        RECT 851.400 723.900 852.450 736.950 ;
        RECT 857.400 724.050 858.450 736.950 ;
        RECT 862.950 729.000 865.050 733.050 ;
        RECT 869.400 729.600 870.450 752.400 ;
        RECT 875.400 730.050 876.450 799.950 ;
        RECT 877.950 799.800 880.050 801.900 ;
        RECT 883.950 799.800 886.050 801.900 ;
        RECT 892.950 799.950 895.050 802.050 ;
        RECT 877.950 793.950 880.050 796.050 ;
        RECT 863.400 727.350 864.600 729.000 ;
        RECT 869.400 727.350 870.600 729.600 ;
        RECT 874.950 727.950 877.050 730.050 ;
        RECT 862.950 724.950 865.050 727.050 ;
        RECT 865.950 724.950 868.050 727.050 ;
        RECT 868.950 724.950 871.050 727.050 ;
        RECT 871.950 724.950 874.050 727.050 ;
        RECT 846.000 721.950 850.050 722.400 ;
        RECT 850.950 721.800 853.050 723.900 ;
        RECT 856.950 721.950 859.050 724.050 ;
        RECT 866.400 722.400 867.600 724.650 ;
        RECT 872.400 723.900 873.600 724.650 ;
        RECT 844.950 718.950 847.050 721.050 ;
        RECT 866.400 720.450 867.450 722.400 ;
        RECT 871.950 721.800 874.050 723.900 ;
        RECT 863.400 719.400 867.450 720.450 ;
        RECT 826.950 685.950 829.050 688.050 ;
        RECT 829.950 685.950 832.050 688.050 ;
        RECT 833.400 684.600 834.450 718.950 ;
        RECT 838.950 694.950 841.050 697.050 ;
        RECT 833.400 682.350 834.600 684.600 ;
        RECT 829.950 679.950 832.050 682.050 ;
        RECT 832.950 679.950 835.050 682.050 ;
        RECT 826.950 676.950 829.050 679.050 ;
        RECT 830.400 678.900 831.600 679.650 ;
        RECT 817.950 673.950 820.050 676.050 ;
        RECT 820.950 673.950 823.050 676.050 ;
        RECT 823.950 673.950 826.050 676.050 ;
        RECT 814.950 661.950 817.050 664.050 ;
        RECT 811.950 655.950 814.050 658.050 ;
        RECT 805.950 650.100 808.050 652.200 ;
        RECT 812.400 651.600 813.450 655.950 ;
        RECT 806.400 649.350 807.600 650.100 ;
        RECT 812.400 649.350 813.600 651.600 ;
        RECT 802.950 646.950 805.050 649.050 ;
        RECT 805.950 646.950 808.050 649.050 ;
        RECT 808.950 646.950 811.050 649.050 ;
        RECT 811.950 646.950 814.050 649.050 ;
        RECT 796.950 643.950 799.050 646.050 ;
        RECT 803.400 645.900 804.600 646.650 ;
        RECT 802.950 643.800 805.050 645.900 ;
        RECT 809.400 645.000 810.600 646.650 ;
        RECT 808.950 640.950 811.050 645.000 ;
        RECT 814.950 643.950 817.050 646.050 ;
        RECT 793.950 637.950 796.050 640.050 ;
        RECT 808.950 637.800 811.050 639.900 ;
        RECT 793.950 634.800 796.050 636.900 ;
        RECT 787.950 613.950 790.050 616.050 ;
        RECT 775.950 605.100 778.050 607.200 ;
        RECT 776.400 604.350 777.600 605.100 ;
        RECT 775.950 601.950 778.050 604.050 ;
        RECT 778.950 601.950 781.050 604.050 ;
        RECT 781.950 601.950 784.050 604.050 ;
        RECT 749.400 599.400 753.600 600.450 ;
        RECT 749.400 595.050 750.450 599.400 ;
        RECT 757.950 598.800 760.050 600.900 ;
        RECT 769.950 598.950 772.050 601.050 ;
        RECT 779.400 599.400 780.600 601.650 ;
        RECT 794.400 600.450 795.450 634.800 ;
        RECT 802.950 605.100 805.050 607.200 ;
        RECT 803.400 604.350 804.600 605.100 ;
        RECT 799.950 601.950 802.050 604.050 ;
        RECT 802.950 601.950 805.050 604.050 ;
        RECT 794.400 599.400 798.450 600.450 ;
        RECT 748.950 592.950 751.050 595.050 ;
        RECT 745.950 586.950 748.050 589.050 ;
        RECT 742.950 583.950 745.050 586.050 ;
        RECT 749.400 580.050 750.450 592.950 ;
        RECT 751.950 580.950 754.050 583.050 ;
        RECT 740.400 578.400 744.450 579.450 ;
        RECT 736.950 572.100 739.050 574.200 ;
        RECT 743.400 573.600 744.450 578.400 ;
        RECT 748.950 577.950 751.050 580.050 ;
        RECT 737.400 571.350 738.600 572.100 ;
        RECT 743.400 571.350 744.600 573.600 ;
        RECT 748.950 571.950 751.050 576.900 ;
        RECT 736.950 568.950 739.050 571.050 ;
        RECT 739.950 568.950 742.050 571.050 ;
        RECT 742.950 568.950 745.050 571.050 ;
        RECT 745.950 568.950 748.050 571.050 ;
        RECT 740.400 566.400 741.600 568.650 ;
        RECT 746.400 567.900 747.600 568.650 ;
        RECT 752.400 567.900 753.450 580.950 ;
        RECT 754.950 572.100 757.050 574.200 ;
        RECT 763.950 572.100 766.050 574.200 ;
        RECT 769.950 572.100 772.050 574.200 ;
        RECT 740.400 547.050 741.450 566.400 ;
        RECT 745.950 565.800 748.050 567.900 ;
        RECT 751.950 565.800 754.050 567.900 ;
        RECT 755.400 547.050 756.450 572.100 ;
        RECT 764.400 571.350 765.600 572.100 ;
        RECT 770.400 571.350 771.600 572.100 ;
        RECT 760.950 568.950 763.050 571.050 ;
        RECT 763.950 568.950 766.050 571.050 ;
        RECT 766.950 568.950 769.050 571.050 ;
        RECT 769.950 568.950 772.050 571.050 ;
        RECT 757.950 565.950 760.050 568.050 ;
        RECT 761.400 566.400 762.600 568.650 ;
        RECT 767.400 567.900 768.600 568.650 ;
        RECT 779.400 567.900 780.450 599.400 ;
        RECT 790.950 580.950 793.050 583.050 ;
        RECT 781.950 571.950 784.050 574.050 ;
        RECT 791.400 573.600 792.450 580.950 ;
        RECT 739.950 544.950 742.050 547.050 ;
        RECT 748.950 544.950 751.050 547.050 ;
        RECT 754.950 544.950 757.050 547.050 ;
        RECT 730.950 541.950 733.050 544.050 ;
        RECT 736.950 541.950 739.050 544.050 ;
        RECT 724.950 538.950 727.050 541.050 ;
        RECT 718.950 526.950 721.050 529.050 ;
        RECT 721.950 528.000 724.050 532.050 ;
        RECT 727.950 528.000 730.050 532.050 ;
        RECT 722.400 526.350 723.600 528.000 ;
        RECT 728.400 526.350 729.600 528.000 ;
        RECT 721.950 523.950 724.050 526.050 ;
        RECT 724.950 523.950 727.050 526.050 ;
        RECT 727.950 523.950 730.050 526.050 ;
        RECT 730.950 523.950 733.050 526.050 ;
        RECT 718.950 520.950 721.050 523.050 ;
        RECT 725.400 521.400 726.600 523.650 ;
        RECT 731.400 522.000 732.600 523.650 ;
        RECT 712.950 517.950 715.050 520.050 ;
        RECT 706.950 511.950 709.050 514.050 ;
        RECT 703.950 510.450 706.050 511.050 ;
        RECT 709.950 510.450 712.050 511.050 ;
        RECT 703.950 509.400 712.050 510.450 ;
        RECT 703.950 508.950 706.050 509.400 ;
        RECT 709.950 508.950 712.050 509.400 ;
        RECT 691.950 502.950 694.050 505.050 ;
        RECT 691.950 496.950 694.050 499.050 ;
        RECT 692.400 489.450 693.450 496.950 ;
        RECT 700.950 494.100 703.050 496.200 ;
        RECT 701.400 493.350 702.600 494.100 ;
        RECT 695.100 490.950 697.200 493.050 ;
        RECT 700.500 490.950 702.600 493.050 ;
        RECT 703.800 490.950 705.900 493.050 ;
        RECT 712.950 490.950 715.050 493.050 ;
        RECT 695.400 489.450 696.600 490.650 ;
        RECT 692.400 488.400 696.600 489.450 ;
        RECT 704.400 488.400 705.600 490.650 ;
        RECT 688.950 484.950 691.050 487.050 ;
        RECT 694.950 484.950 697.050 487.050 ;
        RECT 682.950 475.950 685.050 478.050 ;
        RECT 670.950 469.950 673.050 472.050 ;
        RECT 658.950 442.800 661.050 444.900 ;
        RECT 667.950 442.950 670.050 445.050 ;
        RECT 671.400 442.050 672.450 469.950 ;
        RECT 691.950 466.950 694.050 469.050 ;
        RECT 692.400 457.050 693.450 466.950 ;
        RECT 691.950 454.950 694.050 457.050 ;
        RECT 676.950 449.100 679.050 451.200 ;
        RECT 682.950 449.100 685.050 451.200 ;
        RECT 691.950 449.100 694.050 451.200 ;
        RECT 677.400 448.350 678.600 449.100 ;
        RECT 683.400 448.350 684.600 449.100 ;
        RECT 676.950 445.950 679.050 448.050 ;
        RECT 679.950 445.950 682.050 448.050 ;
        RECT 682.950 445.950 685.050 448.050 ;
        RECT 673.950 442.950 676.050 445.050 ;
        RECT 680.400 444.900 681.600 445.650 ;
        RECT 692.400 445.050 693.450 449.100 ;
        RECT 670.950 439.950 673.050 442.050 ;
        RECT 674.400 436.050 675.450 442.950 ;
        RECT 679.950 442.800 682.050 444.900 ;
        RECT 691.950 442.950 694.050 445.050 ;
        RECT 676.950 439.950 679.050 442.050 ;
        RECT 673.950 433.950 676.050 436.050 ;
        RECT 647.400 415.350 648.600 416.100 ;
        RECT 649.950 415.950 652.050 418.050 ;
        RECT 652.950 415.800 655.050 417.900 ;
        RECT 655.950 415.950 658.050 418.050 ;
        RECT 664.950 416.100 667.050 418.200 ;
        RECT 637.950 412.950 640.050 415.050 ;
        RECT 640.950 412.950 643.050 415.050 ;
        RECT 643.950 412.950 646.050 415.050 ;
        RECT 646.950 412.950 649.050 415.050 ;
        RECT 638.400 411.900 639.600 412.650 ;
        RECT 623.400 406.050 624.450 410.400 ;
        RECT 631.950 409.800 634.050 411.900 ;
        RECT 637.950 409.800 640.050 411.900 ;
        RECT 644.400 410.400 645.600 412.650 ;
        RECT 622.950 403.950 625.050 406.050 ;
        RECT 616.950 397.950 619.050 400.050 ;
        RECT 610.950 376.950 613.050 379.050 ;
        RECT 608.400 370.350 609.600 372.600 ;
        RECT 607.950 367.950 610.050 370.050 ;
        RECT 610.950 367.950 613.050 370.050 ;
        RECT 611.400 366.900 612.600 367.650 ;
        RECT 610.950 364.800 613.050 366.900 ;
        RECT 607.950 361.950 610.050 364.050 ;
        RECT 601.950 355.950 604.050 358.050 ;
        RECT 608.400 355.050 609.450 361.950 ;
        RECT 613.950 355.950 616.050 358.050 ;
        RECT 607.950 352.950 610.050 355.050 ;
        RECT 599.550 345.300 601.650 347.400 ;
        RECT 595.950 340.950 598.050 343.050 ;
        RECT 599.550 332.400 600.750 345.300 ;
        RECT 604.950 339.000 607.050 343.050 ;
        RECT 605.400 337.350 606.600 339.000 ;
        RECT 604.950 334.950 607.050 337.050 ;
        RECT 599.550 330.300 601.650 332.400 ;
        RECT 607.950 331.800 610.050 333.900 ;
        RECT 592.950 322.950 595.050 325.050 ;
        RECT 599.550 323.700 600.750 330.300 ;
        RECT 599.550 321.600 601.650 323.700 ;
        RECT 604.950 322.950 607.050 325.050 ;
        RECT 601.950 316.950 604.050 319.050 ;
        RECT 580.950 310.950 583.050 313.050 ;
        RECT 575.250 296.700 576.450 303.300 ;
        RECT 577.950 301.950 580.050 304.050 ;
        RECT 574.350 294.600 576.450 296.700 ;
        RECT 563.400 292.350 564.600 294.600 ;
        RECT 559.950 289.950 562.050 292.050 ;
        RECT 562.950 289.950 565.050 292.050 ;
        RECT 568.950 289.950 571.050 292.050 ;
        RECT 560.400 288.900 561.600 289.650 ;
        RECT 569.400 288.900 570.600 289.650 ;
        RECT 559.950 286.800 562.050 288.900 ;
        RECT 568.950 286.800 571.050 288.900 ;
        RECT 559.950 283.650 562.050 285.750 ;
        RECT 541.950 277.950 544.050 280.050 ;
        RECT 553.950 277.950 556.050 280.050 ;
        RECT 526.950 274.950 529.050 277.050 ;
        RECT 538.950 274.950 541.050 277.050 ;
        RECT 523.950 271.950 526.050 274.050 ;
        RECT 511.950 268.950 514.050 271.050 ;
        RECT 520.950 268.950 523.050 271.050 ;
        RECT 512.400 261.600 513.450 268.950 ;
        RECT 527.400 265.050 528.450 274.950 ;
        RECT 539.400 271.050 540.450 274.950 ;
        RECT 538.950 268.950 541.050 271.050 ;
        RECT 542.400 268.050 543.450 277.950 ;
        RECT 560.400 277.050 561.450 283.650 ;
        RECT 575.250 281.700 576.450 294.600 ;
        RECT 577.950 289.950 580.050 292.050 ;
        RECT 565.950 277.950 568.050 280.050 ;
        RECT 574.350 279.600 576.450 281.700 ;
        RECT 559.950 274.950 562.050 277.050 ;
        RECT 556.950 271.950 559.050 274.050 ;
        RECT 557.400 268.050 558.450 271.950 ;
        RECT 566.400 268.050 567.450 277.950 ;
        RECT 578.400 277.050 579.450 289.950 ;
        RECT 574.800 276.000 576.900 277.050 ;
        RECT 574.800 274.950 577.050 276.000 ;
        RECT 577.950 274.950 580.050 277.050 ;
        RECT 574.950 273.450 577.050 274.950 ;
        RECT 574.950 273.000 579.450 273.450 ;
        RECT 575.400 272.400 579.450 273.000 ;
        RECT 541.950 265.950 544.050 268.050 ;
        RECT 556.950 265.950 559.050 268.050 ;
        RECT 565.950 265.950 568.050 268.050 ;
        RECT 526.950 262.950 529.050 265.050 ;
        RECT 512.400 259.350 513.600 261.600 ;
        RECT 517.950 260.100 520.050 262.200 ;
        RECT 518.400 259.350 519.600 260.100 ;
        RECT 523.950 259.950 526.050 262.050 ;
        RECT 508.950 256.950 511.050 259.050 ;
        RECT 511.950 256.950 514.050 259.050 ;
        RECT 514.950 256.950 517.050 259.050 ;
        RECT 517.950 256.950 520.050 259.050 ;
        RECT 509.400 255.000 510.600 256.650 ;
        RECT 515.400 255.900 516.600 256.650 ;
        RECT 508.950 250.950 511.050 255.000 ;
        RECT 514.950 253.800 517.050 255.900 ;
        RECT 502.950 247.950 505.050 250.050 ;
        RECT 508.950 247.800 511.050 249.900 ;
        RECT 505.950 238.950 508.050 241.050 ;
        RECT 496.950 235.950 499.050 238.050 ;
        RECT 493.950 223.950 496.050 226.050 ;
        RECT 494.400 220.050 495.450 223.950 ;
        RECT 497.400 223.050 498.450 235.950 ;
        RECT 496.950 220.950 499.050 223.050 ;
        RECT 493.950 217.950 496.050 220.050 ;
        RECT 490.950 215.100 493.050 217.200 ;
        RECT 496.950 216.000 499.050 219.900 ;
        RECT 506.400 216.450 507.450 238.950 ;
        RECT 509.400 237.450 510.450 247.800 ;
        RECT 511.950 244.950 514.050 247.050 ;
        RECT 512.400 241.050 513.450 244.950 ;
        RECT 511.950 238.950 514.050 241.050 ;
        RECT 509.400 236.400 513.450 237.450 ;
        RECT 475.050 201.600 477.150 203.700 ;
        RECT 484.950 202.950 487.050 205.050 ;
        RECT 466.950 193.950 469.050 196.050 ;
        RECT 475.950 193.950 478.050 196.050 ;
        RECT 460.950 190.950 463.050 193.050 ;
        RECT 424.950 187.950 427.050 190.050 ;
        RECT 418.800 181.950 420.900 184.050 ;
        RECT 421.950 181.950 424.050 184.050 ;
        RECT 430.950 182.100 433.050 184.200 ;
        RECT 451.950 182.100 454.050 184.200 ;
        RECT 419.400 175.050 420.450 181.950 ;
        RECT 415.800 172.950 417.900 175.050 ;
        RECT 418.950 172.950 421.050 175.050 ;
        RECT 422.400 145.050 423.450 181.950 ;
        RECT 431.400 181.350 432.600 182.100 ;
        RECT 452.400 181.350 453.600 182.100 ;
        RECT 427.950 178.950 430.050 181.050 ;
        RECT 430.950 178.950 433.050 181.050 ;
        RECT 433.950 178.950 436.050 181.050 ;
        RECT 448.950 178.950 451.050 181.050 ;
        RECT 451.950 178.950 454.050 181.050 ;
        RECT 454.950 178.950 457.050 181.050 ;
        RECT 428.400 177.000 429.600 178.650 ;
        RECT 427.950 172.950 430.050 177.000 ;
        RECT 434.400 176.400 435.600 178.650 ;
        RECT 455.400 177.450 456.600 178.650 ;
        RECT 461.400 177.450 462.450 190.950 ;
        RECT 466.950 181.950 469.050 184.050 ;
        RECT 476.400 183.600 477.450 193.950 ;
        RECT 481.950 190.950 484.050 193.050 ;
        RECT 482.400 183.600 483.450 190.950 ;
        RECT 467.400 177.900 468.450 181.950 ;
        RECT 476.400 181.350 477.600 183.600 ;
        RECT 482.400 181.350 483.600 183.600 ;
        RECT 472.950 178.950 475.050 181.050 ;
        RECT 475.950 178.950 478.050 181.050 ;
        RECT 478.950 178.950 481.050 181.050 ;
        RECT 481.950 178.950 484.050 181.050 ;
        RECT 473.400 177.900 474.600 178.650 ;
        RECT 479.400 177.900 480.600 178.650 ;
        RECT 455.400 176.400 462.450 177.450 ;
        RECT 434.400 154.050 435.450 176.400 ;
        RECT 466.950 175.800 469.050 177.900 ;
        RECT 472.950 175.800 475.050 177.900 ;
        RECT 478.950 175.800 481.050 177.900 ;
        RECT 454.950 157.950 457.050 160.050 ;
        RECT 484.950 157.950 487.050 160.050 ;
        RECT 433.950 151.950 436.050 154.050 ;
        RECT 421.950 142.950 424.050 145.050 ;
        RECT 412.950 137.100 415.050 139.200 ;
        RECT 418.950 137.100 421.050 139.200 ;
        RECT 427.950 137.100 430.050 139.200 ;
        RECT 436.950 137.100 439.050 139.200 ;
        RECT 442.950 137.100 445.050 139.200 ;
        RECT 413.400 136.350 414.600 137.100 ;
        RECT 419.400 136.350 420.600 137.100 ;
        RECT 412.950 133.950 415.050 136.050 ;
        RECT 415.950 133.950 418.050 136.050 ;
        RECT 418.950 133.950 421.050 136.050 ;
        RECT 421.950 133.950 424.050 136.050 ;
        RECT 416.400 131.400 417.600 133.650 ;
        RECT 422.400 131.400 423.600 133.650 ;
        RECT 416.400 130.050 417.450 131.400 ;
        RECT 415.950 127.950 418.050 130.050 ;
        RECT 406.950 115.950 409.050 118.050 ;
        RECT 416.400 112.050 417.450 127.950 ;
        RECT 422.400 112.050 423.450 131.400 ;
        RECT 428.400 130.050 429.450 137.100 ;
        RECT 437.400 136.350 438.600 137.100 ;
        RECT 443.400 136.350 444.600 137.100 ;
        RECT 436.950 133.950 439.050 136.050 ;
        RECT 439.950 133.950 442.050 136.050 ;
        RECT 442.950 133.950 445.050 136.050 ;
        RECT 445.950 133.950 448.050 136.050 ;
        RECT 440.400 132.900 441.600 133.650 ;
        RECT 430.950 130.800 433.050 132.900 ;
        RECT 439.950 130.800 442.050 132.900 ;
        RECT 446.400 131.400 447.600 133.650 ;
        RECT 427.950 127.950 430.050 130.050 ;
        RECT 415.950 109.950 418.050 112.050 ;
        RECT 421.950 109.950 424.050 112.050 ;
        RECT 403.950 105.000 406.050 109.050 ;
        RECT 404.400 103.350 405.600 105.000 ;
        RECT 421.950 104.100 424.050 106.200 ;
        RECT 422.400 103.350 423.600 104.100 ;
        RECT 403.950 100.950 406.050 103.050 ;
        RECT 406.950 100.950 409.050 103.050 ;
        RECT 415.950 100.950 418.050 103.050 ;
        RECT 421.950 100.950 424.050 103.050 ;
        RECT 424.950 100.950 427.050 103.050 ;
        RECT 398.400 98.400 402.450 99.450 ;
        RECT 386.400 82.050 387.450 98.400 ;
        RECT 376.950 79.950 379.050 82.050 ;
        RECT 385.950 79.950 388.050 82.050 ;
        RECT 364.950 67.950 367.050 70.050 ;
        RECT 359.400 58.350 360.600 60.600 ;
        RECT 364.950 59.100 367.050 61.200 ;
        RECT 365.400 58.350 366.600 59.100 ;
        RECT 358.950 55.950 361.050 58.050 ;
        RECT 361.950 55.950 364.050 58.050 ;
        RECT 364.950 55.950 367.050 58.050 ;
        RECT 367.950 55.950 370.050 58.050 ;
        RECT 352.950 52.950 355.050 55.050 ;
        RECT 362.400 53.400 363.600 55.650 ;
        RECT 368.400 53.400 369.600 55.650 ;
        RECT 377.400 54.900 378.450 79.950 ;
        RECT 391.950 73.950 394.050 76.050 ;
        RECT 385.950 59.100 388.050 61.200 ;
        RECT 392.400 60.600 393.450 73.950 ;
        RECT 386.400 58.350 387.600 59.100 ;
        RECT 392.400 58.350 393.600 60.600 ;
        RECT 385.950 55.950 388.050 58.050 ;
        RECT 388.950 55.950 391.050 58.050 ;
        RECT 391.950 55.950 394.050 58.050 ;
        RECT 394.950 55.950 397.050 58.050 ;
        RECT 389.400 54.900 390.600 55.650 ;
        RECT 358.950 46.950 361.050 49.050 ;
        RECT 349.950 31.950 352.050 34.050 ;
        RECT 346.950 27.000 349.050 31.050 ;
        RECT 347.400 25.350 348.600 27.000 ;
        RECT 352.950 26.100 355.050 28.200 ;
        RECT 353.400 25.350 354.600 26.100 ;
        RECT 343.950 22.950 346.050 25.050 ;
        RECT 346.950 22.950 349.050 25.050 ;
        RECT 349.950 22.950 352.050 25.050 ;
        RECT 352.950 22.950 355.050 25.050 ;
        RECT 344.400 21.900 345.600 22.650 ;
        RECT 299.400 16.050 300.450 19.800 ;
        RECT 301.950 16.950 304.050 19.050 ;
        RECT 319.950 16.950 322.050 21.000 ;
        RECT 326.400 20.400 333.450 21.450 ;
        RECT 343.950 19.800 346.050 21.900 ;
        RECT 350.400 20.400 351.600 22.650 ;
        RECT 359.400 21.900 360.450 46.950 ;
        RECT 362.400 46.050 363.450 53.400 ;
        RECT 368.400 46.050 369.450 53.400 ;
        RECT 376.950 52.800 379.050 54.900 ;
        RECT 388.950 52.800 391.050 54.900 ;
        RECT 395.400 53.400 396.600 55.650 ;
        RECT 361.950 43.950 364.050 46.050 ;
        RECT 367.950 43.950 370.050 46.050 ;
        RECT 367.950 31.950 370.050 34.050 ;
        RECT 364.950 25.950 367.050 28.050 ;
        RECT 368.400 27.600 369.450 31.950 ;
        RECT 395.400 30.450 396.450 53.400 ;
        RECT 395.400 29.400 399.450 30.450 ;
        RECT 286.950 13.950 289.050 16.050 ;
        RECT 298.950 13.950 301.050 16.050 ;
        RECT 13.950 10.950 16.050 13.050 ;
        RECT 88.950 10.950 91.050 13.050 ;
        RECT 94.950 10.950 97.050 13.050 ;
        RECT 247.950 10.950 250.050 13.050 ;
        RECT 295.950 12.450 298.050 13.050 ;
        RECT 302.400 12.450 303.450 16.950 ;
        RECT 350.400 16.050 351.450 20.400 ;
        RECT 358.950 19.800 361.050 21.900 ;
        RECT 365.400 16.050 366.450 25.950 ;
        RECT 368.400 25.350 369.600 27.600 ;
        RECT 394.950 26.100 397.050 28.200 ;
        RECT 395.400 25.350 396.600 26.100 ;
        RECT 368.400 22.950 370.500 25.050 ;
        RECT 373.800 22.950 375.900 25.050 ;
        RECT 389.100 22.950 391.200 25.050 ;
        RECT 394.500 22.950 396.600 25.050 ;
        RECT 398.400 21.900 399.450 29.400 ;
        RECT 401.400 28.050 402.450 98.400 ;
        RECT 407.400 98.400 408.600 100.650 ;
        RECT 403.950 73.950 406.050 76.050 ;
        RECT 404.400 54.900 405.450 73.950 ;
        RECT 407.400 61.200 408.450 98.400 ;
        RECT 416.400 88.050 417.450 100.950 ;
        RECT 425.400 99.900 426.600 100.650 ;
        RECT 424.950 97.800 427.050 99.900 ;
        RECT 431.400 99.450 432.450 130.800 ;
        RECT 442.950 127.950 445.050 130.050 ;
        RECT 443.400 105.600 444.450 127.950 ;
        RECT 446.400 127.050 447.450 131.400 ;
        RECT 445.950 124.950 448.050 127.050 ;
        RECT 443.400 103.350 444.600 105.600 ;
        RECT 439.950 100.950 442.050 103.050 ;
        RECT 442.950 100.950 445.050 103.050 ;
        RECT 445.950 100.950 448.050 103.050 ;
        RECT 440.400 99.900 441.600 100.650 ;
        RECT 428.400 98.400 432.450 99.450 ;
        RECT 415.950 85.950 418.050 88.050 ;
        RECT 412.950 67.950 415.050 70.050 ;
        RECT 406.950 59.100 409.050 61.200 ;
        RECT 413.400 60.600 414.450 67.950 ;
        RECT 424.950 61.950 427.050 64.050 ;
        RECT 413.400 58.350 414.600 60.600 ;
        RECT 418.950 59.100 421.050 61.200 ;
        RECT 419.400 58.350 420.600 59.100 ;
        RECT 409.950 55.950 412.050 58.050 ;
        RECT 412.950 55.950 415.050 58.050 ;
        RECT 415.950 55.950 418.050 58.050 ;
        RECT 418.950 55.950 421.050 58.050 ;
        RECT 410.400 54.900 411.600 55.650 ;
        RECT 403.950 52.800 406.050 54.900 ;
        RECT 409.950 52.800 412.050 54.900 ;
        RECT 416.400 54.000 417.600 55.650 ;
        RECT 415.950 49.950 418.050 54.000 ;
        RECT 421.950 52.950 424.050 55.050 ;
        RECT 400.950 25.950 403.050 28.050 ;
        RECT 419.400 27.450 420.600 27.600 ;
        RECT 422.400 27.450 423.450 52.950 ;
        RECT 425.400 46.050 426.450 61.950 ;
        RECT 428.400 54.450 429.450 98.400 ;
        RECT 439.950 97.800 442.050 99.900 ;
        RECT 446.400 98.400 447.600 100.650 ;
        RECT 446.400 94.050 447.450 98.400 ;
        RECT 445.950 91.950 448.050 94.050 ;
        RECT 455.400 82.050 456.450 157.950 ;
        RECT 469.950 142.950 472.050 145.050 ;
        RECT 463.950 137.100 466.050 139.200 ;
        RECT 470.400 138.600 471.450 142.950 ;
        RECT 464.400 136.350 465.600 137.100 ;
        RECT 470.400 136.350 471.600 138.600 ;
        RECT 475.800 137.100 477.900 139.200 ;
        RECT 478.950 137.100 481.050 139.200 ;
        RECT 485.400 138.600 486.450 157.950 ;
        RECT 491.400 145.050 492.450 215.100 ;
        RECT 497.400 214.350 498.600 216.000 ;
        RECT 506.400 215.400 510.450 216.450 ;
        RECT 496.950 211.950 499.050 214.050 ;
        RECT 499.950 211.950 502.050 214.050 ;
        RECT 502.950 211.950 505.050 214.050 ;
        RECT 500.400 209.400 501.600 211.650 ;
        RECT 500.400 208.050 501.450 209.400 ;
        RECT 505.950 208.950 508.050 211.050 ;
        RECT 499.950 205.950 502.050 208.050 ;
        RECT 500.400 186.450 501.450 205.950 ;
        RECT 497.400 185.400 501.450 186.450 ;
        RECT 497.400 184.200 498.450 185.400 ;
        RECT 496.950 182.100 499.050 184.200 ;
        RECT 497.400 181.350 498.600 182.100 ;
        RECT 496.950 178.950 499.050 181.050 ;
        RECT 499.950 178.950 502.050 181.050 ;
        RECT 500.400 176.400 501.600 178.650 ;
        RECT 500.400 151.050 501.450 176.400 ;
        RECT 506.400 154.050 507.450 208.950 ;
        RECT 509.400 160.050 510.450 215.400 ;
        RECT 512.400 211.050 513.450 236.400 ;
        RECT 514.950 229.950 517.050 232.050 ;
        RECT 515.400 223.050 516.450 229.950 ;
        RECT 514.950 220.950 517.050 223.050 ;
        RECT 517.950 215.100 520.050 217.200 ;
        RECT 524.400 217.050 525.450 259.950 ;
        RECT 527.400 256.050 528.450 262.950 ;
        RECT 535.950 261.000 538.050 265.050 ;
        RECT 542.400 262.050 543.450 265.950 ;
        RECT 536.400 259.350 537.600 261.000 ;
        RECT 541.950 259.950 544.050 262.050 ;
        RECT 544.950 259.950 547.050 262.050 ;
        RECT 557.400 261.600 558.450 265.950 ;
        RECT 571.950 262.950 574.050 265.050 ;
        RECT 535.950 256.950 538.050 259.050 ;
        RECT 538.950 256.950 541.050 259.050 ;
        RECT 526.950 253.950 529.050 256.050 ;
        RECT 539.400 255.900 540.600 256.650 ;
        RECT 527.400 250.050 528.450 253.950 ;
        RECT 538.950 253.800 541.050 255.900 ;
        RECT 541.950 250.950 544.050 253.050 ;
        RECT 526.950 247.950 529.050 250.050 ;
        RECT 532.950 241.950 535.050 244.050 ;
        RECT 533.400 232.050 534.450 241.950 ;
        RECT 542.400 238.050 543.450 250.950 ;
        RECT 541.950 235.950 544.050 238.050 ;
        RECT 532.950 229.950 535.050 232.050 ;
        RECT 541.950 226.950 544.050 229.050 ;
        RECT 542.400 220.200 543.450 226.950 ;
        RECT 545.400 226.050 546.450 259.950 ;
        RECT 557.400 259.350 558.600 261.600 ;
        RECT 562.950 260.100 565.050 262.200 ;
        RECT 563.400 259.350 564.600 260.100 ;
        RECT 553.950 256.950 556.050 259.050 ;
        RECT 556.950 256.950 559.050 259.050 ;
        RECT 559.950 256.950 562.050 259.050 ;
        RECT 562.950 256.950 565.050 259.050 ;
        RECT 568.950 256.950 571.050 259.050 ;
        RECT 554.400 256.050 555.600 256.650 ;
        RECT 550.950 254.400 555.600 256.050 ;
        RECT 560.400 255.900 561.600 256.650 ;
        RECT 550.950 253.950 555.450 254.400 ;
        RECT 554.400 238.050 555.450 253.950 ;
        RECT 559.950 253.800 562.050 255.900 ;
        RECT 569.400 250.050 570.450 256.950 ;
        RECT 572.400 256.050 573.450 262.950 ;
        RECT 578.400 261.600 579.450 272.400 ;
        RECT 581.400 265.050 582.450 310.950 ;
        RECT 598.950 304.950 601.050 307.050 ;
        RECT 589.650 301.500 591.750 302.400 ;
        RECT 595.950 301.950 598.050 304.050 ;
        RECT 589.650 300.300 593.850 301.500 ;
        RECT 586.950 293.100 589.050 295.200 ;
        RECT 587.400 292.350 588.600 293.100 ;
        RECT 586.800 289.950 588.900 292.050 ;
        RECT 592.650 281.700 593.850 300.300 ;
        RECT 596.400 294.600 597.450 301.950 ;
        RECT 599.400 301.050 600.450 304.950 ;
        RECT 598.950 298.950 601.050 301.050 ;
        RECT 596.400 292.350 597.600 294.600 ;
        RECT 595.950 289.950 598.050 292.050 ;
        RECT 592.050 279.600 594.150 281.700 ;
        RECT 602.400 280.050 603.450 316.950 ;
        RECT 601.950 277.950 604.050 280.050 ;
        RECT 583.950 265.950 586.050 268.050 ;
        RECT 589.950 265.950 592.050 268.050 ;
        RECT 580.950 262.950 583.050 265.050 ;
        RECT 584.400 261.600 585.450 265.950 ;
        RECT 590.400 262.050 591.450 265.950 ;
        RECT 605.400 265.050 606.450 322.950 ;
        RECT 608.400 310.050 609.450 331.800 ;
        RECT 607.950 307.950 610.050 310.050 ;
        RECT 607.950 304.050 610.050 306.900 ;
        RECT 607.950 303.000 613.050 304.050 ;
        RECT 608.400 302.400 613.050 303.000 ;
        RECT 609.000 301.950 613.050 302.400 ;
        RECT 614.400 294.600 615.450 355.950 ;
        RECT 617.400 334.050 618.450 397.950 ;
        RECT 619.950 376.950 622.050 379.050 ;
        RECT 620.400 366.900 621.450 376.950 ;
        RECT 623.400 376.050 624.450 403.950 ;
        RECT 644.400 400.050 645.450 410.400 ;
        RECT 653.400 406.050 654.450 415.800 ;
        RECT 652.950 403.950 655.050 406.050 ;
        RECT 643.950 397.950 646.050 400.050 ;
        RECT 625.950 391.950 628.050 394.050 ;
        RECT 626.400 382.050 627.450 391.950 ;
        RECT 656.400 391.050 657.450 415.950 ;
        RECT 665.400 415.350 666.600 416.100 ;
        RECT 661.950 412.950 664.050 415.050 ;
        RECT 664.950 412.950 667.050 415.050 ;
        RECT 667.950 412.950 670.050 415.050 ;
        RECT 668.400 411.000 669.600 412.650 ;
        RECT 667.950 406.950 670.050 411.000 ;
        RECT 670.950 409.950 673.050 412.050 ;
        RECT 667.950 403.800 670.050 405.900 ;
        RECT 655.950 388.950 658.050 391.050 ;
        RECT 631.950 385.950 634.050 388.050 ;
        RECT 625.950 379.950 628.050 382.050 ;
        RECT 622.950 373.950 625.050 376.050 ;
        RECT 626.400 372.600 627.450 379.950 ;
        RECT 632.400 372.600 633.450 385.950 ;
        RECT 652.950 379.950 655.050 382.050 ;
        RECT 653.400 372.600 654.450 379.950 ;
        RECT 626.400 370.350 627.600 372.600 ;
        RECT 632.400 370.350 633.600 372.600 ;
        RECT 653.400 370.350 654.600 372.600 ;
        RECT 658.950 371.100 661.050 373.200 ;
        RECT 659.400 370.350 660.600 371.100 ;
        RECT 625.950 367.950 628.050 370.050 ;
        RECT 628.950 367.950 631.050 370.050 ;
        RECT 631.950 367.950 634.050 370.050 ;
        RECT 634.950 367.950 637.050 370.050 ;
        RECT 652.950 367.950 655.050 370.050 ;
        RECT 655.950 367.950 658.050 370.050 ;
        RECT 658.950 367.950 661.050 370.050 ;
        RECT 661.950 367.950 664.050 370.050 ;
        RECT 629.400 366.900 630.600 367.650 ;
        RECT 619.950 364.800 622.050 366.900 ;
        RECT 628.950 364.800 631.050 366.900 ;
        RECT 635.400 365.400 636.600 367.650 ;
        RECT 656.400 365.400 657.600 367.650 ;
        RECT 662.400 365.400 663.600 367.650 ;
        RECT 619.950 346.950 622.050 349.050 ;
        RECT 616.950 331.950 619.050 334.050 ;
        RECT 620.400 319.050 621.450 346.950 ;
        RECT 635.400 343.050 636.450 365.400 ;
        RECT 652.950 358.950 655.050 361.050 ;
        RECT 653.400 355.050 654.450 358.950 ;
        RECT 652.950 352.950 655.050 355.050 ;
        RECT 656.400 346.050 657.450 365.400 ;
        RECT 658.950 358.950 661.050 361.050 ;
        RECT 655.950 343.950 658.050 346.050 ;
        RECT 625.950 339.000 628.050 343.050 ;
        RECT 634.950 340.950 637.050 343.050 ;
        RECT 626.400 337.350 627.600 339.000 ;
        RECT 637.950 337.950 640.050 340.050 ;
        RECT 646.950 339.000 649.050 343.050 ;
        RECT 625.950 334.950 628.050 337.050 ;
        RECT 628.950 334.950 631.050 337.050 ;
        RECT 629.400 333.900 630.600 334.650 ;
        RECT 628.950 331.800 631.050 333.900 ;
        RECT 629.400 328.050 630.450 331.800 ;
        RECT 634.950 328.950 637.050 331.050 ;
        RECT 628.950 325.950 631.050 328.050 ;
        RECT 619.950 316.950 622.050 319.050 ;
        RECT 616.950 313.950 619.050 316.050 ;
        RECT 617.400 298.050 618.450 313.950 ;
        RECT 635.400 310.050 636.450 328.950 ;
        RECT 628.950 307.950 631.050 310.050 ;
        RECT 634.950 307.950 637.050 310.050 ;
        RECT 616.950 295.950 619.050 298.050 ;
        RECT 614.400 292.350 615.600 294.600 ;
        RECT 619.950 293.100 622.050 295.200 ;
        RECT 625.950 294.000 628.050 298.050 ;
        RECT 629.400 295.050 630.450 307.950 ;
        RECT 631.950 295.950 634.050 301.050 ;
        RECT 620.400 292.350 621.600 293.100 ;
        RECT 626.400 292.350 627.600 294.000 ;
        RECT 628.950 292.950 631.050 295.050 ;
        RECT 635.400 294.450 636.450 307.950 ;
        RECT 638.400 295.050 639.450 337.950 ;
        RECT 647.400 337.350 648.600 339.000 ;
        RECT 652.950 338.100 655.050 340.200 ;
        RECT 653.400 337.350 654.600 338.100 ;
        RECT 643.950 334.950 646.050 337.050 ;
        RECT 646.950 334.950 649.050 337.050 ;
        RECT 649.950 334.950 652.050 337.050 ;
        RECT 652.950 334.950 655.050 337.050 ;
        RECT 644.400 333.900 645.600 334.650 ;
        RECT 643.950 331.800 646.050 333.900 ;
        RECT 650.400 333.000 651.600 334.650 ;
        RECT 649.950 328.950 652.050 333.000 ;
        RECT 643.950 325.950 646.050 328.050 ;
        RECT 632.400 293.400 636.450 294.450 ;
        RECT 613.950 289.950 616.050 292.050 ;
        RECT 616.950 289.950 619.050 292.050 ;
        RECT 619.950 289.950 622.050 292.050 ;
        RECT 622.950 289.950 625.050 292.050 ;
        RECT 625.950 289.950 628.050 292.050 ;
        RECT 617.400 288.000 618.600 289.650 ;
        RECT 616.950 283.950 619.050 288.000 ;
        RECT 623.400 287.400 624.600 289.650 ;
        RECT 623.400 283.050 624.450 287.400 ;
        RECT 622.950 280.950 625.050 283.050 ;
        RECT 613.950 277.950 616.050 280.050 ;
        RECT 595.950 262.950 598.050 265.050 ;
        RECT 604.950 262.950 607.050 265.050 ;
        RECT 578.400 259.350 579.600 261.600 ;
        RECT 584.400 259.350 585.600 261.600 ;
        RECT 589.950 259.950 592.050 262.050 ;
        RECT 592.950 259.950 595.050 262.050 ;
        RECT 577.950 256.950 580.050 259.050 ;
        RECT 580.950 256.950 583.050 259.050 ;
        RECT 583.950 256.950 586.050 259.050 ;
        RECT 586.950 256.950 589.050 259.050 ;
        RECT 571.950 253.950 574.050 256.050 ;
        RECT 581.400 255.900 582.600 256.650 ;
        RECT 587.400 255.900 588.600 256.650 ;
        RECT 580.950 253.800 583.050 255.900 ;
        RECT 586.950 253.800 589.050 255.900 ;
        RECT 593.400 253.050 594.450 259.950 ;
        RECT 571.950 250.800 574.050 252.900 ;
        RECT 568.950 247.950 571.050 250.050 ;
        RECT 572.400 241.050 573.450 250.800 ;
        RECT 586.950 250.650 589.050 252.750 ;
        RECT 592.950 250.950 595.050 253.050 ;
        RECT 580.800 241.950 582.900 244.050 ;
        RECT 583.950 241.950 586.050 244.050 ;
        RECT 565.950 238.950 571.050 241.050 ;
        RECT 571.950 238.950 574.050 241.050 ;
        RECT 553.950 235.950 556.050 238.050 ;
        RECT 568.950 235.800 571.050 237.900 ;
        RECT 574.950 235.950 577.050 241.050 ;
        RECT 556.950 229.950 559.050 232.050 ;
        RECT 544.950 223.950 547.050 226.050 ;
        RECT 553.950 223.950 556.050 226.050 ;
        RECT 526.950 217.950 529.050 220.050 ;
        RECT 541.950 218.100 544.050 220.200 ;
        RECT 518.400 214.350 519.600 215.100 ;
        RECT 523.950 214.950 526.050 217.050 ;
        RECT 517.950 211.950 520.050 214.050 ;
        RECT 520.950 211.950 523.050 214.050 ;
        RECT 511.950 208.950 514.050 211.050 ;
        RECT 521.400 210.000 522.600 211.650 ;
        RECT 520.950 205.950 523.050 210.000 ;
        RECT 527.400 202.050 528.450 217.950 ;
        RECT 529.950 214.950 532.050 217.050 ;
        RECT 541.950 214.950 544.050 217.050 ;
        RECT 547.950 215.100 550.050 220.050 ;
        RECT 530.400 208.050 531.450 214.950 ;
        RECT 542.400 214.350 543.600 214.950 ;
        RECT 548.400 214.350 549.600 215.100 ;
        RECT 554.400 214.050 555.450 223.950 ;
        RECT 557.400 223.050 558.450 229.950 ;
        RECT 569.400 226.050 570.450 235.800 ;
        RECT 568.950 223.950 571.050 226.050 ;
        RECT 556.950 220.950 559.050 223.050 ;
        RECT 565.950 220.950 568.050 223.050 ;
        RECT 559.950 214.950 562.050 217.050 ;
        RECT 566.400 216.600 567.450 220.950 ;
        RECT 538.950 211.950 541.050 214.050 ;
        RECT 541.950 211.950 544.050 214.050 ;
        RECT 544.950 211.950 547.050 214.050 ;
        RECT 547.950 211.950 550.050 214.050 ;
        RECT 553.950 211.950 556.050 214.050 ;
        RECT 539.400 209.400 540.600 211.650 ;
        RECT 545.400 209.400 546.600 211.650 ;
        RECT 529.950 205.950 532.050 208.050 ;
        RECT 517.950 199.950 520.050 202.050 ;
        RECT 526.950 199.950 529.050 202.050 ;
        RECT 518.400 183.600 519.450 199.950 ;
        RECT 518.400 181.350 519.600 183.600 ;
        RECT 523.950 182.100 526.050 184.200 ;
        RECT 524.400 181.350 525.600 182.100 ;
        RECT 514.950 178.950 517.050 181.050 ;
        RECT 517.950 178.950 520.050 181.050 ;
        RECT 520.950 178.950 523.050 181.050 ;
        RECT 523.950 178.950 526.050 181.050 ;
        RECT 515.400 177.900 516.600 178.650 ;
        RECT 514.950 175.800 517.050 177.900 ;
        RECT 521.400 177.000 522.600 178.650 ;
        RECT 530.400 177.900 531.450 205.950 ;
        RECT 539.400 190.050 540.450 209.400 ;
        RECT 532.950 187.950 535.050 190.050 ;
        RECT 538.950 187.950 541.050 190.050 ;
        RECT 520.950 172.950 523.050 177.000 ;
        RECT 529.950 175.800 532.050 177.900 ;
        RECT 508.950 157.950 511.050 160.050 ;
        RECT 505.950 151.950 508.050 154.050 ;
        RECT 511.950 151.950 514.050 154.050 ;
        RECT 499.950 148.950 502.050 151.050 ;
        RECT 503.250 145.500 505.350 146.400 ;
        RECT 490.950 142.950 493.050 145.050 ;
        RECT 496.950 142.950 499.050 145.050 ;
        RECT 501.150 144.300 505.350 145.500 ;
        RECT 460.950 133.950 463.050 136.050 ;
        RECT 463.950 133.950 466.050 136.050 ;
        RECT 466.950 133.950 469.050 136.050 ;
        RECT 469.950 133.950 472.050 136.050 ;
        RECT 461.400 131.400 462.600 133.650 ;
        RECT 467.400 132.000 468.600 133.650 ;
        RECT 476.400 133.050 477.450 137.100 ;
        RECT 461.400 127.050 462.450 131.400 ;
        RECT 466.950 127.950 469.050 132.000 ;
        RECT 475.950 130.950 478.050 133.050 ;
        RECT 460.950 124.950 463.050 127.050 ;
        RECT 469.950 115.950 472.050 118.050 ;
        RECT 460.950 109.950 463.050 112.050 ;
        RECT 470.400 111.450 471.450 115.950 ;
        RECT 479.400 112.050 480.450 137.100 ;
        RECT 485.400 136.350 486.600 138.600 ;
        RECT 490.950 137.100 493.050 139.200 ;
        RECT 497.400 138.600 498.450 142.950 ;
        RECT 491.400 136.350 492.600 137.100 ;
        RECT 497.400 136.350 498.600 138.600 ;
        RECT 484.950 133.950 487.050 136.050 ;
        RECT 487.950 133.950 490.050 136.050 ;
        RECT 490.950 133.950 493.050 136.050 ;
        RECT 496.950 133.950 499.050 136.050 ;
        RECT 488.400 132.900 489.600 133.650 ;
        RECT 487.950 130.800 490.050 132.900 ;
        RECT 501.150 125.700 502.350 144.300 ;
        RECT 505.950 137.100 508.050 139.200 ;
        RECT 506.400 136.350 507.600 137.100 ;
        RECT 506.100 133.950 508.200 136.050 ;
        RECT 512.400 127.050 513.450 151.950 ;
        RECT 518.550 147.300 520.650 149.400 ;
        RECT 518.550 140.700 519.750 147.300 ;
        RECT 514.950 137.100 517.050 139.200 ;
        RECT 518.550 138.600 520.650 140.700 ;
        RECT 515.400 130.050 516.450 137.100 ;
        RECT 514.950 127.950 517.050 130.050 ;
        RECT 500.850 123.600 502.950 125.700 ;
        RECT 511.950 124.950 514.050 127.050 ;
        RECT 518.550 125.700 519.750 138.600 ;
        RECT 523.950 133.950 526.050 136.050 ;
        RECT 524.400 131.400 525.600 133.650 ;
        RECT 524.400 127.050 525.450 131.400 ;
        RECT 530.400 130.050 531.450 175.800 ;
        RECT 533.400 175.050 534.450 187.950 ;
        RECT 539.400 183.600 540.450 187.950 ;
        RECT 539.400 181.350 540.600 183.600 ;
        RECT 545.400 183.450 546.450 209.400 ;
        RECT 547.950 202.950 550.050 205.050 ;
        RECT 548.400 196.050 549.450 202.950 ;
        RECT 550.950 196.950 553.050 199.050 ;
        RECT 547.950 193.950 550.050 196.050 ;
        RECT 545.400 182.400 549.450 183.450 ;
        RECT 538.950 178.950 541.050 181.050 ;
        RECT 541.950 178.950 544.050 181.050 ;
        RECT 542.400 176.400 543.600 178.650 ;
        RECT 532.950 172.950 535.050 175.050 ;
        RECT 542.400 166.050 543.450 176.400 ;
        RECT 541.950 163.950 544.050 166.050 ;
        RECT 544.950 160.950 547.050 163.050 ;
        RECT 545.400 141.450 546.450 160.950 ;
        RECT 548.400 145.050 549.450 182.400 ;
        RECT 551.400 160.050 552.450 196.950 ;
        RECT 560.400 190.050 561.450 214.950 ;
        RECT 566.400 214.350 567.600 216.600 ;
        RECT 571.950 216.000 574.050 220.050 ;
        RECT 572.400 214.350 573.600 216.000 ;
        RECT 581.400 214.050 582.450 241.950 ;
        RECT 584.400 226.050 585.450 241.950 ;
        RECT 583.950 223.950 586.050 226.050 ;
        RECT 587.400 220.050 588.450 250.650 ;
        RECT 592.950 247.800 595.050 249.900 ;
        RECT 589.950 229.950 592.050 232.050 ;
        RECT 586.950 217.950 589.050 220.050 ;
        RECT 590.400 216.600 591.450 229.950 ;
        RECT 593.400 223.050 594.450 247.800 ;
        RECT 596.400 234.450 597.450 262.950 ;
        RECT 601.950 260.100 604.050 262.200 ;
        RECT 614.400 262.050 615.450 277.950 ;
        RECT 616.950 274.950 619.050 277.050 ;
        RECT 602.400 259.350 603.600 260.100 ;
        RECT 607.950 259.950 610.050 262.050 ;
        RECT 613.950 259.950 616.050 262.050 ;
        RECT 608.400 259.350 609.600 259.950 ;
        RECT 601.950 256.950 604.050 259.050 ;
        RECT 604.950 256.950 607.050 259.050 ;
        RECT 607.950 256.950 610.050 259.050 ;
        RECT 610.950 256.950 613.050 259.050 ;
        RECT 605.400 255.900 606.600 256.650 ;
        RECT 604.950 253.800 607.050 255.900 ;
        RECT 611.400 255.000 612.600 256.650 ;
        RECT 617.400 256.050 618.450 274.950 ;
        RECT 622.950 268.950 625.050 271.050 ;
        RECT 619.950 256.950 622.050 259.050 ;
        RECT 604.950 250.650 607.050 252.750 ;
        RECT 610.950 250.950 613.050 255.000 ;
        RECT 616.950 253.950 619.050 256.050 ;
        RECT 620.400 252.450 621.450 256.950 ;
        RECT 617.400 251.400 621.450 252.450 ;
        RECT 605.400 244.050 606.450 250.650 ;
        RECT 607.950 247.950 610.050 250.050 ;
        RECT 604.950 241.950 607.050 244.050 ;
        RECT 608.400 241.050 609.450 247.950 ;
        RECT 610.950 241.950 613.050 244.050 ;
        RECT 607.950 238.950 610.050 241.050 ;
        RECT 596.400 233.400 600.450 234.450 ;
        RECT 595.950 229.950 598.050 232.050 ;
        RECT 596.400 226.050 597.450 229.950 ;
        RECT 599.400 226.050 600.450 233.400 ;
        RECT 611.400 226.050 612.450 241.950 ;
        RECT 595.950 223.950 598.050 226.050 ;
        RECT 598.950 225.450 601.050 226.050 ;
        RECT 598.950 224.400 603.450 225.450 ;
        RECT 598.950 223.950 601.050 224.400 ;
        RECT 592.950 220.950 595.050 223.050 ;
        RECT 590.400 214.350 591.600 216.600 ;
        RECT 565.950 211.950 568.050 214.050 ;
        RECT 568.950 211.950 571.050 214.050 ;
        RECT 571.950 211.950 574.050 214.050 ;
        RECT 574.950 211.950 577.050 214.050 ;
        RECT 580.950 211.950 583.050 214.050 ;
        RECT 589.950 211.950 592.050 214.050 ;
        RECT 592.950 211.950 595.050 214.050 ;
        RECT 595.950 211.950 598.050 214.050 ;
        RECT 569.400 210.900 570.600 211.650 ;
        RECT 568.950 208.800 571.050 210.900 ;
        RECT 575.400 209.400 576.600 211.650 ;
        RECT 593.400 209.400 594.600 211.650 ;
        RECT 568.950 202.950 571.050 205.050 ;
        RECT 569.400 196.050 570.450 202.950 ;
        RECT 575.400 196.050 576.450 209.400 ;
        RECT 568.950 193.950 571.050 196.050 ;
        RECT 574.950 193.950 577.050 196.050 ;
        RECT 559.950 187.950 562.050 190.050 ;
        RECT 586.950 187.950 589.050 190.050 ;
        RECT 556.950 182.100 559.050 184.200 ;
        RECT 562.950 183.000 565.050 187.050 ;
        RECT 557.400 181.350 558.600 182.100 ;
        RECT 563.400 181.350 564.600 183.000 ;
        RECT 574.950 181.950 577.050 184.050 ;
        RECT 580.950 182.100 583.050 184.200 ;
        RECT 587.400 183.600 588.450 187.950 ;
        RECT 556.950 178.950 559.050 181.050 ;
        RECT 559.950 178.950 562.050 181.050 ;
        RECT 562.950 178.950 565.050 181.050 ;
        RECT 565.950 178.950 568.050 181.050 ;
        RECT 560.400 176.400 561.600 178.650 ;
        RECT 566.400 176.400 567.600 178.650 ;
        RECT 560.400 160.050 561.450 176.400 ;
        RECT 550.950 157.950 553.050 160.050 ;
        RECT 559.950 157.950 562.050 160.050 ;
        RECT 562.950 148.950 565.050 151.050 ;
        RECT 547.950 142.950 550.050 145.050 ;
        RECT 559.950 142.950 562.050 145.050 ;
        RECT 545.400 140.400 549.450 141.450 ;
        RECT 548.400 138.600 549.450 140.400 ;
        RECT 548.400 136.350 549.600 138.600 ;
        RECT 541.950 133.950 544.050 136.050 ;
        RECT 544.950 133.950 547.050 136.050 ;
        RECT 547.950 133.950 550.050 136.050 ;
        RECT 545.400 131.400 546.600 133.650 ;
        RECT 529.950 127.950 532.050 130.050 ;
        RECT 518.550 123.600 520.650 125.700 ;
        RECT 523.950 124.950 526.050 127.050 ;
        RECT 545.400 121.050 546.450 131.400 ;
        RECT 544.950 118.950 547.050 121.050 ;
        RECT 560.400 118.050 561.450 142.950 ;
        RECT 563.400 138.450 564.450 148.950 ;
        RECT 566.400 148.050 567.450 176.400 ;
        RECT 571.950 163.950 574.050 166.050 ;
        RECT 572.400 154.050 573.450 163.950 ;
        RECT 571.950 151.950 574.050 154.050 ;
        RECT 565.950 145.950 568.050 148.050 ;
        RECT 572.400 138.600 573.450 151.950 ;
        RECT 575.400 145.050 576.450 181.950 ;
        RECT 581.400 181.350 582.600 182.100 ;
        RECT 587.400 181.350 588.600 183.600 ;
        RECT 593.400 183.450 594.450 209.400 ;
        RECT 598.950 196.950 601.050 199.050 ;
        RECT 593.400 182.400 597.450 183.450 ;
        RECT 580.950 178.950 583.050 181.050 ;
        RECT 583.950 178.950 586.050 181.050 ;
        RECT 586.950 178.950 589.050 181.050 ;
        RECT 589.950 178.950 592.050 181.050 ;
        RECT 584.400 177.000 585.600 178.650 ;
        RECT 590.400 177.900 591.600 178.650 ;
        RECT 596.400 177.900 597.450 182.400 ;
        RECT 583.950 172.950 586.050 177.000 ;
        RECT 589.950 175.800 592.050 177.900 ;
        RECT 595.950 175.800 598.050 177.900 ;
        RECT 596.400 169.050 597.450 175.800 ;
        RECT 589.950 166.950 595.050 169.050 ;
        RECT 595.950 166.950 598.050 169.050 ;
        RECT 599.400 163.050 600.450 196.950 ;
        RECT 602.400 175.050 603.450 224.400 ;
        RECT 610.950 223.950 613.050 226.050 ;
        RECT 617.400 217.200 618.450 251.400 ;
        RECT 619.950 229.950 622.050 232.050 ;
        RECT 620.400 223.050 621.450 229.950 ;
        RECT 619.950 220.950 622.050 223.050 ;
        RECT 604.950 215.100 607.050 217.200 ;
        RECT 616.950 215.100 619.050 217.200 ;
        RECT 605.400 199.050 606.450 215.100 ;
        RECT 617.400 214.350 618.600 215.100 ;
        RECT 610.950 211.950 613.050 214.050 ;
        RECT 613.950 211.950 616.050 214.050 ;
        RECT 616.950 211.950 619.050 214.050 ;
        RECT 607.950 208.950 610.050 211.050 ;
        RECT 614.400 210.000 615.600 211.650 ;
        RECT 604.950 196.950 607.050 199.050 ;
        RECT 604.950 181.950 607.050 187.050 ;
        RECT 608.400 183.600 609.450 208.950 ;
        RECT 613.950 205.950 616.050 210.000 ;
        RECT 619.950 193.950 622.050 196.050 ;
        RECT 608.400 181.350 609.600 183.600 ;
        RECT 613.950 182.100 616.050 184.200 ;
        RECT 620.400 184.050 621.450 193.950 ;
        RECT 614.400 181.350 615.600 182.100 ;
        RECT 619.950 181.950 622.050 184.050 ;
        RECT 607.950 178.950 610.050 181.050 ;
        RECT 610.950 178.950 613.050 181.050 ;
        RECT 613.950 178.950 616.050 181.050 ;
        RECT 616.950 178.950 619.050 181.050 ;
        RECT 611.400 177.000 612.600 178.650 ;
        RECT 601.950 172.950 604.050 175.050 ;
        RECT 610.950 172.950 613.050 177.000 ;
        RECT 617.400 176.400 618.600 178.650 ;
        RECT 601.950 163.950 604.050 169.050 ;
        RECT 598.950 160.950 601.050 163.050 ;
        RECT 617.400 154.050 618.450 176.400 ;
        RECT 619.950 175.950 622.050 178.050 ;
        RECT 589.950 151.950 592.050 154.050 ;
        RECT 616.950 151.950 619.050 154.050 ;
        RECT 574.950 142.950 577.050 145.050 ;
        RECT 580.950 142.950 583.050 145.050 ;
        RECT 566.400 138.450 567.600 138.600 ;
        RECT 563.400 137.400 567.600 138.450 ;
        RECT 566.400 136.350 567.600 137.400 ;
        RECT 572.400 136.350 573.600 138.600 ;
        RECT 565.950 133.950 568.050 136.050 ;
        RECT 568.950 133.950 571.050 136.050 ;
        RECT 571.950 133.950 574.050 136.050 ;
        RECT 574.950 133.950 577.050 136.050 ;
        RECT 569.400 132.900 570.600 133.650 ;
        RECT 568.950 127.950 571.050 132.900 ;
        RECT 575.400 131.400 576.600 133.650 ;
        RECT 562.950 121.950 565.050 124.050 ;
        RECT 559.950 115.950 562.050 118.050 ;
        RECT 556.950 112.950 559.050 115.050 ;
        RECT 461.400 105.450 462.450 109.950 ;
        RECT 466.800 108.300 468.900 110.400 ;
        RECT 470.400 109.200 471.600 111.450 ;
        RECT 478.950 109.950 481.050 112.050 ;
        RECT 526.950 109.950 529.050 112.050 ;
        RECT 464.400 105.450 465.600 105.600 ;
        RECT 461.400 104.400 465.600 105.450 ;
        RECT 464.400 103.350 465.600 104.400 ;
        RECT 464.100 100.950 466.200 103.050 ;
        RECT 467.100 102.900 468.000 108.300 ;
        RECT 470.100 106.800 472.200 108.900 ;
        RECT 474.000 105.900 476.100 107.700 ;
        RECT 468.900 104.700 477.600 105.900 ;
        RECT 468.900 103.800 471.000 104.700 ;
        RECT 467.100 101.700 474.000 102.900 ;
        RECT 467.100 94.500 468.300 101.700 ;
        RECT 470.100 97.950 472.200 100.050 ;
        RECT 473.100 99.300 474.000 101.700 ;
        RECT 470.400 95.400 471.600 97.650 ;
        RECT 473.100 97.200 475.200 99.300 ;
        RECT 476.700 95.700 477.600 104.700 ;
        RECT 487.950 104.100 490.050 106.200 ;
        RECT 493.950 104.100 496.050 106.200 ;
        RECT 505.950 104.100 508.050 106.200 ;
        RECT 511.950 104.100 514.050 106.200 ;
        RECT 517.950 104.100 520.050 106.200 ;
        RECT 523.950 104.100 526.050 106.200 ;
        RECT 478.800 100.950 480.900 103.050 ;
        RECT 479.400 99.450 480.600 100.650 ;
        RECT 481.950 99.450 484.050 103.050 ;
        RECT 479.400 99.000 484.050 99.450 ;
        RECT 479.400 98.400 483.450 99.000 ;
        RECT 466.800 92.400 468.900 94.500 ;
        RECT 472.950 91.950 475.050 94.050 ;
        RECT 476.400 93.600 478.500 95.700 ;
        RECT 488.400 94.050 489.450 104.100 ;
        RECT 494.400 103.350 495.600 104.100 ;
        RECT 493.950 100.950 496.050 103.050 ;
        RECT 496.950 100.950 499.050 103.050 ;
        RECT 502.950 100.950 505.050 103.050 ;
        RECT 497.400 99.900 498.600 100.650 ;
        RECT 496.950 97.800 499.050 99.900 ;
        RECT 503.400 97.050 504.450 100.950 ;
        RECT 506.400 100.050 507.450 104.100 ;
        RECT 512.400 103.350 513.600 104.100 ;
        RECT 518.400 103.350 519.600 104.100 ;
        RECT 511.950 100.950 514.050 103.050 ;
        RECT 514.950 100.950 517.050 103.050 ;
        RECT 517.950 100.950 520.050 103.050 ;
        RECT 505.950 97.950 508.050 100.050 ;
        RECT 515.400 99.000 516.600 100.650 ;
        RECT 502.950 94.950 505.050 97.050 ;
        RECT 514.950 94.950 517.050 99.000 ;
        RECT 487.950 91.950 490.050 94.050 ;
        RECT 466.950 85.950 469.050 88.050 ;
        RECT 430.950 79.950 433.050 82.050 ;
        RECT 454.950 79.950 457.050 82.050 ;
        RECT 431.400 61.050 432.450 79.950 ;
        RECT 467.400 79.050 468.450 85.950 ;
        RECT 466.950 76.950 469.050 79.050 ;
        RECT 454.950 73.950 457.050 76.050 ;
        RECT 436.950 67.950 439.050 70.050 ;
        RECT 430.950 58.950 433.050 61.050 ;
        RECT 437.400 60.600 438.450 67.950 ;
        RECT 437.400 58.350 438.600 60.600 ;
        RECT 442.950 59.100 445.050 61.200 ;
        RECT 448.950 59.100 451.050 61.200 ;
        RECT 455.400 61.050 456.450 73.950 ;
        RECT 460.950 67.950 463.050 70.050 ;
        RECT 461.400 64.050 462.450 67.950 ;
        RECT 443.400 58.350 444.600 59.100 ;
        RECT 433.950 55.950 436.050 58.050 ;
        RECT 436.950 55.950 439.050 58.050 ;
        RECT 439.950 55.950 442.050 58.050 ;
        RECT 442.950 55.950 445.050 58.050 ;
        RECT 434.400 54.900 435.600 55.650 ;
        RECT 440.400 54.900 441.600 55.650 ;
        RECT 428.400 53.400 432.450 54.450 ;
        RECT 431.400 49.050 432.450 53.400 ;
        RECT 433.950 52.800 436.050 54.900 ;
        RECT 439.950 52.800 442.050 54.900 ;
        RECT 430.950 46.950 433.050 49.050 ;
        RECT 436.950 46.950 439.050 49.050 ;
        RECT 424.950 43.950 427.050 46.050 ;
        RECT 419.400 26.400 423.450 27.450 ;
        RECT 437.400 27.600 438.450 46.950 ;
        RECT 449.400 43.050 450.450 59.100 ;
        RECT 454.950 58.950 457.050 61.050 ;
        RECT 460.950 60.000 463.050 64.050 ;
        RECT 467.400 60.600 468.450 76.950 ;
        RECT 461.400 58.350 462.600 60.000 ;
        RECT 467.400 58.350 468.600 60.600 ;
        RECT 457.950 55.950 460.050 58.050 ;
        RECT 460.950 55.950 463.050 58.050 ;
        RECT 463.950 55.950 466.050 58.050 ;
        RECT 466.950 55.950 469.050 58.050 ;
        RECT 458.400 53.400 459.600 55.650 ;
        RECT 464.400 54.900 465.600 55.650 ;
        RECT 458.400 49.050 459.450 53.400 ;
        RECT 463.950 49.950 466.050 54.900 ;
        RECT 473.400 52.050 474.450 91.950 ;
        RECT 488.400 73.050 489.450 91.950 ;
        RECT 524.400 73.050 525.450 104.100 ;
        RECT 527.400 99.900 528.450 109.950 ;
        RECT 557.400 109.050 558.450 112.950 ;
        RECT 556.950 106.950 559.050 109.050 ;
        RECT 532.950 104.100 535.050 106.200 ;
        RECT 538.950 104.100 541.050 106.200 ;
        RECT 533.400 103.350 534.600 104.100 ;
        RECT 539.400 103.350 540.600 104.100 ;
        RECT 550.950 103.950 553.050 106.050 ;
        RECT 557.400 105.600 558.450 106.950 ;
        RECT 563.400 106.050 564.450 121.950 ;
        RECT 565.950 115.950 568.050 118.050 ;
        RECT 571.950 115.950 574.050 118.050 ;
        RECT 532.950 100.950 535.050 103.050 ;
        RECT 535.950 100.950 538.050 103.050 ;
        RECT 538.950 100.950 541.050 103.050 ;
        RECT 541.950 100.950 544.050 103.050 ;
        RECT 536.400 99.900 537.600 100.650 ;
        RECT 526.950 97.800 529.050 99.900 ;
        RECT 535.950 97.800 538.050 99.900 ;
        RECT 542.400 98.400 543.600 100.650 ;
        RECT 542.400 94.050 543.450 98.400 ;
        RECT 551.400 94.050 552.450 103.950 ;
        RECT 557.400 103.350 558.600 105.600 ;
        RECT 562.950 103.950 565.050 106.050 ;
        RECT 556.950 100.950 559.050 103.050 ;
        RECT 559.950 100.950 562.050 103.050 ;
        RECT 560.400 99.900 561.600 100.650 ;
        RECT 559.950 97.800 562.050 99.900 ;
        RECT 566.400 97.050 567.450 115.950 ;
        RECT 572.400 112.050 573.450 115.950 ;
        RECT 571.950 109.950 574.050 112.050 ;
        RECT 575.400 109.050 576.450 131.400 ;
        RECT 581.400 118.050 582.450 142.950 ;
        RECT 590.400 138.600 591.450 151.950 ;
        RECT 595.950 148.950 598.050 151.050 ;
        RECT 596.400 138.600 597.450 148.950 ;
        RECT 620.400 142.050 621.450 175.950 ;
        RECT 623.400 172.050 624.450 268.950 ;
        RECT 632.400 261.600 633.450 293.400 ;
        RECT 637.950 292.950 640.050 295.050 ;
        RECT 644.400 294.600 645.450 325.950 ;
        RECT 659.400 322.050 660.450 358.950 ;
        RECT 662.400 355.050 663.450 365.400 ;
        RECT 661.950 352.950 664.050 355.050 ;
        RECT 668.400 340.200 669.450 403.800 ;
        RECT 671.400 388.050 672.450 409.950 ;
        RECT 674.400 406.050 675.450 433.950 ;
        RECT 677.400 409.050 678.450 439.950 ;
        RECT 695.400 430.050 696.450 484.950 ;
        RECT 704.400 481.050 705.450 488.400 ;
        RECT 703.950 478.950 706.050 481.050 ;
        RECT 700.950 466.950 703.050 469.050 ;
        RECT 697.950 463.950 700.050 466.050 ;
        RECT 698.400 454.050 699.450 463.950 ;
        RECT 697.950 451.950 700.050 454.050 ;
        RECT 701.400 450.600 702.450 466.950 ;
        RECT 701.400 448.350 702.600 450.600 ;
        RECT 706.950 449.100 709.050 451.200 ;
        RECT 713.400 451.050 714.450 490.950 ;
        RECT 719.400 489.450 720.450 520.950 ;
        RECT 725.400 505.050 726.450 521.400 ;
        RECT 730.950 517.950 733.050 522.000 ;
        RECT 724.950 502.950 727.050 505.050 ;
        RECT 722.100 490.950 724.200 493.050 ;
        RECT 725.400 490.950 727.500 493.050 ;
        RECT 730.800 490.950 732.900 493.050 ;
        RECT 722.400 489.450 723.600 490.650 ;
        RECT 719.400 488.400 723.600 489.450 ;
        RECT 731.400 489.000 732.600 490.650 ;
        RECT 722.400 465.450 723.450 488.400 ;
        RECT 730.950 484.950 733.050 489.000 ;
        RECT 730.950 478.950 736.050 481.050 ;
        RECT 722.400 464.400 726.450 465.450 ;
        RECT 721.950 460.950 724.050 463.050 ;
        RECT 722.400 451.050 723.450 460.950 ;
        RECT 707.400 448.350 708.600 449.100 ;
        RECT 712.950 448.950 715.050 451.050 ;
        RECT 721.950 448.950 724.050 451.050 ;
        RECT 725.400 450.600 726.450 464.400 ;
        RECT 727.950 460.950 730.050 463.050 ;
        RECT 728.400 454.050 729.450 460.950 ;
        RECT 737.400 454.050 738.450 541.950 ;
        RECT 739.950 529.950 742.050 532.050 ;
        RECT 740.400 522.900 741.450 529.950 ;
        RECT 749.400 528.600 750.450 544.950 ;
        RECT 754.950 538.950 757.050 541.050 ;
        RECT 749.400 526.350 750.600 528.600 ;
        RECT 745.950 523.950 748.050 526.050 ;
        RECT 748.950 523.950 751.050 526.050 ;
        RECT 746.400 522.900 747.600 523.650 ;
        RECT 739.950 520.800 742.050 522.900 ;
        RECT 745.950 520.800 748.050 522.900 ;
        RECT 755.400 517.050 756.450 538.950 ;
        RECT 758.400 538.050 759.450 565.950 ;
        RECT 761.400 559.050 762.450 566.400 ;
        RECT 766.950 565.800 769.050 567.900 ;
        RECT 778.950 565.800 781.050 567.900 ;
        RECT 782.400 567.450 783.450 571.950 ;
        RECT 791.400 571.350 792.600 573.600 ;
        RECT 785.100 568.950 787.200 571.050 ;
        RECT 790.500 568.950 792.600 571.050 ;
        RECT 793.800 568.950 795.900 571.050 ;
        RECT 785.400 567.450 786.600 568.650 ;
        RECT 782.400 566.400 786.600 567.450 ;
        RECT 794.400 567.450 795.600 568.650 ;
        RECT 797.400 567.450 798.450 599.400 ;
        RECT 800.400 599.400 801.600 601.650 ;
        RECT 800.400 595.050 801.450 599.400 ;
        RECT 809.400 598.050 810.450 637.800 ;
        RECT 811.950 604.950 814.050 607.050 ;
        RECT 812.400 600.900 813.450 604.950 ;
        RECT 811.950 598.800 814.050 600.900 ;
        RECT 815.400 600.450 816.450 643.950 ;
        RECT 818.400 637.050 819.450 673.950 ;
        RECT 827.400 672.450 828.450 676.950 ;
        RECT 829.950 676.800 832.050 678.900 ;
        RECT 835.950 675.450 838.050 678.900 ;
        RECT 833.400 675.000 838.050 675.450 ;
        RECT 833.400 674.400 837.450 675.000 ;
        RECT 833.400 672.450 834.450 674.400 ;
        RECT 824.400 671.400 828.450 672.450 ;
        RECT 830.400 671.400 834.450 672.450 ;
        RECT 820.950 661.950 823.050 664.050 ;
        RECT 821.400 645.900 822.450 661.950 ;
        RECT 824.400 652.050 825.450 671.400 ;
        RECT 830.400 670.050 831.450 671.400 ;
        RECT 835.950 670.950 838.050 673.050 ;
        RECT 826.950 668.400 831.450 670.050 ;
        RECT 826.950 667.950 831.000 668.400 ;
        RECT 829.950 664.950 832.050 667.050 ;
        RECT 823.950 649.950 826.050 652.050 ;
        RECT 830.400 651.600 831.450 664.950 ;
        RECT 836.400 651.600 837.450 670.950 ;
        RECT 839.400 658.050 840.450 694.950 ;
        RECT 845.400 684.450 846.450 718.950 ;
        RECT 863.400 715.050 864.450 719.400 ;
        RECT 878.400 718.050 879.450 793.950 ;
        RECT 884.400 763.050 885.450 799.800 ;
        RECT 896.400 796.050 897.450 823.950 ;
        RECT 902.400 820.050 903.450 832.950 ;
        RECT 905.400 826.050 906.450 868.950 ;
        RECT 911.400 841.050 912.450 884.100 ;
        RECT 914.400 871.050 915.450 884.400 ;
        RECT 923.400 883.350 924.600 885.600 ;
        RECT 928.950 884.100 931.050 886.200 ;
        RECT 935.400 886.050 936.450 910.950 ;
        RECT 929.400 883.350 930.600 884.100 ;
        RECT 934.950 883.950 937.050 886.050 ;
        RECT 919.950 880.950 922.050 883.050 ;
        RECT 922.950 880.950 925.050 883.050 ;
        RECT 925.950 880.950 928.050 883.050 ;
        RECT 928.950 880.950 931.050 883.050 ;
        RECT 931.950 880.950 934.050 883.050 ;
        RECT 920.400 878.400 921.600 880.650 ;
        RECT 926.400 878.400 927.600 880.650 ;
        RECT 932.400 879.900 933.600 880.650 ;
        RECT 920.400 874.050 921.450 878.400 ;
        RECT 919.950 871.950 922.050 874.050 ;
        RECT 913.950 868.950 916.050 871.050 ;
        RECT 920.400 856.050 921.450 871.950 ;
        RECT 919.950 853.950 922.050 856.050 ;
        RECT 916.950 844.950 919.050 847.050 ;
        RECT 917.400 841.200 918.450 844.950 ;
        RECT 910.950 838.950 913.050 841.050 ;
        RECT 916.950 839.100 919.050 841.200 ;
        RECT 922.950 839.100 925.050 841.200 ;
        RECT 926.400 841.050 927.450 878.400 ;
        RECT 931.950 877.800 934.050 879.900 ;
        RECT 938.400 874.050 939.450 916.950 ;
        RECT 944.400 898.050 945.450 931.950 ;
        RECT 965.400 928.050 966.450 961.950 ;
        RECT 974.400 961.350 975.600 963.600 ;
        RECT 979.950 962.100 982.050 964.200 ;
        RECT 980.400 961.350 981.600 962.100 ;
        RECT 985.950 961.950 988.050 964.050 ;
        RECT 970.950 958.950 973.050 961.050 ;
        RECT 973.950 958.950 976.050 961.050 ;
        RECT 976.950 958.950 979.050 961.050 ;
        RECT 979.950 958.950 982.050 961.050 ;
        RECT 971.400 957.900 972.600 958.650 ;
        RECT 970.950 955.800 973.050 957.900 ;
        RECT 977.400 956.400 978.600 958.650 ;
        RECT 977.400 954.450 978.450 956.400 ;
        RECT 977.400 953.400 981.450 954.450 ;
        RECT 964.950 925.950 967.050 928.050 ;
        RECT 967.950 922.950 970.050 925.050 ;
        RECT 946.950 918.450 949.050 922.050 ;
        RECT 950.400 918.450 951.600 918.600 ;
        RECT 946.950 918.000 951.600 918.450 ;
        RECT 955.950 918.000 958.050 922.050 ;
        RECT 947.400 917.400 951.600 918.000 ;
        RECT 950.400 916.350 951.600 917.400 ;
        RECT 956.400 916.350 957.600 918.000 ;
        RECT 949.950 913.950 952.050 916.050 ;
        RECT 952.950 913.950 955.050 916.050 ;
        RECT 955.950 913.950 958.050 916.050 ;
        RECT 958.950 913.950 961.050 916.050 ;
        RECT 953.400 912.900 954.600 913.650 ;
        RECT 952.950 910.800 955.050 912.900 ;
        RECT 959.400 911.400 960.600 913.650 ;
        RECT 943.950 895.950 946.050 898.050 ;
        RECT 959.400 889.050 960.450 911.400 ;
        RECT 968.400 910.050 969.450 922.950 ;
        RECT 980.400 922.050 981.450 953.400 ;
        RECT 986.400 925.050 987.450 961.950 ;
        RECT 992.400 943.050 993.450 970.950 ;
        RECT 997.950 962.100 1000.050 964.200 ;
        RECT 1004.400 963.600 1005.450 970.950 ;
        RECT 998.400 961.350 999.600 962.100 ;
        RECT 1004.400 961.350 1005.600 963.600 ;
        RECT 997.950 958.950 1000.050 961.050 ;
        RECT 1000.950 958.950 1003.050 961.050 ;
        RECT 1003.950 958.950 1006.050 961.050 ;
        RECT 1006.950 958.950 1009.050 961.050 ;
        RECT 1001.400 957.900 1002.600 958.650 ;
        RECT 994.950 955.800 997.050 957.900 ;
        RECT 1000.950 955.800 1003.050 957.900 ;
        RECT 1007.400 956.400 1008.600 958.650 ;
        RECT 991.950 940.950 994.050 943.050 ;
        RECT 995.400 934.050 996.450 955.800 ;
        RECT 1007.400 946.050 1008.450 956.400 ;
        RECT 1006.950 943.950 1009.050 946.050 ;
        RECT 1015.950 943.950 1018.050 946.050 ;
        RECT 994.950 931.950 997.050 934.050 ;
        RECT 985.950 922.950 988.050 925.050 ;
        RECT 979.950 919.950 982.050 922.050 ;
        RECT 976.950 917.100 979.050 919.200 ;
        RECT 982.950 918.000 985.050 922.050 ;
        RECT 991.950 919.950 994.050 922.050 ;
        RECT 977.400 916.350 978.600 917.100 ;
        RECT 983.400 916.350 984.600 918.000 ;
        RECT 988.950 916.950 991.050 919.050 ;
        RECT 973.950 913.950 976.050 916.050 ;
        RECT 976.950 913.950 979.050 916.050 ;
        RECT 979.950 913.950 982.050 916.050 ;
        RECT 982.950 913.950 985.050 916.050 ;
        RECT 974.400 911.400 975.600 913.650 ;
        RECT 980.400 912.900 981.600 913.650 ;
        RECT 961.950 907.950 964.050 910.050 ;
        RECT 967.950 907.950 970.050 910.050 ;
        RECT 940.950 883.950 943.050 886.050 ;
        RECT 946.950 884.100 949.050 886.200 ;
        RECT 952.950 885.000 955.050 889.050 ;
        RECT 937.950 871.950 940.050 874.050 ;
        RECT 941.400 844.050 942.450 883.950 ;
        RECT 947.400 883.350 948.600 884.100 ;
        RECT 953.400 883.350 954.600 885.000 ;
        RECT 958.950 883.950 961.050 889.050 ;
        RECT 946.950 880.950 949.050 883.050 ;
        RECT 949.950 880.950 952.050 883.050 ;
        RECT 952.950 880.950 955.050 883.050 ;
        RECT 955.950 880.950 958.050 883.050 ;
        RECT 950.400 879.900 951.600 880.650 ;
        RECT 956.400 879.900 957.600 880.650 ;
        RECT 943.950 877.800 946.050 879.900 ;
        RECT 949.950 877.800 952.050 879.900 ;
        RECT 955.950 877.800 958.050 879.900 ;
        RECT 940.950 841.950 943.050 844.050 ;
        RECT 917.400 838.350 918.600 839.100 ;
        RECT 923.400 838.350 924.600 839.100 ;
        RECT 925.950 838.950 928.050 841.050 ;
        RECT 928.950 839.100 931.050 841.200 ;
        RECT 944.400 841.050 945.450 877.800 ;
        RECT 955.950 847.950 958.050 850.050 ;
        RECT 946.950 844.950 949.050 847.050 ;
        RECT 913.950 835.950 916.050 838.050 ;
        RECT 916.950 835.950 919.050 838.050 ;
        RECT 919.950 835.950 922.050 838.050 ;
        RECT 922.950 835.950 925.050 838.050 ;
        RECT 910.950 832.950 913.050 835.050 ;
        RECT 914.400 833.400 915.600 835.650 ;
        RECT 920.400 833.400 921.600 835.650 ;
        RECT 904.950 823.950 907.050 826.050 ;
        RECT 901.950 817.950 904.050 820.050 ;
        RECT 911.400 808.200 912.450 832.950 ;
        RECT 914.400 817.050 915.450 833.400 ;
        RECT 920.400 823.050 921.450 833.400 ;
        RECT 929.400 826.050 930.450 839.100 ;
        RECT 934.950 838.950 937.050 841.050 ;
        RECT 943.950 838.950 946.050 841.050 ;
        RECT 947.400 840.600 948.450 844.950 ;
        RECT 949.950 841.950 955.050 844.050 ;
        RECT 956.400 840.600 957.450 847.950 ;
        RECT 962.400 846.450 963.450 907.950 ;
        RECT 974.400 907.050 975.450 911.400 ;
        RECT 979.950 910.800 982.050 912.900 ;
        RECT 967.950 904.800 970.050 906.900 ;
        RECT 973.950 904.950 976.050 907.050 ;
        RECT 979.950 904.950 982.050 907.050 ;
        RECT 968.400 886.050 969.450 904.800 ;
        RECT 967.950 883.950 970.050 886.050 ;
        RECT 973.950 884.100 976.050 889.050 ;
        RECT 980.400 885.600 981.450 904.950 ;
        RECT 985.950 901.950 988.050 904.050 ;
        RECT 974.400 883.350 975.600 884.100 ;
        RECT 980.400 883.350 981.600 885.600 ;
        RECT 970.950 880.950 973.050 883.050 ;
        RECT 973.950 880.950 976.050 883.050 ;
        RECT 976.950 880.950 979.050 883.050 ;
        RECT 979.950 880.950 982.050 883.050 ;
        RECT 967.950 877.950 970.050 880.050 ;
        RECT 971.400 878.400 972.600 880.650 ;
        RECT 977.400 878.400 978.600 880.650 ;
        RECT 964.950 868.950 967.050 871.050 ;
        RECT 959.400 845.400 963.450 846.450 ;
        RECT 935.400 832.050 936.450 838.950 ;
        RECT 947.400 838.350 948.600 840.600 ;
        RECT 956.400 838.350 957.600 840.600 ;
        RECT 959.400 838.050 960.450 845.400 ;
        RECT 961.950 841.950 964.050 844.050 ;
        RECT 940.800 835.950 942.900 838.050 ;
        RECT 946.950 835.950 949.050 838.050 ;
        RECT 949.950 835.950 952.050 838.050 ;
        RECT 955.500 835.950 957.600 838.050 ;
        RECT 958.950 835.950 961.050 838.050 ;
        RECT 941.400 834.000 942.600 835.650 ;
        RECT 934.950 829.950 937.050 832.050 ;
        RECT 940.950 829.950 943.050 834.000 ;
        RECT 950.400 833.400 951.600 835.650 ;
        RECT 946.950 829.950 949.050 832.050 ;
        RECT 928.950 823.950 931.050 826.050 ;
        RECT 919.950 820.950 922.050 823.050 ;
        RECT 935.400 817.050 936.450 829.950 ;
        RECT 940.950 823.950 943.050 826.050 ;
        RECT 913.950 814.950 916.050 817.050 ;
        RECT 934.950 814.950 937.050 817.050 ;
        RECT 904.950 806.100 907.050 808.200 ;
        RECT 910.950 806.100 913.050 808.200 ;
        RECT 905.400 805.350 906.600 806.100 ;
        RECT 911.400 805.350 912.600 806.100 ;
        RECT 916.800 805.950 918.900 808.050 ;
        RECT 919.950 805.950 922.050 808.050 ;
        RECT 928.950 806.100 931.050 808.200 ;
        RECT 935.400 807.600 936.450 814.950 ;
        RECT 901.950 802.950 904.050 805.050 ;
        RECT 904.950 802.950 907.050 805.050 ;
        RECT 907.950 802.950 910.050 805.050 ;
        RECT 910.950 802.950 913.050 805.050 ;
        RECT 902.400 800.400 903.600 802.650 ;
        RECT 908.400 800.400 909.600 802.650 ;
        RECT 917.400 801.900 918.450 805.950 ;
        RECT 902.400 798.450 903.450 800.400 ;
        RECT 902.400 797.400 906.450 798.450 ;
        RECT 895.950 793.950 898.050 796.050 ;
        RECT 883.950 760.950 886.050 763.050 ;
        RECT 889.950 762.000 892.050 766.050 ;
        RECT 901.950 763.950 904.050 766.050 ;
        RECT 890.400 760.350 891.600 762.000 ;
        RECT 895.950 761.100 898.050 763.200 ;
        RECT 896.400 760.350 897.600 761.100 ;
        RECT 886.950 757.950 889.050 760.050 ;
        RECT 889.950 757.950 892.050 760.050 ;
        RECT 892.950 757.950 895.050 760.050 ;
        RECT 895.950 757.950 898.050 760.050 ;
        RECT 887.400 756.900 888.600 757.650 ;
        RECT 886.950 754.800 889.050 756.900 ;
        RECT 893.400 755.400 894.600 757.650 ;
        RECT 893.400 753.450 894.450 755.400 ;
        RECT 898.950 754.950 901.050 757.050 ;
        RECT 890.400 752.400 894.450 753.450 ;
        RECT 890.400 730.200 891.450 752.400 ;
        RECT 899.400 738.450 900.450 754.950 ;
        RECT 902.400 748.050 903.450 763.950 ;
        RECT 905.400 757.050 906.450 797.400 ;
        RECT 908.400 781.050 909.450 800.400 ;
        RECT 916.950 799.800 919.050 801.900 ;
        RECT 907.950 778.950 910.050 781.050 ;
        RECT 913.950 769.950 916.050 772.050 ;
        RECT 914.400 762.600 915.450 769.950 ;
        RECT 920.400 766.200 921.450 805.950 ;
        RECT 929.400 805.350 930.600 806.100 ;
        RECT 935.400 805.350 936.600 807.600 ;
        RECT 925.950 802.950 928.050 805.050 ;
        RECT 928.950 802.950 931.050 805.050 ;
        RECT 931.950 802.950 934.050 805.050 ;
        RECT 934.950 802.950 937.050 805.050 ;
        RECT 926.400 800.400 927.600 802.650 ;
        RECT 932.400 801.900 933.600 802.650 ;
        RECT 926.400 793.050 927.450 800.400 ;
        RECT 931.950 799.800 934.050 801.900 ;
        RECT 937.950 799.950 940.050 802.050 ;
        RECT 934.950 796.950 937.050 799.050 ;
        RECT 925.950 790.950 928.050 793.050 ;
        RECT 919.950 764.100 922.050 766.200 ;
        RECT 926.400 763.050 927.450 790.950 ;
        RECT 931.950 772.950 934.050 775.050 ;
        RECT 928.950 763.950 931.050 766.050 ;
        RECT 914.400 760.350 915.600 762.600 ;
        RECT 919.950 760.950 922.050 763.050 ;
        RECT 925.950 760.950 928.050 763.050 ;
        RECT 920.400 760.350 921.600 760.950 ;
        RECT 907.950 757.950 910.050 760.050 ;
        RECT 913.950 757.950 916.050 760.050 ;
        RECT 916.950 757.950 919.050 760.050 ;
        RECT 919.950 757.950 922.050 760.050 ;
        RECT 922.950 757.950 925.050 760.050 ;
        RECT 904.950 754.950 907.050 757.050 ;
        RECT 901.950 745.950 904.050 748.050 ;
        RECT 901.950 738.450 904.050 739.050 ;
        RECT 899.400 737.400 904.050 738.450 ;
        RECT 901.950 736.950 904.050 737.400 ;
        RECT 880.950 728.100 883.050 730.200 ;
        RECT 889.950 728.100 892.050 730.200 ;
        RECT 895.950 728.100 898.050 730.200 ;
        RECT 877.950 715.950 880.050 718.050 ;
        RECT 862.950 712.950 865.050 715.050 ;
        RECT 865.950 708.450 868.050 712.050 ;
        RECT 863.400 708.000 868.050 708.450 ;
        RECT 863.400 707.400 867.450 708.000 ;
        RECT 848.400 684.450 849.600 684.600 ;
        RECT 842.400 683.400 849.600 684.450 ;
        RECT 838.950 655.950 841.050 658.050 ;
        RECT 842.400 652.200 843.450 683.400 ;
        RECT 848.400 682.350 849.600 683.400 ;
        RECT 853.950 683.100 856.050 685.200 ;
        RECT 854.400 682.350 855.600 683.100 ;
        RECT 847.950 679.950 850.050 682.050 ;
        RECT 850.950 679.950 853.050 682.050 ;
        RECT 853.950 679.950 856.050 682.050 ;
        RECT 856.950 679.950 859.050 682.050 ;
        RECT 851.400 677.400 852.600 679.650 ;
        RECT 857.400 679.050 858.600 679.650 ;
        RECT 863.400 679.050 864.450 707.400 ;
        RECT 868.950 706.950 871.050 709.050 ;
        RECT 865.950 683.100 868.050 685.200 ;
        RECT 869.400 685.050 870.450 706.950 ;
        RECT 881.400 697.050 882.450 728.100 ;
        RECT 890.400 727.350 891.600 728.100 ;
        RECT 896.400 727.350 897.600 728.100 ;
        RECT 886.950 724.950 889.050 727.050 ;
        RECT 889.950 724.950 892.050 727.050 ;
        RECT 892.950 724.950 895.050 727.050 ;
        RECT 895.950 724.950 898.050 727.050 ;
        RECT 883.950 721.950 886.050 724.050 ;
        RECT 887.400 723.900 888.600 724.650 ;
        RECT 893.400 723.900 894.600 724.650 ;
        RECT 902.400 723.900 903.450 736.950 ;
        RECT 904.950 727.950 907.050 730.050 ;
        RECT 880.950 694.950 883.050 697.050 ;
        RECT 874.950 688.950 877.050 691.050 ;
        RECT 857.400 677.400 862.050 679.050 ;
        RECT 851.400 664.050 852.450 677.400 ;
        RECT 858.000 676.950 862.050 677.400 ;
        RECT 862.950 676.950 865.050 679.050 ;
        RECT 866.400 666.450 867.450 683.100 ;
        RECT 868.950 682.950 871.050 685.050 ;
        RECT 875.400 684.600 876.450 688.950 ;
        RECT 875.400 682.350 876.600 684.600 ;
        RECT 880.800 683.100 882.900 685.200 ;
        RECT 884.400 685.050 885.450 721.950 ;
        RECT 886.950 721.800 889.050 723.900 ;
        RECT 892.950 721.800 895.050 723.900 ;
        RECT 901.950 721.800 904.050 723.900 ;
        RECT 889.950 718.950 892.050 721.050 ;
        RECT 886.950 715.950 889.050 718.050 ;
        RECT 881.400 682.350 882.600 683.100 ;
        RECT 883.950 682.950 886.050 685.050 ;
        RECT 871.950 679.950 874.050 682.050 ;
        RECT 874.950 679.950 877.050 682.050 ;
        RECT 877.950 679.950 880.050 682.050 ;
        RECT 880.950 679.950 883.050 682.050 ;
        RECT 872.400 678.900 873.600 679.650 ;
        RECT 871.950 676.800 874.050 678.900 ;
        RECT 878.400 677.400 879.600 679.650 ;
        RECT 872.400 670.050 873.450 676.800 ;
        RECT 874.950 673.950 877.050 676.050 ;
        RECT 871.950 667.950 874.050 670.050 ;
        RECT 868.950 666.450 871.050 667.050 ;
        RECT 866.400 665.400 871.050 666.450 ;
        RECT 868.950 664.950 871.050 665.400 ;
        RECT 850.950 663.450 853.050 664.050 ;
        RECT 848.400 662.400 853.050 663.450 ;
        RECT 844.950 658.950 847.050 661.050 ;
        RECT 830.400 649.350 831.600 651.600 ;
        RECT 836.400 649.350 837.600 651.600 ;
        RECT 841.950 650.100 844.050 652.200 ;
        RECT 826.950 646.950 829.050 649.050 ;
        RECT 829.950 646.950 832.050 649.050 ;
        RECT 832.950 646.950 835.050 649.050 ;
        RECT 835.950 646.950 838.050 649.050 ;
        RECT 827.400 645.900 828.600 646.650 ;
        RECT 833.400 645.900 834.600 646.650 ;
        RECT 842.400 645.900 843.450 650.100 ;
        RECT 820.950 643.800 823.050 645.900 ;
        RECT 826.950 643.800 829.050 645.900 ;
        RECT 832.950 643.800 835.050 645.900 ;
        RECT 841.950 643.800 844.050 645.900 ;
        RECT 845.400 637.050 846.450 658.950 ;
        RECT 848.400 645.900 849.450 662.400 ;
        RECT 850.950 661.950 853.050 662.400 ;
        RECT 856.950 650.100 859.050 652.200 ;
        RECT 862.950 650.100 865.050 652.200 ;
        RECT 857.400 649.350 858.600 650.100 ;
        RECT 863.400 649.350 864.600 650.100 ;
        RECT 853.950 646.950 856.050 649.050 ;
        RECT 856.950 646.950 859.050 649.050 ;
        RECT 859.950 646.950 862.050 649.050 ;
        RECT 862.950 646.950 865.050 649.050 ;
        RECT 854.400 645.900 855.600 646.650 ;
        RECT 860.400 645.900 861.600 646.650 ;
        RECT 847.950 643.800 850.050 645.900 ;
        RECT 853.950 643.800 856.050 645.900 ;
        RECT 859.950 643.800 862.050 645.900 ;
        RECT 865.950 643.950 868.050 646.050 ;
        RECT 862.950 640.950 865.050 643.050 ;
        RECT 817.950 634.950 820.050 637.050 ;
        RECT 844.950 634.950 847.050 637.050 ;
        RECT 859.950 622.950 862.050 625.050 ;
        RECT 826.950 619.950 829.050 622.050 ;
        RECT 844.950 619.950 847.050 622.050 ;
        RECT 820.950 613.950 823.050 616.050 ;
        RECT 821.400 606.600 822.450 613.950 ;
        RECT 827.400 606.600 828.450 619.950 ;
        RECT 841.950 613.950 844.050 616.050 ;
        RECT 821.400 604.350 822.600 606.600 ;
        RECT 827.400 604.350 828.600 606.600 ;
        RECT 842.400 606.450 843.450 613.950 ;
        RECT 839.400 605.400 843.450 606.450 ;
        RECT 845.400 606.600 846.450 619.950 ;
        RECT 820.950 601.950 823.050 604.050 ;
        RECT 823.950 601.950 826.050 604.050 ;
        RECT 826.950 601.950 829.050 604.050 ;
        RECT 829.950 601.950 832.050 604.050 ;
        RECT 824.400 600.900 825.600 601.650 ;
        RECT 815.400 599.400 819.450 600.450 ;
        RECT 808.950 595.950 811.050 598.050 ;
        RECT 799.950 592.950 802.050 595.050 ;
        RECT 811.950 572.100 814.050 574.200 ;
        RECT 818.400 573.600 819.450 599.400 ;
        RECT 823.950 598.800 826.050 600.900 ;
        RECT 830.400 600.000 831.600 601.650 ;
        RECT 839.400 600.900 840.450 605.400 ;
        RECT 845.400 604.350 846.600 606.600 ;
        RECT 850.950 605.100 853.050 607.200 ;
        RECT 851.400 604.350 852.600 605.100 ;
        RECT 844.950 601.950 847.050 604.050 ;
        RECT 847.950 601.950 850.050 604.050 ;
        RECT 850.950 601.950 853.050 604.050 ;
        RECT 853.950 601.950 856.050 604.050 ;
        RECT 848.400 600.900 849.600 601.650 ;
        RECT 829.950 595.950 832.050 600.000 ;
        RECT 838.950 598.800 841.050 600.900 ;
        RECT 847.950 598.800 850.050 600.900 ;
        RECT 854.400 599.400 855.600 601.650 ;
        RECT 850.950 595.950 853.050 598.050 ;
        RECT 812.400 571.350 813.600 572.100 ;
        RECT 818.400 571.350 819.600 573.600 ;
        RECT 826.950 572.100 829.050 574.200 ;
        RECT 811.950 568.950 814.050 571.050 ;
        RECT 814.950 568.950 817.050 571.050 ;
        RECT 817.950 568.950 820.050 571.050 ;
        RECT 820.950 568.950 823.050 571.050 ;
        RECT 815.400 567.900 816.600 568.650 ;
        RECT 794.400 566.400 798.450 567.450 ;
        RECT 763.950 562.950 766.050 565.050 ;
        RECT 760.950 556.950 763.050 559.050 ;
        RECT 757.950 535.950 760.050 538.050 ;
        RECT 758.400 523.050 759.450 535.950 ;
        RECT 764.400 535.050 765.450 562.950 ;
        RECT 785.400 556.050 786.450 566.400 ;
        RECT 814.950 565.800 817.050 567.900 ;
        RECT 821.400 566.400 822.600 568.650 ;
        RECT 821.400 556.050 822.450 566.400 ;
        RECT 823.950 565.800 826.050 567.900 ;
        RECT 824.400 562.050 825.450 565.800 ;
        RECT 823.950 559.950 826.050 562.050 ;
        RECT 784.950 553.950 787.050 556.050 ;
        RECT 814.950 553.950 817.050 556.050 ;
        RECT 820.950 553.950 823.050 556.050 ;
        RECT 784.950 541.950 787.050 544.050 ;
        RECT 763.950 532.950 766.050 535.050 ;
        RECT 760.950 527.100 763.050 529.200 ;
        RECT 769.950 527.100 772.050 532.050 ;
        RECT 778.950 529.950 784.050 532.050 ;
        RECT 776.400 528.450 777.600 528.600 ;
        RECT 776.400 527.400 783.450 528.450 ;
        RECT 757.950 520.950 760.050 523.050 ;
        RECT 761.400 520.050 762.450 527.100 ;
        RECT 770.400 526.350 771.600 527.100 ;
        RECT 776.400 526.350 777.600 527.400 ;
        RECT 766.950 523.950 769.050 526.050 ;
        RECT 769.950 523.950 772.050 526.050 ;
        RECT 772.950 523.950 775.050 526.050 ;
        RECT 775.950 523.950 778.050 526.050 ;
        RECT 767.400 523.050 768.600 523.650 ;
        RECT 763.950 521.400 768.600 523.050 ;
        RECT 773.400 522.900 774.600 523.650 ;
        RECT 763.950 520.950 768.000 521.400 ;
        RECT 772.950 520.800 775.050 522.900 ;
        RECT 760.950 517.950 763.050 520.050 ;
        RECT 742.950 514.950 745.050 517.050 ;
        RECT 754.950 514.950 757.050 517.050 ;
        RECT 739.950 502.950 742.050 505.050 ;
        RECT 727.950 451.950 730.050 454.050 ;
        RECT 736.950 451.950 739.050 454.050 ;
        RECT 725.400 448.350 726.600 450.600 ;
        RECT 730.950 449.100 733.050 451.200 ;
        RECT 731.400 448.350 732.600 449.100 ;
        RECT 700.950 445.950 703.050 448.050 ;
        RECT 703.950 445.950 706.050 448.050 ;
        RECT 706.950 445.950 709.050 448.050 ;
        RECT 709.950 445.950 712.050 448.050 ;
        RECT 724.950 445.950 727.050 448.050 ;
        RECT 727.950 445.950 730.050 448.050 ;
        RECT 730.950 445.950 733.050 448.050 ;
        RECT 733.950 445.950 736.050 448.050 ;
        RECT 704.400 443.400 705.600 445.650 ;
        RECT 710.400 444.900 711.600 445.650 ;
        RECT 728.400 444.900 729.600 445.650 ;
        RECT 704.400 433.050 705.450 443.400 ;
        RECT 709.950 442.800 712.050 444.900 ;
        RECT 727.950 442.800 730.050 444.900 ;
        RECT 734.400 443.400 735.600 445.650 ;
        RECT 740.400 445.050 741.450 502.950 ;
        RECT 743.400 484.050 744.450 514.950 ;
        RECT 782.400 511.050 783.450 527.400 ;
        RECT 785.400 523.050 786.450 541.950 ;
        RECT 799.950 538.950 802.050 541.050 ;
        RECT 787.950 535.950 790.050 538.050 ;
        RECT 788.400 529.050 789.450 535.950 ;
        RECT 800.400 535.050 801.450 538.950 ;
        RECT 799.950 532.950 802.050 535.050 ;
        RECT 805.950 532.950 808.050 535.050 ;
        RECT 787.950 526.950 790.050 529.050 ;
        RECT 793.950 528.000 796.050 532.050 ;
        RECT 794.400 526.350 795.600 528.000 ;
        RECT 799.950 527.100 802.050 529.200 ;
        RECT 800.400 526.350 801.600 527.100 ;
        RECT 790.950 523.950 793.050 526.050 ;
        RECT 793.950 523.950 796.050 526.050 ;
        RECT 796.950 523.950 799.050 526.050 ;
        RECT 799.950 523.950 802.050 526.050 ;
        RECT 784.950 520.950 787.050 523.050 ;
        RECT 791.400 522.900 792.600 523.650 ;
        RECT 790.950 520.800 793.050 522.900 ;
        RECT 797.400 521.400 798.600 523.650 ;
        RECT 793.950 517.950 796.050 520.050 ;
        RECT 781.950 508.950 784.050 511.050 ;
        RECT 778.950 505.950 781.050 508.050 ;
        RECT 779.400 502.050 780.450 505.950 ;
        RECT 778.950 499.950 781.050 502.050 ;
        RECT 751.950 494.100 754.050 496.200 ;
        RECT 763.950 494.100 766.050 496.200 ;
        RECT 769.950 494.100 772.050 496.200 ;
        RECT 752.400 493.350 753.600 494.100 ;
        RECT 748.950 490.950 751.050 493.050 ;
        RECT 751.950 490.950 754.050 493.050 ;
        RECT 754.950 490.950 757.050 493.050 ;
        RECT 760.950 490.950 763.050 493.050 ;
        RECT 749.400 489.900 750.600 490.650 ;
        RECT 748.950 487.800 751.050 489.900 ;
        RECT 755.400 488.400 756.600 490.650 ;
        RECT 755.400 484.050 756.450 488.400 ;
        RECT 761.400 487.050 762.450 490.950 ;
        RECT 760.950 484.950 763.050 487.050 ;
        RECT 742.950 481.950 745.050 484.050 ;
        RECT 754.950 481.950 757.050 484.050 ;
        RECT 764.400 483.450 765.450 494.100 ;
        RECT 770.400 493.350 771.600 494.100 ;
        RECT 769.950 490.950 772.050 493.050 ;
        RECT 772.950 490.950 775.050 493.050 ;
        RECT 773.400 489.450 774.600 490.650 ;
        RECT 779.400 489.450 780.450 499.950 ;
        RECT 787.950 494.100 790.050 496.200 ;
        RECT 794.400 495.600 795.450 517.950 ;
        RECT 797.400 517.050 798.450 521.400 ;
        RECT 806.400 517.050 807.450 532.950 ;
        RECT 808.950 527.100 811.050 529.200 ;
        RECT 815.400 528.600 816.450 553.950 ;
        RECT 796.950 514.950 799.050 517.050 ;
        RECT 805.950 514.950 808.050 517.050 ;
        RECT 809.400 511.050 810.450 527.100 ;
        RECT 815.400 526.350 816.600 528.600 ;
        RECT 820.950 527.100 823.050 529.200 ;
        RECT 827.400 529.050 828.450 572.100 ;
        RECT 830.400 559.050 831.450 595.950 ;
        RECT 835.950 573.000 838.050 577.050 ;
        RECT 836.400 571.350 837.600 573.000 ;
        RECT 841.950 572.100 844.050 574.200 ;
        RECT 842.400 571.350 843.600 572.100 ;
        RECT 835.950 568.950 838.050 571.050 ;
        RECT 838.950 568.950 841.050 571.050 ;
        RECT 841.950 568.950 844.050 571.050 ;
        RECT 844.950 568.950 847.050 571.050 ;
        RECT 839.400 567.900 840.600 568.650 ;
        RECT 838.950 565.800 841.050 567.900 ;
        RECT 845.400 566.400 846.600 568.650 ;
        RECT 845.400 562.050 846.450 566.400 ;
        RECT 844.950 559.950 847.050 562.050 ;
        RECT 829.950 556.950 832.050 559.050 ;
        RECT 838.950 553.950 841.050 556.050 ;
        RECT 829.950 544.950 832.050 547.050 ;
        RECT 821.400 526.350 822.600 527.100 ;
        RECT 826.950 526.950 829.050 529.050 ;
        RECT 814.950 523.950 817.050 526.050 ;
        RECT 817.950 523.950 820.050 526.050 ;
        RECT 820.950 523.950 823.050 526.050 ;
        RECT 823.950 523.950 826.050 526.050 ;
        RECT 818.400 522.900 819.600 523.650 ;
        RECT 817.950 520.800 820.050 522.900 ;
        RECT 824.400 521.400 825.600 523.650 ;
        RECT 818.400 514.050 819.450 520.800 ;
        RECT 824.400 514.050 825.450 521.400 ;
        RECT 826.950 520.950 829.050 523.050 ;
        RECT 817.950 511.950 820.050 514.050 ;
        RECT 823.950 511.950 826.050 514.050 ;
        RECT 808.950 508.950 811.050 511.050 ;
        RECT 805.950 499.950 808.050 502.050 ;
        RECT 820.950 499.950 823.050 502.050 ;
        RECT 788.400 493.350 789.600 494.100 ;
        RECT 794.400 493.350 795.600 495.600 ;
        RECT 802.950 494.100 805.050 496.200 ;
        RECT 787.950 490.950 790.050 493.050 ;
        RECT 790.950 490.950 793.050 493.050 ;
        RECT 793.950 490.950 796.050 493.050 ;
        RECT 796.950 490.950 799.050 493.050 ;
        RECT 773.400 488.400 780.450 489.450 ;
        RECT 791.400 488.400 792.600 490.650 ;
        RECT 797.400 489.000 798.600 490.650 ;
        RECT 803.400 489.450 804.450 494.100 ;
        RECT 806.400 489.900 807.450 499.950 ;
        RECT 814.950 494.100 817.050 496.200 ;
        RECT 821.400 495.600 822.450 499.950 ;
        RECT 815.400 493.350 816.600 494.100 ;
        RECT 821.400 493.350 822.600 495.600 ;
        RECT 811.950 490.950 814.050 493.050 ;
        RECT 814.950 490.950 817.050 493.050 ;
        RECT 817.950 490.950 820.050 493.050 ;
        RECT 820.950 490.950 823.050 493.050 ;
        RECT 812.400 489.900 813.600 490.650 ;
        RECT 761.400 482.400 765.450 483.450 ;
        RECT 748.950 480.450 751.050 481.050 ;
        RECT 757.950 480.450 760.050 481.050 ;
        RECT 748.950 479.400 760.050 480.450 ;
        RECT 748.950 478.950 751.050 479.400 ;
        RECT 757.950 478.950 760.050 479.400 ;
        RECT 761.400 469.050 762.450 482.400 ;
        RECT 791.400 481.050 792.450 488.400 ;
        RECT 796.950 484.950 799.050 489.000 ;
        RECT 800.400 488.400 804.450 489.450 ;
        RECT 790.950 478.950 793.050 481.050 ;
        RECT 796.950 472.950 799.050 475.050 ;
        RECT 760.950 466.950 763.050 469.050 ;
        RECT 742.950 449.100 745.050 451.200 ;
        RECT 748.950 450.000 751.050 454.050 ;
        RECT 706.950 439.950 709.050 442.050 ;
        RECT 734.400 441.450 735.450 443.400 ;
        RECT 736.950 442.950 739.050 445.050 ;
        RECT 739.950 442.950 742.050 445.050 ;
        RECT 743.400 444.450 744.450 449.100 ;
        RECT 749.400 448.350 750.600 450.000 ;
        RECT 748.950 445.950 751.050 448.050 ;
        RECT 751.950 445.950 754.050 448.050 ;
        RECT 754.950 445.950 757.050 448.050 ;
        RECT 752.400 444.900 753.600 445.650 ;
        RECT 761.400 445.050 762.450 466.950 ;
        RECT 769.950 454.950 772.050 457.050 ;
        RECT 781.950 454.950 784.050 457.050 ;
        RECT 770.400 450.600 771.450 454.950 ;
        RECT 770.400 448.350 771.600 450.600 ;
        RECT 769.950 445.950 772.050 448.050 ;
        RECT 772.950 445.950 775.050 448.050 ;
        RECT 775.950 445.950 778.050 448.050 ;
        RECT 743.400 443.400 747.450 444.450 ;
        RECT 731.400 440.400 735.450 441.450 ;
        RECT 703.950 430.950 706.050 433.050 ;
        RECT 694.950 427.950 697.050 430.050 ;
        RECT 703.950 427.800 706.050 429.900 ;
        RECT 682.950 412.950 685.050 415.050 ;
        RECT 685.950 412.950 688.050 415.050 ;
        RECT 688.950 412.950 691.050 415.050 ;
        RECT 691.950 412.950 694.050 415.050 ;
        RECT 694.950 412.950 697.050 415.050 ;
        RECT 683.400 410.400 684.600 412.650 ;
        RECT 689.400 410.400 690.600 412.650 ;
        RECT 695.400 410.400 696.600 412.650 ;
        RECT 704.400 412.050 705.450 427.800 ;
        RECT 676.950 406.950 679.050 409.050 ;
        RECT 683.400 406.050 684.450 410.400 ;
        RECT 685.950 406.950 688.050 409.050 ;
        RECT 673.950 403.950 676.050 406.050 ;
        RECT 682.950 403.950 685.050 406.050 ;
        RECT 670.950 385.950 673.050 388.050 ;
        RECT 676.950 379.950 679.050 382.050 ;
        RECT 670.950 370.950 673.050 373.050 ;
        RECT 677.400 372.600 678.450 379.950 ;
        RECT 686.400 379.050 687.450 406.950 ;
        RECT 689.400 385.050 690.450 410.400 ;
        RECT 695.400 408.450 696.450 410.400 ;
        RECT 703.950 409.950 706.050 412.050 ;
        RECT 707.400 409.050 708.450 439.950 ;
        RECT 712.950 412.950 715.050 415.050 ;
        RECT 715.950 412.950 718.050 415.050 ;
        RECT 716.400 410.400 717.600 412.650 ;
        RECT 692.400 407.400 696.450 408.450 ;
        RECT 692.400 394.050 693.450 407.400 ;
        RECT 706.950 406.950 709.050 409.050 ;
        RECT 712.950 406.950 715.050 409.050 ;
        RECT 694.950 403.950 697.050 406.050 ;
        RECT 691.950 391.950 694.050 394.050 ;
        RECT 688.950 382.950 691.050 385.050 ;
        RECT 685.950 376.950 688.050 379.050 ;
        RECT 691.950 376.950 694.050 379.050 ;
        RECT 671.400 364.050 672.450 370.950 ;
        RECT 677.400 370.350 678.600 372.600 ;
        RECT 682.950 372.000 685.050 376.050 ;
        RECT 683.400 370.350 684.600 372.000 ;
        RECT 676.950 367.950 679.050 370.050 ;
        RECT 679.950 367.950 682.050 370.050 ;
        RECT 682.950 367.950 685.050 370.050 ;
        RECT 685.950 367.950 688.050 370.050 ;
        RECT 680.400 365.400 681.600 367.650 ;
        RECT 686.400 365.400 687.600 367.650 ;
        RECT 670.950 361.950 673.050 364.050 ;
        RECT 676.950 355.950 679.050 358.050 ;
        RECT 661.950 337.950 664.050 340.050 ;
        RECT 667.950 338.100 670.050 340.200 ;
        RECT 658.950 319.950 661.050 322.050 ;
        RECT 646.950 310.950 649.050 313.050 ;
        RECT 647.400 304.050 648.450 310.950 ;
        RECT 646.950 301.950 649.050 304.050 ;
        RECT 644.400 292.350 645.600 294.600 ;
        RECT 649.950 294.000 652.050 298.050 ;
        RECT 658.950 295.950 661.050 298.050 ;
        RECT 662.400 297.450 663.450 337.950 ;
        RECT 668.400 337.350 669.600 338.100 ;
        RECT 667.950 334.950 670.050 337.050 ;
        RECT 670.950 334.950 673.050 337.050 ;
        RECT 671.400 332.400 672.600 334.650 ;
        RECT 671.400 328.050 672.450 332.400 ;
        RECT 670.950 325.950 673.050 328.050 ;
        RECT 671.400 313.050 672.450 325.950 ;
        RECT 670.950 310.950 673.050 313.050 ;
        RECT 662.400 296.400 666.450 297.450 ;
        RECT 650.400 292.350 651.600 294.000 ;
        RECT 640.950 289.950 643.050 292.050 ;
        RECT 643.950 289.950 646.050 292.050 ;
        RECT 646.950 289.950 649.050 292.050 ;
        RECT 649.950 289.950 652.050 292.050 ;
        RECT 652.950 289.950 655.050 292.050 ;
        RECT 641.400 287.400 642.600 289.650 ;
        RECT 647.400 288.900 648.600 289.650 ;
        RECT 632.400 259.350 633.600 261.600 ;
        RECT 628.950 256.950 631.050 259.050 ;
        RECT 631.950 256.950 634.050 259.050 ;
        RECT 634.950 256.950 637.050 259.050 ;
        RECT 629.400 255.000 630.600 256.650 ;
        RECT 628.950 250.950 631.050 255.000 ;
        RECT 641.400 250.050 642.450 287.400 ;
        RECT 646.950 286.800 649.050 288.900 ;
        RECT 653.400 287.400 654.600 289.650 ;
        RECT 659.400 288.450 660.450 295.950 ;
        RECT 661.950 292.950 664.050 295.050 ;
        RECT 656.400 287.400 660.450 288.450 ;
        RECT 646.950 271.950 649.050 274.050 ;
        RECT 640.950 247.950 643.050 250.050 ;
        RECT 628.950 229.950 631.050 232.050 ;
        RECT 629.400 217.050 630.450 229.950 ;
        RECT 634.950 223.950 637.050 226.050 ;
        RECT 640.950 223.950 643.050 226.050 ;
        RECT 628.950 214.950 631.050 217.050 ;
        RECT 635.400 216.600 636.450 223.950 ;
        RECT 641.400 216.600 642.450 223.950 ;
        RECT 635.400 214.350 636.600 216.600 ;
        RECT 641.400 214.350 642.600 216.600 ;
        RECT 631.950 211.950 634.050 214.050 ;
        RECT 634.950 211.950 637.050 214.050 ;
        RECT 637.950 211.950 640.050 214.050 ;
        RECT 640.950 211.950 643.050 214.050 ;
        RECT 632.400 209.400 633.600 211.650 ;
        RECT 638.400 210.900 639.600 211.650 ;
        RECT 632.400 183.450 633.450 209.400 ;
        RECT 637.950 208.800 640.050 210.900 ;
        RECT 647.400 205.050 648.450 271.950 ;
        RECT 653.400 271.050 654.450 287.400 ;
        RECT 652.950 268.950 655.050 271.050 ;
        RECT 656.400 261.600 657.450 287.400 ;
        RECT 658.950 277.950 661.050 280.050 ;
        RECT 659.400 271.050 660.450 277.950 ;
        RECT 658.950 268.950 661.050 271.050 ;
        RECT 662.400 262.050 663.450 292.950 ;
        RECT 656.400 259.350 657.600 261.600 ;
        RECT 661.950 259.950 664.050 262.050 ;
        RECT 652.950 256.950 655.050 259.050 ;
        RECT 655.950 256.950 658.050 259.050 ;
        RECT 658.950 256.950 661.050 259.050 ;
        RECT 653.400 254.400 654.600 256.650 ;
        RECT 659.400 254.400 660.600 256.650 ;
        RECT 653.400 250.050 654.450 254.400 ;
        RECT 652.950 247.950 655.050 250.050 ;
        RECT 659.400 241.050 660.450 254.400 ;
        RECT 661.950 253.950 664.050 256.050 ;
        RECT 662.400 247.050 663.450 253.950 ;
        RECT 665.400 253.050 666.450 296.400 ;
        RECT 670.950 294.000 673.050 298.050 ;
        RECT 677.400 294.600 678.450 355.950 ;
        RECT 680.400 346.050 681.450 365.400 ;
        RECT 682.950 361.950 685.050 364.050 ;
        RECT 679.950 343.950 682.050 346.050 ;
        RECT 679.950 340.800 682.050 342.900 ;
        RECT 680.400 313.050 681.450 340.800 ;
        RECT 683.400 328.050 684.450 361.950 ;
        RECT 686.400 343.050 687.450 365.400 ;
        RECT 692.400 346.050 693.450 376.950 ;
        RECT 695.400 366.450 696.450 403.950 ;
        RECT 703.950 376.950 706.050 379.050 ;
        RECT 704.400 372.600 705.450 376.950 ;
        RECT 704.400 370.350 705.600 372.600 ;
        RECT 700.950 367.950 703.050 370.050 ;
        RECT 703.950 367.950 706.050 370.050 ;
        RECT 706.950 367.950 709.050 370.050 ;
        RECT 695.400 365.400 699.450 366.450 ;
        RECT 691.950 343.950 694.050 346.050 ;
        RECT 685.950 340.950 688.050 343.050 ;
        RECT 686.100 334.950 688.200 337.050 ;
        RECT 691.500 334.950 693.600 337.050 ;
        RECT 694.800 334.950 696.900 337.050 ;
        RECT 686.400 332.400 687.600 334.650 ;
        RECT 695.400 333.000 696.600 334.650 ;
        RECT 682.950 325.950 685.050 328.050 ;
        RECT 682.950 322.800 685.050 324.900 ;
        RECT 679.950 310.950 682.050 313.050 ;
        RECT 671.400 292.350 672.600 294.000 ;
        RECT 677.400 292.350 678.600 294.600 ;
        RECT 683.400 294.450 684.450 322.800 ;
        RECT 686.400 319.050 687.450 332.400 ;
        RECT 694.950 328.950 697.050 333.000 ;
        RECT 698.400 325.050 699.450 365.400 ;
        RECT 701.400 365.400 702.600 367.650 ;
        RECT 707.400 366.900 708.600 367.650 ;
        RECT 701.400 352.050 702.450 365.400 ;
        RECT 706.950 364.800 709.050 366.900 ;
        RECT 713.400 358.050 714.450 406.950 ;
        RECT 716.400 403.050 717.450 410.400 ;
        RECT 731.400 409.050 732.450 440.400 ;
        RECT 737.400 430.050 738.450 442.950 ;
        RECT 746.400 439.050 747.450 443.400 ;
        RECT 751.950 442.800 754.050 444.900 ;
        RECT 760.950 442.950 763.050 445.050 ;
        RECT 773.400 444.900 774.600 445.650 ;
        RECT 772.950 442.800 775.050 444.900 ;
        RECT 782.400 442.050 783.450 454.950 ;
        RECT 787.950 451.950 790.050 454.050 ;
        RECT 788.400 445.050 789.450 451.950 ;
        RECT 797.400 450.600 798.450 472.950 ;
        RECT 800.400 463.050 801.450 488.400 ;
        RECT 805.950 487.800 808.050 489.900 ;
        RECT 811.950 487.800 814.050 489.900 ;
        RECT 818.400 489.000 819.600 490.650 ;
        RECT 817.950 484.950 820.050 489.000 ;
        RECT 827.400 475.050 828.450 520.950 ;
        RECT 826.950 472.950 829.050 475.050 ;
        RECT 830.400 463.050 831.450 544.950 ;
        RECT 832.950 538.950 835.050 541.050 ;
        RECT 833.400 511.050 834.450 538.950 ;
        RECT 839.400 528.600 840.450 553.950 ;
        RECT 845.400 547.050 846.450 559.950 ;
        RECT 844.950 544.950 847.050 547.050 ;
        RECT 839.400 526.350 840.600 528.600 ;
        RECT 844.950 527.100 847.050 529.200 ;
        RECT 851.400 529.050 852.450 595.950 ;
        RECT 854.400 577.050 855.450 599.400 ;
        RECT 860.400 595.050 861.450 622.950 ;
        RECT 859.950 592.950 862.050 595.050 ;
        RECT 863.400 586.050 864.450 640.950 ;
        RECT 866.400 607.050 867.450 643.950 ;
        RECT 869.400 643.050 870.450 664.950 ;
        RECT 875.400 652.050 876.450 673.950 ;
        RECT 878.400 658.050 879.450 677.400 ;
        RECT 887.400 675.450 888.450 715.950 ;
        RECT 890.400 678.450 891.450 718.950 ;
        RECT 905.400 697.050 906.450 727.950 ;
        RECT 908.400 712.050 909.450 757.950 ;
        RECT 917.400 756.900 918.600 757.650 ;
        RECT 916.950 754.800 919.050 756.900 ;
        RECT 923.400 755.400 924.600 757.650 ;
        RECT 919.950 748.950 922.050 751.050 ;
        RECT 913.950 728.100 916.050 730.200 ;
        RECT 920.400 729.600 921.450 748.950 ;
        RECT 923.400 748.050 924.450 755.400 ;
        RECT 925.950 754.950 928.050 757.050 ;
        RECT 929.400 756.900 930.450 763.950 ;
        RECT 926.400 751.050 927.450 754.950 ;
        RECT 928.950 754.800 931.050 756.900 ;
        RECT 925.950 748.950 928.050 751.050 ;
        RECT 922.950 745.950 925.050 748.050 ;
        RECT 925.950 739.950 928.050 742.050 ;
        RECT 926.400 733.050 927.450 739.950 ;
        RECT 932.400 736.050 933.450 772.950 ;
        RECT 931.950 733.950 934.050 736.050 ;
        RECT 925.950 730.950 928.050 733.050 ;
        RECT 931.950 730.800 934.050 732.900 ;
        RECT 914.400 727.350 915.600 728.100 ;
        RECT 920.400 727.350 921.600 729.600 ;
        RECT 913.950 724.950 916.050 727.050 ;
        RECT 916.950 724.950 919.050 727.050 ;
        RECT 919.950 724.950 922.050 727.050 ;
        RECT 922.950 724.950 925.050 727.050 ;
        RECT 917.400 722.400 918.600 724.650 ;
        RECT 923.400 722.400 924.600 724.650 ;
        RECT 907.950 709.950 910.050 712.050 ;
        RECT 917.400 709.050 918.450 722.400 ;
        RECT 916.950 706.950 919.050 709.050 ;
        RECT 898.950 694.950 901.050 697.050 ;
        RECT 904.950 694.950 907.050 697.050 ;
        RECT 899.400 691.050 900.450 694.950 ;
        RECT 898.950 688.950 901.050 691.050 ;
        RECT 899.400 684.600 900.450 688.950 ;
        RECT 923.400 688.050 924.450 722.400 ;
        RECT 932.400 700.050 933.450 730.800 ;
        RECT 935.400 730.050 936.450 796.950 ;
        RECT 938.400 769.050 939.450 799.950 ;
        RECT 941.400 799.050 942.450 823.950 ;
        RECT 943.950 811.950 946.050 814.050 ;
        RECT 944.400 802.050 945.450 811.950 ;
        RECT 947.400 808.050 948.450 829.950 ;
        RECT 950.400 826.050 951.450 833.400 ;
        RECT 958.950 832.800 961.050 834.900 ;
        RECT 955.950 826.950 958.050 829.050 ;
        RECT 949.950 823.950 952.050 826.050 ;
        RECT 956.400 811.050 957.450 826.950 ;
        RECT 946.950 805.950 949.050 808.050 ;
        RECT 949.950 806.100 952.050 808.200 ;
        RECT 955.950 806.100 958.050 811.050 ;
        RECT 950.400 805.350 951.600 806.100 ;
        RECT 949.950 802.950 952.050 805.050 ;
        RECT 952.950 802.950 955.050 805.050 ;
        RECT 943.950 799.950 946.050 802.050 ;
        RECT 953.400 801.900 954.600 802.650 ;
        RECT 952.950 799.800 955.050 801.900 ;
        RECT 955.950 799.950 958.050 802.050 ;
        RECT 940.950 796.950 943.050 799.050 ;
        RECT 956.400 793.050 957.450 799.950 ;
        RECT 955.950 790.950 958.050 793.050 ;
        RECT 937.950 766.950 940.050 769.050 ;
        RECT 938.400 762.450 939.450 766.950 ;
        RECT 956.400 763.200 957.450 790.950 ;
        RECT 941.400 762.450 942.600 762.600 ;
        RECT 938.400 761.400 942.600 762.450 ;
        RECT 941.400 760.350 942.600 761.400 ;
        RECT 946.950 761.100 949.050 763.200 ;
        RECT 955.950 761.100 958.050 763.200 ;
        RECT 947.400 760.350 948.600 761.100 ;
        RECT 940.950 757.950 943.050 760.050 ;
        RECT 943.950 757.950 946.050 760.050 ;
        RECT 946.950 757.950 949.050 760.050 ;
        RECT 949.950 757.950 952.050 760.050 ;
        RECT 944.400 756.900 945.600 757.650 ;
        RECT 943.950 751.950 946.050 756.900 ;
        RECT 950.400 755.400 951.600 757.650 ;
        RECT 956.400 756.450 957.450 761.100 ;
        RECT 953.400 755.400 957.450 756.450 ;
        RECT 950.400 751.050 951.450 755.400 ;
        RECT 949.950 748.950 952.050 751.050 ;
        RECT 953.400 747.450 954.450 755.400 ;
        RECT 950.400 746.400 954.450 747.450 ;
        RECT 950.400 742.050 951.450 746.400 ;
        RECT 952.950 742.950 955.050 745.050 ;
        RECT 949.950 739.950 952.050 742.050 ;
        RECT 937.950 736.950 940.050 739.050 ;
        RECT 934.950 727.950 937.050 730.050 ;
        RECT 938.400 729.600 939.450 736.950 ;
        RECT 949.950 730.950 952.050 736.050 ;
        RECT 938.400 727.350 939.600 729.600 ;
        RECT 943.950 728.100 946.050 730.200 ;
        RECT 944.400 727.350 945.600 728.100 ;
        RECT 937.950 724.950 940.050 727.050 ;
        RECT 940.950 724.950 943.050 727.050 ;
        RECT 943.950 724.950 946.050 727.050 ;
        RECT 946.950 724.950 949.050 727.050 ;
        RECT 934.950 721.950 937.050 724.050 ;
        RECT 941.400 722.400 942.600 724.650 ;
        RECT 947.400 722.400 948.600 724.650 ;
        RECT 931.950 697.950 934.050 700.050 ;
        RECT 935.400 691.050 936.450 721.950 ;
        RECT 937.950 718.950 940.050 721.050 ;
        RECT 938.400 703.050 939.450 718.950 ;
        RECT 941.400 715.050 942.450 722.400 ;
        RECT 940.950 712.950 943.050 715.050 ;
        RECT 941.400 706.050 942.450 712.950 ;
        RECT 947.400 712.050 948.450 722.400 ;
        RECT 953.400 718.050 954.450 742.950 ;
        RECT 955.950 736.950 958.050 739.050 ;
        RECT 952.950 715.950 955.050 718.050 ;
        RECT 946.950 709.950 949.050 712.050 ;
        RECT 956.400 706.050 957.450 736.950 ;
        RECT 959.400 736.050 960.450 832.800 ;
        RECT 962.400 829.050 963.450 841.950 ;
        RECT 961.950 826.950 964.050 829.050 ;
        RECT 965.400 825.450 966.450 868.950 ;
        RECT 962.400 824.400 966.450 825.450 ;
        RECT 962.400 796.050 963.450 824.400 ;
        RECT 968.400 814.050 969.450 877.950 ;
        RECT 971.400 868.050 972.450 878.400 ;
        RECT 977.400 871.050 978.450 878.400 ;
        RECT 982.950 877.950 985.050 880.050 ;
        RECT 976.950 868.950 979.050 871.050 ;
        RECT 970.950 865.950 973.050 868.050 ;
        RECT 983.400 865.050 984.450 877.950 ;
        RECT 986.400 865.050 987.450 901.950 ;
        RECT 989.400 879.450 990.450 916.950 ;
        RECT 992.400 904.050 993.450 919.950 ;
        RECT 994.950 917.100 997.050 919.200 ;
        RECT 1000.950 917.100 1003.050 919.200 ;
        RECT 1006.950 918.000 1009.050 922.050 ;
        RECT 995.400 910.050 996.450 917.100 ;
        RECT 1001.400 916.350 1002.600 917.100 ;
        RECT 1007.400 916.350 1008.600 918.000 ;
        RECT 1000.950 913.950 1003.050 916.050 ;
        RECT 1003.950 913.950 1006.050 916.050 ;
        RECT 1006.950 913.950 1009.050 916.050 ;
        RECT 1009.950 913.950 1012.050 916.050 ;
        RECT 1004.400 911.400 1005.600 913.650 ;
        RECT 1010.400 912.450 1011.600 913.650 ;
        RECT 1010.400 911.400 1014.450 912.450 ;
        RECT 994.950 907.950 997.050 910.050 ;
        RECT 1004.400 909.450 1005.450 911.400 ;
        RECT 1004.400 908.400 1008.450 909.450 ;
        RECT 991.950 901.950 994.050 904.050 ;
        RECT 1003.950 901.950 1006.050 904.050 ;
        RECT 997.950 884.100 1000.050 886.200 ;
        RECT 1004.400 885.600 1005.450 901.950 ;
        RECT 1007.400 886.050 1008.450 908.400 ;
        RECT 1009.950 907.950 1012.050 910.050 ;
        RECT 998.400 883.350 999.600 884.100 ;
        RECT 1004.400 883.350 1005.600 885.600 ;
        RECT 1006.950 883.950 1009.050 886.050 ;
        RECT 994.950 880.950 997.050 883.050 ;
        RECT 997.950 880.950 1000.050 883.050 ;
        RECT 1000.950 880.950 1003.050 883.050 ;
        RECT 1003.950 880.950 1006.050 883.050 ;
        RECT 989.400 878.400 993.450 879.450 ;
        RECT 970.950 862.800 973.050 864.900 ;
        RECT 982.800 862.950 984.900 865.050 ;
        RECT 985.950 862.950 988.050 865.050 ;
        RECT 971.400 829.050 972.450 862.800 ;
        RECT 988.950 856.950 991.050 859.050 ;
        RECT 973.950 847.950 976.050 850.050 ;
        RECT 974.400 841.050 975.450 847.950 ;
        RECT 976.950 844.050 979.050 844.200 ;
        RECT 979.950 844.050 982.050 844.200 ;
        RECT 976.950 842.100 982.050 844.050 ;
        RECT 978.000 841.950 981.000 842.100 ;
        RECT 973.950 838.950 976.050 841.050 ;
        RECT 979.950 838.950 982.050 841.050 ;
        RECT 985.950 840.000 988.050 844.050 ;
        RECT 989.400 841.050 990.450 856.950 ;
        RECT 980.400 838.350 981.600 838.950 ;
        RECT 986.400 838.350 987.600 840.000 ;
        RECT 988.950 838.950 991.050 841.050 ;
        RECT 976.950 835.950 979.050 838.050 ;
        RECT 979.950 835.950 982.050 838.050 ;
        RECT 982.950 835.950 985.050 838.050 ;
        RECT 985.950 835.950 988.050 838.050 ;
        RECT 973.950 832.950 976.050 835.050 ;
        RECT 977.400 833.400 978.600 835.650 ;
        RECT 983.400 833.400 984.600 835.650 ;
        RECT 992.400 835.050 993.450 878.400 ;
        RECT 995.400 878.400 996.600 880.650 ;
        RECT 1001.400 878.400 1002.600 880.650 ;
        RECT 1010.400 879.450 1011.450 907.950 ;
        RECT 1013.400 882.450 1014.450 911.400 ;
        RECT 1016.400 886.050 1017.450 943.950 ;
        RECT 1015.950 883.950 1018.050 886.050 ;
        RECT 1013.400 881.400 1017.450 882.450 ;
        RECT 1010.400 878.400 1014.450 879.450 ;
        RECT 995.400 871.050 996.450 878.400 ;
        RECT 994.950 868.950 997.050 871.050 ;
        RECT 1001.400 868.050 1002.450 878.400 ;
        RECT 1009.950 874.950 1012.050 877.050 ;
        RECT 1000.950 865.950 1003.050 868.050 ;
        RECT 997.950 862.950 1000.050 865.050 ;
        RECT 994.950 850.950 997.050 853.050 ;
        RECT 970.950 826.950 973.050 829.050 ;
        RECT 974.400 819.450 975.450 832.950 ;
        RECT 977.400 832.050 978.450 833.400 ;
        RECT 977.400 830.400 982.050 832.050 ;
        RECT 978.000 829.950 982.050 830.400 ;
        RECT 983.400 823.050 984.450 833.400 ;
        RECT 991.950 832.950 994.050 835.050 ;
        RECT 985.950 826.950 988.050 829.050 ;
        RECT 991.950 826.950 994.050 829.050 ;
        RECT 982.950 820.950 985.050 823.050 ;
        RECT 974.400 818.400 978.450 819.450 ;
        RECT 973.950 814.950 976.050 817.050 ;
        RECT 967.950 811.950 970.050 814.050 ;
        RECT 969.000 810.450 973.050 811.050 ;
        RECT 968.400 808.950 973.050 810.450 ;
        RECT 968.400 807.600 969.450 808.950 ;
        RECT 974.400 807.600 975.450 814.950 ;
        RECT 977.400 811.050 978.450 818.400 ;
        RECT 976.950 808.950 979.050 811.050 ;
        RECT 982.950 808.950 985.050 811.050 ;
        RECT 968.400 805.350 969.600 807.600 ;
        RECT 974.400 805.350 975.600 807.600 ;
        RECT 967.950 802.950 970.050 805.050 ;
        RECT 970.950 802.950 973.050 805.050 ;
        RECT 973.950 802.950 976.050 805.050 ;
        RECT 976.950 802.950 979.050 805.050 ;
        RECT 971.400 801.900 972.600 802.650 ;
        RECT 977.400 801.900 978.600 802.650 ;
        RECT 970.950 799.800 973.050 801.900 ;
        RECT 976.950 799.800 979.050 801.900 ;
        RECT 961.950 793.950 964.050 796.050 ;
        RECT 961.950 775.950 964.050 778.050 ;
        RECT 962.400 739.050 963.450 775.950 ;
        RECT 967.950 766.950 970.050 769.050 ;
        RECT 968.400 762.600 969.450 766.950 ;
        RECT 971.400 765.450 972.450 799.800 ;
        RECT 973.950 796.950 976.050 799.050 ;
        RECT 979.950 796.950 982.050 799.050 ;
        RECT 974.400 778.050 975.450 796.950 ;
        RECT 973.950 775.950 976.050 778.050 ;
        RECT 980.400 771.450 981.450 796.950 ;
        RECT 983.400 775.050 984.450 808.950 ;
        RECT 982.950 772.950 985.050 775.050 ;
        RECT 980.400 770.400 984.450 771.450 ;
        RECT 971.400 764.400 975.450 765.450 ;
        RECT 974.400 762.600 975.450 764.400 ;
        RECT 968.400 760.350 969.600 762.600 ;
        RECT 974.400 760.350 975.600 762.600 ;
        RECT 967.950 757.950 970.050 760.050 ;
        RECT 970.950 757.950 973.050 760.050 ;
        RECT 973.950 757.950 976.050 760.050 ;
        RECT 976.950 757.950 979.050 760.050 ;
        RECT 971.400 756.000 972.600 757.650 ;
        RECT 970.950 751.950 973.050 756.000 ;
        RECT 977.400 755.400 978.600 757.650 ;
        RECT 977.400 751.050 978.450 755.400 ;
        RECT 964.950 748.950 967.050 751.050 ;
        RECT 976.950 748.950 979.050 751.050 ;
        RECT 961.950 736.950 964.050 739.050 ;
        RECT 958.950 733.950 961.050 736.050 ;
        RECT 965.400 733.050 966.450 748.950 ;
        RECT 983.400 745.050 984.450 770.400 ;
        RECT 973.950 742.950 976.050 745.050 ;
        RECT 982.950 742.950 985.050 745.050 ;
        RECT 961.950 729.000 964.050 733.050 ;
        RECT 964.950 730.950 967.050 733.050 ;
        RECT 962.400 727.350 963.600 729.000 ;
        RECT 967.950 728.100 970.050 730.200 ;
        RECT 974.400 729.600 975.450 742.950 ;
        RECT 976.950 736.950 979.050 739.050 ;
        RECT 977.400 730.050 978.450 736.950 ;
        RECT 979.800 733.950 981.900 736.050 ;
        RECT 982.950 733.950 985.050 736.050 ;
        RECT 968.400 727.350 969.600 728.100 ;
        RECT 974.400 727.350 975.600 729.600 ;
        RECT 976.950 727.950 979.050 730.050 ;
        RECT 961.950 724.950 964.050 727.050 ;
        RECT 964.950 724.950 967.050 727.050 ;
        RECT 967.950 724.950 970.050 727.050 ;
        RECT 970.950 724.950 973.050 727.050 ;
        RECT 973.950 724.950 976.050 727.050 ;
        RECT 965.400 723.900 966.600 724.650 ;
        RECT 964.950 721.800 967.050 723.900 ;
        RECT 971.400 722.400 972.600 724.650 ;
        RECT 971.400 720.450 972.450 722.400 ;
        RECT 976.950 721.950 979.050 724.050 ;
        RECT 971.400 719.400 975.450 720.450 ;
        RECT 967.950 715.950 970.050 718.050 ;
        RECT 964.950 706.950 967.050 709.050 ;
        RECT 940.950 703.950 943.050 706.050 ;
        RECT 955.950 703.950 958.050 706.050 ;
        RECT 937.950 700.950 940.050 703.050 ;
        RECT 937.950 697.800 940.050 699.900 ;
        RECT 934.950 688.950 937.050 691.050 ;
        RECT 899.400 682.350 900.600 684.600 ;
        RECT 904.950 684.000 907.050 688.050 ;
        RECT 910.950 685.950 913.050 688.050 ;
        RECT 922.950 685.950 925.050 688.050 ;
        RECT 931.950 685.950 934.050 688.050 ;
        RECT 938.400 687.450 939.450 697.800 ;
        RECT 956.400 694.050 957.450 703.950 ;
        RECT 955.950 691.950 958.050 694.050 ;
        RECT 965.400 691.050 966.450 706.950 ;
        RECT 968.400 694.050 969.450 715.950 ;
        RECT 967.950 691.950 970.050 694.050 ;
        RECT 955.950 688.800 958.050 690.900 ;
        RECT 958.950 688.950 961.050 691.050 ;
        RECT 964.950 688.950 967.050 691.050 ;
        RECT 935.400 686.400 939.450 687.450 ;
        RECT 905.400 682.350 906.600 684.000 ;
        RECT 895.950 679.950 898.050 682.050 ;
        RECT 898.950 679.950 901.050 682.050 ;
        RECT 901.950 679.950 904.050 682.050 ;
        RECT 904.950 679.950 907.050 682.050 ;
        RECT 890.400 677.400 894.450 678.450 ;
        RECT 887.400 674.400 891.450 675.450 ;
        RECT 890.400 661.050 891.450 674.400 ;
        RECT 889.950 658.950 892.050 661.050 ;
        RECT 877.950 655.950 880.050 658.050 ;
        RECT 889.950 655.800 892.050 657.900 ;
        RECT 871.950 646.950 874.050 652.050 ;
        RECT 874.950 649.950 877.050 652.050 ;
        RECT 880.950 650.100 883.050 652.200 ;
        RECT 886.950 650.100 889.050 652.200 ;
        RECT 890.400 652.050 891.450 655.800 ;
        RECT 881.400 649.350 882.600 650.100 ;
        RECT 887.400 649.350 888.600 650.100 ;
        RECT 889.950 649.950 892.050 652.050 ;
        RECT 877.950 646.950 880.050 649.050 ;
        RECT 880.950 646.950 883.050 649.050 ;
        RECT 883.950 646.950 886.050 649.050 ;
        RECT 886.950 646.950 889.050 649.050 ;
        RECT 871.950 643.800 874.050 645.900 ;
        RECT 874.950 643.950 877.050 646.050 ;
        RECT 878.400 644.400 879.600 646.650 ;
        RECT 884.400 644.400 885.600 646.650 ;
        RECT 868.950 640.950 871.050 643.050 ;
        RECT 872.400 619.050 873.450 643.800 ;
        RECT 871.950 616.950 874.050 619.050 ;
        RECT 868.950 610.950 871.050 613.050 ;
        RECT 865.950 604.950 868.050 607.050 ;
        RECT 869.400 606.600 870.450 610.950 ;
        RECT 875.400 610.200 876.450 643.950 ;
        RECT 878.400 634.050 879.450 644.400 ;
        RECT 884.400 643.050 885.450 644.400 ;
        RECT 889.950 643.950 892.050 646.050 ;
        RECT 883.950 640.950 886.050 643.050 ;
        RECT 877.950 631.950 880.050 634.050 ;
        RECT 880.950 610.950 883.050 613.050 ;
        RECT 874.950 608.100 877.050 610.200 ;
        RECT 869.400 604.350 870.600 606.600 ;
        RECT 874.950 604.950 877.050 607.050 ;
        RECT 875.400 604.350 876.600 604.950 ;
        RECT 868.950 601.950 871.050 604.050 ;
        RECT 871.950 601.950 874.050 604.050 ;
        RECT 874.950 601.950 877.050 604.050 ;
        RECT 872.400 600.900 873.600 601.650 ;
        RECT 871.950 598.800 874.050 600.900 ;
        RECT 871.950 592.950 874.050 595.050 ;
        RECT 862.950 583.950 865.050 586.050 ;
        RECT 853.950 574.950 856.050 577.050 ;
        RECT 859.950 573.000 862.050 577.050 ;
        RECT 860.400 571.350 861.600 573.000 ;
        RECT 865.950 572.100 868.050 574.200 ;
        RECT 872.400 574.050 873.450 592.950 ;
        RECT 877.950 583.950 880.050 586.050 ;
        RECT 866.400 571.350 867.600 572.100 ;
        RECT 871.950 571.950 874.050 574.050 ;
        RECT 874.950 571.950 877.050 574.050 ;
        RECT 853.950 568.950 856.050 571.050 ;
        RECT 859.950 568.950 862.050 571.050 ;
        RECT 862.950 568.950 865.050 571.050 ;
        RECT 865.950 568.950 868.050 571.050 ;
        RECT 868.950 568.950 871.050 571.050 ;
        RECT 845.400 526.350 846.600 527.100 ;
        RECT 850.950 526.950 853.050 529.050 ;
        RECT 838.950 523.950 841.050 526.050 ;
        RECT 841.950 523.950 844.050 526.050 ;
        RECT 844.950 523.950 847.050 526.050 ;
        RECT 847.950 523.950 850.050 526.050 ;
        RECT 842.400 522.900 843.600 523.650 ;
        RECT 841.950 520.800 844.050 522.900 ;
        RECT 848.400 521.400 849.600 523.650 ;
        RECT 832.950 508.950 835.050 511.050 ;
        RECT 848.400 508.050 849.450 521.400 ;
        RECT 850.950 520.950 853.050 523.050 ;
        RECT 847.950 505.950 850.050 508.050 ;
        RECT 841.950 494.100 844.050 496.200 ;
        RECT 842.400 493.350 843.600 494.100 ;
        RECT 838.950 490.950 841.050 493.050 ;
        RECT 841.950 490.950 844.050 493.050 ;
        RECT 844.950 490.950 847.050 493.050 ;
        RECT 839.400 488.400 840.600 490.650 ;
        RECT 845.400 490.050 846.600 490.650 ;
        RECT 845.400 488.400 850.050 490.050 ;
        RECT 839.400 481.050 840.450 488.400 ;
        RECT 846.000 487.950 850.050 488.400 ;
        RECT 851.400 487.050 852.450 520.950 ;
        RECT 844.950 484.950 847.050 487.050 ;
        RECT 850.950 484.950 853.050 487.050 ;
        RECT 838.950 478.950 841.050 481.050 ;
        RECT 839.400 466.050 840.450 478.950 ;
        RECT 841.950 472.950 844.050 475.050 ;
        RECT 838.950 463.950 841.050 466.050 ;
        RECT 799.950 460.950 802.050 463.050 ;
        RECT 829.950 460.950 832.050 463.050 ;
        RECT 823.950 454.950 826.050 457.050 ;
        RECT 832.950 454.950 835.050 457.050 ;
        RECT 797.400 448.350 798.600 450.600 ;
        RECT 817.950 449.100 820.050 451.200 ;
        RECT 824.400 450.600 825.450 454.950 ;
        RECT 818.400 448.350 819.600 449.100 ;
        RECT 824.400 448.350 825.600 450.600 ;
        RECT 793.950 445.950 796.050 448.050 ;
        RECT 796.950 445.950 799.050 448.050 ;
        RECT 808.950 445.950 811.050 448.050 ;
        RECT 814.950 445.950 817.050 448.050 ;
        RECT 817.950 445.950 820.050 448.050 ;
        RECT 820.950 445.950 823.050 448.050 ;
        RECT 823.950 445.950 826.050 448.050 ;
        RECT 787.950 442.950 790.050 445.050 ;
        RECT 794.400 443.400 795.600 445.650 ;
        RECT 775.950 439.950 778.050 442.050 ;
        RECT 781.950 439.950 784.050 442.050 ;
        RECT 745.950 436.950 748.050 439.050 ;
        RECT 736.950 427.950 739.050 430.050 ;
        RECT 734.100 412.950 736.200 415.050 ;
        RECT 737.400 412.950 739.500 415.050 ;
        RECT 742.800 412.950 744.900 415.050 ;
        RECT 734.400 410.400 735.600 412.650 ;
        RECT 743.400 411.900 744.600 412.650 ;
        RECT 730.950 406.950 733.050 409.050 ;
        RECT 715.950 400.950 718.050 403.050 ;
        RECT 716.400 366.900 717.450 400.950 ;
        RECT 734.400 400.050 735.450 410.400 ;
        RECT 742.950 409.800 745.050 411.900 ;
        RECT 739.950 406.950 742.050 409.050 ;
        RECT 733.950 397.950 736.050 400.050 ;
        RECT 727.950 388.950 730.050 391.050 ;
        RECT 728.400 372.600 729.450 388.950 ;
        RECT 734.400 372.600 735.450 397.950 ;
        RECT 728.400 370.350 729.600 372.600 ;
        RECT 734.400 370.350 735.600 372.600 ;
        RECT 724.950 367.950 727.050 370.050 ;
        RECT 727.950 367.950 730.050 370.050 ;
        RECT 730.950 367.950 733.050 370.050 ;
        RECT 733.950 367.950 736.050 370.050 ;
        RECT 715.950 364.800 718.050 366.900 ;
        RECT 721.950 364.950 724.050 367.050 ;
        RECT 725.400 365.400 726.600 367.650 ;
        RECT 731.400 365.400 732.600 367.650 ;
        RECT 722.400 361.050 723.450 364.950 ;
        RECT 721.950 358.950 724.050 361.050 ;
        RECT 703.950 355.950 706.050 358.050 ;
        RECT 712.950 355.950 715.050 358.050 ;
        RECT 700.950 349.950 703.050 352.050 ;
        RECT 704.400 331.050 705.450 355.950 ;
        RECT 715.950 352.950 718.050 355.050 ;
        RECT 716.400 339.600 717.450 352.950 ;
        RECT 716.400 337.350 717.600 339.600 ;
        RECT 712.950 334.950 715.050 337.050 ;
        RECT 715.950 334.950 718.050 337.050 ;
        RECT 718.950 334.950 721.050 337.050 ;
        RECT 706.950 331.800 709.050 333.900 ;
        RECT 713.400 333.000 714.600 334.650 ;
        RECT 719.400 333.900 720.600 334.650 ;
        RECT 703.950 328.950 706.050 331.050 ;
        RECT 697.950 322.950 700.050 325.050 ;
        RECT 697.950 319.800 700.050 321.900 ;
        RECT 685.950 316.950 688.050 319.050 ;
        RECT 686.400 298.050 687.450 316.950 ;
        RECT 691.950 304.950 694.050 307.050 ;
        RECT 688.950 298.950 691.050 301.050 ;
        RECT 685.950 295.950 688.050 298.050 ;
        RECT 683.400 293.400 687.450 294.450 ;
        RECT 670.950 289.950 673.050 292.050 ;
        RECT 673.950 289.950 676.050 292.050 ;
        RECT 676.950 289.950 679.050 292.050 ;
        RECT 679.950 289.950 682.050 292.050 ;
        RECT 674.400 288.900 675.600 289.650 ;
        RECT 680.400 289.050 681.600 289.650 ;
        RECT 673.950 286.800 676.050 288.900 ;
        RECT 680.400 287.400 685.050 289.050 ;
        RECT 681.000 286.950 685.050 287.400 ;
        RECT 681.000 285.900 684.000 286.050 ;
        RECT 681.000 285.450 685.050 285.900 ;
        RECT 680.400 283.950 685.050 285.450 ;
        RECT 670.950 280.950 673.050 283.050 ;
        RECT 667.950 259.950 670.050 262.050 ;
        RECT 664.950 250.950 667.050 253.050 ;
        RECT 668.400 250.050 669.450 259.950 ;
        RECT 667.950 247.950 670.050 250.050 ;
        RECT 661.950 244.950 664.050 247.050 ;
        RECT 671.400 244.050 672.450 280.950 ;
        RECT 680.400 274.050 681.450 283.950 ;
        RECT 682.950 283.800 685.050 283.950 ;
        RECT 686.400 283.050 687.450 293.400 ;
        RECT 689.400 289.050 690.450 298.950 ;
        RECT 692.400 295.050 693.450 304.950 ;
        RECT 698.400 301.050 699.450 319.800 ;
        RECT 697.950 298.950 700.050 301.050 ;
        RECT 703.950 298.950 706.050 301.050 ;
        RECT 691.950 292.950 694.050 295.050 ;
        RECT 697.950 294.000 700.050 297.900 ;
        RECT 704.400 295.050 705.450 298.950 ;
        RECT 698.400 292.350 699.600 294.000 ;
        RECT 703.950 292.950 706.050 295.050 ;
        RECT 694.950 289.950 697.050 292.050 ;
        RECT 697.950 289.950 700.050 292.050 ;
        RECT 700.950 289.950 703.050 292.050 ;
        RECT 688.950 286.950 691.050 289.050 ;
        RECT 695.400 287.400 696.600 289.650 ;
        RECT 701.400 288.900 702.600 289.650 ;
        RECT 695.400 283.050 696.450 287.400 ;
        RECT 700.950 286.800 703.050 288.900 ;
        RECT 703.950 286.950 706.050 289.050 ;
        RECT 685.950 280.950 688.050 283.050 ;
        RECT 694.950 280.950 697.050 283.050 ;
        RECT 685.950 274.950 688.050 277.050 ;
        RECT 679.950 271.950 682.050 274.050 ;
        RECT 680.400 261.600 681.450 271.950 ;
        RECT 680.400 259.350 681.600 261.600 ;
        RECT 676.950 256.950 679.050 259.050 ;
        RECT 679.950 256.950 682.050 259.050 ;
        RECT 677.400 255.900 678.600 256.650 ;
        RECT 686.400 255.900 687.450 274.950 ;
        RECT 688.950 271.950 691.050 274.050 ;
        RECT 676.950 253.800 679.050 255.900 ;
        RECT 685.950 253.800 688.050 255.900 ;
        RECT 676.950 250.650 679.050 252.750 ;
        RECT 670.950 241.950 673.050 244.050 ;
        RECT 652.950 238.950 655.050 241.050 ;
        RECT 658.950 238.950 661.050 241.050 ;
        RECT 673.950 238.950 676.050 241.050 ;
        RECT 649.950 226.950 652.050 229.050 ;
        RECT 650.400 208.050 651.450 226.950 ;
        RECT 649.950 205.950 652.050 208.050 ;
        RECT 646.950 202.950 649.050 205.050 ;
        RECT 653.400 202.050 654.450 238.950 ;
        RECT 667.950 226.950 670.050 229.050 ;
        RECT 661.950 215.100 664.050 217.200 ;
        RECT 668.400 216.600 669.450 226.950 ;
        RECT 662.400 214.350 663.600 215.100 ;
        RECT 668.400 214.350 669.600 216.600 ;
        RECT 658.950 211.950 661.050 214.050 ;
        RECT 661.950 211.950 664.050 214.050 ;
        RECT 664.950 211.950 667.050 214.050 ;
        RECT 667.950 211.950 670.050 214.050 ;
        RECT 659.400 209.400 660.600 211.650 ;
        RECT 665.400 210.900 666.600 211.650 ;
        RECT 674.400 211.050 675.450 238.950 ;
        RECT 655.950 202.950 658.050 205.050 ;
        RECT 652.950 199.950 655.050 202.050 ;
        RECT 640.950 187.950 643.050 190.050 ;
        RECT 652.950 187.950 655.050 190.050 ;
        RECT 634.950 183.450 637.050 184.200 ;
        RECT 632.400 182.400 637.050 183.450 ;
        RECT 634.950 182.100 637.050 182.400 ;
        RECT 641.400 183.600 642.450 187.950 ;
        RECT 635.400 181.350 636.600 182.100 ;
        RECT 641.400 181.350 642.600 183.600 ;
        RECT 646.950 182.100 649.050 184.200 ;
        RECT 647.400 181.350 648.600 182.100 ;
        RECT 634.950 178.950 637.050 181.050 ;
        RECT 637.950 178.950 640.050 181.050 ;
        RECT 640.950 178.950 643.050 181.050 ;
        RECT 643.950 178.950 646.050 181.050 ;
        RECT 646.950 178.950 649.050 181.050 ;
        RECT 638.400 177.000 639.600 178.650 ;
        RECT 644.400 177.000 645.600 178.650 ;
        RECT 637.950 172.950 640.050 177.000 ;
        RECT 643.950 172.950 646.050 177.000 ;
        RECT 649.950 175.950 652.050 178.050 ;
        RECT 622.950 169.950 625.050 172.050 ;
        RECT 644.400 160.050 645.450 172.950 ;
        RECT 650.400 166.050 651.450 175.950 ;
        RECT 649.950 163.950 652.050 166.050 ;
        RECT 653.400 160.050 654.450 187.950 ;
        RECT 656.400 184.200 657.450 202.950 ;
        RECT 659.400 199.050 660.450 209.400 ;
        RECT 664.950 208.800 667.050 210.900 ;
        RECT 673.950 205.950 676.050 211.050 ;
        RECT 658.950 196.950 661.050 199.050 ;
        RECT 658.950 190.950 661.050 193.050 ;
        RECT 655.950 178.950 658.050 184.200 ;
        RECT 655.950 172.950 658.050 177.900 ;
        RECT 659.400 177.450 660.450 190.950 ;
        RECT 677.400 190.050 678.450 250.650 ;
        RECT 686.400 235.050 687.450 253.800 ;
        RECT 685.950 232.950 688.050 235.050 ;
        RECT 679.950 226.950 682.050 229.050 ;
        RECT 676.950 189.450 679.050 190.050 ;
        RECT 674.400 188.400 679.050 189.450 ;
        RECT 674.400 181.050 675.450 188.400 ;
        RECT 676.950 187.950 679.050 188.400 ;
        RECT 680.400 184.200 681.450 226.950 ;
        RECT 689.400 217.200 690.450 271.950 ;
        RECT 701.400 270.450 702.450 286.800 ;
        RECT 704.400 274.050 705.450 286.950 ;
        RECT 703.950 271.950 706.050 274.050 ;
        RECT 701.400 269.400 705.450 270.450 ;
        RECT 697.950 260.100 700.050 262.200 ;
        RECT 698.400 259.350 699.600 260.100 ;
        RECT 694.950 256.950 697.050 259.050 ;
        RECT 697.950 256.950 700.050 259.050 ;
        RECT 695.400 254.400 696.600 256.650 ;
        RECT 695.400 232.050 696.450 254.400 ;
        RECT 700.950 253.950 703.050 256.050 ;
        RECT 701.400 250.050 702.450 253.950 ;
        RECT 697.950 247.950 700.050 250.050 ;
        RECT 700.950 247.950 703.050 250.050 ;
        RECT 698.400 241.050 699.450 247.950 ;
        RECT 697.950 238.950 700.050 241.050 ;
        RECT 704.400 238.050 705.450 269.400 ;
        RECT 707.400 253.050 708.450 331.800 ;
        RECT 712.950 328.950 715.050 333.000 ;
        RECT 718.950 331.800 721.050 333.900 ;
        RECT 718.950 325.950 721.050 330.750 ;
        RECT 725.400 328.050 726.450 365.400 ;
        RECT 731.400 358.050 732.450 365.400 ;
        RECT 730.950 355.950 733.050 358.050 ;
        RECT 736.950 346.950 739.050 349.050 ;
        RECT 727.950 343.950 730.050 346.050 ;
        RECT 724.950 325.950 727.050 328.050 ;
        RECT 728.400 319.050 729.450 343.950 ;
        RECT 737.400 339.600 738.450 346.950 ;
        RECT 740.400 343.050 741.450 406.950 ;
        RECT 743.400 399.450 744.450 409.800 ;
        RECT 746.400 403.050 747.450 436.950 ;
        RECT 769.950 427.950 772.050 430.050 ;
        RECT 758.100 412.950 760.200 415.050 ;
        RECT 763.500 412.950 765.600 415.050 ;
        RECT 766.800 412.950 768.900 415.050 ;
        RECT 758.400 410.400 759.600 412.650 ;
        RECT 767.400 411.900 768.600 412.650 ;
        RECT 745.950 400.950 748.050 403.050 ;
        RECT 743.400 398.400 747.450 399.450 ;
        RECT 742.950 376.950 745.050 379.050 ;
        RECT 743.400 364.050 744.450 376.950 ;
        RECT 746.400 373.050 747.450 398.400 ;
        RECT 758.400 394.050 759.450 410.400 ;
        RECT 766.950 409.800 769.050 411.900 ;
        RECT 757.950 391.950 760.050 394.050 ;
        RECT 745.950 370.950 748.050 373.050 ;
        RECT 751.950 371.100 754.050 373.200 ;
        RECT 758.400 372.450 759.600 372.600 ;
        RECT 758.400 371.400 765.450 372.450 ;
        RECT 752.400 370.350 753.600 371.100 ;
        RECT 758.400 370.350 759.600 371.400 ;
        RECT 748.950 367.950 751.050 370.050 ;
        RECT 751.950 367.950 754.050 370.050 ;
        RECT 754.950 367.950 757.050 370.050 ;
        RECT 757.950 367.950 760.050 370.050 ;
        RECT 749.400 365.400 750.600 367.650 ;
        RECT 755.400 365.400 756.600 367.650 ;
        RECT 742.950 361.950 745.050 364.050 ;
        RECT 749.400 363.450 750.450 365.400 ;
        RECT 749.400 362.400 753.450 363.450 ;
        RECT 748.950 358.950 751.050 361.050 ;
        RECT 739.950 340.950 742.050 343.050 ;
        RECT 745.950 340.950 748.050 343.050 ;
        RECT 737.400 337.350 738.600 339.600 ;
        RECT 733.950 334.950 736.050 337.050 ;
        RECT 736.950 334.950 739.050 337.050 ;
        RECT 739.950 334.950 742.050 337.050 ;
        RECT 734.400 333.000 735.600 334.650 ;
        RECT 733.950 330.450 736.050 333.000 ;
        RECT 731.400 329.400 736.050 330.450 ;
        RECT 727.950 316.950 730.050 319.050 ;
        RECT 724.950 313.950 727.050 316.050 ;
        RECT 725.400 310.050 726.450 313.950 ;
        RECT 724.950 307.950 727.050 310.050 ;
        RECT 728.400 301.050 729.450 316.950 ;
        RECT 727.950 298.950 730.050 301.050 ;
        RECT 712.950 295.950 715.050 298.050 ;
        RECT 709.950 293.100 712.050 295.200 ;
        RECT 710.400 283.050 711.450 293.100 ;
        RECT 709.950 280.950 712.050 283.050 ;
        RECT 710.400 262.050 711.450 280.950 ;
        RECT 713.400 280.050 714.450 295.950 ;
        RECT 721.950 293.100 724.050 295.200 ;
        RECT 727.950 294.000 730.050 297.900 ;
        RECT 731.400 295.050 732.450 329.400 ;
        RECT 733.950 328.950 736.050 329.400 ;
        RECT 733.950 325.800 736.050 327.900 ;
        RECT 722.400 292.350 723.600 293.100 ;
        RECT 728.400 292.350 729.600 294.000 ;
        RECT 730.950 292.950 733.050 295.050 ;
        RECT 718.950 289.950 721.050 292.050 ;
        RECT 721.950 289.950 724.050 292.050 ;
        RECT 724.950 289.950 727.050 292.050 ;
        RECT 727.950 289.950 730.050 292.050 ;
        RECT 719.400 288.900 720.600 289.650 ;
        RECT 718.950 286.800 721.050 288.900 ;
        RECT 725.400 287.400 726.600 289.650 ;
        RECT 734.400 288.450 735.450 325.800 ;
        RECT 736.950 322.950 739.050 325.050 ;
        RECT 737.400 310.050 738.450 322.950 ;
        RECT 746.400 315.450 747.450 340.950 ;
        RECT 743.400 314.400 747.450 315.450 ;
        RECT 736.950 307.950 739.050 310.050 ;
        RECT 736.950 295.950 739.050 301.050 ;
        RECT 743.400 300.450 744.450 314.400 ;
        RECT 745.950 307.950 748.050 310.050 ;
        RECT 740.400 299.400 744.450 300.450 ;
        RECT 740.400 295.050 741.450 299.400 ;
        RECT 746.400 298.050 747.450 307.950 ;
        RECT 745.950 295.950 748.050 298.050 ;
        RECT 736.950 292.800 739.050 294.900 ;
        RECT 739.950 292.950 742.050 295.050 ;
        RECT 746.400 294.600 747.450 295.950 ;
        RECT 749.400 295.050 750.450 358.950 ;
        RECT 752.400 340.050 753.450 362.400 ;
        RECT 755.400 361.050 756.450 365.400 ;
        RECT 760.950 364.950 763.050 367.050 ;
        RECT 754.950 358.950 757.050 361.050 ;
        RECT 754.950 346.950 757.050 349.050 ;
        RECT 751.950 337.950 754.050 340.050 ;
        RECT 755.400 339.600 756.450 346.950 ;
        RECT 761.400 340.050 762.450 364.950 ;
        RECT 755.400 337.350 756.600 339.600 ;
        RECT 760.950 337.950 763.050 340.050 ;
        RECT 754.950 334.950 757.050 337.050 ;
        RECT 757.950 334.950 760.050 337.050 ;
        RECT 751.950 331.950 754.050 334.050 ;
        RECT 758.400 332.400 759.600 334.650 ;
        RECT 752.400 316.050 753.450 331.950 ;
        RECT 758.400 322.050 759.450 332.400 ;
        RECT 757.950 319.950 760.050 322.050 ;
        RECT 751.950 313.950 754.050 316.050 ;
        RECT 752.400 295.050 753.450 313.950 ;
        RECT 764.400 313.050 765.450 371.400 ;
        RECT 766.950 364.800 769.050 366.900 ;
        RECT 767.400 358.050 768.450 364.800 ;
        RECT 766.950 355.950 769.050 358.050 ;
        RECT 770.400 357.450 771.450 427.950 ;
        RECT 776.400 394.050 777.450 439.950 ;
        RECT 784.950 424.950 787.050 427.050 ;
        RECT 785.400 417.600 786.450 424.950 ;
        RECT 785.400 415.350 786.600 417.600 ;
        RECT 781.950 412.950 784.050 415.050 ;
        RECT 784.950 412.950 787.050 415.050 ;
        RECT 787.950 412.950 790.050 415.050 ;
        RECT 782.400 411.900 783.600 412.650 ;
        RECT 781.950 409.800 784.050 411.900 ;
        RECT 788.400 410.400 789.600 412.650 ;
        RECT 775.950 391.950 778.050 394.050 ;
        RECT 775.950 376.950 778.050 379.050 ;
        RECT 776.400 372.600 777.450 376.950 ;
        RECT 782.400 372.600 783.450 409.800 ;
        RECT 788.400 400.050 789.450 410.400 ;
        RECT 794.400 400.050 795.450 443.400 ;
        RECT 809.400 439.050 810.450 445.950 ;
        RECT 815.400 443.400 816.600 445.650 ;
        RECT 821.400 443.400 822.600 445.650 ;
        RECT 833.400 444.900 834.450 454.950 ;
        RECT 842.400 450.600 843.450 472.950 ;
        RECT 845.400 472.050 846.450 484.950 ;
        RECT 844.950 469.950 847.050 472.050 ;
        RECT 854.400 457.050 855.450 568.950 ;
        RECT 863.400 567.900 864.600 568.650 ;
        RECT 862.950 565.800 865.050 567.900 ;
        RECT 869.400 566.400 870.600 568.650 ;
        RECT 869.400 556.050 870.450 566.400 ;
        RECT 868.950 553.950 871.050 556.050 ;
        RECT 875.400 535.050 876.450 571.950 ;
        RECT 868.950 532.950 871.050 535.050 ;
        RECT 874.950 532.950 877.050 535.050 ;
        RECT 856.950 527.100 859.050 529.200 ;
        RECT 862.950 527.100 865.050 529.200 ;
        RECT 869.400 528.600 870.450 532.950 ;
        RECT 857.400 487.050 858.450 527.100 ;
        RECT 863.400 526.350 864.600 527.100 ;
        RECT 869.400 526.350 870.600 528.600 ;
        RECT 862.950 523.950 865.050 526.050 ;
        RECT 865.950 523.950 868.050 526.050 ;
        RECT 868.950 523.950 871.050 526.050 ;
        RECT 871.950 523.950 874.050 526.050 ;
        RECT 866.400 521.400 867.600 523.650 ;
        RECT 872.400 523.050 873.600 523.650 ;
        RECT 872.400 521.400 877.050 523.050 ;
        RECT 866.400 514.050 867.450 521.400 ;
        RECT 873.000 520.950 877.050 521.400 ;
        RECT 874.950 517.800 877.050 519.900 ;
        RECT 868.950 514.950 871.050 517.050 ;
        RECT 865.950 511.950 868.050 514.050 ;
        RECT 869.400 508.050 870.450 514.950 ;
        RECT 871.950 508.950 874.050 511.050 ;
        RECT 868.950 505.950 871.050 508.050 ;
        RECT 872.400 502.050 873.450 508.950 ;
        RECT 875.400 502.050 876.450 517.800 ;
        RECT 878.400 517.050 879.450 583.950 ;
        RECT 881.400 523.050 882.450 610.950 ;
        RECT 884.400 607.050 885.450 640.950 ;
        RECT 890.400 634.050 891.450 643.950 ;
        RECT 893.400 643.050 894.450 677.400 ;
        RECT 896.400 677.400 897.600 679.650 ;
        RECT 902.400 677.400 903.600 679.650 ;
        RECT 911.400 678.450 912.450 685.950 ;
        RECT 913.950 682.950 916.050 685.050 ;
        RECT 919.950 683.100 922.050 685.200 ;
        RECT 928.950 683.100 931.050 685.200 ;
        RECT 908.400 677.400 912.450 678.450 ;
        RECT 896.400 670.050 897.450 677.400 ;
        RECT 895.950 667.950 898.050 670.050 ;
        RECT 895.950 658.950 898.050 661.050 ;
        RECT 892.950 640.950 895.050 643.050 ;
        RECT 889.950 631.950 892.050 634.050 ;
        RECT 890.400 610.200 891.450 631.950 ;
        RECT 896.400 625.050 897.450 658.950 ;
        RECT 902.400 658.050 903.450 677.400 ;
        RECT 904.950 658.950 907.050 661.050 ;
        RECT 901.950 655.950 904.050 658.050 ;
        RECT 898.950 649.950 901.050 652.050 ;
        RECT 905.400 651.600 906.450 658.950 ;
        RECT 908.400 655.050 909.450 677.400 ;
        RECT 914.400 675.450 915.450 682.950 ;
        RECT 920.400 682.350 921.600 683.100 ;
        RECT 919.950 679.950 922.050 682.050 ;
        RECT 922.950 679.950 925.050 682.050 ;
        RECT 923.400 678.900 924.600 679.650 ;
        RECT 922.950 676.800 925.050 678.900 ;
        RECT 925.950 676.950 928.050 679.050 ;
        RECT 914.400 674.400 921.450 675.450 ;
        RECT 916.950 670.950 919.050 673.050 ;
        RECT 910.950 655.950 913.050 658.050 ;
        RECT 907.950 652.950 910.050 655.050 ;
        RECT 911.400 651.600 912.450 655.950 ;
        RECT 917.400 652.050 918.450 670.950 ;
        RECT 920.400 669.450 921.450 674.400 ;
        RECT 923.400 673.050 924.450 676.800 ;
        RECT 922.950 670.950 925.050 673.050 ;
        RECT 926.400 669.450 927.450 676.950 ;
        RECT 920.400 668.400 927.450 669.450 ;
        RECT 929.400 667.050 930.450 683.100 ;
        RECT 932.400 679.050 933.450 685.950 ;
        RECT 935.400 682.050 936.450 686.400 ;
        RECT 940.950 683.100 943.050 685.200 ;
        RECT 946.950 684.000 949.050 688.050 ;
        RECT 941.400 682.350 942.600 683.100 ;
        RECT 947.400 682.350 948.600 684.000 ;
        RECT 934.950 679.950 937.050 682.050 ;
        RECT 940.950 679.950 943.050 682.050 ;
        RECT 943.950 679.950 946.050 682.050 ;
        RECT 946.950 679.950 949.050 682.050 ;
        RECT 949.950 679.950 952.050 682.050 ;
        RECT 931.950 676.950 934.050 679.050 ;
        RECT 934.950 675.450 937.050 678.900 ;
        RECT 932.400 675.000 937.050 675.450 ;
        RECT 944.400 677.400 945.600 679.650 ;
        RECT 950.400 679.050 951.600 679.650 ;
        RECT 950.400 677.400 955.050 679.050 ;
        RECT 932.400 674.400 936.450 675.000 ;
        RECT 919.950 664.950 922.050 667.050 ;
        RECT 928.950 664.950 931.050 667.050 ;
        RECT 899.400 631.050 900.450 649.950 ;
        RECT 905.400 649.350 906.600 651.600 ;
        RECT 911.400 649.350 912.600 651.600 ;
        RECT 916.950 649.950 919.050 652.050 ;
        RECT 904.950 646.950 907.050 649.050 ;
        RECT 907.950 646.950 910.050 649.050 ;
        RECT 910.950 646.950 913.050 649.050 ;
        RECT 913.950 646.950 916.050 649.050 ;
        RECT 908.400 645.000 909.600 646.650 ;
        RECT 914.400 645.900 915.600 646.650 ;
        RECT 907.950 640.950 910.050 645.000 ;
        RECT 913.950 643.800 916.050 645.900 ;
        RECT 916.950 642.450 919.050 643.050 ;
        RECT 920.400 642.450 921.450 664.950 ;
        RECT 932.400 663.450 933.450 674.400 ;
        RECT 929.400 662.400 933.450 663.450 ;
        RECT 922.950 658.950 925.050 661.050 ;
        RECT 916.950 641.400 921.450 642.450 ;
        RECT 916.950 640.950 919.050 641.400 ;
        RECT 907.950 637.800 910.050 639.900 ;
        RECT 898.950 628.950 901.050 631.050 ;
        RECT 895.950 622.950 898.050 625.050 ;
        RECT 889.950 608.100 892.050 610.200 ;
        RECT 883.950 604.950 886.050 607.050 ;
        RECT 889.950 604.950 892.050 607.050 ;
        RECT 895.950 606.000 898.050 610.050 ;
        RECT 884.400 601.050 885.450 604.950 ;
        RECT 890.400 604.350 891.600 604.950 ;
        RECT 896.400 604.350 897.600 606.000 ;
        RECT 889.950 601.950 892.050 604.050 ;
        RECT 892.950 601.950 895.050 604.050 ;
        RECT 895.950 601.950 898.050 604.050 ;
        RECT 898.950 601.950 901.050 604.050 ;
        RECT 904.950 601.950 907.050 604.050 ;
        RECT 883.950 598.950 886.050 601.050 ;
        RECT 886.950 595.950 889.050 601.050 ;
        RECT 893.400 600.000 894.600 601.650 ;
        RECT 899.400 600.450 900.600 601.650 ;
        RECT 892.950 595.950 895.050 600.000 ;
        RECT 899.400 599.400 903.450 600.450 ;
        RECT 898.950 595.950 901.050 598.050 ;
        RECT 889.950 577.950 892.050 580.050 ;
        RECT 890.400 573.600 891.450 577.950 ;
        RECT 890.400 571.350 891.600 573.600 ;
        RECT 886.950 568.950 889.050 571.050 ;
        RECT 889.950 568.950 892.050 571.050 ;
        RECT 892.950 568.950 895.050 571.050 ;
        RECT 883.950 565.950 886.050 568.050 ;
        RECT 887.400 567.900 888.600 568.650 ;
        RECT 884.400 529.050 885.450 565.950 ;
        RECT 886.950 565.800 889.050 567.900 ;
        RECT 893.400 566.400 894.600 568.650 ;
        RECT 899.400 568.050 900.450 595.950 ;
        RECT 902.400 589.050 903.450 599.400 ;
        RECT 905.400 598.050 906.450 601.950 ;
        RECT 904.950 595.950 907.050 598.050 ;
        RECT 901.950 586.950 904.050 589.050 ;
        RECT 908.400 583.050 909.450 637.800 ;
        RECT 910.950 631.950 913.050 634.050 ;
        RECT 911.400 592.050 912.450 631.950 ;
        RECT 913.950 616.950 916.050 619.050 ;
        RECT 914.400 597.450 915.450 616.950 ;
        RECT 917.400 606.600 918.450 640.950 ;
        RECT 923.400 616.050 924.450 658.950 ;
        RECT 929.400 655.050 930.450 662.400 ;
        RECT 934.950 658.950 937.050 661.050 ;
        RECT 931.950 655.950 934.050 658.050 ;
        RECT 928.950 652.950 931.050 655.050 ;
        RECT 932.400 651.600 933.450 655.950 ;
        RECT 935.400 655.050 936.450 658.950 ;
        RECT 944.400 658.050 945.450 677.400 ;
        RECT 951.000 676.950 955.050 677.400 ;
        RECT 946.950 673.950 949.050 676.050 ;
        RECT 943.950 655.950 946.050 658.050 ;
        RECT 934.950 652.950 937.050 655.050 ;
        RECT 932.400 649.350 933.600 651.600 ;
        RECT 937.950 650.100 940.050 652.200 ;
        RECT 938.400 649.350 939.600 650.100 ;
        RECT 943.950 649.950 946.050 652.050 ;
        RECT 928.950 646.950 931.050 649.050 ;
        RECT 931.950 646.950 934.050 649.050 ;
        RECT 934.950 646.950 937.050 649.050 ;
        RECT 937.950 646.950 940.050 649.050 ;
        RECT 925.950 643.950 928.050 646.050 ;
        RECT 929.400 645.900 930.600 646.650 ;
        RECT 926.400 640.050 927.450 643.950 ;
        RECT 928.950 643.800 931.050 645.900 ;
        RECT 935.400 645.000 936.600 646.650 ;
        RECT 934.950 640.950 937.050 645.000 ;
        RECT 940.950 643.950 943.050 646.050 ;
        RECT 937.950 640.950 940.050 643.050 ;
        RECT 925.950 637.950 928.050 640.050 ;
        RECT 931.950 625.950 934.050 628.050 ;
        RECT 922.950 613.950 925.050 616.050 ;
        RECT 928.950 613.950 931.050 616.050 ;
        RECT 925.950 610.950 928.050 613.050 ;
        RECT 926.400 606.600 927.450 610.950 ;
        RECT 917.400 604.350 918.600 606.600 ;
        RECT 926.400 604.350 927.600 606.600 ;
        RECT 917.100 601.950 919.200 604.050 ;
        RECT 920.400 601.950 922.500 604.050 ;
        RECT 925.800 601.950 927.900 604.050 ;
        RECT 920.400 600.000 921.600 601.650 ;
        RECT 914.400 596.400 918.450 597.450 ;
        RECT 910.950 589.950 913.050 592.050 ;
        RECT 901.950 580.950 904.050 583.050 ;
        RECT 907.950 580.950 910.050 583.050 ;
        RECT 887.400 532.050 888.450 565.800 ;
        RECT 889.950 538.950 892.050 541.050 ;
        RECT 886.950 529.950 889.050 532.050 ;
        RECT 883.950 526.950 886.050 529.050 ;
        RECT 890.400 528.600 891.450 538.950 ;
        RECT 893.400 532.050 894.450 566.400 ;
        RECT 898.950 565.950 901.050 568.050 ;
        RECT 902.400 567.450 903.450 580.950 ;
        RECT 910.950 572.100 913.050 574.200 ;
        RECT 911.400 571.350 912.600 572.100 ;
        RECT 907.950 568.950 910.050 571.050 ;
        RECT 910.950 568.950 913.050 571.050 ;
        RECT 902.400 566.400 906.450 567.450 ;
        RECT 905.400 532.050 906.450 566.400 ;
        RECT 908.400 566.400 909.600 568.650 ;
        RECT 908.400 556.050 909.450 566.400 ;
        RECT 913.950 565.950 916.050 568.050 ;
        RECT 914.400 562.050 915.450 565.950 ;
        RECT 913.950 559.950 916.050 562.050 ;
        RECT 907.950 553.950 910.050 556.050 ;
        RECT 908.400 541.050 909.450 553.950 ;
        RECT 917.400 553.050 918.450 596.400 ;
        RECT 919.950 595.950 922.050 600.000 ;
        RECT 929.400 595.050 930.450 613.950 ;
        RECT 928.950 592.950 931.050 595.050 ;
        RECT 919.950 589.950 922.050 592.050 ;
        RECT 920.400 565.050 921.450 589.950 ;
        RECT 922.950 586.950 925.050 589.050 ;
        RECT 923.400 574.050 924.450 586.950 ;
        RECT 922.950 571.950 925.050 574.050 ;
        RECT 929.400 573.600 930.450 592.950 ;
        RECT 932.400 580.050 933.450 625.950 ;
        RECT 938.400 616.050 939.450 640.950 ;
        RECT 941.400 628.050 942.450 643.950 ;
        RECT 944.400 642.450 945.450 649.950 ;
        RECT 947.400 646.050 948.450 673.950 ;
        RECT 952.950 667.950 955.050 670.050 ;
        RECT 949.950 664.950 952.050 667.050 ;
        RECT 946.950 643.950 949.050 646.050 ;
        RECT 944.400 641.400 948.450 642.450 ;
        RECT 943.950 634.950 946.050 640.050 ;
        RECT 940.950 625.950 943.050 628.050 ;
        RECT 937.950 613.950 940.050 616.050 ;
        RECT 947.400 610.200 948.450 641.400 ;
        RECT 950.400 640.050 951.450 664.950 ;
        RECT 953.400 652.050 954.450 667.950 ;
        RECT 956.400 661.050 957.450 688.800 ;
        RECT 959.400 682.050 960.450 688.950 ;
        RECT 968.400 684.600 969.450 691.950 ;
        RECT 968.400 682.350 969.600 684.600 ;
        RECT 958.950 679.950 961.050 682.050 ;
        RECT 964.950 679.950 967.050 682.050 ;
        RECT 967.950 679.950 970.050 682.050 ;
        RECT 958.950 676.800 961.050 678.900 ;
        RECT 965.400 677.400 966.600 679.650 ;
        RECT 974.400 679.050 975.450 719.400 ;
        RECT 959.400 667.050 960.450 676.800 ;
        RECT 958.950 664.950 961.050 667.050 ;
        RECT 955.950 658.950 958.050 661.050 ;
        RECT 952.950 649.950 955.050 652.050 ;
        RECT 959.400 651.600 960.450 664.950 ;
        RECT 965.400 664.050 966.450 677.400 ;
        RECT 973.950 676.950 976.050 679.050 ;
        RECT 970.950 673.950 973.050 676.050 ;
        RECT 971.400 664.050 972.450 673.950 ;
        RECT 973.950 670.950 976.050 673.050 ;
        RECT 964.950 661.950 967.050 664.050 ;
        RECT 970.950 661.950 973.050 664.050 ;
        RECT 966.000 660.600 970.050 661.050 ;
        RECT 965.400 658.950 970.050 660.600 ;
        RECT 965.400 655.050 966.450 658.950 ;
        RECT 967.950 655.800 970.050 657.900 ;
        RECT 959.400 649.350 960.600 651.600 ;
        RECT 964.950 651.000 967.050 655.050 ;
        RECT 968.400 652.050 969.450 655.800 ;
        RECT 965.400 649.350 966.600 651.000 ;
        RECT 967.950 649.950 970.050 652.050 ;
        RECT 955.950 646.950 958.050 649.050 ;
        RECT 958.950 646.950 961.050 649.050 ;
        RECT 961.950 646.950 964.050 649.050 ;
        RECT 964.950 646.950 967.050 649.050 ;
        RECT 952.950 643.950 955.050 646.050 ;
        RECT 956.400 645.000 957.600 646.650 ;
        RECT 953.400 640.050 954.450 643.950 ;
        RECT 955.950 640.950 958.050 645.000 ;
        RECT 962.400 644.400 963.600 646.650 ;
        RECT 958.950 640.950 961.050 643.050 ;
        RECT 962.400 642.450 963.450 644.400 ;
        RECT 962.400 641.400 966.450 642.450 ;
        RECT 949.950 637.950 952.050 640.050 ;
        RECT 952.950 637.950 955.050 640.050 ;
        RECT 949.950 631.950 952.050 636.900 ;
        RECT 959.400 636.450 960.450 640.950 ;
        RECT 956.400 635.400 960.450 636.450 ;
        RECT 934.950 607.950 937.050 610.050 ;
        RECT 946.950 608.100 949.050 610.200 ;
        RECT 935.400 580.050 936.450 607.950 ;
        RECT 940.950 605.100 943.050 607.200 ;
        RECT 941.400 604.350 942.600 605.100 ;
        RECT 946.950 604.950 949.050 607.050 ;
        RECT 947.400 604.350 948.600 604.950 ;
        RECT 940.950 601.950 943.050 604.050 ;
        RECT 943.950 601.950 946.050 604.050 ;
        RECT 946.950 601.950 949.050 604.050 ;
        RECT 949.950 601.950 952.050 604.050 ;
        RECT 937.950 598.950 940.050 601.050 ;
        RECT 944.400 599.400 945.600 601.650 ;
        RECT 950.400 599.400 951.600 601.650 ;
        RECT 956.400 601.050 957.450 635.400 ;
        RECT 961.950 631.950 964.050 634.050 ;
        RECT 958.950 628.950 961.050 631.050 ;
        RECT 938.400 589.050 939.450 598.950 ;
        RECT 944.400 597.450 945.450 599.400 ;
        RECT 941.400 597.000 945.450 597.450 ;
        RECT 940.950 596.400 945.450 597.000 ;
        RECT 940.950 595.050 943.050 596.400 ;
        RECT 940.800 594.000 943.050 595.050 ;
        RECT 940.800 592.950 942.900 594.000 ;
        RECT 943.950 592.950 946.050 595.050 ;
        RECT 937.950 586.950 940.050 589.050 ;
        RECT 931.800 577.950 933.900 580.050 ;
        RECT 934.950 577.950 937.050 580.050 ;
        RECT 940.950 577.950 943.050 580.050 ;
        RECT 929.400 571.350 930.600 573.600 ;
        RECT 934.950 572.100 937.050 574.200 ;
        RECT 935.400 571.350 936.600 572.100 ;
        RECT 925.950 568.950 928.050 571.050 ;
        RECT 928.950 568.950 931.050 571.050 ;
        RECT 931.950 568.950 934.050 571.050 ;
        RECT 934.950 568.950 937.050 571.050 ;
        RECT 926.400 567.900 927.600 568.650 ;
        RECT 925.950 565.800 928.050 567.900 ;
        RECT 932.400 566.400 933.600 568.650 ;
        RECT 932.400 565.050 933.450 566.400 ;
        RECT 937.950 565.950 940.050 568.050 ;
        RECT 919.950 562.950 922.050 565.050 ;
        RECT 931.950 562.950 934.050 565.050 ;
        RECT 932.400 559.050 933.450 562.950 ;
        RECT 938.400 561.450 939.450 565.950 ;
        RECT 935.400 560.400 939.450 561.450 ;
        RECT 925.950 556.950 928.050 559.050 ;
        RECT 931.950 556.950 934.050 559.050 ;
        RECT 916.950 550.950 919.050 553.050 ;
        RECT 907.950 538.950 910.050 541.050 ;
        RECT 913.950 538.950 916.050 541.050 ;
        RECT 892.950 529.950 895.050 532.050 ;
        RECT 904.950 529.950 907.050 532.050 ;
        RECT 890.400 526.350 891.600 528.600 ;
        RECT 895.950 527.100 898.050 529.200 ;
        RECT 901.950 527.100 904.050 529.200 ;
        RECT 914.400 528.600 915.450 538.950 ;
        RECT 896.400 526.350 897.600 527.100 ;
        RECT 886.950 523.950 889.050 526.050 ;
        RECT 889.950 523.950 892.050 526.050 ;
        RECT 892.950 523.950 895.050 526.050 ;
        RECT 895.950 523.950 898.050 526.050 ;
        RECT 880.950 520.950 883.050 523.050 ;
        RECT 887.400 522.900 888.600 523.650 ;
        RECT 893.400 522.900 894.600 523.650 ;
        RECT 886.950 520.800 889.050 522.900 ;
        RECT 892.950 517.950 895.050 522.900 ;
        RECT 898.950 520.950 901.050 523.050 ;
        RECT 877.950 514.950 880.050 517.050 ;
        RECT 883.950 514.950 886.050 517.050 ;
        RECT 880.950 511.950 883.050 514.050 ;
        RECT 859.950 499.950 862.050 502.050 ;
        RECT 871.950 499.950 874.050 502.050 ;
        RECT 874.950 499.950 877.050 502.050 ;
        RECT 877.950 499.950 880.050 502.050 ;
        RECT 860.400 490.050 861.450 499.950 ;
        RECT 869.400 497.400 876.450 498.450 ;
        RECT 869.400 495.600 870.450 497.400 ;
        RECT 869.400 493.350 870.600 495.600 ;
        RECT 863.100 490.950 865.200 493.050 ;
        RECT 868.500 490.950 870.600 493.050 ;
        RECT 871.800 490.950 873.900 493.050 ;
        RECT 859.950 489.450 862.050 490.050 ;
        RECT 863.400 489.450 864.600 490.650 ;
        RECT 859.950 488.400 864.600 489.450 ;
        RECT 872.400 488.400 873.600 490.650 ;
        RECT 859.950 487.950 862.050 488.400 ;
        RECT 856.950 484.950 859.050 487.050 ;
        RECT 859.950 484.800 862.050 486.900 ;
        RECT 865.950 484.950 868.050 487.050 ;
        RECT 853.950 454.950 856.050 457.050 ;
        RECT 842.400 448.350 843.600 450.600 ;
        RECT 847.950 449.100 850.050 451.200 ;
        RECT 853.950 449.100 856.050 451.200 ;
        RECT 848.400 448.350 849.600 449.100 ;
        RECT 838.950 445.950 841.050 448.050 ;
        RECT 841.950 445.950 844.050 448.050 ;
        RECT 844.950 445.950 847.050 448.050 ;
        RECT 847.950 445.950 850.050 448.050 ;
        RECT 839.400 444.900 840.600 445.650 ;
        RECT 845.400 444.900 846.600 445.650 ;
        RECT 808.950 436.950 811.050 439.050 ;
        RECT 815.400 436.050 816.450 443.400 ;
        RECT 811.950 433.950 814.050 436.050 ;
        RECT 814.950 433.950 817.050 436.050 ;
        RECT 805.950 416.100 808.050 418.200 ;
        RECT 812.400 417.600 813.450 433.950 ;
        RECT 821.400 430.050 822.450 443.400 ;
        RECT 832.950 442.800 835.050 444.900 ;
        RECT 838.950 442.800 841.050 444.900 ;
        RECT 844.950 442.800 847.050 444.900 ;
        RECT 854.400 433.050 855.450 449.100 ;
        RECT 860.400 433.050 861.450 484.800 ;
        RECT 862.950 466.950 865.050 469.050 ;
        RECT 838.950 430.950 841.050 433.050 ;
        RECT 847.950 430.950 850.050 433.050 ;
        RECT 853.950 430.950 856.050 433.050 ;
        RECT 859.950 430.950 862.050 433.050 ;
        RECT 820.950 427.950 823.050 430.050 ;
        RECT 835.950 424.950 838.050 427.050 ;
        RECT 806.400 415.350 807.600 416.100 ;
        RECT 812.400 415.350 813.600 417.600 ;
        RECT 814.950 417.450 819.000 418.050 ;
        RECT 814.950 415.950 819.450 417.450 ;
        RECT 820.950 416.100 823.050 418.200 ;
        RECT 826.950 416.100 829.050 418.200 ;
        RECT 802.950 412.950 805.050 415.050 ;
        RECT 805.950 412.950 808.050 415.050 ;
        RECT 808.950 412.950 811.050 415.050 ;
        RECT 811.950 412.950 814.050 415.050 ;
        RECT 803.400 411.900 804.600 412.650 ;
        RECT 802.950 409.800 805.050 411.900 ;
        RECT 809.400 410.400 810.600 412.650 ;
        RECT 809.400 403.050 810.450 410.400 ;
        RECT 808.950 400.950 811.050 403.050 ;
        RECT 787.950 397.950 790.050 400.050 ;
        RECT 793.950 397.950 796.050 400.050 ;
        RECT 787.950 391.950 790.050 394.050 ;
        RECT 776.400 370.350 777.600 372.600 ;
        RECT 782.400 370.350 783.600 372.600 ;
        RECT 775.950 367.950 778.050 370.050 ;
        RECT 778.950 367.950 781.050 370.050 ;
        RECT 781.950 367.950 784.050 370.050 ;
        RECT 779.400 365.400 780.600 367.650 ;
        RECT 788.400 367.050 789.450 391.950 ;
        RECT 796.950 385.950 799.050 388.050 ;
        RECT 790.950 376.950 793.050 379.050 ;
        RECT 791.400 367.050 792.450 376.950 ;
        RECT 797.400 372.600 798.450 385.950 ;
        RECT 811.950 382.950 814.050 385.050 ;
        RECT 797.400 370.350 798.600 372.600 ;
        RECT 802.950 371.100 805.050 373.200 ;
        RECT 803.400 370.350 804.600 371.100 ;
        RECT 796.950 367.950 799.050 370.050 ;
        RECT 799.950 367.950 802.050 370.050 ;
        RECT 802.950 367.950 805.050 370.050 ;
        RECT 805.950 367.950 808.050 370.050 ;
        RECT 770.400 356.400 774.450 357.450 ;
        RECT 769.950 352.950 772.050 355.050 ;
        RECT 766.950 337.950 769.050 340.050 ;
        RECT 767.400 325.050 768.450 337.950 ;
        RECT 770.400 333.900 771.450 352.950 ;
        RECT 773.400 340.050 774.450 356.400 ;
        RECT 779.400 355.050 780.450 365.400 ;
        RECT 787.950 364.950 790.050 367.050 ;
        RECT 790.950 364.950 793.050 367.050 ;
        RECT 793.950 364.950 796.050 367.050 ;
        RECT 800.400 366.900 801.600 367.650 ;
        RECT 781.950 355.950 784.050 358.050 ;
        RECT 778.950 352.950 781.050 355.050 ;
        RECT 782.400 351.450 783.450 355.950 ;
        RECT 779.400 350.400 783.450 351.450 ;
        RECT 772.950 337.950 775.050 340.050 ;
        RECT 779.400 339.600 780.450 350.400 ;
        RECT 784.950 346.950 787.050 349.050 ;
        RECT 785.400 340.200 786.450 346.950 ;
        RECT 790.950 340.950 793.050 343.050 ;
        RECT 779.400 337.350 780.600 339.600 ;
        RECT 784.950 338.100 787.050 340.200 ;
        RECT 785.400 337.350 786.600 338.100 ;
        RECT 775.950 334.950 778.050 337.050 ;
        RECT 778.950 334.950 781.050 337.050 ;
        RECT 781.950 334.950 784.050 337.050 ;
        RECT 784.950 334.950 787.050 337.050 ;
        RECT 769.950 331.800 772.050 333.900 ;
        RECT 772.950 331.950 775.050 334.050 ;
        RECT 776.400 333.900 777.600 334.650 ;
        RECT 766.950 322.950 769.050 325.050 ;
        RECT 754.950 310.950 757.050 313.050 ;
        RECT 763.950 310.950 766.050 313.050 ;
        RECT 731.400 287.400 735.450 288.450 ;
        RECT 712.950 277.950 715.050 280.050 ;
        RECT 725.400 271.050 726.450 287.400 ;
        RECT 731.400 285.450 732.450 287.400 ;
        RECT 728.400 284.400 732.450 285.450 ;
        RECT 724.950 268.950 727.050 271.050 ;
        RECT 709.950 259.950 712.050 262.050 ;
        RECT 715.950 260.100 718.050 262.200 ;
        RECT 724.950 260.100 727.050 262.200 ;
        RECT 716.400 259.350 717.600 260.100 ;
        RECT 712.950 256.950 715.050 259.050 ;
        RECT 715.950 256.950 718.050 259.050 ;
        RECT 713.400 255.900 714.600 256.650 ;
        RECT 712.950 253.800 715.050 255.900 ;
        RECT 706.950 250.950 709.050 253.050 ;
        RECT 703.950 235.950 706.050 238.050 ;
        RECT 694.950 229.950 697.050 232.050 ;
        RECT 697.950 226.050 700.050 229.050 ;
        RECT 707.400 226.050 708.450 250.950 ;
        RECT 709.950 247.950 712.050 253.050 ;
        RECT 712.950 235.950 715.050 238.050 ;
        RECT 697.800 225.000 700.050 226.050 ;
        RECT 697.800 223.950 699.900 225.000 ;
        RECT 706.950 223.950 709.050 226.050 ;
        RECT 688.950 215.100 691.050 217.200 ;
        RECT 694.950 216.000 697.050 220.050 ;
        RECT 706.950 217.950 712.050 220.050 ;
        RECT 689.400 214.350 690.600 215.100 ;
        RECT 695.400 214.350 696.600 216.000 ;
        RECT 703.950 214.950 706.050 217.050 ;
        RECT 713.400 216.600 714.450 235.950 ;
        RECT 685.950 211.950 688.050 214.050 ;
        RECT 688.950 211.950 691.050 214.050 ;
        RECT 691.950 211.950 694.050 214.050 ;
        RECT 694.950 211.950 697.050 214.050 ;
        RECT 686.400 211.050 687.600 211.650 ;
        RECT 682.950 209.400 687.600 211.050 ;
        RECT 692.400 210.900 693.600 211.650 ;
        RECT 682.950 208.950 687.000 209.400 ;
        RECT 691.950 208.800 694.050 210.900 ;
        RECT 694.950 196.950 697.050 199.050 ;
        RECT 679.950 182.100 682.050 184.200 ;
        RECT 685.950 182.100 688.050 184.200 ;
        RECT 686.400 181.350 687.600 182.100 ;
        RECT 662.100 178.950 664.200 181.050 ;
        RECT 667.500 178.950 669.600 181.050 ;
        RECT 670.800 178.950 672.900 181.050 ;
        RECT 673.950 178.950 676.050 181.050 ;
        RECT 685.950 178.950 688.050 181.050 ;
        RECT 688.950 178.950 691.050 181.050 ;
        RECT 662.400 177.450 663.600 178.650 ;
        RECT 659.400 176.400 663.600 177.450 ;
        RECT 671.400 176.400 672.600 178.650 ;
        RECT 689.400 176.400 690.600 178.650 ;
        RECT 655.950 169.800 658.050 171.900 ;
        RECT 643.950 157.950 646.050 160.050 ;
        RECT 652.950 157.950 655.050 160.050 ;
        RECT 656.400 157.050 657.450 169.800 ;
        RECT 661.950 160.950 664.050 163.050 ;
        RECT 655.950 154.950 658.050 157.050 ;
        RECT 649.950 145.950 652.050 148.050 ;
        RECT 619.950 139.950 622.050 142.050 ;
        RECT 620.400 138.600 621.450 139.950 ;
        RECT 590.400 136.350 591.600 138.600 ;
        RECT 596.400 136.350 597.600 138.600 ;
        RECT 614.400 138.450 615.600 138.600 ;
        RECT 608.400 137.400 615.600 138.450 ;
        RECT 589.950 133.950 592.050 136.050 ;
        RECT 592.950 133.950 595.050 136.050 ;
        RECT 595.950 133.950 598.050 136.050 ;
        RECT 598.950 133.950 601.050 136.050 ;
        RECT 593.400 132.900 594.600 133.650 ;
        RECT 592.950 130.800 595.050 132.900 ;
        RECT 599.400 131.400 600.600 133.650 ;
        RECT 592.950 124.950 595.050 127.050 ;
        RECT 580.950 115.950 583.050 118.050 ;
        RECT 568.950 106.950 571.050 109.050 ;
        RECT 574.950 106.950 577.050 109.050 ;
        RECT 569.400 99.900 570.450 106.950 ;
        RECT 571.950 103.950 574.050 106.050 ;
        RECT 580.950 105.000 583.050 112.050 ;
        RECT 568.950 97.800 571.050 99.900 ;
        RECT 565.950 94.950 568.050 97.050 ;
        RECT 541.950 91.950 544.050 94.050 ;
        RECT 550.950 91.950 553.050 94.050 ;
        RECT 526.950 76.950 529.050 79.050 ;
        RECT 478.950 70.950 481.050 73.050 ;
        RECT 487.950 70.950 490.050 73.050 ;
        RECT 523.950 70.950 526.050 73.050 ;
        RECT 472.950 49.950 475.050 52.050 ;
        RECT 457.950 46.950 460.050 49.050 ;
        RECT 448.950 40.950 451.050 43.050 ;
        RECT 457.950 31.950 460.050 34.050 ;
        RECT 458.400 27.600 459.450 31.950 ;
        RECT 419.400 25.350 420.600 26.400 ;
        RECT 437.400 25.350 438.600 27.600 ;
        RECT 458.400 25.350 459.600 27.600 ;
        RECT 463.950 26.100 466.050 28.200 ;
        RECT 469.950 26.100 472.050 28.200 ;
        RECT 479.400 27.600 480.450 70.950 ;
        RECT 490.950 67.950 493.050 70.050 ;
        RECT 508.950 67.950 511.050 70.050 ;
        RECT 484.950 59.100 487.050 61.200 ;
        RECT 491.400 60.600 492.450 67.950 ;
        RECT 485.400 58.350 486.600 59.100 ;
        RECT 491.400 58.350 492.600 60.600 ;
        RECT 496.950 59.100 499.050 61.200 ;
        RECT 509.400 60.600 510.450 67.950 ;
        RECT 484.950 55.950 487.050 58.050 ;
        RECT 487.950 55.950 490.050 58.050 ;
        RECT 490.950 55.950 493.050 58.050 ;
        RECT 488.400 54.000 489.600 55.650 ;
        RECT 497.400 55.050 498.450 59.100 ;
        RECT 509.400 58.350 510.600 60.600 ;
        RECT 517.950 59.100 520.050 61.200 ;
        RECT 518.400 58.350 519.600 59.100 ;
        RECT 527.400 58.050 528.450 76.950 ;
        RECT 538.950 70.950 541.050 73.050 ;
        RECT 532.950 59.100 535.050 61.200 ;
        RECT 539.400 60.600 540.450 70.950 ;
        RECT 572.400 61.200 573.450 103.950 ;
        RECT 581.400 103.350 582.600 105.000 ;
        RECT 586.950 104.100 589.050 106.200 ;
        RECT 587.400 103.350 588.600 104.100 ;
        RECT 577.950 100.950 580.050 103.050 ;
        RECT 580.950 100.950 583.050 103.050 ;
        RECT 583.950 100.950 586.050 103.050 ;
        RECT 586.950 100.950 589.050 103.050 ;
        RECT 578.400 99.000 579.600 100.650 ;
        RECT 584.400 99.900 585.600 100.650 ;
        RECT 577.950 94.950 580.050 99.000 ;
        RECT 583.950 97.800 586.050 99.900 ;
        RECT 589.950 96.450 592.050 97.050 ;
        RECT 593.400 96.450 594.450 124.950 ;
        RECT 599.400 124.050 600.450 131.400 ;
        RECT 595.800 121.950 597.900 124.050 ;
        RECT 598.950 121.950 601.050 124.050 ;
        RECT 596.400 118.050 597.450 121.950 ;
        RECT 595.950 115.950 598.050 118.050 ;
        RECT 604.950 109.950 607.050 112.050 ;
        RECT 605.400 106.200 606.450 109.950 ;
        RECT 608.400 109.050 609.450 137.400 ;
        RECT 614.400 136.350 615.600 137.400 ;
        RECT 620.400 136.350 621.600 138.600 ;
        RECT 631.950 137.100 634.050 139.200 ;
        RECT 640.950 138.000 643.050 142.050 ;
        RECT 613.950 133.950 616.050 136.050 ;
        RECT 616.950 133.950 619.050 136.050 ;
        RECT 619.950 133.950 622.050 136.050 ;
        RECT 622.950 133.950 625.050 136.050 ;
        RECT 617.400 131.400 618.600 133.650 ;
        RECT 623.400 131.400 624.600 133.650 ;
        RECT 632.400 132.450 633.450 137.100 ;
        RECT 641.400 136.350 642.600 138.000 ;
        RECT 646.800 137.100 648.900 139.200 ;
        RECT 650.400 139.050 651.450 145.950 ;
        RECT 647.400 136.350 648.600 137.100 ;
        RECT 649.950 136.950 652.050 139.050 ;
        RECT 662.400 138.600 663.450 160.950 ;
        RECT 671.400 154.050 672.450 176.400 ;
        RECT 689.400 166.050 690.450 176.400 ;
        RECT 688.950 163.950 691.050 166.050 ;
        RECT 695.400 154.050 696.450 196.950 ;
        RECT 704.400 196.050 705.450 214.950 ;
        RECT 713.400 214.350 714.600 216.600 ;
        RECT 712.950 211.950 715.050 214.050 ;
        RECT 715.950 211.950 718.050 214.050 ;
        RECT 716.400 210.000 717.600 211.650 ;
        RECT 715.950 205.950 718.050 210.000 ;
        RECT 725.400 205.050 726.450 260.100 ;
        RECT 728.400 235.050 729.450 284.400 ;
        RECT 737.400 265.050 738.450 292.800 ;
        RECT 746.400 292.350 747.600 294.600 ;
        RECT 748.950 292.950 751.050 295.050 ;
        RECT 751.950 292.950 754.050 295.050 ;
        RECT 742.950 289.950 745.050 292.050 ;
        RECT 745.950 289.950 748.050 292.050 ;
        RECT 743.400 288.900 744.600 289.650 ;
        RECT 742.950 286.800 745.050 288.900 ;
        RECT 748.950 286.950 751.050 289.050 ;
        RECT 736.950 262.950 739.050 265.050 ;
        RECT 731.100 256.950 733.200 259.050 ;
        RECT 734.400 256.950 736.500 259.050 ;
        RECT 739.800 256.950 741.900 259.050 ;
        RECT 731.400 254.400 732.600 256.650 ;
        RECT 740.400 255.900 741.600 256.650 ;
        RECT 731.400 253.050 732.450 254.400 ;
        RECT 739.950 253.800 742.050 255.900 ;
        RECT 730.950 250.950 733.050 253.050 ;
        RECT 727.950 232.950 730.050 235.050 ;
        RECT 731.400 228.450 732.450 250.950 ;
        RECT 743.400 244.050 744.450 286.800 ;
        RECT 745.950 283.950 748.050 286.050 ;
        RECT 746.400 255.900 747.450 283.950 ;
        RECT 745.950 253.800 748.050 255.900 ;
        RECT 742.950 241.950 745.050 244.050 ;
        RECT 746.400 235.050 747.450 253.800 ;
        RECT 745.950 232.950 748.050 235.050 ;
        RECT 728.400 227.400 732.450 228.450 ;
        RECT 728.400 216.450 729.450 227.400 ;
        RECT 742.950 217.950 745.050 220.050 ;
        RECT 731.400 216.450 732.600 216.600 ;
        RECT 728.400 215.400 732.600 216.450 ;
        RECT 731.400 214.350 732.600 215.400 ;
        RECT 736.950 215.100 739.050 217.200 ;
        RECT 737.400 214.350 738.600 215.100 ;
        RECT 730.950 211.950 733.050 214.050 ;
        RECT 733.950 211.950 736.050 214.050 ;
        RECT 736.950 211.950 739.050 214.050 ;
        RECT 734.400 209.400 735.600 211.650 ;
        RECT 724.950 202.950 727.050 205.050 ;
        RECT 697.950 193.950 700.050 196.050 ;
        RECT 703.950 193.950 706.050 196.050 ;
        RECT 698.400 177.900 699.450 193.950 ;
        RECT 703.950 187.950 706.050 190.050 ;
        RECT 704.400 183.600 705.450 187.950 ;
        RECT 734.400 187.050 735.450 209.400 ;
        RECT 743.400 193.050 744.450 217.950 ;
        RECT 745.950 202.950 748.050 205.050 ;
        RECT 742.950 190.950 745.050 193.050 ;
        RECT 733.950 184.950 736.050 187.050 ;
        RECT 704.400 181.350 705.600 183.600 ;
        RECT 709.950 182.100 712.050 184.200 ;
        RECT 721.950 182.100 724.050 184.200 ;
        RECT 730.950 182.100 733.050 184.200 ;
        RECT 736.950 182.100 739.050 184.200 ;
        RECT 710.400 181.350 711.600 182.100 ;
        RECT 703.950 178.950 706.050 181.050 ;
        RECT 706.950 178.950 709.050 181.050 ;
        RECT 709.950 178.950 712.050 181.050 ;
        RECT 712.950 178.950 715.050 181.050 ;
        RECT 707.400 177.900 708.600 178.650 ;
        RECT 697.950 175.800 700.050 177.900 ;
        RECT 706.950 175.800 709.050 177.900 ;
        RECT 713.400 177.000 714.600 178.650 ;
        RECT 712.950 172.950 715.050 177.000 ;
        RECT 712.950 169.800 715.050 171.900 ;
        RECT 670.950 151.950 673.050 154.050 ;
        RECT 694.950 151.950 697.050 154.050 ;
        RECT 671.400 145.050 672.450 151.950 ;
        RECT 670.950 142.950 673.050 145.050 ;
        RECT 694.950 142.950 697.050 145.050 ;
        RECT 662.400 136.350 663.600 138.600 ;
        RECT 670.950 137.100 673.050 139.200 ;
        RECT 688.950 137.100 691.050 139.200 ;
        RECT 695.400 138.600 696.450 142.950 ;
        RECT 671.400 136.350 672.600 137.100 ;
        RECT 689.400 136.350 690.600 137.100 ;
        RECT 695.400 136.350 696.600 138.600 ;
        RECT 706.950 137.100 709.050 139.200 ;
        RECT 713.400 138.600 714.450 169.800 ;
        RECT 722.400 160.050 723.450 182.100 ;
        RECT 731.400 181.350 732.600 182.100 ;
        RECT 737.400 181.350 738.600 182.100 ;
        RECT 742.950 181.950 745.050 184.050 ;
        RECT 727.950 178.950 730.050 181.050 ;
        RECT 730.950 178.950 733.050 181.050 ;
        RECT 733.950 178.950 736.050 181.050 ;
        RECT 736.950 178.950 739.050 181.050 ;
        RECT 728.400 176.400 729.600 178.650 ;
        RECT 734.400 177.900 735.600 178.650 ;
        RECT 728.400 166.050 729.450 176.400 ;
        RECT 733.950 175.800 736.050 177.900 ;
        RECT 730.950 172.950 733.050 175.050 ;
        RECT 727.950 163.950 730.050 166.050 ;
        RECT 721.950 157.950 724.050 160.050 ;
        RECT 637.950 133.950 640.050 136.050 ;
        RECT 640.950 133.950 643.050 136.050 ;
        RECT 643.950 133.950 646.050 136.050 ;
        RECT 646.950 133.950 649.050 136.050 ;
        RECT 662.100 133.950 664.200 136.050 ;
        RECT 667.500 133.950 669.600 136.050 ;
        RECT 670.800 133.950 672.900 136.050 ;
        RECT 688.950 133.950 691.050 136.050 ;
        RECT 691.950 133.950 694.050 136.050 ;
        RECT 694.950 133.950 697.050 136.050 ;
        RECT 632.400 131.400 636.450 132.450 ;
        RECT 617.400 115.050 618.450 131.400 ;
        RECT 623.400 124.050 624.450 131.400 ;
        RECT 628.950 124.800 631.050 126.900 ;
        RECT 622.950 121.950 625.050 124.050 ;
        RECT 622.950 115.950 625.050 118.050 ;
        RECT 616.950 112.950 619.050 115.050 ;
        RECT 607.950 106.950 610.050 109.050 ;
        RECT 595.950 103.950 598.050 106.050 ;
        RECT 604.950 104.100 607.050 106.200 ;
        RECT 623.400 106.050 624.450 115.950 ;
        RECT 612.000 105.600 616.050 106.050 ;
        RECT 589.950 95.400 594.450 96.450 ;
        RECT 589.950 94.950 592.050 95.400 ;
        RECT 578.400 91.050 579.450 94.950 ;
        RECT 590.400 91.050 591.450 94.950 ;
        RECT 596.400 91.050 597.450 103.950 ;
        RECT 605.400 103.350 606.600 104.100 ;
        RECT 611.400 103.950 616.050 105.600 ;
        RECT 622.950 103.950 625.050 106.050 ;
        RECT 629.400 105.600 630.450 124.800 ;
        RECT 635.400 118.050 636.450 131.400 ;
        RECT 638.400 131.400 639.600 133.650 ;
        RECT 644.400 131.400 645.600 133.650 ;
        RECT 692.400 132.900 693.600 133.650 ;
        RECT 707.400 133.050 708.450 137.100 ;
        RECT 713.400 136.350 714.600 138.600 ;
        RECT 718.950 137.100 721.050 139.200 ;
        RECT 719.400 136.350 720.600 137.100 ;
        RECT 727.950 136.950 730.050 139.050 ;
        RECT 712.950 133.950 715.050 136.050 ;
        RECT 715.950 133.950 718.050 136.050 ;
        RECT 718.950 133.950 721.050 136.050 ;
        RECT 721.950 133.950 724.050 136.050 ;
        RECT 638.400 124.050 639.450 131.400 ;
        RECT 637.950 121.950 640.050 124.050 ;
        RECT 634.950 115.950 637.050 118.050 ;
        RECT 640.950 112.950 643.050 115.050 ;
        RECT 611.400 103.350 612.600 103.950 ;
        RECT 629.400 103.350 630.600 105.600 ;
        RECT 634.950 104.100 637.050 106.200 ;
        RECT 635.400 103.350 636.600 104.100 ;
        RECT 601.950 100.950 604.050 103.050 ;
        RECT 604.950 100.950 607.050 103.050 ;
        RECT 607.950 100.950 610.050 103.050 ;
        RECT 610.950 100.950 613.050 103.050 ;
        RECT 625.950 100.950 628.050 103.050 ;
        RECT 628.950 100.950 631.050 103.050 ;
        RECT 631.950 100.950 634.050 103.050 ;
        RECT 634.950 100.950 637.050 103.050 ;
        RECT 602.400 99.900 603.600 100.650 ;
        RECT 601.950 97.800 604.050 99.900 ;
        RECT 608.400 99.000 609.600 100.650 ;
        RECT 607.950 94.950 610.050 99.000 ;
        RECT 622.950 97.950 625.050 100.050 ;
        RECT 626.400 99.900 627.600 100.650 ;
        RECT 632.400 99.900 633.600 100.650 ;
        RECT 577.950 88.950 580.050 91.050 ;
        RECT 589.950 88.950 592.050 91.050 ;
        RECT 595.950 88.950 598.050 91.050 ;
        RECT 601.950 82.950 604.050 85.050 ;
        RECT 574.950 79.950 577.050 82.050 ;
        RECT 592.950 79.950 595.050 82.050 ;
        RECT 533.400 58.350 534.600 59.100 ;
        RECT 539.400 58.350 540.600 60.600 ;
        RECT 545.400 60.450 546.600 60.600 ;
        RECT 560.400 60.450 561.600 60.600 ;
        RECT 545.400 59.400 552.450 60.450 ;
        RECT 545.400 58.350 546.600 59.400 ;
        RECT 509.100 55.950 511.200 58.050 ;
        RECT 514.500 55.950 516.600 58.050 ;
        RECT 517.800 55.950 519.900 58.050 ;
        RECT 526.950 55.950 529.050 58.050 ;
        RECT 532.950 55.950 535.050 58.050 ;
        RECT 535.950 55.950 538.050 58.050 ;
        RECT 538.950 55.950 541.050 58.050 ;
        RECT 541.950 55.950 544.050 58.050 ;
        RECT 544.950 55.950 547.050 58.050 ;
        RECT 487.950 49.950 490.050 54.000 ;
        RECT 496.950 52.950 499.050 55.050 ;
        RECT 515.400 54.900 516.600 55.650 ;
        RECT 536.400 54.900 537.600 55.650 ;
        RECT 542.400 54.900 543.600 55.650 ;
        RECT 514.950 52.800 517.050 54.900 ;
        RECT 535.950 52.800 538.050 54.900 ;
        RECT 541.950 52.800 544.050 54.900 ;
        RECT 541.950 49.650 544.050 51.750 ;
        RECT 484.950 46.950 487.050 49.050 ;
        RECT 485.400 34.050 486.450 46.950 ;
        RECT 542.400 46.050 543.450 49.650 ;
        RECT 551.400 49.050 552.450 59.400 ;
        RECT 557.400 59.400 561.600 60.450 ;
        RECT 557.400 52.050 558.450 59.400 ;
        RECT 560.400 58.350 561.600 59.400 ;
        RECT 569.400 60.450 570.600 60.600 ;
        RECT 571.950 60.450 574.050 61.200 ;
        RECT 569.400 59.400 574.050 60.450 ;
        RECT 569.400 58.350 570.600 59.400 ;
        RECT 571.950 59.100 574.050 59.400 ;
        RECT 560.100 55.950 562.200 58.050 ;
        RECT 563.400 55.950 565.500 58.050 ;
        RECT 568.800 55.950 570.900 58.050 ;
        RECT 563.400 54.900 564.600 55.650 ;
        RECT 575.400 54.900 576.450 79.950 ;
        RECT 580.950 70.950 583.050 73.050 ;
        RECT 577.950 64.950 580.050 67.050 ;
        RECT 562.950 52.800 565.050 54.900 ;
        RECT 574.950 52.800 577.050 54.900 ;
        RECT 556.950 49.950 559.050 52.050 ;
        RECT 550.950 46.950 553.050 49.050 ;
        RECT 541.950 43.950 544.050 46.050 ;
        RECT 551.400 43.050 552.450 46.950 ;
        RECT 496.950 40.950 499.050 43.050 ;
        RECT 550.950 40.950 553.050 43.050 ;
        RECT 574.950 40.950 577.050 43.050 ;
        RECT 484.950 31.950 487.050 34.050 ;
        RECT 485.400 27.600 486.450 31.950 ;
        RECT 464.400 25.350 465.600 26.100 ;
        RECT 413.100 22.950 415.200 25.050 ;
        RECT 418.500 22.950 420.600 25.050 ;
        RECT 433.950 22.950 436.050 25.050 ;
        RECT 436.950 22.950 439.050 25.050 ;
        RECT 454.950 22.950 457.050 25.050 ;
        RECT 457.950 22.950 460.050 25.050 ;
        RECT 460.950 22.950 463.050 25.050 ;
        RECT 463.950 22.950 466.050 25.050 ;
        RECT 397.950 19.800 400.050 21.900 ;
        RECT 434.400 20.400 435.600 22.650 ;
        RECT 455.400 21.900 456.600 22.650 ;
        RECT 349.950 13.950 352.050 16.050 ;
        RECT 364.950 13.950 367.050 16.050 ;
        RECT 434.400 13.050 435.450 20.400 ;
        RECT 454.950 19.800 457.050 21.900 ;
        RECT 461.400 21.000 462.600 22.650 ;
        RECT 460.950 16.950 463.050 21.000 ;
        RECT 295.950 11.400 303.450 12.450 ;
        RECT 295.950 10.950 298.050 11.400 ;
        RECT 433.950 10.950 436.050 13.050 ;
        RECT 470.400 7.050 471.450 26.100 ;
        RECT 479.400 25.350 480.600 27.600 ;
        RECT 485.400 25.350 486.600 27.600 ;
        RECT 493.950 25.950 496.050 28.050 ;
        RECT 478.950 22.950 481.050 25.050 ;
        RECT 481.950 22.950 484.050 25.050 ;
        RECT 484.950 22.950 487.050 25.050 ;
        RECT 487.950 22.950 490.050 25.050 ;
        RECT 482.400 20.400 483.600 22.650 ;
        RECT 488.400 22.050 489.600 22.650 ;
        RECT 488.400 20.400 493.050 22.050 ;
        RECT 482.400 13.050 483.450 20.400 ;
        RECT 489.000 19.950 493.050 20.400 ;
        RECT 494.400 19.050 495.450 25.950 ;
        RECT 497.400 22.050 498.450 40.950 ;
        RECT 535.800 37.950 537.900 40.050 ;
        RECT 538.950 37.950 541.050 40.050 ;
        RECT 536.400 31.050 537.450 37.950 ;
        RECT 535.950 28.950 538.050 31.050 ;
        RECT 502.950 26.100 505.050 28.200 ;
        RECT 508.950 26.100 511.050 28.200 ;
        RECT 532.950 26.100 535.050 28.200 ;
        RECT 539.400 27.600 540.450 37.950 ;
        RECT 547.950 28.950 550.050 31.050 ;
        RECT 503.400 25.350 504.600 26.100 ;
        RECT 509.400 25.350 510.600 26.100 ;
        RECT 533.400 25.350 534.600 26.100 ;
        RECT 539.400 25.350 540.600 27.600 ;
        RECT 544.950 25.950 547.050 28.050 ;
        RECT 502.950 22.950 505.050 25.050 ;
        RECT 505.950 22.950 508.050 25.050 ;
        RECT 508.950 22.950 511.050 25.050 ;
        RECT 511.950 22.950 514.050 25.050 ;
        RECT 529.950 22.950 532.050 25.050 ;
        RECT 532.950 22.950 535.050 25.050 ;
        RECT 535.950 22.950 538.050 25.050 ;
        RECT 538.950 22.950 541.050 25.050 ;
        RECT 496.950 19.950 499.050 22.050 ;
        RECT 506.400 20.400 507.600 22.650 ;
        RECT 512.400 21.900 513.600 22.650 ;
        RECT 493.950 16.950 496.050 19.050 ;
        RECT 506.400 13.050 507.450 20.400 ;
        RECT 511.950 19.800 514.050 21.900 ;
        RECT 530.400 20.400 531.600 22.650 ;
        RECT 536.400 21.900 537.600 22.650 ;
        RECT 530.400 13.050 531.450 20.400 ;
        RECT 535.950 16.950 538.050 21.900 ;
        RECT 545.400 19.050 546.450 25.950 ;
        RECT 548.400 21.900 549.450 28.950 ;
        RECT 556.950 26.100 559.050 28.200 ;
        RECT 562.950 27.000 565.050 31.050 ;
        RECT 557.400 25.350 558.600 26.100 ;
        RECT 563.400 25.350 564.600 27.000 ;
        RECT 553.950 22.950 556.050 25.050 ;
        RECT 556.950 22.950 559.050 25.050 ;
        RECT 559.950 22.950 562.050 25.050 ;
        RECT 562.950 22.950 565.050 25.050 ;
        RECT 554.400 21.900 555.600 22.650 ;
        RECT 560.400 21.900 561.600 22.650 ;
        RECT 575.400 21.900 576.450 40.950 ;
        RECT 578.400 40.050 579.450 64.950 ;
        RECT 581.400 43.050 582.450 70.950 ;
        RECT 586.950 59.100 589.050 61.200 ;
        RECT 593.400 60.600 594.450 79.950 ;
        RECT 587.400 58.350 588.600 59.100 ;
        RECT 593.400 58.350 594.600 60.600 ;
        RECT 586.950 55.950 589.050 58.050 ;
        RECT 589.950 55.950 592.050 58.050 ;
        RECT 592.950 55.950 595.050 58.050 ;
        RECT 598.950 55.950 601.050 58.050 ;
        RECT 590.400 53.400 591.600 55.650 ;
        RECT 586.950 49.950 589.050 52.050 ;
        RECT 580.950 40.950 583.050 43.050 ;
        RECT 577.950 37.950 580.050 40.050 ;
        RECT 580.950 27.000 583.050 31.050 ;
        RECT 587.400 27.600 588.450 49.950 ;
        RECT 590.400 37.050 591.450 53.400 ;
        RECT 589.950 34.950 592.050 37.050 ;
        RECT 599.400 31.050 600.450 55.950 ;
        RECT 602.400 54.900 603.450 82.950 ;
        RECT 623.400 79.050 624.450 97.950 ;
        RECT 625.950 97.800 628.050 99.900 ;
        RECT 631.950 97.800 634.050 99.900 ;
        RECT 637.950 91.950 640.050 97.050 ;
        RECT 636.000 90.900 639.000 91.050 ;
        RECT 634.950 88.950 640.050 90.900 ;
        RECT 634.950 88.800 637.050 88.950 ;
        RECT 637.950 88.800 640.050 88.950 ;
        RECT 622.950 76.950 625.050 79.050 ;
        RECT 613.950 73.950 616.050 76.050 ;
        RECT 607.950 64.950 610.050 67.050 ;
        RECT 608.400 60.600 609.450 64.950 ;
        RECT 614.400 60.600 615.450 73.950 ;
        RECT 641.400 64.050 642.450 112.950 ;
        RECT 644.400 109.050 645.450 131.400 ;
        RECT 691.950 130.800 694.050 132.900 ;
        RECT 706.950 130.950 709.050 133.050 ;
        RECT 716.400 132.900 717.600 133.650 ;
        RECT 715.950 130.800 718.050 132.900 ;
        RECT 722.400 131.400 723.600 133.650 ;
        RECT 728.400 132.900 729.450 136.950 ;
        RECT 709.950 124.950 712.050 127.050 ;
        RECT 655.950 112.950 658.050 115.050 ;
        RECT 685.950 112.950 688.050 115.050 ;
        RECT 656.400 109.050 657.450 112.950 ;
        RECT 673.950 109.950 676.050 112.050 ;
        RECT 643.950 106.950 646.050 109.050 ;
        RECT 643.950 103.800 646.050 105.900 ;
        RECT 655.950 105.000 658.050 109.050 ;
        RECT 640.950 61.950 643.050 64.050 ;
        RECT 608.400 58.350 609.600 60.600 ;
        RECT 614.400 58.350 615.600 60.600 ;
        RECT 634.950 59.100 637.050 61.200 ;
        RECT 641.400 60.600 642.450 61.950 ;
        RECT 635.400 58.350 636.600 59.100 ;
        RECT 641.400 58.350 642.600 60.600 ;
        RECT 644.400 60.450 645.450 103.800 ;
        RECT 656.400 103.350 657.600 105.000 ;
        RECT 661.950 104.100 664.050 106.200 ;
        RECT 662.400 103.350 663.600 104.100 ;
        RECT 667.800 103.950 669.900 106.050 ;
        RECT 670.950 103.950 673.050 106.050 ;
        RECT 652.950 100.950 655.050 103.050 ;
        RECT 655.950 100.950 658.050 103.050 ;
        RECT 658.950 100.950 661.050 103.050 ;
        RECT 661.950 100.950 664.050 103.050 ;
        RECT 653.400 99.450 654.600 100.650 ;
        RECT 659.400 99.900 660.600 100.650 ;
        RECT 650.400 99.000 654.600 99.450 ;
        RECT 650.400 98.400 655.050 99.000 ;
        RECT 646.950 88.950 649.050 94.050 ;
        RECT 650.400 79.050 651.450 98.400 ;
        RECT 652.950 94.950 655.050 98.400 ;
        RECT 658.950 97.800 661.050 99.900 ;
        RECT 655.950 91.950 658.050 97.050 ;
        RECT 652.950 90.450 655.050 91.050 ;
        RECT 658.950 90.450 661.050 91.050 ;
        RECT 652.950 89.400 661.050 90.450 ;
        RECT 652.950 88.950 655.050 89.400 ;
        RECT 658.950 88.950 661.050 89.400 ;
        RECT 655.950 85.950 658.050 88.050 ;
        RECT 649.950 76.950 652.050 79.050 ;
        RECT 649.950 64.950 652.050 67.050 ;
        RECT 644.400 59.400 648.450 60.450 ;
        RECT 607.950 55.950 610.050 58.050 ;
        RECT 610.950 55.950 613.050 58.050 ;
        RECT 613.950 55.950 616.050 58.050 ;
        RECT 616.950 55.950 619.050 58.050 ;
        RECT 631.950 55.950 634.050 58.050 ;
        RECT 634.950 55.950 637.050 58.050 ;
        RECT 637.950 55.950 640.050 58.050 ;
        RECT 640.950 55.950 643.050 58.050 ;
        RECT 611.400 54.900 612.600 55.650 ;
        RECT 601.950 52.800 604.050 54.900 ;
        RECT 610.950 52.800 613.050 54.900 ;
        RECT 617.400 53.400 618.600 55.650 ;
        RECT 632.400 54.900 633.600 55.650 ;
        RECT 617.400 49.050 618.450 53.400 ;
        RECT 631.950 52.800 634.050 54.900 ;
        RECT 638.400 54.000 639.600 55.650 ;
        RECT 637.950 49.950 640.050 54.000 ;
        RECT 647.400 52.050 648.450 59.400 ;
        RECT 650.400 52.050 651.450 64.950 ;
        RECT 656.400 61.200 657.450 85.950 ;
        RECT 668.400 73.050 669.450 103.950 ;
        RECT 667.950 70.950 670.050 73.050 ;
        RECT 658.950 64.950 664.050 67.050 ;
        RECT 671.400 64.050 672.450 103.950 ;
        RECT 674.400 99.900 675.450 109.950 ;
        RECT 679.950 104.100 682.050 106.200 ;
        RECT 686.400 105.600 687.450 112.950 ;
        RECT 680.400 103.350 681.600 104.100 ;
        RECT 686.400 103.350 687.600 105.600 ;
        RECT 703.950 104.100 706.050 106.200 ;
        RECT 710.400 105.600 711.450 124.950 ;
        RECT 704.400 103.350 705.600 104.100 ;
        RECT 710.400 103.350 711.600 105.600 ;
        RECT 718.950 104.100 721.050 106.200 ;
        RECT 679.950 100.950 682.050 103.050 ;
        RECT 682.950 100.950 685.050 103.050 ;
        RECT 685.950 100.950 688.050 103.050 ;
        RECT 688.950 100.950 691.050 103.050 ;
        RECT 703.950 100.950 706.050 103.050 ;
        RECT 706.950 100.950 709.050 103.050 ;
        RECT 709.950 100.950 712.050 103.050 ;
        RECT 712.950 100.950 715.050 103.050 ;
        RECT 683.400 99.900 684.600 100.650 ;
        RECT 673.950 97.800 676.050 99.900 ;
        RECT 682.950 97.800 685.050 99.900 ;
        RECT 689.400 99.000 690.600 100.650 ;
        RECT 707.400 99.900 708.600 100.650 ;
        RECT 685.950 91.950 688.050 97.050 ;
        RECT 688.950 94.950 691.050 99.000 ;
        RECT 700.950 97.800 703.050 99.900 ;
        RECT 706.950 97.800 709.050 99.900 ;
        RECT 713.400 99.000 714.600 100.650 ;
        RECT 701.400 91.050 702.450 97.800 ;
        RECT 706.950 94.650 709.050 96.750 ;
        RECT 712.950 94.950 715.050 99.000 ;
        RECT 707.400 91.050 708.450 94.650 ;
        RECT 700.950 88.950 703.050 91.050 ;
        RECT 706.950 88.950 709.050 91.050 ;
        RECT 719.400 88.050 720.450 104.100 ;
        RECT 722.400 97.050 723.450 131.400 ;
        RECT 727.950 130.800 730.050 132.900 ;
        RECT 731.400 121.050 732.450 172.950 ;
        RECT 733.950 166.950 736.050 169.050 ;
        RECT 734.400 132.900 735.450 166.950 ;
        RECT 743.400 142.050 744.450 181.950 ;
        RECT 746.400 166.050 747.450 202.950 ;
        RECT 749.400 184.050 750.450 286.950 ;
        RECT 755.400 264.450 756.450 310.950 ;
        RECT 760.950 304.950 763.050 307.050 ;
        RECT 761.400 294.600 762.450 304.950 ;
        RECT 761.400 292.350 762.600 294.600 ;
        RECT 760.950 289.950 763.050 292.050 ;
        RECT 763.950 289.950 766.050 292.050 ;
        RECT 764.400 288.450 765.600 289.650 ;
        RECT 764.400 287.400 768.450 288.450 ;
        RECT 767.400 280.050 768.450 287.400 ;
        RECT 769.950 280.950 772.050 283.050 ;
        RECT 766.950 277.950 769.050 280.050 ;
        RECT 755.400 263.400 759.450 264.450 ;
        RECT 758.400 261.600 759.450 263.400 ;
        RECT 763.950 262.950 766.050 265.050 ;
        RECT 758.400 259.350 759.600 261.600 ;
        RECT 754.950 256.950 757.050 259.050 ;
        RECT 757.950 256.950 760.050 259.050 ;
        RECT 755.400 255.900 756.600 256.650 ;
        RECT 754.950 253.800 757.050 255.900 ;
        RECT 760.950 247.950 763.050 250.050 ;
        RECT 761.400 244.050 762.450 247.950 ;
        RECT 760.950 241.950 763.050 244.050 ;
        RECT 760.950 219.450 763.050 220.050 ;
        RECT 764.400 219.450 765.450 262.950 ;
        RECT 760.950 218.400 765.450 219.450 ;
        RECT 760.950 217.950 763.050 218.400 ;
        RECT 751.950 215.100 754.050 217.200 ;
        RECT 761.400 216.600 762.450 217.950 ;
        RECT 752.400 214.350 753.600 215.100 ;
        RECT 761.400 214.350 762.600 216.600 ;
        RECT 763.950 214.950 766.050 217.050 ;
        RECT 752.100 211.950 754.200 214.050 ;
        RECT 755.400 211.950 757.500 214.050 ;
        RECT 760.800 211.950 762.900 214.050 ;
        RECT 757.950 202.950 760.050 205.050 ;
        RECT 751.950 199.950 754.050 202.050 ;
        RECT 748.950 181.950 751.050 184.050 ;
        RECT 752.400 183.600 753.450 199.950 ;
        RECT 758.400 183.600 759.450 202.950 ;
        RECT 764.400 183.600 765.450 214.950 ;
        RECT 767.400 202.050 768.450 277.950 ;
        RECT 770.400 277.050 771.450 280.950 ;
        RECT 773.400 280.050 774.450 331.950 ;
        RECT 775.950 331.800 778.050 333.900 ;
        RECT 782.400 332.400 783.600 334.650 ;
        RECT 782.400 328.050 783.450 332.400 ;
        RECT 781.950 325.950 784.050 328.050 ;
        RECT 791.400 322.050 792.450 340.950 ;
        RECT 790.950 319.950 793.050 322.050 ;
        RECT 791.400 316.050 792.450 319.950 ;
        RECT 790.950 313.950 793.050 316.050 ;
        RECT 775.950 292.950 778.050 295.050 ;
        RECT 787.950 294.000 790.050 298.050 ;
        RECT 772.950 277.950 775.050 280.050 ;
        RECT 769.950 274.950 772.050 277.050 ;
        RECT 773.400 261.600 774.450 277.950 ;
        RECT 776.400 268.050 777.450 292.950 ;
        RECT 788.400 292.350 789.600 294.000 ;
        RECT 781.950 289.950 784.050 292.050 ;
        RECT 784.950 289.950 787.050 292.050 ;
        RECT 787.950 289.950 790.050 292.050 ;
        RECT 785.400 288.900 786.600 289.650 ;
        RECT 784.950 286.800 787.050 288.900 ;
        RECT 775.950 265.950 778.050 268.050 ;
        RECT 787.950 265.950 790.050 268.050 ;
        RECT 773.400 259.350 774.600 261.600 ;
        RECT 778.950 260.100 781.050 262.200 ;
        RECT 779.400 259.350 780.600 260.100 ;
        RECT 772.950 256.950 775.050 259.050 ;
        RECT 775.950 256.950 778.050 259.050 ;
        RECT 778.950 256.950 781.050 259.050 ;
        RECT 781.950 256.950 784.050 259.050 ;
        RECT 776.400 255.900 777.600 256.650 ;
        RECT 782.400 255.900 783.600 256.650 ;
        RECT 788.400 255.900 789.450 265.950 ;
        RECT 775.950 253.800 778.050 255.900 ;
        RECT 781.950 253.800 784.050 255.900 ;
        RECT 787.950 253.800 790.050 255.900 ;
        RECT 769.950 244.950 772.050 247.050 ;
        RECT 770.400 205.050 771.450 244.950 ;
        RECT 794.400 244.050 795.450 364.950 ;
        RECT 799.950 364.800 802.050 366.900 ;
        RECT 806.400 365.400 807.600 367.650 ;
        RECT 806.400 355.050 807.450 365.400 ;
        RECT 805.950 352.950 808.050 355.050 ;
        RECT 812.400 346.050 813.450 382.950 ;
        RECT 818.400 373.200 819.450 415.950 ;
        RECT 821.400 388.050 822.450 416.100 ;
        RECT 827.400 415.350 828.600 416.100 ;
        RECT 826.950 412.950 829.050 415.050 ;
        RECT 829.950 412.950 832.050 415.050 ;
        RECT 830.400 410.400 831.600 412.650 ;
        RECT 836.400 411.900 837.450 424.950 ;
        RECT 830.400 406.050 831.450 410.400 ;
        RECT 835.950 409.800 838.050 411.900 ;
        RECT 829.950 403.950 832.050 406.050 ;
        RECT 839.400 391.050 840.450 430.950 ;
        RECT 841.950 416.100 844.050 418.200 ;
        RECT 848.400 417.600 849.450 430.950 ;
        RECT 842.400 406.050 843.450 416.100 ;
        RECT 848.400 415.350 849.600 417.600 ;
        RECT 853.950 416.100 856.050 418.200 ;
        RECT 854.400 415.350 855.600 416.100 ;
        RECT 847.950 412.950 850.050 415.050 ;
        RECT 850.950 412.950 853.050 415.050 ;
        RECT 853.950 412.950 856.050 415.050 ;
        RECT 856.950 412.950 859.050 415.050 ;
        RECT 851.400 411.900 852.600 412.650 ;
        RECT 857.400 411.900 858.600 412.650 ;
        RECT 850.950 406.950 853.050 411.900 ;
        RECT 856.950 409.800 859.050 411.900 ;
        RECT 841.950 403.950 844.050 406.050 ;
        RECT 838.950 388.950 841.050 391.050 ;
        RECT 820.950 385.950 823.050 388.050 ;
        RECT 826.950 385.950 829.050 388.050 ;
        RECT 820.950 376.950 823.050 379.050 ;
        RECT 817.950 372.450 820.050 373.200 ;
        RECT 815.400 371.400 820.050 372.450 ;
        RECT 815.400 366.900 816.450 371.400 ;
        RECT 817.950 371.100 820.050 371.400 ;
        RECT 821.400 372.600 822.450 376.950 ;
        RECT 827.400 372.600 828.450 385.950 ;
        RECT 835.950 382.950 838.050 385.050 ;
        RECT 821.400 370.350 822.600 372.600 ;
        RECT 827.400 370.350 828.600 372.600 ;
        RECT 820.950 367.950 823.050 370.050 ;
        RECT 823.950 367.950 826.050 370.050 ;
        RECT 826.950 367.950 829.050 370.050 ;
        RECT 829.950 367.950 832.050 370.050 ;
        RECT 824.400 366.900 825.600 367.650 ;
        RECT 814.950 364.800 817.050 366.900 ;
        RECT 823.950 364.800 826.050 366.900 ;
        RECT 830.400 366.000 831.600 367.650 ;
        RECT 829.950 361.950 832.050 366.000 ;
        RECT 836.400 349.050 837.450 382.950 ;
        RECT 839.400 379.050 840.450 388.950 ;
        RECT 838.950 376.950 841.050 379.050 ;
        RECT 844.950 376.950 847.050 379.050 ;
        RECT 845.400 372.600 846.450 376.950 ;
        RECT 845.400 370.350 846.600 372.600 ;
        RECT 850.950 371.100 853.050 373.200 ;
        RECT 851.400 370.350 852.600 371.100 ;
        RECT 859.950 370.950 862.050 376.050 ;
        RECT 844.950 367.950 847.050 370.050 ;
        RECT 847.950 367.950 850.050 370.050 ;
        RECT 850.950 367.950 853.050 370.050 ;
        RECT 853.950 367.950 856.050 370.050 ;
        RECT 841.950 364.950 844.050 367.050 ;
        RECT 848.400 365.400 849.600 367.650 ;
        RECT 854.400 366.900 855.600 367.650 ;
        RECT 842.400 358.050 843.450 364.950 ;
        RECT 841.950 355.950 844.050 358.050 ;
        RECT 848.400 355.050 849.450 365.400 ;
        RECT 853.950 364.800 856.050 366.900 ;
        RECT 863.400 361.050 864.450 466.950 ;
        RECT 866.400 450.600 867.450 484.950 ;
        RECT 872.400 475.050 873.450 488.400 ;
        RECT 875.400 481.050 876.450 497.400 ;
        RECT 878.400 490.050 879.450 499.950 ;
        RECT 877.950 487.950 880.050 490.050 ;
        RECT 877.950 484.800 880.050 486.900 ;
        RECT 874.950 478.950 877.050 481.050 ;
        RECT 871.950 472.950 874.050 475.050 ;
        RECT 866.400 448.350 867.600 450.600 ;
        RECT 874.950 449.100 877.050 451.200 ;
        RECT 875.400 448.350 876.600 449.100 ;
        RECT 866.100 445.950 868.200 448.050 ;
        RECT 869.400 445.950 871.500 448.050 ;
        RECT 874.800 445.950 876.900 448.050 ;
        RECT 869.400 443.400 870.600 445.650 ;
        RECT 865.950 427.950 868.050 430.050 ;
        RECT 866.400 411.900 867.450 427.950 ;
        RECT 869.400 427.050 870.450 443.400 ;
        RECT 878.400 442.050 879.450 484.800 ;
        RECT 881.400 445.050 882.450 511.950 ;
        RECT 884.400 508.050 885.450 514.950 ;
        RECT 889.950 508.950 892.050 511.050 ;
        RECT 883.950 505.950 886.050 508.050 ;
        RECT 890.400 495.600 891.450 508.950 ;
        RECT 899.400 504.450 900.450 520.950 ;
        RECT 902.400 514.050 903.450 527.100 ;
        RECT 914.400 526.350 915.600 528.600 ;
        RECT 919.950 527.100 922.050 529.200 ;
        RECT 920.400 526.350 921.600 527.100 ;
        RECT 910.950 523.950 913.050 526.050 ;
        RECT 913.950 523.950 916.050 526.050 ;
        RECT 916.950 523.950 919.050 526.050 ;
        RECT 919.950 523.950 922.050 526.050 ;
        RECT 911.400 521.400 912.600 523.650 ;
        RECT 917.400 522.900 918.600 523.650 ;
        RECT 901.950 511.950 904.050 514.050 ;
        RECT 907.950 511.950 910.050 514.050 ;
        RECT 899.400 503.400 903.450 504.450 ;
        RECT 890.400 493.350 891.600 495.600 ;
        RECT 895.950 494.100 898.050 496.200 ;
        RECT 896.400 493.350 897.600 494.100 ;
        RECT 902.400 493.050 903.450 503.400 ;
        RECT 904.950 499.950 907.050 502.050 ;
        RECT 886.950 490.950 889.050 493.050 ;
        RECT 889.950 490.950 892.050 493.050 ;
        RECT 892.950 490.950 895.050 493.050 ;
        RECT 895.950 490.950 898.050 493.050 ;
        RECT 901.950 490.950 904.050 493.050 ;
        RECT 887.400 489.900 888.600 490.650 ;
        RECT 886.950 487.800 889.050 489.900 ;
        RECT 893.400 488.400 894.600 490.650 ;
        RECT 883.950 484.950 886.050 487.050 ;
        RECT 880.950 442.950 883.050 445.050 ;
        RECT 877.950 439.950 880.050 442.050 ;
        RECT 884.400 430.050 885.450 484.950 ;
        RECT 887.400 481.050 888.450 487.800 ;
        RECT 886.950 478.950 889.050 481.050 ;
        RECT 893.400 478.050 894.450 488.400 ;
        RECT 901.950 487.800 904.050 489.900 ;
        RECT 892.950 475.950 895.050 478.050 ;
        RECT 893.400 469.050 894.450 475.950 ;
        RECT 895.950 469.950 898.050 472.050 ;
        RECT 892.950 466.950 895.050 469.050 ;
        RECT 886.950 460.950 889.050 463.050 ;
        RECT 887.400 451.050 888.450 460.950 ;
        RECT 889.950 454.950 892.050 457.050 ;
        RECT 886.950 448.950 889.050 451.050 ;
        RECT 890.400 450.600 891.450 454.950 ;
        RECT 896.400 451.200 897.450 469.950 ;
        RECT 902.400 463.050 903.450 487.800 ;
        RECT 901.950 460.950 904.050 463.050 ;
        RECT 890.400 448.350 891.600 450.600 ;
        RECT 895.950 449.100 898.050 451.200 ;
        RECT 896.400 448.350 897.600 449.100 ;
        RECT 889.950 445.950 892.050 448.050 ;
        RECT 892.950 445.950 895.050 448.050 ;
        RECT 895.950 445.950 898.050 448.050 ;
        RECT 898.950 445.950 901.050 448.050 ;
        RECT 886.950 442.950 889.050 445.050 ;
        RECT 893.400 444.000 894.600 445.650 ;
        RECT 874.950 427.950 877.050 430.050 ;
        RECT 883.950 427.950 886.050 430.050 ;
        RECT 868.950 424.950 871.050 427.050 ;
        RECT 875.400 417.600 876.450 427.950 ;
        RECT 875.400 415.350 876.600 417.600 ;
        RECT 880.950 416.100 883.050 418.200 ;
        RECT 881.400 415.350 882.600 416.100 ;
        RECT 871.950 412.950 874.050 415.050 ;
        RECT 874.950 412.950 877.050 415.050 ;
        RECT 877.950 412.950 880.050 415.050 ;
        RECT 880.950 412.950 883.050 415.050 ;
        RECT 865.950 409.800 868.050 411.900 ;
        RECT 872.400 411.000 873.600 412.650 ;
        RECT 871.950 406.950 874.050 411.000 ;
        RECT 878.400 410.400 879.600 412.650 ;
        RECT 887.400 411.450 888.450 442.950 ;
        RECT 889.950 439.950 892.050 442.050 ;
        RECT 892.950 439.950 895.050 444.000 ;
        RECT 899.400 443.400 900.600 445.650 ;
        RECT 905.400 444.900 906.450 499.950 ;
        RECT 908.400 496.050 909.450 511.950 ;
        RECT 911.400 502.050 912.450 521.400 ;
        RECT 916.950 520.800 919.050 522.900 ;
        RECT 922.950 520.950 925.050 523.050 ;
        RECT 926.400 522.900 927.450 556.950 ;
        RECT 928.950 541.950 931.050 544.050 ;
        RECT 916.950 505.950 919.050 508.050 ;
        RECT 910.950 499.950 913.050 502.050 ;
        RECT 907.950 493.950 910.050 496.050 ;
        RECT 910.950 494.100 913.050 496.200 ;
        RECT 917.400 495.600 918.450 505.950 ;
        RECT 923.400 496.050 924.450 520.950 ;
        RECT 925.950 520.800 928.050 522.900 ;
        RECT 926.400 511.050 927.450 520.800 ;
        RECT 925.950 508.950 928.050 511.050 ;
        RECT 926.400 505.050 927.450 508.950 ;
        RECT 925.950 502.950 928.050 505.050 ;
        RECT 925.950 496.950 928.050 499.050 ;
        RECT 911.400 493.350 912.600 494.100 ;
        RECT 917.400 493.350 918.600 495.600 ;
        RECT 922.950 493.950 925.050 496.050 ;
        RECT 910.950 490.950 913.050 493.050 ;
        RECT 913.950 490.950 916.050 493.050 ;
        RECT 916.950 490.950 919.050 493.050 ;
        RECT 919.950 490.950 922.050 493.050 ;
        RECT 907.950 487.950 910.050 490.050 ;
        RECT 914.400 489.000 915.600 490.650 ;
        RECT 920.400 489.900 921.600 490.650 ;
        RECT 926.400 490.050 927.450 496.950 ;
        RECT 908.400 472.050 909.450 487.950 ;
        RECT 913.950 484.950 916.050 489.000 ;
        RECT 919.950 487.800 922.050 489.900 ;
        RECT 925.950 487.950 928.050 490.050 ;
        RECT 920.400 472.050 921.450 487.800 ;
        RECT 925.950 484.800 928.050 486.900 ;
        RECT 907.950 469.950 910.050 472.050 ;
        RECT 919.950 469.950 922.050 472.050 ;
        RECT 907.950 460.950 910.050 463.050 ;
        RECT 884.400 410.400 888.450 411.450 ;
        RECT 878.400 406.050 879.450 410.400 ;
        RECT 877.950 403.950 880.050 406.050 ;
        RECT 868.950 388.950 871.050 391.050 ;
        RECT 865.950 379.950 868.050 382.050 ;
        RECT 866.400 376.050 867.450 379.950 ;
        RECT 865.950 373.950 868.050 376.050 ;
        RECT 869.400 372.600 870.450 388.950 ;
        RECT 874.950 382.950 877.050 385.050 ;
        RECT 871.950 373.950 874.050 379.050 ;
        RECT 875.400 372.600 876.450 382.950 ;
        RECT 869.400 370.350 870.600 372.600 ;
        RECT 875.400 370.350 876.600 372.600 ;
        RECT 868.950 367.950 871.050 370.050 ;
        RECT 871.950 367.950 874.050 370.050 ;
        RECT 874.950 367.950 877.050 370.050 ;
        RECT 877.950 367.950 880.050 370.050 ;
        RECT 872.400 365.400 873.600 367.650 ;
        RECT 878.400 365.400 879.600 367.650 ;
        RECT 865.950 361.950 868.050 364.050 ;
        RECT 862.950 358.950 865.050 361.050 ;
        RECT 866.400 357.450 867.450 361.950 ;
        RECT 863.400 356.400 867.450 357.450 ;
        RECT 847.950 352.950 850.050 355.050 ;
        RECT 835.950 346.950 838.050 349.050 ;
        RECT 859.950 346.950 862.050 349.050 ;
        RECT 811.950 343.950 814.050 346.050 ;
        RECT 802.950 339.000 805.050 343.050 ;
        RECT 803.400 337.350 804.600 339.000 ;
        RECT 808.950 338.100 811.050 340.200 ;
        RECT 809.400 337.350 810.600 338.100 ;
        RECT 820.950 337.950 823.050 340.050 ;
        RECT 829.950 338.100 832.050 340.200 ;
        RECT 837.000 339.600 841.050 340.050 ;
        RECT 799.950 334.950 802.050 337.050 ;
        RECT 802.950 334.950 805.050 337.050 ;
        RECT 805.950 334.950 808.050 337.050 ;
        RECT 808.950 334.950 811.050 337.050 ;
        RECT 800.400 332.400 801.600 334.650 ;
        RECT 806.400 333.900 807.600 334.650 ;
        RECT 800.400 310.050 801.450 332.400 ;
        RECT 805.950 331.800 808.050 333.900 ;
        RECT 799.950 307.950 802.050 310.050 ;
        RECT 817.950 307.950 820.050 310.050 ;
        RECT 805.950 298.950 808.050 301.050 ;
        RECT 806.400 294.600 807.450 298.950 ;
        RECT 806.400 292.350 807.600 294.600 ;
        RECT 811.950 293.100 814.050 295.200 ;
        RECT 812.400 292.350 813.600 293.100 ;
        RECT 802.950 289.950 805.050 292.050 ;
        RECT 805.950 289.950 808.050 292.050 ;
        RECT 808.950 289.950 811.050 292.050 ;
        RECT 811.950 289.950 814.050 292.050 ;
        RECT 803.400 287.400 804.600 289.650 ;
        RECT 809.400 288.000 810.600 289.650 ;
        RECT 803.400 283.050 804.450 287.400 ;
        RECT 808.950 283.950 811.050 288.000 ;
        RECT 818.400 286.050 819.450 307.950 ;
        RECT 821.400 307.050 822.450 337.950 ;
        RECT 830.400 337.350 831.600 338.100 ;
        RECT 836.400 337.950 841.050 339.600 ;
        RECT 841.950 338.100 844.050 340.200 ;
        RECT 836.400 337.350 837.600 337.950 ;
        RECT 826.950 334.950 829.050 337.050 ;
        RECT 829.950 334.950 832.050 337.050 ;
        RECT 832.950 334.950 835.050 337.050 ;
        RECT 835.950 334.950 838.050 337.050 ;
        RECT 827.400 333.900 828.600 334.650 ;
        RECT 826.950 331.800 829.050 333.900 ;
        RECT 833.400 332.400 834.600 334.650 ;
        RECT 826.950 325.950 829.050 328.050 ;
        RECT 827.400 322.050 828.450 325.950 ;
        RECT 833.400 322.050 834.450 332.400 ;
        RECT 838.950 331.950 841.050 334.050 ;
        RECT 835.950 328.950 838.050 331.050 ;
        RECT 826.950 319.950 829.050 322.050 ;
        RECT 832.950 319.950 835.050 322.050 ;
        RECT 820.950 304.950 823.050 307.050 ;
        RECT 827.400 294.600 828.450 319.950 ;
        RECT 836.400 316.050 837.450 328.950 ;
        RECT 835.950 313.950 838.050 316.050 ;
        RECT 839.400 301.050 840.450 331.950 ;
        RECT 842.400 310.050 843.450 338.100 ;
        RECT 844.950 337.950 847.050 340.050 ;
        RECT 853.950 338.100 856.050 340.200 ;
        RECT 860.400 339.600 861.450 346.950 ;
        RECT 863.400 342.450 864.450 356.400 ;
        RECT 872.400 355.050 873.450 365.400 ;
        RECT 871.950 352.950 874.050 355.050 ;
        RECT 871.950 349.800 874.050 351.900 ;
        RECT 865.950 343.950 871.050 346.050 ;
        RECT 872.400 343.050 873.450 349.800 ;
        RECT 874.950 343.950 877.050 349.050 ;
        RECT 878.400 348.450 879.450 365.400 ;
        RECT 880.950 364.950 883.050 367.050 ;
        RECT 881.400 358.050 882.450 364.950 ;
        RECT 880.950 355.950 883.050 358.050 ;
        RECT 884.400 352.050 885.450 410.400 ;
        RECT 886.950 406.950 889.050 409.050 ;
        RECT 887.400 364.050 888.450 406.950 ;
        RECT 890.400 397.050 891.450 439.950 ;
        RECT 892.950 430.950 895.050 433.050 ;
        RECT 893.400 409.050 894.450 430.950 ;
        RECT 899.400 421.050 900.450 443.400 ;
        RECT 904.950 442.800 907.050 444.900 ;
        RECT 908.400 424.050 909.450 460.950 ;
        RECT 919.950 454.950 922.050 457.050 ;
        RECT 913.950 449.100 916.050 451.200 ;
        RECT 920.400 450.600 921.450 454.950 ;
        RECT 926.400 451.050 927.450 484.800 ;
        RECT 914.400 448.350 915.600 449.100 ;
        RECT 920.400 448.350 921.600 450.600 ;
        RECT 925.950 448.950 928.050 451.050 ;
        RECT 913.950 445.950 916.050 448.050 ;
        RECT 916.950 445.950 919.050 448.050 ;
        RECT 919.950 445.950 922.050 448.050 ;
        RECT 922.950 445.950 925.050 448.050 ;
        RECT 917.400 444.900 918.600 445.650 ;
        RECT 923.400 444.900 924.600 445.650 ;
        RECT 916.950 442.800 919.050 444.900 ;
        RECT 922.950 442.800 925.050 444.900 ;
        RECT 929.400 439.050 930.450 541.950 ;
        RECT 931.950 527.100 934.050 529.200 ;
        RECT 935.400 529.050 936.450 560.400 ;
        RECT 941.400 544.050 942.450 577.950 ;
        RECT 944.400 568.050 945.450 592.950 ;
        RECT 950.400 586.050 951.450 599.400 ;
        RECT 952.950 598.950 955.050 601.050 ;
        RECT 955.950 598.950 958.050 601.050 ;
        RECT 959.400 600.900 960.450 628.950 ;
        RECT 949.950 583.950 952.050 586.050 ;
        RECT 953.400 582.450 954.450 598.950 ;
        RECT 958.950 598.800 961.050 600.900 ;
        RECT 962.400 586.050 963.450 631.950 ;
        RECT 965.400 631.050 966.450 641.400 ;
        RECT 967.950 637.950 970.050 640.050 ;
        RECT 964.950 628.950 967.050 631.050 ;
        RECT 968.400 625.050 969.450 637.950 ;
        RECT 971.400 634.050 972.450 661.950 ;
        RECT 970.950 631.950 973.050 634.050 ;
        RECT 974.400 631.050 975.450 670.950 ;
        RECT 977.400 670.050 978.450 721.950 ;
        RECT 980.400 709.050 981.450 733.950 ;
        RECT 983.400 723.900 984.450 733.950 ;
        RECT 986.400 730.050 987.450 826.950 ;
        RECT 988.950 811.950 991.050 814.050 ;
        RECT 989.400 772.050 990.450 811.950 ;
        RECT 992.400 808.050 993.450 826.950 ;
        RECT 995.400 814.050 996.450 850.950 ;
        RECT 998.400 817.050 999.450 862.950 ;
        RECT 1003.950 850.950 1006.050 853.050 ;
        RECT 1004.400 840.600 1005.450 850.950 ;
        RECT 1010.400 841.050 1011.450 874.950 ;
        RECT 1004.400 838.350 1005.600 840.600 ;
        RECT 1009.950 838.950 1012.050 841.050 ;
        RECT 1003.950 835.950 1006.050 838.050 ;
        RECT 1006.950 835.950 1009.050 838.050 ;
        RECT 1007.400 833.400 1008.600 835.650 ;
        RECT 1007.400 829.050 1008.450 833.400 ;
        RECT 1009.950 832.950 1012.050 835.050 ;
        RECT 1006.950 826.950 1009.050 829.050 ;
        RECT 1010.400 825.450 1011.450 832.950 ;
        RECT 1007.400 824.400 1011.450 825.450 ;
        RECT 997.950 814.950 1000.050 817.050 ;
        RECT 994.950 811.950 997.050 814.050 ;
        RECT 998.400 810.450 999.450 814.950 ;
        RECT 998.400 809.400 1002.450 810.450 ;
        RECT 991.950 805.950 994.050 808.050 ;
        RECT 994.950 806.100 997.050 808.200 ;
        RECT 1001.400 807.600 1002.450 809.400 ;
        RECT 1007.400 808.050 1008.450 824.400 ;
        RECT 1009.950 820.950 1012.050 823.050 ;
        RECT 995.400 805.350 996.600 806.100 ;
        RECT 1001.400 805.350 1002.600 807.600 ;
        RECT 1006.950 805.950 1009.050 808.050 ;
        RECT 994.950 802.950 997.050 805.050 ;
        RECT 997.950 802.950 1000.050 805.050 ;
        RECT 1000.950 802.950 1003.050 805.050 ;
        RECT 1003.950 802.950 1006.050 805.050 ;
        RECT 991.950 799.950 994.050 802.050 ;
        RECT 998.400 800.400 999.600 802.650 ;
        RECT 1004.400 801.000 1005.600 802.650 ;
        RECT 988.950 769.950 991.050 772.050 ;
        RECT 992.400 769.050 993.450 799.950 ;
        RECT 998.400 793.050 999.450 800.400 ;
        RECT 1003.950 796.950 1006.050 801.000 ;
        RECT 1006.950 799.950 1009.050 802.050 ;
        RECT 1007.400 793.050 1008.450 799.950 ;
        RECT 1010.400 799.050 1011.450 820.950 ;
        RECT 1009.950 796.950 1012.050 799.050 ;
        RECT 1013.400 795.450 1014.450 878.400 ;
        RECT 1010.400 794.400 1014.450 795.450 ;
        RECT 997.950 790.950 1000.050 793.050 ;
        RECT 1006.950 790.950 1009.050 793.050 ;
        RECT 1006.950 769.950 1009.050 772.050 ;
        RECT 991.950 766.950 994.050 769.050 ;
        RECT 997.950 766.950 1000.050 769.050 ;
        RECT 991.950 761.100 994.050 763.200 ;
        RECT 998.400 762.600 999.450 766.950 ;
        RECT 992.400 760.350 993.600 761.100 ;
        RECT 998.400 760.350 999.600 762.600 ;
        RECT 991.950 757.950 994.050 760.050 ;
        RECT 994.950 757.950 997.050 760.050 ;
        RECT 997.950 757.950 1000.050 760.050 ;
        RECT 1000.950 757.950 1003.050 760.050 ;
        RECT 995.400 755.400 996.600 757.650 ;
        RECT 1001.400 755.400 1002.600 757.650 ;
        RECT 995.400 736.050 996.450 755.400 ;
        RECT 1001.400 751.050 1002.450 755.400 ;
        RECT 1003.950 754.950 1006.050 757.050 ;
        RECT 1000.950 748.950 1003.050 751.050 ;
        RECT 1000.950 742.950 1003.050 745.050 ;
        RECT 994.950 733.950 997.050 736.050 ;
        RECT 985.950 727.950 988.050 730.050 ;
        RECT 991.950 728.100 994.050 730.200 ;
        RECT 992.400 727.350 993.600 728.100 ;
        RECT 997.950 727.950 1000.050 733.050 ;
        RECT 988.950 724.950 991.050 727.050 ;
        RECT 991.950 724.950 994.050 727.050 ;
        RECT 994.950 724.950 997.050 727.050 ;
        RECT 982.950 721.800 985.050 723.900 ;
        RECT 985.950 721.950 988.050 724.050 ;
        RECT 989.400 723.000 990.600 724.650 ;
        RECT 995.400 723.900 996.600 724.650 ;
        RECT 979.950 706.950 982.050 709.050 ;
        RECT 986.400 703.050 987.450 721.950 ;
        RECT 988.950 718.950 991.050 723.000 ;
        RECT 994.800 721.800 996.900 723.900 ;
        RECT 997.950 721.950 1000.050 724.050 ;
        RECT 989.400 712.050 990.450 718.950 ;
        RECT 994.950 718.650 997.050 720.750 ;
        RECT 995.400 715.050 996.450 718.650 ;
        RECT 994.950 712.950 997.050 715.050 ;
        RECT 988.950 709.950 991.050 712.050 ;
        RECT 979.950 700.950 982.050 703.050 ;
        RECT 985.950 700.950 988.050 703.050 ;
        RECT 980.400 685.050 981.450 700.950 ;
        RECT 988.950 691.950 991.050 694.050 ;
        RECT 979.800 682.950 981.900 685.050 ;
        RECT 982.950 683.100 985.050 685.200 ;
        RECT 989.400 684.600 990.450 691.950 ;
        RECT 983.400 682.350 984.600 683.100 ;
        RECT 989.400 682.350 990.600 684.600 ;
        RECT 982.950 679.950 985.050 682.050 ;
        RECT 985.950 679.950 988.050 682.050 ;
        RECT 988.950 679.950 991.050 682.050 ;
        RECT 991.950 679.950 994.050 682.050 ;
        RECT 979.950 676.950 982.050 679.050 ;
        RECT 986.400 678.900 987.600 679.650 ;
        RECT 980.400 673.050 981.450 676.950 ;
        RECT 985.950 676.800 988.050 678.900 ;
        RECT 992.400 678.450 993.600 679.650 ;
        RECT 998.400 678.450 999.450 721.950 ;
        RECT 992.400 677.400 999.450 678.450 ;
        RECT 985.950 673.650 988.050 675.750 ;
        RECT 988.950 673.950 991.050 676.050 ;
        RECT 991.950 673.950 994.050 676.050 ;
        RECT 997.950 673.950 1000.050 676.050 ;
        RECT 979.950 670.950 982.050 673.050 ;
        RECT 976.950 667.950 979.050 670.050 ;
        RECT 976.950 658.950 979.050 661.050 ;
        RECT 977.400 652.050 978.450 658.950 ;
        RECT 982.950 655.950 985.050 658.050 ;
        RECT 976.950 649.950 979.050 652.050 ;
        RECT 983.400 651.600 984.450 655.950 ;
        RECT 986.400 655.050 987.450 673.650 ;
        RECT 989.400 667.050 990.450 673.950 ;
        RECT 988.950 664.950 991.050 667.050 ;
        RECT 992.400 661.050 993.450 673.950 ;
        RECT 994.950 670.950 997.050 673.050 ;
        RECT 991.950 658.950 994.050 661.050 ;
        RECT 985.950 652.950 988.050 655.050 ;
        RECT 983.400 649.350 984.600 651.600 ;
        RECT 988.950 650.100 991.050 652.200 ;
        RECT 989.400 649.350 990.600 650.100 ;
        RECT 979.950 646.950 982.050 649.050 ;
        RECT 982.950 646.950 985.050 649.050 ;
        RECT 985.950 646.950 988.050 649.050 ;
        RECT 988.950 646.950 991.050 649.050 ;
        RECT 980.400 645.900 981.600 646.650 ;
        RECT 979.950 643.800 982.050 645.900 ;
        RECT 986.400 644.400 987.600 646.650 ;
        RECT 995.400 645.450 996.450 670.950 ;
        RECT 992.400 644.400 996.450 645.450 ;
        RECT 998.400 645.450 999.450 673.950 ;
        RECT 1001.400 652.050 1002.450 742.950 ;
        RECT 1004.400 724.050 1005.450 754.950 ;
        RECT 1003.950 721.950 1006.050 724.050 ;
        RECT 1003.950 703.950 1006.050 706.050 ;
        RECT 1004.400 676.050 1005.450 703.950 ;
        RECT 1003.950 673.950 1006.050 676.050 ;
        RECT 1007.400 655.050 1008.450 769.950 ;
        RECT 1010.400 673.050 1011.450 794.400 ;
        RECT 1012.950 790.950 1015.050 793.050 ;
        RECT 1013.400 691.050 1014.450 790.950 ;
        RECT 1012.950 688.950 1015.050 691.050 ;
        RECT 1009.950 670.950 1012.050 673.050 ;
        RECT 1009.950 664.950 1012.050 667.050 ;
        RECT 1006.950 652.950 1009.050 655.050 ;
        RECT 1000.950 649.950 1003.050 652.050 ;
        RECT 1003.950 650.100 1006.050 652.200 ;
        RECT 1010.400 651.600 1011.450 664.950 ;
        RECT 1016.400 652.050 1017.450 881.400 ;
        RECT 1004.400 649.350 1005.600 650.100 ;
        RECT 1010.400 649.350 1011.600 651.600 ;
        RECT 1015.950 649.950 1018.050 652.050 ;
        RECT 1003.950 646.950 1006.050 649.050 ;
        RECT 1006.950 646.950 1009.050 649.050 ;
        RECT 1009.950 646.950 1012.050 649.050 ;
        RECT 1012.950 646.950 1015.050 649.050 ;
        RECT 1007.400 645.900 1008.600 646.650 ;
        RECT 998.400 644.400 1002.450 645.450 ;
        RECT 979.950 640.650 982.050 642.750 ;
        RECT 982.950 640.950 985.050 643.050 ;
        RECT 973.950 628.950 976.050 631.050 ;
        RECT 967.950 622.950 970.050 625.050 ;
        RECT 980.400 622.050 981.450 640.650 ;
        RECT 970.950 619.950 973.050 622.050 ;
        RECT 979.950 619.950 982.050 622.050 ;
        RECT 971.400 606.600 972.450 619.950 ;
        RECT 979.950 613.950 982.050 616.050 ;
        RECT 971.400 604.350 972.600 606.600 ;
        RECT 976.950 605.100 979.050 607.200 ;
        RECT 980.400 607.050 981.450 613.950 ;
        RECT 977.400 604.350 978.600 605.100 ;
        RECT 979.950 604.950 982.050 607.050 ;
        RECT 967.950 601.950 970.050 604.050 ;
        RECT 970.950 601.950 973.050 604.050 ;
        RECT 973.950 601.950 976.050 604.050 ;
        RECT 976.950 601.950 979.050 604.050 ;
        RECT 964.950 598.950 967.050 601.050 ;
        RECT 968.400 600.900 969.600 601.650 ;
        RECT 965.400 595.050 966.450 598.950 ;
        RECT 967.950 598.800 970.050 600.900 ;
        RECT 974.400 599.400 975.600 601.650 ;
        RECT 970.950 595.950 973.050 598.050 ;
        RECT 964.950 592.950 967.050 595.050 ;
        RECT 967.950 589.950 970.050 592.050 ;
        RECT 961.950 583.950 964.050 586.050 ;
        RECT 950.400 581.400 954.450 582.450 ;
        RECT 950.400 574.050 951.450 581.400 ;
        RECT 946.950 571.950 949.050 574.050 ;
        RECT 949.950 571.950 952.050 574.050 ;
        RECT 952.950 572.100 955.050 574.200 ;
        RECT 958.950 573.000 961.050 577.050 ;
        RECT 943.950 565.950 946.050 568.050 ;
        RECT 947.400 565.050 948.450 571.950 ;
        RECT 953.400 571.350 954.600 572.100 ;
        RECT 959.400 571.350 960.600 573.000 ;
        RECT 952.950 568.950 955.050 571.050 ;
        RECT 955.950 568.950 958.050 571.050 ;
        RECT 958.950 568.950 961.050 571.050 ;
        RECT 961.950 568.950 964.050 571.050 ;
        RECT 949.950 565.950 952.050 568.050 ;
        RECT 956.400 566.400 957.600 568.650 ;
        RECT 962.400 567.900 963.600 568.650 ;
        RECT 946.950 562.950 949.050 565.050 ;
        RECT 946.950 550.950 949.050 553.050 ;
        RECT 940.950 541.950 943.050 544.050 ;
        RECT 943.950 535.950 946.050 538.050 ;
        RECT 940.950 532.950 943.050 535.050 ;
        RECT 932.400 496.050 933.450 527.100 ;
        RECT 934.950 526.950 937.050 529.050 ;
        RECT 941.400 528.600 942.450 532.950 ;
        RECT 944.400 529.050 945.450 535.950 ;
        RECT 941.400 526.350 942.600 528.600 ;
        RECT 943.950 526.950 946.050 529.050 ;
        RECT 937.950 523.950 940.050 526.050 ;
        RECT 940.950 523.950 943.050 526.050 ;
        RECT 938.400 521.400 939.600 523.650 ;
        RECT 947.400 523.050 948.450 550.950 ;
        RECT 938.400 519.450 939.450 521.400 ;
        RECT 943.950 520.950 946.050 523.050 ;
        RECT 946.950 520.950 949.050 523.050 ;
        RECT 938.400 518.400 942.450 519.450 ;
        RECT 937.950 502.950 940.050 505.050 ;
        RECT 931.950 493.950 934.050 496.050 ;
        RECT 938.400 495.600 939.450 502.950 ;
        RECT 941.400 499.050 942.450 518.400 ;
        RECT 944.400 502.050 945.450 520.950 ;
        RECT 950.400 514.050 951.450 565.950 ;
        RECT 952.950 550.950 955.050 553.050 ;
        RECT 953.400 529.050 954.450 550.950 ;
        RECT 956.400 550.050 957.450 566.400 ;
        RECT 961.950 562.950 964.050 567.900 ;
        RECT 968.400 562.050 969.450 589.950 ;
        RECT 967.950 559.950 970.050 562.050 ;
        RECT 967.950 556.800 970.050 558.900 ;
        RECT 955.950 547.950 958.050 550.050 ;
        RECT 958.950 532.950 961.050 535.050 ;
        RECT 964.950 532.950 967.050 535.050 ;
        RECT 952.950 526.950 955.050 529.050 ;
        RECT 959.400 528.600 960.450 532.950 ;
        RECT 965.400 528.600 966.450 532.950 ;
        RECT 968.400 529.050 969.450 556.800 ;
        RECT 959.400 526.350 960.600 528.600 ;
        RECT 965.400 526.350 966.600 528.600 ;
        RECT 967.950 526.950 970.050 529.050 ;
        RECT 955.950 523.950 958.050 526.050 ;
        RECT 958.950 523.950 961.050 526.050 ;
        RECT 961.950 523.950 964.050 526.050 ;
        RECT 964.950 523.950 967.050 526.050 ;
        RECT 956.400 523.050 957.600 523.650 ;
        RECT 952.950 521.400 957.600 523.050 ;
        RECT 962.400 521.400 963.600 523.650 ;
        RECT 952.950 520.950 957.000 521.400 ;
        RECT 955.950 517.950 958.050 520.050 ;
        RECT 949.950 511.950 952.050 514.050 ;
        RECT 949.950 505.950 952.050 508.050 ;
        RECT 943.950 499.950 946.050 502.050 ;
        RECT 940.950 498.450 943.050 499.050 ;
        RECT 940.950 497.400 945.450 498.450 ;
        RECT 940.950 496.950 943.050 497.400 ;
        RECT 944.400 495.600 945.450 497.400 ;
        RECT 938.400 493.350 939.600 495.600 ;
        RECT 944.400 493.350 945.600 495.600 ;
        RECT 934.950 490.950 937.050 493.050 ;
        RECT 937.950 490.950 940.050 493.050 ;
        RECT 940.950 490.950 943.050 493.050 ;
        RECT 943.950 490.950 946.050 493.050 ;
        RECT 935.400 488.400 936.600 490.650 ;
        RECT 941.400 489.900 942.600 490.650 ;
        RECT 950.400 490.050 951.450 505.950 ;
        RECT 952.950 496.950 955.050 499.050 ;
        RECT 935.400 478.050 936.450 488.400 ;
        RECT 940.950 487.800 943.050 489.900 ;
        RECT 946.950 487.950 949.050 490.050 ;
        RECT 949.950 487.950 952.050 490.050 ;
        RECT 941.400 481.050 942.450 487.800 ;
        RECT 940.950 478.950 943.050 481.050 ;
        RECT 934.950 475.950 937.050 478.050 ;
        RECT 947.400 457.050 948.450 487.950 ;
        RECT 953.400 463.050 954.450 496.950 ;
        RECT 956.400 496.050 957.450 517.950 ;
        RECT 962.400 502.050 963.450 521.400 ;
        RECT 971.400 520.050 972.450 595.950 ;
        RECT 974.400 577.050 975.450 599.400 ;
        RECT 983.400 598.050 984.450 640.950 ;
        RECT 986.400 631.050 987.450 644.400 ;
        RECT 985.950 628.950 988.050 631.050 ;
        RECT 992.400 628.050 993.450 644.400 ;
        RECT 997.950 640.950 1000.050 643.050 ;
        RECT 994.950 637.950 997.050 640.050 ;
        RECT 985.950 625.800 988.050 627.900 ;
        RECT 991.950 625.950 994.050 628.050 ;
        RECT 982.950 595.950 985.050 598.050 ;
        RECT 986.400 592.050 987.450 625.800 ;
        RECT 995.400 624.450 996.450 637.950 ;
        RECT 998.400 633.450 999.450 640.950 ;
        RECT 1001.400 637.050 1002.450 644.400 ;
        RECT 1006.950 643.800 1009.050 645.900 ;
        RECT 1013.400 644.400 1014.600 646.650 ;
        RECT 1007.400 642.450 1008.450 643.800 ;
        RECT 1004.400 641.400 1008.450 642.450 ;
        RECT 1000.950 634.950 1003.050 637.050 ;
        RECT 998.400 632.400 1002.450 633.450 ;
        RECT 997.950 624.450 1000.050 625.050 ;
        RECT 995.400 623.400 1000.050 624.450 ;
        RECT 997.950 622.950 1000.050 623.400 ;
        RECT 991.950 610.950 994.050 613.050 ;
        RECT 992.400 607.200 993.450 610.950 ;
        RECT 991.950 605.100 994.050 607.200 ;
        RECT 998.400 606.600 999.450 622.950 ;
        RECT 1001.400 609.450 1002.450 632.400 ;
        RECT 1004.400 613.050 1005.450 641.400 ;
        RECT 1009.950 640.950 1012.050 643.050 ;
        RECT 1006.950 634.950 1009.050 637.050 ;
        RECT 1003.950 610.950 1006.050 613.050 ;
        RECT 1001.400 609.000 1005.450 609.450 ;
        RECT 1001.400 608.400 1006.050 609.000 ;
        RECT 992.400 604.350 993.600 605.100 ;
        RECT 998.400 604.350 999.600 606.600 ;
        RECT 1003.950 604.950 1006.050 608.400 ;
        RECT 991.950 601.950 994.050 604.050 ;
        RECT 994.950 601.950 997.050 604.050 ;
        RECT 997.950 601.950 1000.050 604.050 ;
        RECT 1000.950 601.950 1003.050 604.050 ;
        RECT 988.950 597.450 991.050 601.050 ;
        RECT 995.400 599.400 996.600 601.650 ;
        RECT 1001.400 599.400 1002.600 601.650 ;
        RECT 988.950 597.000 993.450 597.450 ;
        RECT 989.400 596.400 993.450 597.000 ;
        RECT 985.950 589.950 988.050 592.050 ;
        RECT 988.950 586.950 991.050 589.050 ;
        RECT 976.950 580.950 979.050 583.050 ;
        RECT 973.950 574.950 976.050 577.050 ;
        RECT 977.400 573.600 978.450 580.950 ;
        RECT 977.400 571.350 978.600 573.600 ;
        RECT 982.950 573.000 985.050 577.050 ;
        RECT 989.400 574.050 990.450 586.950 ;
        RECT 983.400 571.350 984.600 573.000 ;
        RECT 988.950 571.950 991.050 574.050 ;
        RECT 976.950 568.950 979.050 571.050 ;
        RECT 979.950 568.950 982.050 571.050 ;
        RECT 982.950 568.950 985.050 571.050 ;
        RECT 985.950 568.950 988.050 571.050 ;
        RECT 980.400 567.900 981.600 568.650 ;
        RECT 979.950 565.800 982.050 567.900 ;
        RECT 986.400 566.400 987.600 568.650 ;
        RECT 992.400 567.450 993.450 596.400 ;
        RECT 995.400 586.050 996.450 599.400 ;
        RECT 997.950 595.950 1000.050 598.050 ;
        RECT 994.950 583.950 997.050 586.050 ;
        RECT 998.400 582.450 999.450 595.950 ;
        RECT 989.400 566.400 993.450 567.450 ;
        RECT 995.400 581.400 999.450 582.450 ;
        RECT 986.400 564.450 987.450 566.400 ;
        RECT 983.400 563.400 987.450 564.450 ;
        RECT 973.950 559.950 976.050 562.050 ;
        RECT 970.950 517.950 973.050 520.050 ;
        RECT 961.950 499.950 964.050 502.050 ;
        RECT 964.950 499.950 967.050 502.050 ;
        RECT 955.950 493.950 958.050 496.050 ;
        RECT 958.950 495.000 961.050 499.050 ;
        RECT 965.400 495.600 966.450 499.950 ;
        RECT 959.400 493.350 960.600 495.000 ;
        RECT 965.400 493.350 966.600 495.600 ;
        RECT 958.950 490.950 961.050 493.050 ;
        RECT 961.950 490.950 964.050 493.050 ;
        RECT 964.950 490.950 967.050 493.050 ;
        RECT 967.950 490.950 970.050 493.050 ;
        RECT 955.950 487.950 958.050 490.050 ;
        RECT 962.400 488.400 963.600 490.650 ;
        RECT 968.400 489.900 969.600 490.650 ;
        RECT 952.950 460.950 955.050 463.050 ;
        RECT 931.950 454.950 934.050 457.050 ;
        RECT 937.950 454.950 940.050 457.050 ;
        RECT 940.950 454.950 943.050 457.050 ;
        RECT 946.950 454.950 949.050 457.050 ;
        RECT 932.400 445.050 933.450 454.950 ;
        RECT 934.950 451.950 937.050 454.050 ;
        RECT 931.950 442.950 934.050 445.050 ;
        RECT 932.400 439.050 933.450 442.950 ;
        RECT 935.400 442.050 936.450 451.950 ;
        RECT 938.400 451.050 939.450 454.950 ;
        RECT 937.950 448.950 940.050 451.050 ;
        RECT 941.400 450.600 942.450 454.950 ;
        RECT 941.400 448.350 942.600 450.600 ;
        RECT 946.950 449.100 949.050 453.900 ;
        RECT 947.400 448.350 948.600 449.100 ;
        RECT 940.950 445.950 943.050 448.050 ;
        RECT 943.950 445.950 946.050 448.050 ;
        RECT 946.950 445.950 949.050 448.050 ;
        RECT 949.950 445.950 952.050 448.050 ;
        RECT 937.950 442.950 940.050 445.050 ;
        RECT 944.400 443.400 945.600 445.650 ;
        RECT 950.400 444.900 951.600 445.650 ;
        RECT 956.400 445.050 957.450 487.950 ;
        RECT 962.400 475.050 963.450 488.400 ;
        RECT 967.950 487.800 970.050 489.900 ;
        RECT 961.950 472.950 964.050 475.050 ;
        RECT 968.400 472.050 969.450 487.800 ;
        RECT 974.400 487.050 975.450 559.950 ;
        RECT 983.400 550.050 984.450 563.400 ;
        RECT 989.400 553.050 990.450 566.400 ;
        RECT 991.950 562.950 994.050 565.050 ;
        RECT 992.400 556.050 993.450 562.950 ;
        RECT 991.950 553.950 994.050 556.050 ;
        RECT 988.950 550.950 991.050 553.050 ;
        RECT 982.950 547.950 985.050 550.050 ;
        RECT 976.950 529.950 979.050 532.050 ;
        RECT 973.950 484.950 976.050 487.050 ;
        RECT 967.950 469.950 970.050 472.050 ;
        RECT 970.950 466.950 973.050 469.050 ;
        RECT 958.950 457.950 961.050 460.050 ;
        RECT 964.950 457.950 967.050 460.050 ;
        RECT 934.950 439.950 937.050 442.050 ;
        RECT 922.950 436.050 925.050 439.050 ;
        RECT 928.800 436.950 930.900 439.050 ;
        RECT 931.950 436.950 934.050 439.050 ;
        RECT 910.950 433.950 913.050 436.050 ;
        RECT 919.950 435.000 925.050 436.050 ;
        RECT 919.950 434.400 924.450 435.000 ;
        RECT 919.950 433.950 924.000 434.400 ;
        RECT 907.950 421.950 910.050 424.050 ;
        RECT 898.950 418.950 901.050 421.050 ;
        RECT 899.400 417.600 900.450 418.950 ;
        RECT 899.400 415.350 900.600 417.600 ;
        RECT 904.950 416.100 907.050 418.200 ;
        RECT 911.400 418.050 912.450 433.950 ;
        RECT 919.950 427.950 922.050 430.050 ;
        RECT 913.950 421.950 916.050 424.050 ;
        RECT 905.400 415.350 906.600 416.100 ;
        RECT 910.950 415.950 913.050 418.050 ;
        RECT 898.950 412.950 901.050 415.050 ;
        RECT 901.950 412.950 904.050 415.050 ;
        RECT 904.950 412.950 907.050 415.050 ;
        RECT 907.950 412.950 910.050 415.050 ;
        RECT 895.950 409.950 898.050 412.050 ;
        RECT 902.400 410.400 903.600 412.650 ;
        RECT 908.400 411.000 909.600 412.650 ;
        RECT 892.950 406.950 895.050 409.050 ;
        RECT 889.950 394.950 892.050 397.050 ;
        RECT 896.400 376.050 897.450 409.950 ;
        RECT 902.400 403.050 903.450 410.400 ;
        RECT 907.950 406.950 910.050 411.000 ;
        RECT 910.950 409.950 913.050 412.050 ;
        RECT 914.400 411.900 915.450 421.950 ;
        RECT 920.400 418.050 921.450 427.950 ;
        RECT 938.400 427.050 939.450 442.950 ;
        RECT 940.950 439.950 943.050 442.050 ;
        RECT 937.950 424.950 940.050 427.050 ;
        RECT 916.950 415.950 919.050 418.050 ;
        RECT 919.950 415.950 922.050 418.050 ;
        RECT 922.950 417.000 925.050 421.050 ;
        RECT 928.950 417.000 931.050 421.050 ;
        RECT 901.950 400.950 904.050 403.050 ;
        RECT 904.950 394.950 907.050 397.050 ;
        RECT 895.950 373.950 898.050 376.050 ;
        RECT 889.950 372.600 894.000 373.050 ;
        RECT 889.950 370.950 894.600 372.600 ;
        RECT 898.950 371.100 901.050 376.050 ;
        RECT 905.400 372.450 906.450 394.950 ;
        RECT 911.400 390.450 912.450 409.950 ;
        RECT 913.950 409.800 916.050 411.900 ;
        RECT 914.400 403.050 915.450 409.800 ;
        RECT 913.950 400.950 916.050 403.050 ;
        RECT 917.400 391.050 918.450 415.950 ;
        RECT 923.400 415.350 924.600 417.000 ;
        RECT 929.400 415.350 930.600 417.000 ;
        RECT 922.950 412.950 925.050 415.050 ;
        RECT 925.950 412.950 928.050 415.050 ;
        RECT 928.950 412.950 931.050 415.050 ;
        RECT 931.950 412.950 934.050 415.050 ;
        RECT 937.950 412.950 940.050 415.050 ;
        RECT 919.950 409.950 922.050 412.050 ;
        RECT 926.400 411.900 927.600 412.650 ;
        RECT 920.400 406.050 921.450 409.950 ;
        RECT 925.950 409.800 928.050 411.900 ;
        RECT 932.400 411.000 933.600 412.650 ;
        RECT 931.950 406.950 934.050 411.000 ;
        RECT 938.400 409.050 939.450 412.950 ;
        RECT 941.400 409.050 942.450 439.950 ;
        RECT 944.400 436.050 945.450 443.400 ;
        RECT 949.950 442.800 952.050 444.900 ;
        RECT 955.950 442.950 958.050 445.050 ;
        RECT 959.400 436.050 960.450 457.950 ;
        RECT 965.400 450.600 966.450 457.950 ;
        RECT 971.400 454.200 972.450 466.950 ;
        RECT 977.400 463.050 978.450 529.950 ;
        RECT 983.400 528.600 984.450 547.950 ;
        RECT 985.950 544.950 988.050 547.050 ;
        RECT 986.400 532.050 987.450 544.950 ;
        RECT 991.950 532.950 994.050 535.050 ;
        RECT 985.950 529.950 988.050 532.050 ;
        RECT 983.400 526.350 984.600 528.600 ;
        RECT 982.950 523.950 985.050 526.050 ;
        RECT 985.950 523.950 988.050 526.050 ;
        RECT 986.400 522.900 987.600 523.650 ;
        RECT 985.950 520.800 988.050 522.900 ;
        RECT 986.400 519.450 987.450 520.800 ;
        RECT 983.400 518.400 987.450 519.450 ;
        RECT 983.400 496.050 984.450 518.400 ;
        RECT 992.400 502.050 993.450 532.950 ;
        RECT 995.400 523.050 996.450 581.400 ;
        RECT 1001.400 576.450 1002.450 599.400 ;
        RECT 1003.950 598.950 1006.050 601.050 ;
        RECT 1004.400 589.050 1005.450 598.950 ;
        RECT 1003.950 586.950 1006.050 589.050 ;
        RECT 1003.950 580.950 1006.050 583.050 ;
        RECT 998.400 576.000 1002.450 576.450 ;
        RECT 997.950 575.400 1002.450 576.000 ;
        RECT 997.950 571.950 1000.050 575.400 ;
        RECT 1004.400 573.600 1005.450 580.950 ;
        RECT 1007.400 576.450 1008.450 634.950 ;
        RECT 1010.400 633.450 1011.450 640.950 ;
        RECT 1013.400 640.050 1014.450 644.400 ;
        RECT 1015.950 643.950 1018.050 646.050 ;
        RECT 1012.950 637.950 1015.050 640.050 ;
        RECT 1010.400 632.400 1014.450 633.450 ;
        RECT 1009.950 628.950 1012.050 631.050 ;
        RECT 1010.400 580.050 1011.450 628.950 ;
        RECT 1009.950 577.950 1012.050 580.050 ;
        RECT 1007.400 575.400 1011.450 576.450 ;
        RECT 1010.400 573.600 1011.450 575.400 ;
        RECT 1013.400 574.050 1014.450 632.400 ;
        RECT 1004.400 571.350 1005.600 573.600 ;
        RECT 1010.400 571.350 1011.600 573.600 ;
        RECT 1012.950 571.950 1015.050 574.050 ;
        RECT 1000.950 568.950 1003.050 571.050 ;
        RECT 1003.950 568.950 1006.050 571.050 ;
        RECT 1006.950 568.950 1009.050 571.050 ;
        RECT 1009.950 568.950 1012.050 571.050 ;
        RECT 997.950 565.800 1000.050 567.900 ;
        RECT 1001.400 567.000 1002.600 568.650 ;
        RECT 1007.400 567.900 1008.600 568.650 ;
        RECT 998.400 529.050 999.450 565.800 ;
        RECT 1000.950 562.950 1003.050 567.000 ;
        RECT 1006.950 565.800 1009.050 567.900 ;
        RECT 1012.950 565.950 1015.050 568.050 ;
        RECT 1009.950 553.950 1012.050 556.050 ;
        RECT 1003.950 532.950 1006.050 535.050 ;
        RECT 997.950 526.950 1000.050 529.050 ;
        RECT 1004.400 528.600 1005.450 532.950 ;
        RECT 1010.400 529.200 1011.450 553.950 ;
        RECT 1004.400 526.350 1005.600 528.600 ;
        RECT 1009.800 527.100 1011.900 529.200 ;
        RECT 1013.400 529.050 1014.450 565.950 ;
        RECT 1016.400 547.050 1017.450 643.950 ;
        RECT 1015.950 544.950 1018.050 547.050 ;
        RECT 1015.950 532.950 1018.050 535.050 ;
        RECT 1010.400 526.350 1011.600 527.100 ;
        RECT 1012.950 526.950 1015.050 529.050 ;
        RECT 1000.950 523.950 1003.050 526.050 ;
        RECT 1003.950 523.950 1006.050 526.050 ;
        RECT 1006.950 523.950 1009.050 526.050 ;
        RECT 1009.950 523.950 1012.050 526.050 ;
        RECT 994.950 520.950 997.050 523.050 ;
        RECT 1001.400 521.400 1002.600 523.650 ;
        RECT 1007.400 522.900 1008.600 523.650 ;
        RECT 997.950 517.950 1000.050 520.050 ;
        RECT 998.400 505.050 999.450 517.950 ;
        RECT 1001.400 508.050 1002.450 521.400 ;
        RECT 1006.950 520.800 1009.050 522.900 ;
        RECT 1016.400 522.450 1017.450 532.950 ;
        RECT 1013.400 521.400 1017.450 522.450 ;
        RECT 1003.950 517.950 1006.050 520.050 ;
        RECT 1009.800 517.950 1011.900 520.050 ;
        RECT 1004.400 510.450 1005.450 517.950 ;
        RECT 1004.400 509.400 1008.450 510.450 ;
        RECT 1000.950 505.950 1003.050 508.050 ;
        RECT 997.950 502.950 1000.050 505.050 ;
        RECT 1003.950 502.950 1006.050 505.050 ;
        RECT 991.950 499.950 994.050 502.050 ;
        RECT 1000.950 499.950 1003.050 502.050 ;
        RECT 982.950 493.950 985.050 496.050 ;
        RECT 988.950 495.000 991.050 499.050 ;
        RECT 989.400 493.350 990.600 495.000 ;
        RECT 994.950 494.100 997.050 496.200 ;
        RECT 995.400 493.350 996.600 494.100 ;
        RECT 979.950 490.950 982.050 493.050 ;
        RECT 985.950 490.950 988.050 493.050 ;
        RECT 988.950 490.950 991.050 493.050 ;
        RECT 991.950 490.950 994.050 493.050 ;
        RECT 994.950 490.950 997.050 493.050 ;
        RECT 976.950 460.950 979.050 463.050 ;
        RECT 980.400 460.050 981.450 490.950 ;
        RECT 982.950 487.950 985.050 490.050 ;
        RECT 986.400 489.900 987.600 490.650 ;
        RECT 979.950 457.950 982.050 460.050 ;
        RECT 976.950 454.950 979.050 457.050 ;
        RECT 970.950 452.100 973.050 454.200 ;
        RECT 977.400 451.200 978.450 454.950 ;
        RECT 979.950 451.950 982.050 454.050 ;
        RECT 965.400 448.350 966.600 450.600 ;
        RECT 970.950 448.950 973.050 451.050 ;
        RECT 976.950 449.100 979.050 451.200 ;
        RECT 971.400 448.350 972.600 448.950 ;
        RECT 964.950 445.950 967.050 448.050 ;
        RECT 967.950 445.950 970.050 448.050 ;
        RECT 970.950 445.950 973.050 448.050 ;
        RECT 973.950 445.950 976.050 448.050 ;
        RECT 961.950 442.950 964.050 445.050 ;
        RECT 968.400 443.400 969.600 445.650 ;
        RECT 974.400 443.400 975.600 445.650 ;
        RECT 943.950 433.950 946.050 436.050 ;
        RECT 952.950 433.950 955.050 436.050 ;
        RECT 958.950 433.950 961.050 436.050 ;
        RECT 943.950 417.600 948.000 418.050 ;
        RECT 953.400 417.600 954.450 433.950 ;
        RECT 943.950 415.950 948.600 417.600 ;
        RECT 947.400 415.350 948.600 415.950 ;
        RECT 953.400 415.350 954.600 417.600 ;
        RECT 946.950 412.950 949.050 415.050 ;
        RECT 949.950 412.950 952.050 415.050 ;
        RECT 952.950 412.950 955.050 415.050 ;
        RECT 955.950 412.950 958.050 415.050 ;
        RECT 943.950 409.950 946.050 412.050 ;
        RECT 950.400 411.900 951.600 412.650 ;
        RECT 934.950 406.950 937.050 409.050 ;
        RECT 937.950 406.950 940.050 409.050 ;
        RECT 940.950 406.950 943.050 409.050 ;
        RECT 919.950 403.950 922.050 406.050 ;
        RECT 911.400 389.400 915.450 390.450 ;
        RECT 910.950 385.950 913.050 388.050 ;
        RECT 907.950 382.950 910.050 385.050 ;
        RECT 908.400 379.050 909.450 382.950 ;
        RECT 907.950 376.950 910.050 379.050 ;
        RECT 905.400 371.400 909.450 372.450 ;
        RECT 893.400 370.350 894.600 370.950 ;
        RECT 899.400 370.350 900.600 371.100 ;
        RECT 892.950 367.950 895.050 370.050 ;
        RECT 895.950 367.950 898.050 370.050 ;
        RECT 898.950 367.950 901.050 370.050 ;
        RECT 901.950 367.950 904.050 370.050 ;
        RECT 896.400 365.400 897.600 367.650 ;
        RECT 902.400 366.900 903.600 367.650 ;
        RECT 886.950 361.950 889.050 364.050 ;
        RECT 883.950 349.950 886.050 352.050 ;
        RECT 878.400 347.400 882.450 348.450 ;
        RECT 863.400 341.400 867.450 342.450 ;
        RECT 845.400 331.050 846.450 337.950 ;
        RECT 854.400 337.350 855.600 338.100 ;
        RECT 860.400 337.350 861.600 339.600 ;
        RECT 850.950 334.950 853.050 337.050 ;
        RECT 853.950 334.950 856.050 337.050 ;
        RECT 856.950 334.950 859.050 337.050 ;
        RECT 859.950 334.950 862.050 337.050 ;
        RECT 851.400 333.000 852.600 334.650 ;
        RECT 844.950 328.950 847.050 331.050 ;
        RECT 850.950 328.950 853.050 333.000 ;
        RECT 857.400 332.400 858.600 334.650 ;
        RECT 853.950 330.450 856.050 331.050 ;
        RECT 857.400 330.450 858.450 332.400 ;
        RECT 853.950 329.400 858.450 330.450 ;
        RECT 853.950 328.950 856.050 329.400 ;
        RECT 844.950 310.950 847.050 313.050 ;
        RECT 841.950 307.950 844.050 310.050 ;
        RECT 838.950 298.950 841.050 301.050 ;
        RECT 827.400 292.350 828.600 294.600 ;
        RECT 835.950 294.450 838.050 295.200 ;
        RECT 835.950 293.400 840.450 294.450 ;
        RECT 835.950 293.100 838.050 293.400 ;
        RECT 836.400 292.350 837.600 293.100 ;
        RECT 827.100 289.950 829.200 292.050 ;
        RECT 830.400 289.950 832.500 292.050 ;
        RECT 835.800 289.950 837.900 292.050 ;
        RECT 830.400 288.900 831.600 289.650 ;
        RECT 829.950 286.800 832.050 288.900 ;
        RECT 839.400 286.050 840.450 293.400 ;
        RECT 817.950 283.950 820.050 286.050 ;
        RECT 838.950 283.950 841.050 286.050 ;
        RECT 802.950 280.950 805.050 283.050 ;
        RECT 799.950 277.950 802.050 280.050 ;
        RECT 800.400 261.600 801.450 277.950 ;
        RECT 817.950 265.950 820.050 268.050 ;
        RECT 800.400 259.350 801.600 261.600 ;
        RECT 808.950 259.950 811.050 262.050 ;
        RECT 818.400 261.600 819.450 265.950 ;
        RECT 845.400 262.200 846.450 310.950 ;
        RECT 854.400 294.600 855.450 328.950 ;
        RECT 854.400 292.350 855.600 294.600 ;
        RECT 850.950 289.950 853.050 292.050 ;
        RECT 853.950 289.950 856.050 292.050 ;
        RECT 856.950 289.950 859.050 292.050 ;
        RECT 851.400 287.400 852.600 289.650 ;
        RECT 857.400 288.900 858.600 289.650 ;
        RECT 851.400 286.050 852.450 287.400 ;
        RECT 856.950 286.800 859.050 288.900 ;
        RECT 866.400 286.050 867.450 341.400 ;
        RECT 871.950 340.950 874.050 343.050 ;
        RECT 872.400 333.900 873.450 340.950 ;
        RECT 881.400 339.600 882.450 347.400 ;
        RECT 896.400 342.450 897.450 365.400 ;
        RECT 901.950 364.800 904.050 366.900 ;
        RECT 908.400 358.050 909.450 371.400 ;
        RECT 911.400 361.050 912.450 385.950 ;
        RECT 914.400 373.050 915.450 389.400 ;
        RECT 916.950 388.950 919.050 391.050 ;
        RECT 931.950 379.950 934.050 382.050 ;
        RECT 925.950 376.950 928.050 379.050 ;
        RECT 913.950 370.950 916.050 373.050 ;
        RECT 919.950 372.000 922.050 376.050 ;
        RECT 926.400 372.600 927.450 376.950 ;
        RECT 920.400 370.350 921.600 372.000 ;
        RECT 926.400 370.350 927.600 372.600 ;
        RECT 916.950 367.950 919.050 370.050 ;
        RECT 919.950 367.950 922.050 370.050 ;
        RECT 922.950 367.950 925.050 370.050 ;
        RECT 925.950 367.950 928.050 370.050 ;
        RECT 913.950 364.950 916.050 367.050 ;
        RECT 917.400 366.900 918.600 367.650 ;
        RECT 910.950 358.950 913.050 361.050 ;
        RECT 898.950 355.950 901.050 358.050 ;
        RECT 907.950 355.950 910.050 358.050 ;
        RECT 893.400 341.400 897.450 342.450 ;
        RECT 881.400 337.350 882.600 339.600 ;
        RECT 886.950 338.100 889.050 340.200 ;
        RECT 887.400 337.350 888.600 338.100 ;
        RECT 877.950 334.950 880.050 337.050 ;
        RECT 880.950 334.950 883.050 337.050 ;
        RECT 883.950 334.950 886.050 337.050 ;
        RECT 886.950 334.950 889.050 337.050 ;
        RECT 878.400 333.900 879.600 334.650 ;
        RECT 871.950 331.800 874.050 333.900 ;
        RECT 877.950 331.800 880.050 333.900 ;
        RECT 884.400 333.000 885.600 334.650 ;
        RECT 883.950 328.950 886.050 333.000 ;
        RECT 889.950 331.950 892.050 334.050 ;
        RECT 874.950 304.950 877.050 307.050 ;
        RECT 875.400 295.200 876.450 304.950 ;
        RECT 880.950 298.950 883.050 301.050 ;
        RECT 874.950 293.100 877.050 295.200 ;
        RECT 881.400 294.600 882.450 298.950 ;
        RECT 875.400 292.350 876.600 293.100 ;
        RECT 881.400 292.350 882.600 294.600 ;
        RECT 874.950 289.950 877.050 292.050 ;
        RECT 877.950 289.950 880.050 292.050 ;
        RECT 880.950 289.950 883.050 292.050 ;
        RECT 878.400 287.400 879.600 289.650 ;
        RECT 850.950 285.450 853.050 286.050 ;
        RECT 850.950 284.400 855.450 285.450 ;
        RECT 850.950 283.950 853.050 284.400 ;
        RECT 799.950 256.950 802.050 259.050 ;
        RECT 802.950 256.950 805.050 259.050 ;
        RECT 803.400 255.900 804.600 256.650 ;
        RECT 802.950 253.800 805.050 255.900 ;
        RECT 809.400 244.050 810.450 259.950 ;
        RECT 818.400 259.350 819.600 261.600 ;
        RECT 832.950 259.950 835.050 262.050 ;
        RECT 838.950 260.100 841.050 262.200 ;
        RECT 844.950 260.100 847.050 262.200 ;
        RECT 817.950 256.950 820.050 259.050 ;
        RECT 820.950 256.950 823.050 259.050 ;
        RECT 829.950 256.950 832.050 259.050 ;
        RECT 821.400 255.000 822.600 256.650 ;
        RECT 820.950 250.950 823.050 255.000 ;
        RECT 830.400 250.050 831.450 256.950 ;
        RECT 829.950 247.950 832.050 250.050 ;
        RECT 793.950 241.950 796.050 244.050 ;
        RECT 808.950 241.950 811.050 244.050 ;
        RECT 802.950 238.950 805.050 241.050 ;
        RECT 796.950 223.950 799.050 226.050 ;
        RECT 778.950 215.100 781.050 217.200 ;
        RECT 797.400 216.600 798.450 223.950 ;
        RECT 803.400 220.050 804.450 238.950 ;
        RECT 814.950 232.950 817.050 235.050 ;
        RECT 811.950 220.950 814.050 223.050 ;
        RECT 802.950 217.950 805.050 220.050 ;
        RECT 803.400 216.600 804.450 217.950 ;
        RECT 779.400 214.350 780.600 215.100 ;
        RECT 797.400 214.350 798.600 216.600 ;
        RECT 803.400 214.350 804.600 216.600 ;
        RECT 778.950 211.950 781.050 214.050 ;
        RECT 781.950 211.950 784.050 214.050 ;
        RECT 796.950 211.950 799.050 214.050 ;
        RECT 799.950 211.950 802.050 214.050 ;
        RECT 802.950 211.950 805.050 214.050 ;
        RECT 805.950 211.950 808.050 214.050 ;
        RECT 782.400 209.400 783.600 211.650 ;
        RECT 800.400 209.400 801.600 211.650 ;
        RECT 806.400 210.000 807.600 211.650 ;
        RECT 772.950 205.950 775.050 208.050 ;
        RECT 769.950 202.950 772.050 205.050 ;
        RECT 766.950 199.950 769.050 202.050 ;
        RECT 773.400 184.050 774.450 205.950 ;
        RECT 782.400 199.050 783.450 209.400 ;
        RECT 781.950 196.950 784.050 199.050 ;
        RECT 790.950 196.950 793.050 199.050 ;
        RECT 752.400 181.350 753.600 183.600 ;
        RECT 758.400 181.350 759.600 183.600 ;
        RECT 764.400 181.350 765.600 183.600 ;
        RECT 772.950 181.950 775.050 184.050 ;
        RECT 781.950 182.100 784.050 184.200 ;
        RECT 782.400 181.350 783.600 182.100 ;
        RECT 751.950 178.950 754.050 181.050 ;
        RECT 754.950 178.950 757.050 181.050 ;
        RECT 757.950 178.950 760.050 181.050 ;
        RECT 760.950 178.950 763.050 181.050 ;
        RECT 763.950 178.950 766.050 181.050 ;
        RECT 779.100 178.950 781.200 181.050 ;
        RECT 782.400 178.950 784.500 181.050 ;
        RECT 787.800 178.950 789.900 181.050 ;
        RECT 755.400 176.400 756.600 178.650 ;
        RECT 761.400 177.900 762.600 178.650 ;
        RECT 779.400 177.900 780.600 178.650 ;
        RECT 788.400 177.900 789.600 178.650 ;
        RECT 755.400 166.050 756.450 176.400 ;
        RECT 760.950 175.800 763.050 177.900 ;
        RECT 778.950 175.800 781.050 177.900 ;
        RECT 787.950 175.800 790.050 177.900 ;
        RECT 757.950 172.950 760.050 175.050 ;
        RECT 745.950 163.950 748.050 166.050 ;
        RECT 754.950 163.950 757.050 166.050 ;
        RECT 758.400 151.050 759.450 172.950 ;
        RECT 791.400 169.050 792.450 196.950 ;
        RECT 793.950 182.100 796.050 184.200 ;
        RECT 800.400 183.450 801.450 209.400 ;
        RECT 805.950 205.950 808.050 210.000 ;
        RECT 812.400 202.050 813.450 220.950 ;
        RECT 805.950 199.950 808.050 202.050 ;
        RECT 811.950 199.950 814.050 202.050 ;
        RECT 797.400 182.400 801.450 183.450 ;
        RECT 806.400 183.600 807.450 199.950 ;
        RECT 790.950 166.950 793.050 169.050 ;
        RECT 763.950 157.950 766.050 160.050 ;
        RECT 790.950 157.950 793.050 160.050 ;
        RECT 764.400 154.050 765.450 157.950 ;
        RECT 763.950 151.950 766.050 154.050 ;
        RECT 757.950 148.950 760.050 151.050 ;
        RECT 742.950 139.950 745.050 142.050 ;
        RECT 748.950 139.950 751.050 142.050 ;
        RECT 739.950 137.100 742.050 139.200 ;
        RECT 740.400 136.350 741.600 137.100 ;
        RECT 739.950 133.950 742.050 136.050 ;
        RECT 742.950 133.950 745.050 136.050 ;
        RECT 743.400 132.900 744.600 133.650 ;
        RECT 733.950 130.800 736.050 132.900 ;
        RECT 742.950 130.800 745.050 132.900 ;
        RECT 742.950 121.950 745.050 124.050 ;
        RECT 730.950 118.950 733.050 121.050 ;
        RECT 736.950 118.950 739.050 121.050 ;
        RECT 730.950 104.100 733.050 106.200 ;
        RECT 737.400 105.600 738.450 118.950 ;
        RECT 731.400 103.350 732.600 104.100 ;
        RECT 737.400 103.350 738.600 105.600 ;
        RECT 727.950 100.950 730.050 103.050 ;
        RECT 730.950 100.950 733.050 103.050 ;
        RECT 733.950 100.950 736.050 103.050 ;
        RECT 736.950 100.950 739.050 103.050 ;
        RECT 724.950 97.950 727.050 100.050 ;
        RECT 728.400 99.000 729.600 100.650 ;
        RECT 734.400 99.900 735.600 100.650 ;
        RECT 743.400 99.900 744.450 121.950 ;
        RECT 745.950 106.950 748.050 109.050 ;
        RECT 721.950 94.950 724.050 97.050 ;
        RECT 718.950 85.950 721.050 88.050 ;
        RECT 697.950 82.950 700.050 85.050 ;
        RECT 655.950 59.100 658.050 61.200 ;
        RECT 661.950 60.000 664.050 63.900 ;
        RECT 670.950 61.950 673.050 64.050 ;
        RECT 656.400 58.350 657.600 59.100 ;
        RECT 662.400 58.350 663.600 60.000 ;
        RECT 655.950 55.950 658.050 58.050 ;
        RECT 658.950 55.950 661.050 58.050 ;
        RECT 661.950 55.950 664.050 58.050 ;
        RECT 664.950 55.950 667.050 58.050 ;
        RECT 659.400 54.900 660.600 55.650 ;
        RECT 643.950 49.950 646.050 52.050 ;
        RECT 646.950 49.950 649.050 52.050 ;
        RECT 649.950 49.950 652.050 52.050 ;
        RECT 652.950 49.950 655.050 54.900 ;
        RECT 658.950 52.800 661.050 54.900 ;
        RECT 665.400 53.400 666.600 55.650 ;
        RECT 616.950 46.950 619.050 49.050 ;
        RECT 619.950 42.450 622.050 43.050 ;
        RECT 614.400 41.400 622.050 42.450 ;
        RECT 614.400 34.050 615.450 41.400 ;
        RECT 619.950 40.950 622.050 41.400 ;
        RECT 616.950 37.950 619.050 40.050 ;
        RECT 613.950 31.950 616.050 34.050 ;
        RECT 598.950 28.950 601.050 31.050 ;
        RECT 581.400 25.350 582.600 27.000 ;
        RECT 587.400 25.350 588.600 27.600 ;
        RECT 604.950 26.100 607.050 28.200 ;
        RECT 610.950 27.000 613.050 31.050 ;
        RECT 617.400 28.050 618.450 37.950 ;
        RECT 634.950 34.950 637.050 37.050 ;
        RECT 619.950 28.950 622.050 31.050 ;
        RECT 605.400 25.350 606.600 26.100 ;
        RECT 611.400 25.350 612.600 27.000 ;
        RECT 616.950 25.950 619.050 28.050 ;
        RECT 620.400 25.050 621.450 28.950 ;
        RECT 622.950 25.950 625.050 28.050 ;
        RECT 628.950 26.100 631.050 28.200 ;
        RECT 635.400 27.600 636.450 34.950 ;
        RECT 580.950 22.950 583.050 25.050 ;
        RECT 583.950 22.950 586.050 25.050 ;
        RECT 586.950 22.950 589.050 25.050 ;
        RECT 589.950 22.950 592.050 25.050 ;
        RECT 604.950 22.950 607.050 25.050 ;
        RECT 607.950 22.950 610.050 25.050 ;
        RECT 610.950 22.950 613.050 25.050 ;
        RECT 613.950 22.950 616.050 25.050 ;
        RECT 619.950 22.950 622.050 25.050 ;
        RECT 584.400 21.900 585.600 22.650 ;
        RECT 547.950 19.800 550.050 21.900 ;
        RECT 553.950 19.800 556.050 21.900 ;
        RECT 559.950 19.800 562.050 21.900 ;
        RECT 574.950 19.800 577.050 21.900 ;
        RECT 583.950 19.800 586.050 21.900 ;
        RECT 590.400 20.400 591.600 22.650 ;
        RECT 608.400 20.400 609.600 22.650 ;
        RECT 614.400 21.900 615.600 22.650 ;
        RECT 544.950 16.950 547.050 19.050 ;
        RECT 590.400 16.050 591.450 20.400 ;
        RECT 608.400 16.050 609.450 20.400 ;
        RECT 613.950 19.800 616.050 21.900 ;
        RECT 589.950 13.950 592.050 16.050 ;
        RECT 607.950 13.950 610.050 16.050 ;
        RECT 481.950 10.950 484.050 13.050 ;
        RECT 505.950 10.950 508.050 13.050 ;
        RECT 529.950 10.950 532.050 13.050 ;
        RECT 623.400 7.050 624.450 25.950 ;
        RECT 629.400 25.350 630.600 26.100 ;
        RECT 635.400 25.350 636.600 27.600 ;
        RECT 628.950 22.950 631.050 25.050 ;
        RECT 631.950 22.950 634.050 25.050 ;
        RECT 634.950 22.950 637.050 25.050 ;
        RECT 637.950 22.950 640.050 25.050 ;
        RECT 632.400 21.900 633.600 22.650 ;
        RECT 631.950 19.800 634.050 21.900 ;
        RECT 638.400 21.000 639.600 22.650 ;
        RECT 637.950 16.950 640.050 21.000 ;
        RECT 644.400 19.050 645.450 49.950 ;
        RECT 658.800 40.950 660.900 43.050 ;
        RECT 661.950 40.950 664.050 43.050 ;
        RECT 659.400 34.050 660.450 40.950 ;
        RECT 658.950 31.950 661.050 34.050 ;
        RECT 646.950 28.950 649.050 31.050 ;
        RECT 643.950 16.950 646.050 19.050 ;
        RECT 647.400 13.050 648.450 28.950 ;
        RECT 652.950 27.000 655.050 31.050 ;
        RECT 653.400 25.350 654.600 27.000 ;
        RECT 652.950 22.950 655.050 25.050 ;
        RECT 655.950 22.950 658.050 25.050 ;
        RECT 656.400 21.900 657.600 22.650 ;
        RECT 655.950 19.800 658.050 21.900 ;
        RECT 658.950 16.950 661.050 22.050 ;
        RECT 662.400 21.900 663.450 40.950 ;
        RECT 665.400 40.050 666.450 53.400 ;
        RECT 671.400 43.050 672.450 61.950 ;
        RECT 673.950 59.100 676.050 61.200 ;
        RECT 679.950 59.100 682.050 61.200 ;
        RECT 685.950 60.000 688.050 64.050 ;
        RECT 670.950 40.950 673.050 43.050 ;
        RECT 674.400 40.050 675.450 59.100 ;
        RECT 680.400 58.350 681.600 59.100 ;
        RECT 686.400 58.350 687.600 60.000 ;
        RECT 679.950 55.950 682.050 58.050 ;
        RECT 682.950 55.950 685.050 58.050 ;
        RECT 685.950 55.950 688.050 58.050 ;
        RECT 688.950 55.950 691.050 58.050 ;
        RECT 683.400 53.400 684.600 55.650 ;
        RECT 689.400 53.400 690.600 55.650 ;
        RECT 698.400 54.450 699.450 82.950 ;
        RECT 722.400 82.050 723.450 94.950 ;
        RECT 721.950 79.950 724.050 82.050 ;
        RECT 725.400 70.050 726.450 97.950 ;
        RECT 727.950 94.950 730.050 99.000 ;
        RECT 733.950 97.800 736.050 99.900 ;
        RECT 742.950 97.800 745.050 99.900 ;
        RECT 746.400 94.050 747.450 106.950 ;
        RECT 745.950 91.950 748.050 94.050 ;
        RECT 724.950 67.950 727.050 70.050 ;
        RECT 706.950 64.950 709.050 67.050 ;
        RECT 707.400 61.200 708.450 64.950 ;
        RECT 706.950 59.100 709.050 61.200 ;
        RECT 712.950 59.100 715.050 61.200 ;
        RECT 725.400 60.450 726.450 67.950 ;
        RECT 730.500 63.300 732.600 65.400 ;
        RECT 740.100 64.500 742.200 66.600 ;
        RECT 728.400 60.450 729.600 60.600 ;
        RECT 725.400 59.400 729.600 60.450 ;
        RECT 707.400 58.350 708.600 59.100 ;
        RECT 713.400 58.350 714.600 59.100 ;
        RECT 728.400 58.350 729.600 59.400 ;
        RECT 703.950 55.950 706.050 58.050 ;
        RECT 706.950 55.950 709.050 58.050 ;
        RECT 709.950 55.950 712.050 58.050 ;
        RECT 712.950 55.950 715.050 58.050 ;
        RECT 724.950 55.950 727.050 58.050 ;
        RECT 728.100 55.950 730.200 58.050 ;
        RECT 704.400 54.450 705.600 55.650 ;
        RECT 698.400 53.400 705.600 54.450 ;
        RECT 710.400 53.400 711.600 55.650 ;
        RECT 664.950 37.950 667.050 40.050 ;
        RECT 673.950 37.950 676.050 40.050 ;
        RECT 664.950 31.950 667.050 34.050 ;
        RECT 661.950 19.800 664.050 21.900 ;
        RECT 665.400 19.050 666.450 31.950 ;
        RECT 667.950 25.950 670.050 31.050 ;
        RECT 674.400 27.600 675.450 37.950 ;
        RECT 683.400 34.050 684.450 53.400 ;
        RECT 689.400 34.050 690.450 53.400 ;
        RECT 700.950 49.950 703.050 52.050 ;
        RECT 682.950 31.950 685.050 34.050 ;
        RECT 688.950 31.950 691.050 34.050 ;
        RECT 674.400 25.350 675.600 27.600 ;
        RECT 679.950 26.100 682.050 28.200 ;
        RECT 680.400 25.350 681.600 26.100 ;
        RECT 691.950 25.950 694.050 28.050 ;
        RECT 701.400 27.600 702.450 49.950 ;
        RECT 706.950 34.950 709.050 37.050 ;
        RECT 707.400 27.600 708.450 34.950 ;
        RECT 710.400 28.050 711.450 53.400 ;
        RECT 715.950 34.950 718.050 37.050 ;
        RECT 670.950 22.950 673.050 25.050 ;
        RECT 673.950 22.950 676.050 25.050 ;
        RECT 676.950 22.950 679.050 25.050 ;
        RECT 679.950 22.950 682.050 25.050 ;
        RECT 671.400 21.900 672.600 22.650 ;
        RECT 670.950 19.800 673.050 21.900 ;
        RECT 677.400 21.000 678.600 22.650 ;
        RECT 664.950 16.950 667.050 19.050 ;
        RECT 676.950 16.950 679.050 21.000 ;
        RECT 692.400 16.050 693.450 25.950 ;
        RECT 701.400 25.350 702.600 27.600 ;
        RECT 707.400 25.350 708.600 27.600 ;
        RECT 709.950 25.950 712.050 28.050 ;
        RECT 697.950 22.950 700.050 25.050 ;
        RECT 700.950 22.950 703.050 25.050 ;
        RECT 703.950 22.950 706.050 25.050 ;
        RECT 706.950 22.950 709.050 25.050 ;
        RECT 698.400 21.900 699.600 22.650 ;
        RECT 704.400 21.900 705.600 22.650 ;
        RECT 697.950 19.800 700.050 21.900 ;
        RECT 703.950 19.800 706.050 21.900 ;
        RECT 716.400 16.050 717.450 34.950 ;
        RECT 725.400 34.050 726.450 55.950 ;
        RECT 731.400 54.300 732.300 63.300 ;
        RECT 733.800 59.700 735.900 61.800 ;
        RECT 737.400 61.350 738.600 63.600 ;
        RECT 735.000 57.300 735.900 59.700 ;
        RECT 736.800 58.950 738.900 61.050 ;
        RECT 740.700 57.300 741.900 64.500 ;
        RECT 749.400 61.200 750.450 139.950 ;
        RECT 758.400 139.200 759.450 148.950 ;
        RECT 751.950 136.950 754.050 139.050 ;
        RECT 757.950 137.100 760.050 139.200 ;
        RECT 764.400 138.600 765.450 151.950 ;
        RECT 791.400 138.600 792.450 157.950 ;
        RECT 752.400 132.900 753.450 136.950 ;
        RECT 758.400 136.350 759.600 137.100 ;
        RECT 764.400 136.350 765.600 138.600 ;
        RECT 782.400 138.450 783.600 138.600 ;
        RECT 779.400 137.400 783.600 138.450 ;
        RECT 757.950 133.950 760.050 136.050 ;
        RECT 760.950 133.950 763.050 136.050 ;
        RECT 763.950 133.950 766.050 136.050 ;
        RECT 751.950 130.800 754.050 132.900 ;
        RECT 761.400 131.400 762.600 133.650 ;
        RECT 754.950 105.000 757.050 109.050 ;
        RECT 761.400 105.450 762.450 131.400 ;
        RECT 775.950 112.950 778.050 115.050 ;
        RECT 766.950 106.950 769.050 112.050 ;
        RECT 755.400 103.350 756.600 105.000 ;
        RECT 761.400 104.400 765.450 105.450 ;
        RECT 754.950 100.950 757.050 103.050 ;
        RECT 757.950 100.950 760.050 103.050 ;
        RECT 758.400 98.400 759.600 100.650 ;
        RECT 758.400 97.050 759.450 98.400 ;
        RECT 758.400 95.400 763.050 97.050 ;
        RECT 759.000 94.950 763.050 95.400 ;
        RECT 764.400 88.050 765.450 104.400 ;
        RECT 767.400 99.900 768.450 106.950 ;
        RECT 776.400 105.600 777.450 112.950 ;
        RECT 779.400 109.050 780.450 137.400 ;
        RECT 782.400 136.350 783.600 137.400 ;
        RECT 791.400 136.350 792.600 138.600 ;
        RECT 782.100 133.950 784.200 136.050 ;
        RECT 785.400 133.950 787.500 136.050 ;
        RECT 790.800 133.950 792.900 136.050 ;
        RECT 785.400 132.900 786.600 133.650 ;
        RECT 784.950 130.800 787.050 132.900 ;
        RECT 778.950 106.950 781.050 109.050 ;
        RECT 776.400 103.350 777.600 105.600 ;
        RECT 781.950 104.100 784.050 106.200 ;
        RECT 794.400 106.050 795.450 182.100 ;
        RECT 797.400 160.050 798.450 182.400 ;
        RECT 806.400 181.350 807.600 183.600 ;
        RECT 802.950 178.950 805.050 181.050 ;
        RECT 805.950 178.950 808.050 181.050 ;
        RECT 808.950 178.950 811.050 181.050 ;
        RECT 803.400 177.900 804.600 178.650 ;
        RECT 802.950 175.800 805.050 177.900 ;
        RECT 809.400 176.400 810.600 178.650 ;
        RECT 799.950 163.950 802.050 166.050 ;
        RECT 796.950 157.950 799.050 160.050 ;
        RECT 796.950 151.950 799.050 154.050 ;
        RECT 782.400 103.350 783.600 104.100 ;
        RECT 787.950 103.950 790.050 106.050 ;
        RECT 793.950 103.950 796.050 106.050 ;
        RECT 797.400 105.600 798.450 151.950 ;
        RECT 800.400 118.050 801.450 163.950 ;
        RECT 803.400 163.050 804.450 175.800 ;
        RECT 809.400 169.050 810.450 176.400 ;
        RECT 808.950 166.950 811.050 169.050 ;
        RECT 802.950 160.950 805.050 163.050 ;
        RECT 815.400 138.600 816.450 232.950 ;
        RECT 833.400 229.050 834.450 259.950 ;
        RECT 839.400 259.350 840.600 260.100 ;
        RECT 845.400 259.350 846.600 260.100 ;
        RECT 838.950 256.950 841.050 259.050 ;
        RECT 841.950 256.950 844.050 259.050 ;
        RECT 844.950 256.950 847.050 259.050 ;
        RECT 847.950 256.950 850.050 259.050 ;
        RECT 842.400 255.000 843.600 256.650 ;
        RECT 841.950 250.950 844.050 255.000 ;
        RECT 848.400 254.400 849.600 256.650 ;
        RECT 848.400 253.050 849.450 254.400 ;
        RECT 847.950 247.950 850.050 253.050 ;
        RECT 841.950 229.950 844.050 232.050 ;
        RECT 817.950 226.950 820.050 229.050 ;
        RECT 832.950 226.950 835.050 229.050 ;
        RECT 818.400 205.050 819.450 226.950 ;
        RECT 838.950 223.950 841.050 226.050 ;
        RECT 826.950 216.000 829.050 220.050 ;
        RECT 827.400 214.350 828.600 216.000 ;
        RECT 832.950 215.100 835.050 217.200 ;
        RECT 833.400 214.350 834.600 215.100 ;
        RECT 823.950 211.950 826.050 214.050 ;
        RECT 826.950 211.950 829.050 214.050 ;
        RECT 829.950 211.950 832.050 214.050 ;
        RECT 832.950 211.950 835.050 214.050 ;
        RECT 824.400 209.400 825.600 211.650 ;
        RECT 830.400 209.400 831.600 211.650 ;
        RECT 824.400 205.050 825.450 209.400 ;
        RECT 817.950 202.950 820.050 205.050 ;
        RECT 823.950 202.950 826.050 205.050 ;
        RECT 817.950 199.800 820.050 201.900 ;
        RECT 818.400 139.050 819.450 199.800 ;
        RECT 830.400 187.050 831.450 209.400 ;
        RECT 839.400 208.050 840.450 223.950 ;
        RECT 838.950 205.950 841.050 208.050 ;
        RECT 838.950 193.950 841.050 196.050 ;
        RECT 832.950 187.950 835.050 190.050 ;
        RECT 829.950 186.450 832.050 187.050 ;
        RECT 827.400 185.400 832.050 186.450 ;
        RECT 827.400 183.600 828.450 185.400 ;
        RECT 829.950 184.950 832.050 185.400 ;
        RECT 833.400 183.600 834.450 187.950 ;
        RECT 827.400 181.350 828.600 183.600 ;
        RECT 833.400 181.350 834.600 183.600 ;
        RECT 823.950 178.950 826.050 181.050 ;
        RECT 826.950 178.950 829.050 181.050 ;
        RECT 829.950 178.950 832.050 181.050 ;
        RECT 832.950 178.950 835.050 181.050 ;
        RECT 824.400 176.400 825.600 178.650 ;
        RECT 830.400 177.000 831.600 178.650 ;
        RECT 824.400 172.050 825.450 176.400 ;
        RECT 829.950 172.950 832.050 177.000 ;
        RECT 823.950 169.950 826.050 172.050 ;
        RECT 839.400 169.050 840.450 193.950 ;
        RECT 842.400 177.900 843.450 229.950 ;
        RECT 854.400 223.050 855.450 284.400 ;
        RECT 856.950 283.650 859.050 285.750 ;
        RECT 865.950 283.950 868.050 286.050 ;
        RECT 857.400 255.450 858.450 283.650 ;
        RECT 878.400 277.050 879.450 287.400 ;
        RECT 890.400 283.050 891.450 331.950 ;
        RECT 893.400 331.050 894.450 341.400 ;
        RECT 899.400 340.050 900.450 355.950 ;
        RECT 914.400 348.450 915.450 364.950 ;
        RECT 916.950 364.800 919.050 366.900 ;
        RECT 923.400 365.400 924.600 367.650 ;
        RECT 923.400 361.050 924.450 365.400 ;
        RECT 928.950 364.950 931.050 367.050 ;
        RECT 922.950 358.950 925.050 361.050 ;
        RECT 916.950 349.950 919.050 352.050 ;
        RECT 911.400 347.400 915.450 348.450 ;
        RECT 901.950 343.950 904.050 346.050 ;
        RECT 895.950 337.950 898.050 340.050 ;
        RECT 898.950 337.950 901.050 340.050 ;
        RECT 902.400 339.600 903.450 343.950 ;
        RECT 892.950 328.950 895.050 331.050 ;
        RECT 896.400 322.050 897.450 337.950 ;
        RECT 902.400 337.350 903.600 339.600 ;
        RECT 907.950 338.100 910.050 340.200 ;
        RECT 911.400 340.050 912.450 347.400 ;
        RECT 913.950 343.950 916.050 346.050 ;
        RECT 908.400 337.350 909.600 338.100 ;
        RECT 910.950 337.950 913.050 340.050 ;
        RECT 901.950 334.950 904.050 337.050 ;
        RECT 904.950 334.950 907.050 337.050 ;
        RECT 907.950 334.950 910.050 337.050 ;
        RECT 905.400 332.400 906.600 334.650 ;
        RECT 905.400 328.050 906.450 332.400 ;
        RECT 904.950 325.950 907.050 328.050 ;
        RECT 895.950 319.950 898.050 322.050 ;
        RECT 895.950 298.950 898.050 301.050 ;
        RECT 904.950 300.450 907.050 301.050 ;
        RECT 904.950 299.400 909.450 300.450 ;
        RECT 904.950 298.950 907.050 299.400 ;
        RECT 892.950 292.950 895.050 295.050 ;
        RECT 896.400 294.600 897.450 298.950 ;
        RECT 905.400 294.600 906.450 298.950 ;
        RECT 893.400 288.900 894.450 292.950 ;
        RECT 896.400 292.350 897.600 294.600 ;
        RECT 905.400 292.350 906.600 294.600 ;
        RECT 896.100 289.950 898.200 292.050 ;
        RECT 901.500 289.950 903.600 292.050 ;
        RECT 904.800 289.950 906.900 292.050 ;
        RECT 902.400 288.900 903.600 289.650 ;
        RECT 892.950 286.800 895.050 288.900 ;
        RECT 901.950 286.800 904.050 288.900 ;
        RECT 889.950 280.950 892.050 283.050 ;
        RECT 901.950 280.950 904.050 283.050 ;
        RECT 877.950 276.450 880.050 277.050 ;
        RECT 877.950 275.400 882.450 276.450 ;
        RECT 877.950 274.950 880.050 275.400 ;
        RECT 877.950 265.950 880.050 268.050 ;
        RECT 865.950 260.100 868.050 262.200 ;
        RECT 871.950 260.100 874.050 262.200 ;
        RECT 866.400 259.350 867.600 260.100 ;
        RECT 872.400 259.350 873.600 260.100 ;
        RECT 862.950 256.950 865.050 259.050 ;
        RECT 865.950 256.950 868.050 259.050 ;
        RECT 868.950 256.950 871.050 259.050 ;
        RECT 871.950 256.950 874.050 259.050 ;
        RECT 857.400 254.400 861.450 255.450 ;
        RECT 863.400 255.000 864.600 256.650 ;
        RECT 869.400 255.000 870.600 256.650 ;
        RECT 856.950 232.950 859.050 235.050 ;
        RECT 853.950 220.950 856.050 223.050 ;
        RECT 850.950 215.100 853.050 217.200 ;
        RECT 851.400 214.350 852.600 215.100 ;
        RECT 847.950 211.950 850.050 214.050 ;
        RECT 850.950 211.950 853.050 214.050 ;
        RECT 848.400 210.000 849.600 211.650 ;
        RECT 847.950 205.950 850.050 210.000 ;
        RECT 857.400 202.050 858.450 232.950 ;
        RECT 850.950 199.950 853.050 202.050 ;
        RECT 856.950 199.950 859.050 202.050 ;
        RECT 851.400 187.050 852.450 199.950 ;
        RECT 850.950 183.000 853.050 187.050 ;
        RECT 851.400 181.350 852.600 183.000 ;
        RECT 856.950 182.100 859.050 184.200 ;
        RECT 860.400 184.050 861.450 254.400 ;
        RECT 862.950 250.950 865.050 255.000 ;
        RECT 868.950 250.950 871.050 255.000 ;
        RECT 874.950 253.950 877.050 256.050 ;
        RECT 868.950 215.100 871.050 217.200 ;
        RECT 875.400 216.600 876.450 253.950 ;
        RECT 878.400 235.050 879.450 265.950 ;
        RECT 877.950 232.950 880.050 235.050 ;
        RECT 869.400 214.350 870.600 215.100 ;
        RECT 875.400 214.350 876.600 216.600 ;
        RECT 865.950 211.950 868.050 214.050 ;
        RECT 868.950 211.950 871.050 214.050 ;
        RECT 871.950 211.950 874.050 214.050 ;
        RECT 874.950 211.950 877.050 214.050 ;
        RECT 866.400 209.400 867.600 211.650 ;
        RECT 872.400 210.900 873.600 211.650 ;
        RECT 866.400 205.050 867.450 209.400 ;
        RECT 871.950 208.800 874.050 210.900 ;
        RECT 865.950 202.950 868.050 205.050 ;
        RECT 862.950 199.950 865.050 202.050 ;
        RECT 857.400 181.350 858.600 182.100 ;
        RECT 859.950 181.950 862.050 184.050 ;
        RECT 847.950 178.950 850.050 181.050 ;
        RECT 850.950 178.950 853.050 181.050 ;
        RECT 853.950 178.950 856.050 181.050 ;
        RECT 856.950 178.950 859.050 181.050 ;
        RECT 841.950 175.800 844.050 177.900 ;
        RECT 848.400 176.400 849.600 178.650 ;
        RECT 854.400 177.900 855.600 178.650 ;
        RECT 848.400 172.050 849.450 176.400 ;
        RECT 853.950 175.800 856.050 177.900 ;
        RECT 859.950 175.950 862.050 178.050 ;
        RECT 847.950 169.950 850.050 172.050 ;
        RECT 838.950 166.950 841.050 169.050 ;
        RECT 860.400 166.050 861.450 175.950 ;
        RECT 863.400 172.050 864.450 199.950 ;
        RECT 881.400 196.050 882.450 275.400 ;
        RECT 895.950 271.950 898.050 274.050 ;
        RECT 896.400 268.050 897.450 271.950 ;
        RECT 895.950 265.950 898.050 268.050 ;
        RECT 889.950 260.100 892.050 262.200 ;
        RECT 896.400 261.600 897.450 265.950 ;
        RECT 890.400 259.350 891.600 260.100 ;
        RECT 896.400 259.350 897.600 261.600 ;
        RECT 886.950 256.950 889.050 259.050 ;
        RECT 889.950 256.950 892.050 259.050 ;
        RECT 892.950 256.950 895.050 259.050 ;
        RECT 895.950 256.950 898.050 259.050 ;
        RECT 887.400 254.400 888.600 256.650 ;
        RECT 893.400 254.400 894.600 256.650 ;
        RECT 887.400 253.050 888.450 254.400 ;
        RECT 886.950 250.950 889.050 253.050 ;
        RECT 883.950 241.950 886.050 244.050 ;
        RECT 884.400 214.050 885.450 241.950 ;
        RECT 887.400 226.050 888.450 250.950 ;
        RECT 893.400 244.050 894.450 254.400 ;
        RECT 892.950 241.950 895.050 244.050 ;
        RECT 902.400 241.050 903.450 280.950 ;
        RECT 908.400 261.450 909.450 299.400 ;
        RECT 914.400 271.050 915.450 343.950 ;
        RECT 917.400 307.050 918.450 349.950 ;
        RECT 922.950 339.000 925.050 343.050 ;
        RECT 929.400 340.050 930.450 364.950 ;
        RECT 932.400 364.050 933.450 379.950 ;
        RECT 931.950 361.950 934.050 364.050 ;
        RECT 931.950 358.800 934.050 360.900 ;
        RECT 923.400 337.350 924.600 339.000 ;
        RECT 928.950 337.950 931.050 340.050 ;
        RECT 922.950 334.950 925.050 337.050 ;
        RECT 925.950 334.950 928.050 337.050 ;
        RECT 919.950 331.950 922.050 334.050 ;
        RECT 926.400 333.900 927.600 334.650 ;
        RECT 932.400 334.050 933.450 358.800 ;
        RECT 916.950 304.950 919.050 307.050 ;
        RECT 920.400 304.050 921.450 331.950 ;
        RECT 925.950 331.800 928.050 333.900 ;
        RECT 931.950 331.950 934.050 334.050 ;
        RECT 931.950 328.800 934.050 330.900 ;
        RECT 932.400 322.050 933.450 328.800 ;
        RECT 935.400 325.050 936.450 406.950 ;
        RECT 938.400 361.050 939.450 406.950 ;
        RECT 944.400 379.050 945.450 409.950 ;
        RECT 949.950 409.800 952.050 411.900 ;
        RECT 956.400 411.000 957.600 412.650 ;
        RECT 955.950 406.950 958.050 411.000 ;
        RECT 958.950 409.950 961.050 412.050 ;
        RECT 952.950 405.900 957.000 406.050 ;
        RECT 952.950 403.950 958.050 405.900 ;
        RECT 955.950 403.800 958.050 403.950 ;
        RECT 949.950 385.950 952.050 388.050 ;
        RECT 943.950 376.950 946.050 379.050 ;
        RECT 943.950 371.100 946.050 373.200 ;
        RECT 950.400 372.600 951.450 385.950 ;
        RECT 944.400 370.350 945.600 371.100 ;
        RECT 950.400 370.350 951.600 372.600 ;
        RECT 943.950 367.950 946.050 370.050 ;
        RECT 946.950 367.950 949.050 370.050 ;
        RECT 949.950 367.950 952.050 370.050 ;
        RECT 952.950 367.950 955.050 370.050 ;
        RECT 947.400 366.000 948.600 367.650 ;
        RECT 946.950 361.950 949.050 366.000 ;
        RECT 953.400 365.400 954.600 367.650 ;
        RECT 937.950 358.950 940.050 361.050 ;
        RECT 946.950 352.950 949.050 355.050 ;
        RECT 943.950 349.950 946.050 352.050 ;
        RECT 944.400 339.600 945.450 349.950 ;
        RECT 947.400 346.050 948.450 352.950 ;
        RECT 953.400 349.050 954.450 365.400 ;
        RECT 959.400 355.050 960.450 409.950 ;
        RECT 962.400 400.050 963.450 442.950 ;
        RECT 964.950 439.950 967.050 442.050 ;
        RECT 965.400 412.050 966.450 439.950 ;
        RECT 968.400 436.050 969.450 443.400 ;
        RECT 974.400 439.050 975.450 443.400 ;
        RECT 980.400 439.050 981.450 451.950 ;
        RECT 983.400 442.050 984.450 487.950 ;
        RECT 985.950 487.800 988.050 489.900 ;
        RECT 992.400 488.400 993.600 490.650 ;
        RECT 985.950 484.650 988.050 486.750 ;
        RECT 982.950 439.950 985.050 442.050 ;
        RECT 973.950 436.950 976.050 439.050 ;
        RECT 979.950 436.950 982.050 439.050 ;
        RECT 967.950 433.950 970.050 436.050 ;
        RECT 968.400 418.050 969.450 433.950 ;
        RECT 979.950 433.800 982.050 435.900 ;
        RECT 970.950 427.950 973.050 430.050 ;
        RECT 971.400 421.050 972.450 427.950 ;
        RECT 973.950 421.950 976.050 424.050 ;
        RECT 970.950 418.950 973.050 421.050 ;
        RECT 974.400 418.200 975.450 421.950 ;
        RECT 967.950 415.950 970.050 418.050 ;
        RECT 973.950 416.100 976.050 418.200 ;
        RECT 974.400 415.350 975.600 416.100 ;
        RECT 970.950 412.950 973.050 415.050 ;
        RECT 973.950 412.950 976.050 415.050 ;
        RECT 964.950 409.950 967.050 412.050 ;
        RECT 971.400 411.900 972.600 412.650 ;
        RECT 970.950 409.800 973.050 411.900 ;
        RECT 964.950 400.950 967.050 406.050 ;
        RECT 961.950 397.950 964.050 400.050 ;
        RECT 961.950 388.950 964.050 391.050 ;
        RECT 962.400 364.050 963.450 388.950 ;
        RECT 970.950 376.950 973.050 379.050 ;
        RECT 971.400 373.200 972.450 376.950 ;
        RECT 976.950 375.450 979.050 376.050 ;
        RECT 980.400 375.450 981.450 433.800 ;
        RECT 986.400 430.050 987.450 484.650 ;
        RECT 992.400 475.050 993.450 488.400 ;
        RECT 1001.400 475.050 1002.450 499.950 ;
        RECT 991.950 472.950 994.050 475.050 ;
        RECT 1000.950 472.950 1003.050 475.050 ;
        RECT 997.950 454.950 1000.050 457.050 ;
        RECT 991.950 449.100 994.050 451.200 ;
        RECT 998.400 450.600 999.450 454.950 ;
        RECT 1004.400 451.050 1005.450 502.950 ;
        RECT 992.400 448.350 993.600 449.100 ;
        RECT 998.400 448.350 999.600 450.600 ;
        RECT 1003.950 448.950 1006.050 451.050 ;
        RECT 991.950 445.950 994.050 448.050 ;
        RECT 994.950 445.950 997.050 448.050 ;
        RECT 997.950 445.950 1000.050 448.050 ;
        RECT 1000.950 445.950 1003.050 448.050 ;
        RECT 988.950 442.950 991.050 445.050 ;
        RECT 995.400 443.400 996.600 445.650 ;
        RECT 1001.400 443.400 1002.600 445.650 ;
        RECT 1007.400 444.450 1008.450 509.400 ;
        RECT 1010.400 508.050 1011.450 517.950 ;
        RECT 1009.950 505.950 1012.050 508.050 ;
        RECT 1009.950 502.800 1012.050 504.900 ;
        RECT 1004.400 443.400 1008.450 444.450 ;
        RECT 985.950 429.450 988.050 430.050 ;
        RECT 976.950 374.400 981.450 375.450 ;
        RECT 983.400 428.400 988.050 429.450 ;
        RECT 970.950 371.100 973.050 373.200 ;
        RECT 976.950 372.000 979.050 374.400 ;
        RECT 971.400 370.350 972.600 371.100 ;
        RECT 977.400 370.350 978.600 372.000 ;
        RECT 967.950 367.950 970.050 370.050 ;
        RECT 970.950 367.950 973.050 370.050 ;
        RECT 973.950 367.950 976.050 370.050 ;
        RECT 976.950 367.950 979.050 370.050 ;
        RECT 964.950 364.950 967.050 367.050 ;
        RECT 968.400 365.400 969.600 367.650 ;
        RECT 974.400 366.000 975.600 367.650 ;
        RECT 961.950 361.950 964.050 364.050 ;
        RECT 958.950 352.950 961.050 355.050 ;
        RECT 955.950 349.950 958.050 352.050 ;
        RECT 952.950 348.450 955.050 349.050 ;
        RECT 950.400 347.400 955.050 348.450 ;
        RECT 946.950 343.950 949.050 346.050 ;
        RECT 950.400 340.050 951.450 347.400 ;
        RECT 952.950 346.950 955.050 347.400 ;
        RECT 956.400 342.450 957.450 349.950 ;
        RECT 965.400 346.050 966.450 364.950 ;
        RECT 964.950 343.950 967.050 346.050 ;
        RECT 968.400 343.200 969.450 365.400 ;
        RECT 973.950 361.950 976.050 366.000 ;
        RECT 979.950 363.450 982.050 367.050 ;
        RECT 977.400 363.000 982.050 363.450 ;
        RECT 977.400 362.400 981.450 363.000 ;
        RECT 953.400 341.400 957.450 342.450 ;
        RECT 944.400 337.350 945.600 339.600 ;
        RECT 949.950 337.950 952.050 340.050 ;
        RECT 940.950 334.950 943.050 337.050 ;
        RECT 943.950 334.950 946.050 337.050 ;
        RECT 946.950 334.950 949.050 337.050 ;
        RECT 937.950 331.950 940.050 334.050 ;
        RECT 941.400 333.000 942.600 334.650 ;
        RECT 947.400 333.900 948.600 334.650 ;
        RECT 953.400 333.900 954.450 341.400 ;
        RECT 967.950 341.100 970.050 343.200 ;
        RECT 955.950 337.950 958.050 340.050 ;
        RECT 961.950 338.100 964.050 340.200 ;
        RECT 974.400 340.050 975.450 361.950 ;
        RECT 934.950 322.950 937.050 325.050 ;
        RECT 931.950 319.950 934.050 322.050 ;
        RECT 919.950 301.950 922.050 304.050 ;
        RECT 916.950 293.100 919.050 295.200 ;
        RECT 925.950 293.100 928.050 295.200 ;
        RECT 931.950 293.100 934.050 295.200 ;
        RECT 917.400 288.450 918.450 293.100 ;
        RECT 926.400 292.350 927.600 293.100 ;
        RECT 932.400 292.350 933.600 293.100 ;
        RECT 922.950 289.950 925.050 292.050 ;
        RECT 925.950 289.950 928.050 292.050 ;
        RECT 928.950 289.950 931.050 292.050 ;
        RECT 931.950 289.950 934.050 292.050 ;
        RECT 917.400 287.400 921.450 288.450 ;
        RECT 913.950 268.950 916.050 271.050 ;
        RECT 905.400 260.400 909.450 261.450 ;
        RECT 901.950 238.950 904.050 241.050 ;
        RECT 905.400 232.050 906.450 260.400 ;
        RECT 913.950 260.100 916.050 262.200 ;
        RECT 920.400 261.600 921.450 287.400 ;
        RECT 923.400 287.400 924.600 289.650 ;
        RECT 929.400 288.900 930.600 289.650 ;
        RECT 923.400 277.050 924.450 287.400 ;
        RECT 928.950 286.800 931.050 288.900 ;
        RECT 938.400 286.050 939.450 331.950 ;
        RECT 940.950 328.950 943.050 333.000 ;
        RECT 946.950 331.800 949.050 333.900 ;
        RECT 952.950 331.800 955.050 333.900 ;
        RECT 943.950 325.950 946.050 328.050 ;
        RECT 940.950 322.950 943.050 325.050 ;
        RECT 941.400 289.050 942.450 322.950 ;
        RECT 940.950 286.950 943.050 289.050 ;
        RECT 937.950 283.950 940.050 286.050 ;
        RECT 922.950 274.950 925.050 277.050 ;
        RECT 928.950 268.950 931.050 271.050 ;
        RECT 914.400 259.350 915.600 260.100 ;
        RECT 920.400 259.350 921.600 261.600 ;
        RECT 925.950 259.950 928.050 262.050 ;
        RECT 910.950 256.950 913.050 259.050 ;
        RECT 913.950 256.950 916.050 259.050 ;
        RECT 916.950 256.950 919.050 259.050 ;
        RECT 919.950 256.950 922.050 259.050 ;
        RECT 911.400 254.400 912.600 256.650 ;
        RECT 917.400 255.000 918.600 256.650 ;
        RECT 911.400 244.050 912.450 254.400 ;
        RECT 916.950 250.950 919.050 255.000 ;
        RECT 910.950 241.950 913.050 244.050 ;
        RECT 910.950 232.950 913.050 235.050 ;
        RECT 904.950 229.950 907.050 232.050 ;
        RECT 886.950 223.950 889.050 226.050 ;
        RECT 895.950 223.950 898.050 226.050 ;
        RECT 896.400 216.600 897.450 223.950 ;
        RECT 907.950 220.950 910.050 223.050 ;
        RECT 896.400 214.350 897.600 216.600 ;
        RECT 901.950 215.100 904.050 217.200 ;
        RECT 902.400 214.350 903.600 215.100 ;
        RECT 883.950 211.950 886.050 214.050 ;
        RECT 892.950 211.950 895.050 214.050 ;
        RECT 895.950 211.950 898.050 214.050 ;
        RECT 898.950 211.950 901.050 214.050 ;
        RECT 901.950 211.950 904.050 214.050 ;
        RECT 893.400 209.400 894.600 211.650 ;
        RECT 899.400 210.900 900.600 211.650 ;
        RECT 908.400 210.900 909.450 220.950 ;
        RECT 886.950 202.950 889.050 205.050 ;
        RECT 874.950 193.950 877.050 196.050 ;
        RECT 880.950 193.950 883.050 196.050 ;
        RECT 865.950 187.950 868.050 190.050 ;
        RECT 862.950 169.950 865.050 172.050 ;
        RECT 859.950 163.950 862.050 166.050 ;
        RECT 859.950 151.950 862.050 154.050 ;
        RECT 841.950 145.950 844.050 148.050 ;
        RECT 815.400 136.350 816.600 138.600 ;
        RECT 817.950 136.950 820.050 139.050 ;
        RECT 823.950 137.100 826.050 139.200 ;
        RECT 833.400 138.450 834.600 138.600 ;
        RECT 827.400 137.400 834.600 138.450 ;
        RECT 808.950 133.950 811.050 136.050 ;
        RECT 811.950 133.950 814.050 136.050 ;
        RECT 814.950 133.950 817.050 136.050 ;
        RECT 812.400 132.900 813.600 133.650 ;
        RECT 824.400 133.050 825.450 137.100 ;
        RECT 811.950 130.800 814.050 132.900 ;
        RECT 823.950 130.950 826.050 133.050 ;
        RECT 827.400 124.050 828.450 137.400 ;
        RECT 833.400 136.350 834.600 137.400 ;
        RECT 832.950 133.950 835.050 136.050 ;
        RECT 835.950 133.950 838.050 136.050 ;
        RECT 836.400 132.900 837.600 133.650 ;
        RECT 842.400 132.900 843.450 145.950 ;
        RECT 853.950 137.100 856.050 139.200 ;
        RECT 860.400 138.600 861.450 151.950 ;
        RECT 854.400 136.350 855.600 137.100 ;
        RECT 860.400 136.350 861.600 138.600 ;
        RECT 850.950 133.950 853.050 136.050 ;
        RECT 853.950 133.950 856.050 136.050 ;
        RECT 856.950 133.950 859.050 136.050 ;
        RECT 859.950 133.950 862.050 136.050 ;
        RECT 835.950 130.800 838.050 132.900 ;
        RECT 841.950 130.800 844.050 132.900 ;
        RECT 851.400 131.400 852.600 133.650 ;
        RECT 857.400 132.900 858.600 133.650 ;
        RECT 838.950 124.950 841.050 127.050 ;
        RECT 826.950 121.950 829.050 124.050 ;
        RECT 799.950 115.950 802.050 118.050 ;
        RECT 829.950 115.950 832.050 118.050 ;
        RECT 772.950 100.950 775.050 103.050 ;
        RECT 775.950 100.950 778.050 103.050 ;
        RECT 778.950 100.950 781.050 103.050 ;
        RECT 781.950 100.950 784.050 103.050 ;
        RECT 773.400 99.900 774.600 100.650 ;
        RECT 766.950 97.800 769.050 99.900 ;
        RECT 772.950 97.800 775.050 99.900 ;
        RECT 779.400 99.000 780.600 100.650 ;
        RECT 778.950 94.950 781.050 99.000 ;
        RECT 784.950 97.800 787.050 99.900 ;
        RECT 785.400 91.050 786.450 97.800 ;
        RECT 788.400 94.050 789.450 103.950 ;
        RECT 797.400 103.350 798.600 105.600 ;
        RECT 802.950 104.100 805.050 106.200 ;
        RECT 811.950 104.100 814.050 106.200 ;
        RECT 823.950 104.100 826.050 106.200 ;
        RECT 830.400 105.600 831.450 115.950 ;
        RECT 803.400 103.350 804.600 104.100 ;
        RECT 796.950 100.950 799.050 103.050 ;
        RECT 799.950 100.950 802.050 103.050 ;
        RECT 802.950 100.950 805.050 103.050 ;
        RECT 805.950 100.950 808.050 103.050 ;
        RECT 800.400 99.900 801.600 100.650 ;
        RECT 799.950 97.800 802.050 99.900 ;
        RECT 806.400 98.400 807.600 100.650 ;
        RECT 806.400 97.050 807.450 98.400 ;
        RECT 812.400 97.050 813.450 104.100 ;
        RECT 824.400 103.350 825.600 104.100 ;
        RECT 830.400 103.350 831.600 105.600 ;
        RECT 820.950 100.950 823.050 103.050 ;
        RECT 823.950 100.950 826.050 103.050 ;
        RECT 826.950 100.950 829.050 103.050 ;
        RECT 829.950 100.950 832.050 103.050 ;
        RECT 821.400 99.000 822.600 100.650 ;
        RECT 827.400 99.000 828.600 100.650 ;
        RECT 839.400 99.900 840.450 124.950 ;
        RECT 851.400 124.050 852.450 131.400 ;
        RECT 856.950 130.800 859.050 132.900 ;
        RECT 859.950 127.950 862.050 130.050 ;
        RECT 850.950 121.950 853.050 124.050 ;
        RECT 853.950 115.950 856.050 118.050 ;
        RECT 847.950 104.100 850.050 106.200 ;
        RECT 854.400 105.600 855.450 115.950 ;
        RECT 848.400 103.350 849.600 104.100 ;
        RECT 854.400 103.350 855.600 105.600 ;
        RECT 844.950 100.950 847.050 103.050 ;
        RECT 847.950 100.950 850.050 103.050 ;
        RECT 850.950 100.950 853.050 103.050 ;
        RECT 853.950 100.950 856.050 103.050 ;
        RECT 845.400 99.900 846.600 100.650 ;
        RECT 851.400 99.900 852.600 100.650 ;
        RECT 805.950 94.950 808.050 97.050 ;
        RECT 811.950 94.950 814.050 97.050 ;
        RECT 820.950 94.950 823.050 99.000 ;
        RECT 826.950 94.950 829.050 99.000 ;
        RECT 838.950 97.800 841.050 99.900 ;
        RECT 844.950 97.800 847.050 99.900 ;
        RECT 850.950 97.800 853.050 99.900 ;
        RECT 787.950 91.950 790.050 94.050 ;
        RECT 784.950 88.950 787.050 91.050 ;
        RECT 763.950 85.950 766.050 88.050 ;
        RECT 806.400 85.050 807.450 94.950 ;
        RECT 808.950 88.950 811.050 94.050 ;
        RECT 805.950 82.950 808.050 85.050 ;
        RECT 812.400 79.050 813.450 94.950 ;
        RECT 825.000 93.900 828.000 94.050 ;
        RECT 823.950 91.950 829.050 93.900 ;
        RECT 823.950 91.800 826.050 91.950 ;
        RECT 826.950 91.800 829.050 91.950 ;
        RECT 814.950 82.950 817.050 85.050 ;
        RECT 790.950 76.950 793.050 79.050 ;
        RECT 811.950 76.950 814.050 79.050 ;
        RECT 775.950 67.950 778.050 70.050 ;
        RECT 745.950 58.950 748.050 61.050 ;
        RECT 748.950 59.100 751.050 61.200 ;
        RECT 754.950 60.600 759.000 61.050 ;
        RECT 776.400 60.600 777.450 67.950 ;
        RECT 735.000 56.100 741.900 57.300 ;
        RECT 738.000 54.300 740.100 55.200 ;
        RECT 731.400 53.100 740.100 54.300 ;
        RECT 732.900 51.300 735.000 53.100 ;
        RECT 736.800 50.100 738.900 52.200 ;
        RECT 741.000 50.700 741.900 56.100 ;
        RECT 742.800 55.950 744.900 58.050 ;
        RECT 743.400 54.450 744.600 55.650 ;
        RECT 746.400 54.450 747.450 58.950 ;
        RECT 749.400 54.900 750.450 59.100 ;
        RECT 754.950 58.950 759.600 60.600 ;
        RECT 758.400 58.350 759.600 58.950 ;
        RECT 776.400 58.350 777.600 60.600 ;
        RECT 781.950 59.100 784.050 61.200 ;
        RECT 782.400 58.350 783.600 59.100 ;
        RECT 757.950 55.950 760.050 58.050 ;
        RECT 760.950 55.950 763.050 58.050 ;
        RECT 775.950 55.950 778.050 58.050 ;
        RECT 778.950 55.950 781.050 58.050 ;
        RECT 781.950 55.950 784.050 58.050 ;
        RECT 761.400 54.900 762.600 55.650 ;
        RECT 743.400 53.400 747.450 54.450 ;
        RECT 748.950 52.800 751.050 54.900 ;
        RECT 760.950 52.800 763.050 54.900 ;
        RECT 779.400 53.400 780.600 55.650 ;
        RECT 737.400 47.550 738.600 49.800 ;
        RECT 740.100 48.600 742.200 50.700 ;
        RECT 724.950 31.950 727.050 34.050 ;
        RECT 733.950 31.950 736.050 34.050 ;
        RECT 725.400 27.600 726.450 31.950 ;
        RECT 725.400 25.350 726.600 27.600 ;
        RECT 721.950 22.950 724.050 25.050 ;
        RECT 724.950 22.950 727.050 25.050 ;
        RECT 722.400 21.900 723.600 22.650 ;
        RECT 734.400 21.900 735.450 31.950 ;
        RECT 737.400 28.200 738.450 47.550 ;
        RECT 769.950 46.950 772.050 49.050 ;
        RECT 748.950 31.950 751.050 34.050 ;
        RECT 736.950 26.100 739.050 28.200 ;
        RECT 742.950 26.100 745.050 28.200 ;
        RECT 749.400 27.600 750.450 31.950 ;
        RECT 770.400 27.600 771.450 46.950 ;
        RECT 779.400 40.050 780.450 53.400 ;
        RECT 791.400 43.050 792.450 76.950 ;
        RECT 793.950 59.100 796.050 61.200 ;
        RECT 799.950 59.100 802.050 61.200 ;
        RECT 805.950 60.000 808.050 64.050 ;
        RECT 794.400 49.050 795.450 59.100 ;
        RECT 800.400 58.350 801.600 59.100 ;
        RECT 806.400 58.350 807.600 60.000 ;
        RECT 799.950 55.950 802.050 58.050 ;
        RECT 802.950 55.950 805.050 58.050 ;
        RECT 805.950 55.950 808.050 58.050 ;
        RECT 808.950 55.950 811.050 58.050 ;
        RECT 803.400 54.000 804.600 55.650 ;
        RECT 809.400 54.900 810.600 55.650 ;
        RECT 802.950 49.950 805.050 54.000 ;
        RECT 808.950 52.800 811.050 54.900 ;
        RECT 811.950 52.950 814.050 55.050 ;
        RECT 793.950 46.950 796.050 49.050 ;
        RECT 812.400 48.450 813.450 52.950 ;
        RECT 815.400 52.050 816.450 82.950 ;
        RECT 826.950 59.100 829.050 61.200 ;
        RECT 844.950 59.100 847.050 64.050 ;
        RECT 850.950 59.100 853.050 61.200 ;
        RECT 827.400 58.350 828.600 59.100 ;
        RECT 845.400 58.350 846.600 59.100 ;
        RECT 851.400 58.350 852.600 59.100 ;
        RECT 823.950 55.950 826.050 58.050 ;
        RECT 826.950 55.950 829.050 58.050 ;
        RECT 841.950 55.950 844.050 58.050 ;
        RECT 844.950 55.950 847.050 58.050 ;
        RECT 847.950 55.950 850.050 58.050 ;
        RECT 850.950 55.950 853.050 58.050 ;
        RECT 824.400 53.400 825.600 55.650 ;
        RECT 842.400 54.900 843.600 55.650 ;
        RECT 814.950 49.950 817.050 52.050 ;
        RECT 812.400 47.400 816.450 48.450 ;
        RECT 796.950 43.950 799.050 46.050 ;
        RECT 790.950 40.950 793.050 43.050 ;
        RECT 778.950 37.950 781.050 40.050 ;
        RECT 781.950 31.950 784.050 34.050 ;
        RECT 743.400 25.350 744.600 26.100 ;
        RECT 749.400 25.350 750.600 27.600 ;
        RECT 770.400 25.350 771.600 27.600 ;
        RECT 742.950 22.950 745.050 25.050 ;
        RECT 745.950 22.950 748.050 25.050 ;
        RECT 748.950 22.950 751.050 25.050 ;
        RECT 751.950 22.950 754.050 25.050 ;
        RECT 769.950 22.950 772.050 25.050 ;
        RECT 772.950 22.950 775.050 25.050 ;
        RECT 721.950 19.800 724.050 21.900 ;
        RECT 733.950 19.800 736.050 21.900 ;
        RECT 746.400 21.000 747.600 22.650 ;
        RECT 752.400 21.900 753.600 22.650 ;
        RECT 773.400 21.900 774.600 22.650 ;
        RECT 745.950 16.950 748.050 21.000 ;
        RECT 751.950 19.800 754.050 21.900 ;
        RECT 772.950 19.800 775.050 21.900 ;
        RECT 691.950 13.950 694.050 16.050 ;
        RECT 715.950 13.950 718.050 16.050 ;
        RECT 646.950 10.950 649.050 13.050 ;
        RECT 782.400 7.050 783.450 31.950 ;
        RECT 797.400 30.450 798.450 43.950 ;
        RECT 799.950 40.950 802.050 43.050 ;
        RECT 794.400 29.400 798.450 30.450 ;
        RECT 794.400 27.600 795.450 29.400 ;
        RECT 800.400 27.600 801.450 40.950 ;
        RECT 808.950 37.950 811.050 40.050 ;
        RECT 805.950 31.950 808.050 34.050 ;
        RECT 794.400 25.350 795.600 27.600 ;
        RECT 800.400 25.350 801.600 27.600 ;
        RECT 790.950 22.950 793.050 25.050 ;
        RECT 793.950 22.950 796.050 25.050 ;
        RECT 796.950 22.950 799.050 25.050 ;
        RECT 799.950 22.950 802.050 25.050 ;
        RECT 791.400 21.900 792.600 22.650 ;
        RECT 797.400 21.900 798.600 22.650 ;
        RECT 806.400 21.900 807.450 31.950 ;
        RECT 809.400 21.900 810.450 37.950 ;
        RECT 815.400 27.600 816.450 47.400 ;
        RECT 824.400 40.050 825.450 53.400 ;
        RECT 841.950 52.800 844.050 54.900 ;
        RECT 848.400 54.000 849.600 55.650 ;
        RECT 844.950 49.950 847.050 52.050 ;
        RECT 847.950 49.950 850.050 54.000 ;
        RECT 853.800 52.950 855.900 55.050 ;
        RECT 845.400 46.050 846.450 49.950 ;
        RECT 854.400 49.050 855.450 52.950 ;
        RECT 856.950 49.950 859.050 55.050 ;
        RECT 853.950 46.950 856.050 49.050 ;
        RECT 860.400 46.050 861.450 127.950 ;
        RECT 866.400 105.450 867.450 187.950 ;
        RECT 875.400 183.600 876.450 193.950 ;
        RECT 875.400 181.350 876.600 183.600 ;
        RECT 880.950 183.000 883.050 187.050 ;
        RECT 881.400 181.350 882.600 183.000 ;
        RECT 871.950 178.950 874.050 181.050 ;
        RECT 874.950 178.950 877.050 181.050 ;
        RECT 877.950 178.950 880.050 181.050 ;
        RECT 880.950 178.950 883.050 181.050 ;
        RECT 868.950 175.800 871.050 177.900 ;
        RECT 872.400 176.400 873.600 178.650 ;
        RECT 878.400 177.000 879.600 178.650 ;
        RECT 869.400 145.050 870.450 175.800 ;
        RECT 868.950 142.950 871.050 145.050 ;
        RECT 869.400 133.050 870.450 142.950 ;
        RECT 868.950 130.950 871.050 133.050 ;
        RECT 872.400 130.050 873.450 176.400 ;
        RECT 877.950 172.950 880.050 177.000 ;
        RECT 887.400 151.050 888.450 202.950 ;
        RECT 889.950 193.950 892.050 196.050 ;
        RECT 886.950 148.950 889.050 151.050 ;
        RECT 880.950 137.100 883.050 139.200 ;
        RECT 886.950 138.000 889.050 142.050 ;
        RECT 890.400 139.200 891.450 193.950 ;
        RECT 893.400 184.050 894.450 209.400 ;
        RECT 898.950 208.800 901.050 210.900 ;
        RECT 907.950 208.800 910.050 210.900 ;
        RECT 911.400 202.050 912.450 232.950 ;
        RECT 926.400 223.050 927.450 259.950 ;
        RECT 929.400 226.050 930.450 268.950 ;
        RECT 944.400 265.050 945.450 325.950 ;
        RECT 956.400 301.050 957.450 337.950 ;
        RECT 962.400 337.350 963.600 338.100 ;
        RECT 967.950 337.950 970.050 340.050 ;
        RECT 973.950 337.950 976.050 340.050 ;
        RECT 968.400 337.350 969.600 337.950 ;
        RECT 961.950 334.950 964.050 337.050 ;
        RECT 964.950 334.950 967.050 337.050 ;
        RECT 967.950 334.950 970.050 337.050 ;
        RECT 970.950 334.950 973.050 337.050 ;
        RECT 965.400 333.900 966.600 334.650 ;
        RECT 964.950 331.800 967.050 333.900 ;
        RECT 971.400 332.400 972.600 334.650 ;
        RECT 977.400 334.050 978.450 362.400 ;
        RECT 979.950 340.950 982.050 343.050 ;
        RECT 971.400 313.050 972.450 332.400 ;
        RECT 976.950 331.950 979.050 334.050 ;
        RECT 970.950 310.950 973.050 313.050 ;
        RECT 980.400 310.050 981.450 340.950 ;
        RECT 979.950 307.950 982.050 310.050 ;
        RECT 964.950 306.450 969.000 307.050 ;
        RECT 964.950 304.950 969.450 306.450 ;
        RECT 961.950 301.950 964.050 304.050 ;
        RECT 949.950 298.950 952.050 301.050 ;
        RECT 955.950 298.950 958.050 301.050 ;
        RECT 950.400 294.600 951.450 298.950 ;
        RECT 962.400 298.050 963.450 301.950 ;
        RECT 964.950 298.950 967.050 301.050 ;
        RECT 961.950 295.950 964.050 298.050 ;
        RECT 950.400 292.350 951.600 294.600 ;
        RECT 955.950 293.100 958.050 295.200 ;
        RECT 956.400 292.350 957.600 293.100 ;
        RECT 949.950 289.950 952.050 292.050 ;
        RECT 952.950 289.950 955.050 292.050 ;
        RECT 955.950 289.950 958.050 292.050 ;
        RECT 958.950 289.950 961.050 292.050 ;
        RECT 946.950 286.800 949.050 288.900 ;
        RECT 953.400 287.400 954.600 289.650 ;
        RECT 959.400 287.400 960.600 289.650 ;
        RECT 947.400 277.050 948.450 286.800 ;
        RECT 946.950 274.950 949.050 277.050 ;
        RECT 943.950 262.950 946.050 265.050 ;
        RECT 949.950 262.950 952.050 265.050 ;
        RECT 937.950 260.100 940.050 262.200 ;
        RECT 945.000 261.600 949.050 262.050 ;
        RECT 938.400 259.350 939.600 260.100 ;
        RECT 944.400 259.950 949.050 261.600 ;
        RECT 944.400 259.350 945.600 259.950 ;
        RECT 934.950 256.950 937.050 259.050 ;
        RECT 937.950 256.950 940.050 259.050 ;
        RECT 940.950 256.950 943.050 259.050 ;
        RECT 943.950 256.950 946.050 259.050 ;
        RECT 935.400 254.400 936.600 256.650 ;
        RECT 941.400 255.900 942.600 256.650 ;
        RECT 935.400 229.050 936.450 254.400 ;
        RECT 940.950 253.800 943.050 255.900 ;
        RECT 940.950 238.950 943.050 241.050 ;
        RECT 934.950 226.950 937.050 229.050 ;
        RECT 928.950 223.950 931.050 226.050 ;
        RECT 913.950 220.950 916.050 223.050 ;
        RECT 925.950 220.950 928.050 223.050 ;
        RECT 914.400 208.050 915.450 220.950 ;
        RECT 929.400 217.200 930.450 223.950 ;
        RECT 934.950 220.950 937.050 223.050 ;
        RECT 922.950 215.100 925.050 217.200 ;
        RECT 928.950 215.100 931.050 217.200 ;
        RECT 923.400 214.350 924.600 215.100 ;
        RECT 929.400 214.350 930.600 215.100 ;
        RECT 919.950 211.950 922.050 214.050 ;
        RECT 922.950 211.950 925.050 214.050 ;
        RECT 925.950 211.950 928.050 214.050 ;
        RECT 928.950 211.950 931.050 214.050 ;
        RECT 920.400 209.400 921.600 211.650 ;
        RECT 926.400 210.000 927.600 211.650 ;
        RECT 913.950 205.950 916.050 208.050 ;
        RECT 910.950 199.950 913.050 202.050 ;
        RECT 920.400 193.050 921.450 209.400 ;
        RECT 925.950 205.950 928.050 210.000 ;
        RECT 922.950 199.950 925.050 202.050 ;
        RECT 910.950 190.950 913.050 193.050 ;
        RECT 919.950 190.950 922.050 193.050 ;
        RECT 901.950 189.450 904.050 190.050 ;
        RECT 896.400 189.000 904.050 189.450 ;
        RECT 895.950 188.400 904.050 189.000 ;
        RECT 895.950 187.050 898.050 188.400 ;
        RECT 901.950 187.950 904.050 188.400 ;
        RECT 895.800 186.000 898.050 187.050 ;
        RECT 895.800 184.950 897.900 186.000 ;
        RECT 892.950 181.950 895.050 184.050 ;
        RECT 898.950 183.000 901.050 187.050 ;
        RECT 899.400 181.350 900.600 183.000 ;
        RECT 907.950 181.950 910.050 184.050 ;
        RECT 895.950 178.950 898.050 181.050 ;
        RECT 898.950 178.950 901.050 181.050 ;
        RECT 901.950 178.950 904.050 181.050 ;
        RECT 896.400 177.900 897.600 178.650 ;
        RECT 895.950 175.800 898.050 177.900 ;
        RECT 902.400 177.000 903.600 178.650 ;
        RECT 901.950 172.950 904.050 177.000 ;
        RECT 904.950 175.950 907.050 178.050 ;
        RECT 892.950 163.950 895.050 166.050 ;
        RECT 881.400 136.350 882.600 137.100 ;
        RECT 887.400 136.350 888.600 138.000 ;
        RECT 889.950 137.100 892.050 139.200 ;
        RECT 877.950 133.950 880.050 136.050 ;
        RECT 880.950 133.950 883.050 136.050 ;
        RECT 883.950 133.950 886.050 136.050 ;
        RECT 886.950 133.950 889.050 136.050 ;
        RECT 878.400 131.400 879.600 133.650 ;
        RECT 884.400 132.900 885.600 133.650 ;
        RECT 871.950 127.950 874.050 130.050 ;
        RECT 878.400 118.050 879.450 131.400 ;
        RECT 883.950 130.800 886.050 132.900 ;
        RECT 893.400 132.450 894.450 163.950 ;
        RECT 895.950 148.950 898.050 151.050 ;
        RECT 896.400 132.900 897.450 148.950 ;
        RECT 905.400 148.050 906.450 175.950 ;
        RECT 908.400 163.050 909.450 181.950 ;
        RECT 911.400 177.900 912.450 190.950 ;
        RECT 916.950 182.100 919.050 184.200 ;
        RECT 923.400 183.600 924.450 199.950 ;
        RECT 928.950 187.950 931.050 190.050 ;
        RECT 929.400 184.050 930.450 187.950 ;
        RECT 917.400 181.350 918.600 182.100 ;
        RECT 923.400 181.350 924.600 183.600 ;
        RECT 928.950 181.950 931.050 184.050 ;
        RECT 916.950 178.950 919.050 181.050 ;
        RECT 919.950 178.950 922.050 181.050 ;
        RECT 922.950 178.950 925.050 181.050 ;
        RECT 925.950 178.950 928.050 181.050 ;
        RECT 920.400 177.900 921.600 178.650 ;
        RECT 910.950 175.800 913.050 177.900 ;
        RECT 919.950 175.800 922.050 177.900 ;
        RECT 926.400 176.400 927.600 178.650 ;
        RECT 926.400 174.450 927.450 176.400 ;
        RECT 935.400 175.050 936.450 220.950 ;
        RECT 937.950 215.100 940.050 217.200 ;
        RECT 938.400 193.050 939.450 215.100 ;
        RECT 941.400 210.450 942.450 238.950 ;
        RECT 950.400 223.050 951.450 262.950 ;
        RECT 953.400 235.050 954.450 287.400 ;
        RECT 959.400 286.050 960.450 287.400 ;
        RECT 955.950 284.400 960.450 286.050 ;
        RECT 955.950 283.950 960.000 284.400 ;
        RECT 965.400 277.050 966.450 298.950 ;
        RECT 968.400 280.050 969.450 304.950 ;
        RECT 983.400 301.050 984.450 428.400 ;
        RECT 985.950 427.950 988.050 428.400 ;
        RECT 989.400 424.050 990.450 442.950 ;
        RECT 995.400 432.450 996.450 443.400 ;
        RECT 997.950 439.950 1000.050 442.050 ;
        RECT 992.400 431.400 996.450 432.450 ;
        RECT 998.400 432.450 999.450 439.950 ;
        RECT 1001.400 436.050 1002.450 443.400 ;
        RECT 1000.950 433.950 1003.050 436.050 ;
        RECT 998.400 431.400 1002.450 432.450 ;
        RECT 992.400 427.050 993.450 431.400 ;
        RECT 994.950 427.950 997.050 430.050 ;
        RECT 991.950 424.950 994.050 427.050 ;
        RECT 988.950 421.950 991.050 424.050 ;
        RECT 990.000 420.450 994.050 421.050 ;
        RECT 989.400 418.950 994.050 420.450 ;
        RECT 989.400 417.600 990.450 418.950 ;
        RECT 995.400 417.600 996.450 427.950 ;
        RECT 989.400 415.350 990.600 417.600 ;
        RECT 995.400 415.350 996.600 417.600 ;
        RECT 1001.400 417.450 1002.450 431.400 ;
        RECT 1004.400 421.050 1005.450 443.400 ;
        RECT 1006.950 439.950 1009.050 442.050 ;
        RECT 1003.950 418.950 1006.050 421.050 ;
        RECT 1001.400 416.400 1005.450 417.450 ;
        RECT 988.950 412.950 991.050 415.050 ;
        RECT 991.950 412.950 994.050 415.050 ;
        RECT 994.950 412.950 997.050 415.050 ;
        RECT 997.950 412.950 1000.050 415.050 ;
        RECT 992.400 411.900 993.600 412.650 ;
        RECT 991.950 409.800 994.050 411.900 ;
        RECT 998.400 410.400 999.600 412.650 ;
        RECT 998.400 408.450 999.450 410.400 ;
        RECT 1000.950 409.950 1003.050 412.050 ;
        RECT 995.400 407.400 999.450 408.450 ;
        RECT 995.400 403.050 996.450 407.400 ;
        RECT 997.950 403.950 1000.050 406.050 ;
        RECT 994.950 400.950 997.050 403.050 ;
        RECT 995.400 376.050 996.450 400.950 ;
        RECT 998.400 385.050 999.450 403.950 ;
        RECT 997.950 382.950 1000.050 385.050 ;
        RECT 997.950 379.800 1000.050 381.900 ;
        RECT 985.950 373.950 988.050 376.050 ;
        RECT 994.950 373.950 997.050 376.050 ;
        RECT 986.400 352.050 987.450 373.950 ;
        RECT 988.950 372.600 993.000 373.050 ;
        RECT 998.400 372.600 999.450 379.800 ;
        RECT 1001.400 373.050 1002.450 409.950 ;
        RECT 988.950 370.950 993.600 372.600 ;
        RECT 992.400 370.350 993.600 370.950 ;
        RECT 998.400 370.350 999.600 372.600 ;
        RECT 1000.950 370.950 1003.050 373.050 ;
        RECT 991.950 367.950 994.050 370.050 ;
        RECT 994.950 367.950 997.050 370.050 ;
        RECT 997.950 367.950 1000.050 370.050 ;
        RECT 988.950 364.950 991.050 367.050 ;
        RECT 995.400 366.000 996.600 367.650 ;
        RECT 985.950 349.950 988.050 352.050 ;
        RECT 989.400 348.450 990.450 364.950 ;
        RECT 994.950 361.950 997.050 366.000 ;
        RECT 1000.950 364.950 1003.050 367.050 ;
        RECT 991.950 348.450 994.050 349.050 ;
        RECT 989.400 347.400 994.050 348.450 ;
        RECT 991.950 346.950 994.050 347.400 ;
        RECT 992.400 339.600 993.450 346.950 ;
        RECT 997.950 343.950 1000.050 346.050 ;
        RECT 992.400 337.350 993.600 339.600 ;
        RECT 986.100 334.950 988.200 337.050 ;
        RECT 991.500 334.950 993.600 337.050 ;
        RECT 994.800 334.950 996.900 337.050 ;
        RECT 986.400 332.400 987.600 334.650 ;
        RECT 995.400 333.900 996.600 334.650 ;
        RECT 986.400 322.050 987.450 332.400 ;
        RECT 994.950 331.800 997.050 333.900 ;
        RECT 985.950 319.950 988.050 322.050 ;
        RECT 985.950 307.950 988.050 310.050 ;
        RECT 982.950 298.950 985.050 301.050 ;
        RECT 982.950 295.800 985.050 297.900 ;
        RECT 973.950 293.100 976.050 295.200 ;
        RECT 974.400 292.350 975.600 293.100 ;
        RECT 973.950 289.950 976.050 292.050 ;
        RECT 976.950 289.950 979.050 292.050 ;
        RECT 977.400 288.900 978.600 289.650 ;
        RECT 976.950 286.800 979.050 288.900 ;
        RECT 983.400 286.050 984.450 295.800 ;
        RECT 982.950 283.950 985.050 286.050 ;
        RECT 982.950 280.800 985.050 282.900 ;
        RECT 967.950 277.950 970.050 280.050 ;
        RECT 976.950 277.950 979.050 280.050 ;
        RECT 955.950 274.950 958.050 277.050 ;
        RECT 964.950 274.950 967.050 277.050 ;
        RECT 956.400 255.900 957.450 274.950 ;
        RECT 964.950 268.950 967.050 271.050 ;
        RECT 958.950 259.950 961.050 265.050 ;
        RECT 965.400 261.600 966.450 268.950 ;
        RECT 965.400 259.350 966.600 261.600 ;
        RECT 970.950 261.450 973.050 262.200 ;
        RECT 973.950 261.450 976.050 265.050 ;
        RECT 970.950 261.000 976.050 261.450 ;
        RECT 970.950 260.400 975.450 261.000 ;
        RECT 970.950 260.100 973.050 260.400 ;
        RECT 971.400 259.350 972.600 260.100 ;
        RECT 961.950 256.950 964.050 259.050 ;
        RECT 964.950 256.950 967.050 259.050 ;
        RECT 967.950 256.950 970.050 259.050 ;
        RECT 970.950 256.950 973.050 259.050 ;
        RECT 955.950 253.800 958.050 255.900 ;
        RECT 962.400 254.400 963.600 256.650 ;
        RECT 968.400 255.900 969.600 256.650 ;
        RECT 955.950 238.950 958.050 241.050 ;
        RECT 952.950 232.950 955.050 235.050 ;
        RECT 949.950 220.950 952.050 223.050 ;
        RECT 949.950 216.000 952.050 219.900 ;
        RECT 956.400 217.200 957.450 238.950 ;
        RECT 962.400 220.050 963.450 254.400 ;
        RECT 967.950 253.800 970.050 255.900 ;
        RECT 977.400 238.050 978.450 277.950 ;
        RECT 979.950 262.950 982.050 265.050 ;
        RECT 980.400 241.050 981.450 262.950 ;
        RECT 983.400 262.050 984.450 280.800 ;
        RECT 986.400 265.050 987.450 307.950 ;
        RECT 991.950 301.950 994.050 304.050 ;
        RECT 992.400 294.600 993.450 301.950 ;
        RECT 995.400 298.050 996.450 331.800 ;
        RECT 998.400 313.050 999.450 343.950 ;
        RECT 997.950 310.950 1000.050 313.050 ;
        RECT 1001.400 304.050 1002.450 364.950 ;
        RECT 1004.400 364.050 1005.450 416.400 ;
        RECT 1007.400 406.050 1008.450 439.950 ;
        RECT 1006.950 403.950 1009.050 406.050 ;
        RECT 1006.950 397.950 1009.050 400.050 ;
        RECT 1003.950 361.950 1006.050 364.050 ;
        RECT 1003.950 358.800 1006.050 360.900 ;
        RECT 1000.950 301.950 1003.050 304.050 ;
        RECT 997.950 298.950 1000.050 301.050 ;
        RECT 994.950 295.950 997.050 298.050 ;
        RECT 998.400 294.600 999.450 298.950 ;
        RECT 1004.400 295.050 1005.450 358.800 ;
        RECT 992.400 292.350 993.600 294.600 ;
        RECT 998.400 292.350 999.600 294.600 ;
        RECT 1003.950 292.950 1006.050 295.050 ;
        RECT 991.950 289.950 994.050 292.050 ;
        RECT 994.950 289.950 997.050 292.050 ;
        RECT 997.950 289.950 1000.050 292.050 ;
        RECT 1000.950 289.950 1003.050 292.050 ;
        RECT 995.400 288.900 996.600 289.650 ;
        RECT 994.950 286.800 997.050 288.900 ;
        RECT 1001.400 287.400 1002.600 289.650 ;
        RECT 997.950 283.950 1000.050 286.050 ;
        RECT 994.950 274.950 997.050 277.050 ;
        RECT 988.950 268.950 991.050 271.050 ;
        RECT 985.950 262.950 988.050 265.050 ;
        RECT 982.950 259.950 985.050 262.050 ;
        RECT 989.400 261.600 990.450 268.950 ;
        RECT 991.950 262.950 994.050 268.050 ;
        RECT 995.400 261.600 996.450 274.950 ;
        RECT 998.400 262.050 999.450 283.950 ;
        RECT 1001.400 283.050 1002.450 287.400 ;
        RECT 1003.950 286.950 1006.050 289.050 ;
        RECT 1000.950 280.950 1003.050 283.050 ;
        RECT 1000.950 268.950 1003.050 271.050 ;
        RECT 989.400 259.350 990.600 261.600 ;
        RECT 995.400 259.350 996.600 261.600 ;
        RECT 997.950 259.950 1000.050 262.050 ;
        RECT 985.950 256.950 988.050 259.050 ;
        RECT 988.950 256.950 991.050 259.050 ;
        RECT 991.950 256.950 994.050 259.050 ;
        RECT 994.950 256.950 997.050 259.050 ;
        RECT 982.950 253.950 985.050 256.050 ;
        RECT 986.400 254.400 987.600 256.650 ;
        RECT 992.400 255.900 993.600 256.650 ;
        RECT 979.950 238.950 982.050 241.050 ;
        RECT 976.950 235.950 979.050 238.050 ;
        RECT 964.950 232.950 967.050 235.050 ;
        RECT 965.400 220.050 966.450 232.950 ;
        RECT 973.950 226.950 976.050 229.050 ;
        RECT 961.800 217.950 963.900 220.050 ;
        RECT 964.950 217.950 967.050 220.050 ;
        RECT 950.400 214.350 951.600 216.000 ;
        RECT 955.950 215.100 958.050 217.200 ;
        RECT 956.400 214.350 957.600 215.100 ;
        RECT 946.950 211.950 949.050 214.050 ;
        RECT 949.950 211.950 952.050 214.050 ;
        RECT 952.950 211.950 955.050 214.050 ;
        RECT 955.950 211.950 958.050 214.050 ;
        RECT 947.400 210.900 948.600 211.650 ;
        RECT 941.400 209.400 945.450 210.450 ;
        RECT 940.950 199.950 943.050 202.050 ;
        RECT 941.400 196.050 942.450 199.950 ;
        RECT 940.950 193.950 943.050 196.050 ;
        RECT 937.950 190.950 940.050 193.050 ;
        RECT 938.400 187.050 939.450 190.950 ;
        RECT 944.400 190.050 945.450 209.400 ;
        RECT 946.950 208.800 949.050 210.900 ;
        RECT 953.400 209.400 954.600 211.650 ;
        RECT 962.400 210.450 963.450 217.950 ;
        RECT 974.400 217.200 975.450 226.950 ;
        RECT 980.400 226.050 981.450 238.950 ;
        RECT 979.950 223.950 982.050 226.050 ;
        RECT 964.950 214.800 967.050 216.900 ;
        RECT 973.950 215.100 976.050 217.200 ;
        RECT 980.400 216.450 981.600 216.600 ;
        RECT 983.400 216.450 984.450 253.950 ;
        RECT 986.400 241.050 987.450 254.400 ;
        RECT 991.950 253.800 994.050 255.900 ;
        RECT 1001.400 244.050 1002.450 268.950 ;
        RECT 988.950 241.950 991.050 244.050 ;
        RECT 1000.950 241.950 1003.050 244.050 ;
        RECT 985.950 238.950 988.050 241.050 ;
        RECT 980.400 215.400 987.450 216.450 ;
        RECT 959.400 209.400 963.450 210.450 ;
        RECT 953.400 202.050 954.450 209.400 ;
        RECT 952.950 199.950 955.050 202.050 ;
        RECT 943.950 187.950 946.050 190.050 ;
        RECT 955.950 187.950 958.050 190.050 ;
        RECT 937.950 184.950 940.050 187.050 ;
        RECT 939.000 183.900 942.000 184.050 ;
        RECT 937.950 183.600 942.000 183.900 ;
        RECT 937.950 181.950 942.600 183.600 ;
        RECT 946.950 182.100 949.050 184.200 ;
        RECT 937.950 181.800 940.050 181.950 ;
        RECT 941.400 181.350 942.600 181.950 ;
        RECT 947.400 181.350 948.600 182.100 ;
        RECT 940.950 178.950 943.050 181.050 ;
        RECT 943.950 178.950 946.050 181.050 ;
        RECT 946.950 178.950 949.050 181.050 ;
        RECT 949.950 178.950 952.050 181.050 ;
        RECT 944.400 176.400 945.600 178.650 ;
        RECT 950.400 177.900 951.600 178.650 ;
        RECT 923.400 173.400 927.450 174.450 ;
        RECT 907.950 160.950 910.050 163.050 ;
        RECT 910.950 157.950 913.050 160.050 ;
        RECT 898.950 145.950 901.050 148.050 ;
        RECT 904.950 145.950 907.050 148.050 ;
        RECT 890.400 131.400 894.450 132.450 ;
        RECT 868.950 115.950 871.050 118.050 ;
        RECT 877.950 115.950 880.050 118.050 ;
        RECT 863.400 104.400 867.450 105.450 ;
        RECT 869.400 105.600 870.450 115.950 ;
        RECT 890.400 112.050 891.450 131.400 ;
        RECT 895.950 130.800 898.050 132.900 ;
        RECT 892.950 112.950 895.050 115.050 ;
        RECT 874.950 109.950 877.050 112.050 ;
        RECT 889.950 109.950 892.050 112.050 ;
        RECT 875.400 105.600 876.450 109.950 ;
        RECT 863.400 99.900 864.450 104.400 ;
        RECT 869.400 103.350 870.600 105.600 ;
        RECT 875.400 103.350 876.600 105.600 ;
        RECT 886.950 103.950 889.050 106.050 ;
        RECT 893.400 105.600 894.450 112.950 ;
        RECT 899.400 106.200 900.450 145.950 ;
        RECT 911.400 142.050 912.450 157.950 ;
        RECT 910.950 139.950 913.050 142.050 ;
        RECT 904.950 137.100 907.050 139.200 ;
        RECT 911.400 138.600 912.450 139.950 ;
        RECT 905.400 136.350 906.600 137.100 ;
        RECT 911.400 136.350 912.600 138.600 ;
        RECT 919.950 137.100 922.050 139.200 ;
        RECT 904.950 133.950 907.050 136.050 ;
        RECT 907.950 133.950 910.050 136.050 ;
        RECT 910.950 133.950 913.050 136.050 ;
        RECT 913.950 133.950 916.050 136.050 ;
        RECT 908.400 132.900 909.600 133.650 ;
        RECT 914.400 132.900 915.600 133.650 ;
        RECT 907.950 130.800 910.050 132.900 ;
        RECT 913.950 130.800 916.050 132.900 ;
        RECT 868.950 100.950 871.050 103.050 ;
        RECT 871.950 100.950 874.050 103.050 ;
        RECT 874.950 100.950 877.050 103.050 ;
        RECT 877.950 100.950 880.050 103.050 ;
        RECT 872.400 99.900 873.600 100.650 ;
        RECT 862.950 97.800 865.050 99.900 ;
        RECT 871.950 97.800 874.050 99.900 ;
        RECT 878.400 98.400 879.600 100.650 ;
        RECT 878.400 94.050 879.450 98.400 ;
        RECT 877.950 91.950 880.050 94.050 ;
        RECT 887.400 70.050 888.450 103.950 ;
        RECT 893.400 103.350 894.600 105.600 ;
        RECT 898.950 104.100 901.050 106.200 ;
        RECT 899.400 103.350 900.600 104.100 ;
        RECT 907.950 103.950 910.050 106.050 ;
        RECT 914.400 105.450 915.450 130.800 ;
        RECT 920.400 127.050 921.450 137.100 ;
        RECT 923.400 130.050 924.450 173.400 ;
        RECT 934.950 172.950 937.050 175.050 ;
        RECT 944.400 163.050 945.450 176.400 ;
        RECT 949.950 175.800 952.050 177.900 ;
        RECT 946.950 172.950 949.050 175.050 ;
        RECT 943.950 160.950 946.050 163.050 ;
        RECT 928.950 145.950 931.050 148.050 ;
        RECT 929.400 138.600 930.450 145.950 ;
        RECT 947.400 139.200 948.450 172.950 ;
        RECT 956.400 154.050 957.450 187.950 ;
        RECT 959.400 169.050 960.450 209.400 ;
        RECT 965.400 199.050 966.450 214.800 ;
        RECT 974.400 214.350 975.600 215.100 ;
        RECT 980.400 214.350 981.600 215.400 ;
        RECT 970.950 211.950 973.050 214.050 ;
        RECT 973.950 211.950 976.050 214.050 ;
        RECT 976.950 211.950 979.050 214.050 ;
        RECT 979.950 211.950 982.050 214.050 ;
        RECT 971.400 211.050 972.600 211.650 ;
        RECT 967.950 209.400 972.600 211.050 ;
        RECT 977.400 210.900 978.600 211.650 ;
        RECT 967.950 208.950 972.450 209.400 ;
        RECT 964.950 196.950 967.050 199.050 ;
        RECT 964.950 193.800 967.050 195.900 ;
        RECT 965.400 183.600 966.450 193.800 ;
        RECT 971.400 184.200 972.450 208.950 ;
        RECT 976.950 208.800 979.050 210.900 ;
        RECT 982.950 208.950 985.050 211.050 ;
        RECT 979.950 196.950 982.050 199.050 ;
        RECT 965.400 181.350 966.600 183.600 ;
        RECT 970.950 182.100 973.050 184.200 ;
        RECT 971.400 181.350 972.600 182.100 ;
        RECT 964.950 178.950 967.050 181.050 ;
        RECT 967.950 178.950 970.050 181.050 ;
        RECT 970.950 178.950 973.050 181.050 ;
        RECT 973.950 178.950 976.050 181.050 ;
        RECT 968.400 177.900 969.600 178.650 ;
        RECT 967.950 175.800 970.050 177.900 ;
        RECT 974.400 177.450 975.600 178.650 ;
        RECT 974.400 177.000 978.450 177.450 ;
        RECT 974.400 176.400 979.050 177.000 ;
        RECT 958.950 166.950 961.050 169.050 ;
        RECT 974.400 163.050 975.450 176.400 ;
        RECT 976.950 172.950 979.050 176.400 ;
        RECT 973.950 160.950 976.050 163.050 ;
        RECT 955.950 151.950 958.050 154.050 ;
        RECT 970.950 151.950 973.050 154.050 ;
        RECT 949.950 142.950 952.050 145.050 ;
        RECT 929.400 136.350 930.600 138.600 ;
        RECT 934.950 137.100 937.050 139.200 ;
        RECT 946.950 137.100 949.050 139.200 ;
        RECT 935.400 136.350 936.600 137.100 ;
        RECT 928.950 133.950 931.050 136.050 ;
        RECT 931.950 133.950 934.050 136.050 ;
        RECT 934.950 133.950 937.050 136.050 ;
        RECT 937.950 133.950 940.050 136.050 ;
        RECT 932.400 132.900 933.600 133.650 ;
        RECT 931.950 130.800 934.050 132.900 ;
        RECT 938.400 131.400 939.600 133.650 ;
        RECT 950.400 132.450 951.450 142.950 ;
        RECT 956.100 142.500 958.200 144.600 ;
        RECT 953.100 133.950 955.200 136.050 ;
        RECT 956.100 135.900 957.000 142.500 ;
        RECT 965.100 142.200 967.200 144.300 ;
        RECT 959.400 139.350 960.600 141.600 ;
        RECT 958.800 136.950 960.900 139.050 ;
        RECT 963.000 135.900 965.100 136.200 ;
        RECT 956.100 135.000 965.100 135.900 ;
        RECT 953.400 132.900 954.600 133.650 ;
        RECT 952.950 132.450 955.050 132.900 ;
        RECT 950.400 131.400 955.050 132.450 ;
        RECT 922.950 127.950 925.050 130.050 ;
        RECT 934.950 127.950 937.050 130.050 ;
        RECT 919.950 124.950 922.050 127.050 ;
        RECT 911.400 104.400 915.450 105.450 ;
        RECT 920.400 105.600 921.450 124.950 ;
        RECT 931.950 112.950 934.050 115.050 ;
        RECT 892.950 100.950 895.050 103.050 ;
        RECT 895.950 100.950 898.050 103.050 ;
        RECT 898.950 100.950 901.050 103.050 ;
        RECT 901.950 100.950 904.050 103.050 ;
        RECT 896.400 98.400 897.600 100.650 ;
        RECT 902.400 99.900 903.600 100.650 ;
        RECT 896.400 94.050 897.450 98.400 ;
        RECT 901.950 97.800 904.050 99.900 ;
        RECT 908.400 97.050 909.450 103.950 ;
        RECT 911.400 99.900 912.450 104.400 ;
        RECT 920.400 103.350 921.600 105.600 ;
        RECT 925.950 104.100 928.050 106.200 ;
        RECT 926.400 103.350 927.600 104.100 ;
        RECT 916.950 100.950 919.050 103.050 ;
        RECT 919.950 100.950 922.050 103.050 ;
        RECT 922.950 100.950 925.050 103.050 ;
        RECT 925.950 100.950 928.050 103.050 ;
        RECT 917.400 99.900 918.600 100.650 ;
        RECT 910.950 97.800 913.050 99.900 ;
        RECT 916.950 97.800 919.050 99.900 ;
        RECT 923.400 99.000 924.600 100.650 ;
        RECT 907.950 94.950 910.050 97.050 ;
        RECT 922.950 94.950 925.050 99.000 ;
        RECT 895.950 91.950 898.050 94.050 ;
        RECT 886.950 67.950 889.050 70.050 ;
        RECT 925.950 67.950 928.050 70.050 ;
        RECT 862.950 59.100 865.050 61.200 ;
        RECT 871.950 59.100 874.050 61.200 ;
        RECT 877.950 60.000 880.050 64.050 ;
        RECT 863.400 54.450 864.450 59.100 ;
        RECT 872.400 58.350 873.600 59.100 ;
        RECT 878.400 58.350 879.600 60.000 ;
        RECT 886.950 59.100 889.050 61.200 ;
        RECT 895.950 59.100 898.050 61.200 ;
        RECT 901.950 60.000 904.050 64.050 ;
        RECT 868.950 55.950 871.050 58.050 ;
        RECT 871.950 55.950 874.050 58.050 ;
        RECT 874.950 55.950 877.050 58.050 ;
        RECT 877.950 55.950 880.050 58.050 ;
        RECT 863.400 53.400 867.450 54.450 ;
        RECT 862.950 49.950 865.050 52.050 ;
        RECT 844.950 43.950 847.050 46.050 ;
        RECT 859.950 43.950 862.050 46.050 ;
        RECT 826.950 40.950 829.050 43.050 ;
        RECT 838.950 40.950 841.050 43.050 ;
        RECT 823.950 37.950 826.050 40.050 ;
        RECT 827.400 34.050 828.450 40.950 ;
        RECT 826.950 31.950 829.050 34.050 ;
        RECT 832.950 31.950 835.050 34.050 ;
        RECT 815.400 25.350 816.600 27.600 ;
        RECT 820.950 26.100 823.050 28.200 ;
        RECT 821.400 25.350 822.600 26.100 ;
        RECT 814.950 22.950 817.050 25.050 ;
        RECT 817.950 22.950 820.050 25.050 ;
        RECT 820.950 22.950 823.050 25.050 ;
        RECT 823.950 22.950 826.050 25.050 ;
        RECT 818.400 21.900 819.600 22.650 ;
        RECT 824.400 21.900 825.600 22.650 ;
        RECT 833.400 21.900 834.450 31.950 ;
        RECT 839.400 27.600 840.450 40.950 ;
        RECT 853.950 37.950 856.050 40.050 ;
        RECT 839.400 25.350 840.600 27.600 ;
        RECT 844.950 26.100 847.050 28.200 ;
        RECT 845.400 25.350 846.600 26.100 ;
        RECT 838.950 22.950 841.050 25.050 ;
        RECT 841.950 22.950 844.050 25.050 ;
        RECT 844.950 22.950 847.050 25.050 ;
        RECT 847.950 22.950 850.050 25.050 ;
        RECT 842.400 21.900 843.600 22.650 ;
        RECT 790.950 19.800 793.050 21.900 ;
        RECT 796.950 19.800 799.050 21.900 ;
        RECT 805.800 19.800 807.900 21.900 ;
        RECT 808.950 19.800 811.050 21.900 ;
        RECT 817.950 19.800 820.050 21.900 ;
        RECT 823.950 19.800 826.050 21.900 ;
        RECT 832.950 19.800 835.050 21.900 ;
        RECT 841.950 19.800 844.050 21.900 ;
        RECT 848.400 21.450 849.600 22.650 ;
        RECT 854.400 21.450 855.450 37.950 ;
        RECT 863.400 27.600 864.450 49.950 ;
        RECT 866.400 37.050 867.450 53.400 ;
        RECT 869.400 53.400 870.600 55.650 ;
        RECT 875.400 53.400 876.600 55.650 ;
        RECT 869.400 46.050 870.450 53.400 ;
        RECT 875.400 49.050 876.450 53.400 ;
        RECT 887.400 49.050 888.450 59.100 ;
        RECT 896.400 58.350 897.600 59.100 ;
        RECT 902.400 58.350 903.600 60.000 ;
        RECT 919.950 59.100 922.050 61.200 ;
        RECT 926.400 60.600 927.450 67.950 ;
        RECT 920.400 58.350 921.600 59.100 ;
        RECT 926.400 58.350 927.600 60.600 ;
        RECT 892.950 55.950 895.050 58.050 ;
        RECT 895.950 55.950 898.050 58.050 ;
        RECT 898.950 55.950 901.050 58.050 ;
        RECT 901.950 55.950 904.050 58.050 ;
        RECT 916.950 55.950 919.050 58.050 ;
        RECT 919.950 55.950 922.050 58.050 ;
        RECT 922.950 55.950 925.050 58.050 ;
        RECT 925.950 55.950 928.050 58.050 ;
        RECT 893.400 54.900 894.600 55.650 ;
        RECT 892.950 52.800 895.050 54.900 ;
        RECT 899.400 54.000 900.600 55.650 ;
        RECT 898.950 49.950 901.050 54.000 ;
        RECT 917.400 53.400 918.600 55.650 ;
        RECT 923.400 54.900 924.600 55.650 ;
        RECT 932.400 54.900 933.450 112.950 ;
        RECT 935.400 94.050 936.450 127.950 ;
        RECT 938.400 126.450 939.450 131.400 ;
        RECT 952.950 130.800 955.050 131.400 ;
        RECT 956.100 129.900 957.000 135.000 ;
        RECT 963.000 134.100 965.100 135.000 ;
        RECT 957.900 133.200 960.000 134.100 ;
        RECT 957.900 132.000 965.100 133.200 ;
        RECT 963.000 131.100 965.100 132.000 ;
        RECT 955.500 127.800 957.600 129.900 ;
        RECT 958.800 128.100 960.900 130.200 ;
        RECT 966.000 129.600 966.900 142.200 ;
        RECT 967.950 137.100 970.050 139.200 ;
        RECT 968.400 136.350 969.600 137.100 ;
        RECT 967.800 133.950 969.900 136.050 ;
        RECT 938.400 125.400 942.450 126.450 ;
        RECT 941.400 105.600 942.450 125.400 ;
        RECT 946.950 124.950 949.050 127.050 ;
        RECT 959.400 125.550 960.600 127.800 ;
        RECT 965.400 127.500 967.500 129.600 ;
        RECT 947.400 105.600 948.450 124.950 ;
        RECT 941.400 103.350 942.600 105.600 ;
        RECT 947.400 103.350 948.600 105.600 ;
        RECT 955.950 103.950 958.050 106.050 ;
        RECT 940.950 100.950 943.050 103.050 ;
        RECT 943.950 100.950 946.050 103.050 ;
        RECT 946.950 100.950 949.050 103.050 ;
        RECT 949.950 100.950 952.050 103.050 ;
        RECT 944.400 98.400 945.600 100.650 ;
        RECT 950.400 99.900 951.600 100.650 ;
        RECT 956.400 99.900 957.450 103.950 ;
        RECT 934.950 91.950 937.050 94.050 ;
        RECT 944.400 91.050 945.450 98.400 ;
        RECT 949.950 97.800 952.050 99.900 ;
        RECT 955.950 97.800 958.050 99.900 ;
        RECT 943.950 90.450 946.050 91.050 ;
        RECT 941.400 89.400 946.050 90.450 ;
        RECT 941.400 61.200 942.450 89.400 ;
        RECT 943.950 88.950 946.050 89.400 ;
        RECT 946.950 67.950 949.050 70.050 ;
        RECT 940.950 59.100 943.050 61.200 ;
        RECT 947.400 60.600 948.450 67.950 ;
        RECT 941.400 58.350 942.600 59.100 ;
        RECT 947.400 58.350 948.600 60.600 ;
        RECT 940.950 55.950 943.050 58.050 ;
        RECT 943.950 55.950 946.050 58.050 ;
        RECT 946.950 55.950 949.050 58.050 ;
        RECT 949.950 55.950 952.050 58.050 ;
        RECT 944.400 54.900 945.600 55.650 ;
        RECT 874.950 46.950 877.050 49.050 ;
        RECT 886.950 46.950 889.050 49.050 ;
        RECT 910.950 46.950 913.050 49.050 ;
        RECT 868.950 43.950 871.050 46.050 ;
        RECT 892.950 40.950 895.050 43.050 ;
        RECT 865.950 34.950 868.050 37.050 ;
        RECT 871.950 34.950 874.050 37.050 ;
        RECT 863.400 25.350 864.600 27.600 ;
        RECT 862.950 22.950 865.050 25.050 ;
        RECT 865.950 22.950 868.050 25.050 ;
        RECT 866.400 21.900 867.600 22.650 ;
        RECT 872.400 22.050 873.450 34.950 ;
        RECT 886.950 26.100 889.050 28.200 ;
        RECT 893.400 27.600 894.450 40.950 ;
        RECT 898.950 34.950 901.050 37.050 ;
        RECT 887.400 25.350 888.600 26.100 ;
        RECT 893.400 25.350 894.600 27.600 ;
        RECT 883.950 22.950 886.050 25.050 ;
        RECT 886.950 22.950 889.050 25.050 ;
        RECT 889.950 22.950 892.050 25.050 ;
        RECT 892.950 22.950 895.050 25.050 ;
        RECT 848.400 20.400 855.450 21.450 ;
        RECT 865.950 19.800 868.050 21.900 ;
        RECT 871.950 19.950 874.050 22.050 ;
        RECT 884.400 20.400 885.600 22.650 ;
        RECT 890.400 21.900 891.600 22.650 ;
        RECT 899.400 22.050 900.450 34.950 ;
        RECT 911.400 27.600 912.450 46.950 ;
        RECT 917.400 45.450 918.450 53.400 ;
        RECT 922.950 52.800 925.050 54.900 ;
        RECT 931.950 52.800 934.050 54.900 ;
        RECT 943.950 52.800 946.050 54.900 ;
        RECT 950.400 53.400 951.600 55.650 ;
        RECT 914.400 44.400 918.450 45.450 ;
        RECT 914.400 37.050 915.450 44.400 ;
        RECT 916.950 40.950 919.050 43.050 ;
        RECT 934.950 40.950 937.050 43.050 ;
        RECT 913.950 34.950 916.050 37.050 ;
        RECT 917.400 27.600 918.450 40.950 ;
        RECT 935.400 37.050 936.450 40.950 ;
        RECT 934.950 34.950 937.050 37.050 ;
        RECT 931.950 31.950 934.050 34.050 ;
        RECT 932.400 27.600 933.450 31.950 ;
        RECT 911.400 25.350 912.600 27.600 ;
        RECT 917.400 25.350 918.600 27.600 ;
        RECT 932.400 25.350 933.600 27.600 ;
        RECT 937.950 26.100 940.050 28.200 ;
        RECT 938.400 25.350 939.600 26.100 ;
        RECT 907.950 22.950 910.050 25.050 ;
        RECT 910.950 22.950 913.050 25.050 ;
        RECT 913.950 22.950 916.050 25.050 ;
        RECT 916.950 22.950 919.050 25.050 ;
        RECT 931.950 22.950 934.050 25.050 ;
        RECT 934.950 22.950 937.050 25.050 ;
        RECT 937.950 22.950 940.050 25.050 ;
        RECT 940.950 22.950 943.050 25.050 ;
        RECT 884.400 7.050 885.450 20.400 ;
        RECT 889.950 19.800 892.050 21.900 ;
        RECT 898.950 19.950 901.050 22.050 ;
        RECT 904.800 19.950 906.900 22.050 ;
        RECT 908.400 21.900 909.600 22.650 ;
        RECT 898.950 13.950 901.050 18.900 ;
        RECT 905.400 16.050 906.450 19.950 ;
        RECT 907.950 16.950 910.050 21.900 ;
        RECT 914.400 20.400 915.600 22.650 ;
        RECT 935.400 21.900 936.600 22.650 ;
        RECT 941.400 22.050 942.600 22.650 ;
        RECT 950.400 22.050 951.450 53.400 ;
        RECT 956.400 46.050 957.450 97.800 ;
        RECT 959.400 91.050 960.450 125.550 ;
        RECT 964.950 104.100 967.050 106.200 ;
        RECT 971.400 106.050 972.450 151.950 ;
        RECT 980.400 127.050 981.450 196.950 ;
        RECT 983.400 175.050 984.450 208.950 ;
        RECT 986.400 208.050 987.450 215.400 ;
        RECT 985.950 205.950 988.050 208.050 ;
        RECT 986.400 202.050 987.450 205.950 ;
        RECT 985.950 199.950 988.050 202.050 ;
        RECT 989.400 192.450 990.450 241.950 ;
        RECT 991.950 238.950 994.050 241.050 ;
        RECT 992.400 211.050 993.450 238.950 ;
        RECT 1004.400 235.050 1005.450 286.950 ;
        RECT 1007.400 262.050 1008.450 397.950 ;
        RECT 1010.400 277.050 1011.450 502.800 ;
        RECT 1009.950 274.950 1012.050 277.050 ;
        RECT 1006.950 259.950 1009.050 262.050 ;
        RECT 1009.950 259.950 1012.050 262.050 ;
        RECT 1003.950 232.950 1006.050 235.050 ;
        RECT 1000.950 226.950 1003.050 229.050 ;
        RECT 997.950 223.950 1000.050 226.050 ;
        RECT 998.400 220.050 999.450 223.950 ;
        RECT 997.950 217.950 1000.050 220.050 ;
        RECT 1001.400 216.600 1002.450 226.950 ;
        RECT 1001.400 214.350 1002.600 216.600 ;
        RECT 1006.950 216.000 1009.050 220.050 ;
        RECT 1010.400 217.050 1011.450 259.950 ;
        RECT 1007.400 214.350 1008.600 216.000 ;
        RECT 1009.950 214.950 1012.050 217.050 ;
        RECT 997.950 211.950 1000.050 214.050 ;
        RECT 1000.950 211.950 1003.050 214.050 ;
        RECT 1003.950 211.950 1006.050 214.050 ;
        RECT 1006.950 211.950 1009.050 214.050 ;
        RECT 991.950 208.950 994.050 211.050 ;
        RECT 998.400 210.900 999.600 211.650 ;
        RECT 997.950 208.800 1000.050 210.900 ;
        RECT 1004.400 210.000 1005.600 211.650 ;
        RECT 1013.400 211.050 1014.450 521.400 ;
        RECT 1015.950 517.950 1018.050 520.050 ;
        RECT 1016.400 469.050 1017.450 517.950 ;
        RECT 1015.950 466.950 1018.050 469.050 ;
        RECT 1015.950 460.950 1018.050 463.050 ;
        RECT 1016.400 265.050 1017.450 460.950 ;
        RECT 1015.950 262.950 1018.050 265.050 ;
        RECT 1015.950 235.950 1018.050 238.050 ;
        RECT 1003.950 205.950 1006.050 210.000 ;
        RECT 1009.950 208.950 1012.050 211.050 ;
        RECT 1012.950 208.950 1015.050 211.050 ;
        RECT 986.400 191.400 990.450 192.450 ;
        RECT 986.400 184.050 987.450 191.400 ;
        RECT 988.950 187.950 991.050 190.050 ;
        RECT 985.950 181.950 988.050 184.050 ;
        RECT 989.400 183.600 990.450 187.950 ;
        RECT 989.400 181.350 990.600 183.600 ;
        RECT 988.950 178.950 991.050 181.050 ;
        RECT 991.950 178.950 994.050 181.050 ;
        RECT 992.400 177.000 993.600 178.650 ;
        RECT 982.950 172.950 985.050 175.050 ;
        RECT 991.950 172.950 994.050 177.000 ;
        RECT 982.950 166.950 985.050 169.050 ;
        RECT 979.950 124.950 982.050 127.050 ;
        RECT 983.400 123.450 984.450 166.950 ;
        RECT 988.800 142.500 990.900 144.600 ;
        RECT 986.100 133.950 988.200 136.050 ;
        RECT 989.100 135.300 990.300 142.500 ;
        RECT 992.400 139.350 993.600 141.600 ;
        RECT 998.400 141.300 1000.500 143.400 ;
        RECT 992.100 136.950 994.200 139.050 ;
        RECT 995.100 137.700 997.200 139.800 ;
        RECT 995.100 135.300 996.000 137.700 ;
        RECT 989.100 134.100 996.000 135.300 ;
        RECT 986.400 132.900 987.600 133.650 ;
        RECT 985.950 130.800 988.050 132.900 ;
        RECT 989.100 128.700 990.000 134.100 ;
        RECT 990.900 132.300 993.000 133.200 ;
        RECT 998.700 132.300 999.600 141.300 ;
        RECT 1000.950 137.100 1003.050 139.200 ;
        RECT 1001.400 136.350 1002.600 137.100 ;
        RECT 1000.800 133.950 1002.900 136.050 ;
        RECT 990.900 131.100 999.600 132.300 ;
        RECT 988.800 126.600 990.900 128.700 ;
        RECT 992.100 128.100 994.200 130.200 ;
        RECT 996.000 129.300 998.100 131.100 ;
        RECT 992.400 125.550 993.600 127.800 ;
        RECT 983.400 122.400 987.450 123.450 ;
        RECT 979.950 109.950 982.050 112.050 ;
        RECT 965.400 103.350 966.600 104.100 ;
        RECT 970.950 103.950 973.050 106.050 ;
        RECT 964.950 100.950 967.050 103.050 ;
        RECT 967.950 100.950 970.050 103.050 ;
        RECT 968.400 100.050 969.600 100.650 ;
        RECT 968.400 99.900 972.000 100.050 ;
        RECT 968.400 98.400 973.050 99.900 ;
        RECT 969.000 97.950 973.050 98.400 ;
        RECT 970.950 97.800 973.050 97.950 ;
        RECT 958.950 88.950 961.050 91.050 ;
        RECT 958.950 59.100 961.050 61.200 ;
        RECT 964.950 59.100 967.050 61.200 ;
        RECT 970.950 60.000 973.050 64.050 ;
        RECT 980.400 61.200 981.450 109.950 ;
        RECT 986.400 105.600 987.450 122.400 ;
        RECT 992.400 115.050 993.450 125.550 ;
        RECT 991.950 112.950 994.050 115.050 ;
        RECT 1000.950 112.950 1003.050 115.050 ;
        RECT 988.950 108.450 991.050 112.050 ;
        RECT 988.950 108.000 993.450 108.450 ;
        RECT 989.400 107.400 993.450 108.000 ;
        RECT 992.400 105.600 993.450 107.400 ;
        RECT 986.400 103.350 987.600 105.600 ;
        RECT 992.400 103.350 993.600 105.600 ;
        RECT 985.950 100.950 988.050 103.050 ;
        RECT 988.950 100.950 991.050 103.050 ;
        RECT 991.950 100.950 994.050 103.050 ;
        RECT 994.950 100.950 997.050 103.050 ;
        RECT 989.400 99.900 990.600 100.650 ;
        RECT 988.950 97.800 991.050 99.900 ;
        RECT 995.400 99.000 996.600 100.650 ;
        RECT 994.950 96.450 997.050 99.000 ;
        RECT 1001.400 97.050 1002.450 112.950 ;
        RECT 992.400 95.400 997.050 96.450 ;
        RECT 982.950 91.950 985.050 94.050 ;
        RECT 959.400 52.050 960.450 59.100 ;
        RECT 965.400 58.350 966.600 59.100 ;
        RECT 971.400 58.350 972.600 60.000 ;
        RECT 979.950 59.100 982.050 61.200 ;
        RECT 964.950 55.950 967.050 58.050 ;
        RECT 967.950 55.950 970.050 58.050 ;
        RECT 970.950 55.950 973.050 58.050 ;
        RECT 973.950 55.950 976.050 58.050 ;
        RECT 968.400 54.900 969.600 55.650 ;
        RECT 967.950 52.800 970.050 54.900 ;
        RECT 974.400 53.400 975.600 55.650 ;
        RECT 983.400 55.050 984.450 91.950 ;
        RECT 992.400 60.600 993.450 95.400 ;
        RECT 994.950 94.950 997.050 95.400 ;
        RECT 1000.950 94.950 1003.050 97.050 ;
        RECT 992.400 58.350 993.600 60.600 ;
        RECT 997.950 59.100 1000.050 61.200 ;
        RECT 998.400 58.350 999.600 59.100 ;
        RECT 988.950 55.950 991.050 58.050 ;
        RECT 991.950 55.950 994.050 58.050 ;
        RECT 994.950 55.950 997.050 58.050 ;
        RECT 997.950 55.950 1000.050 58.050 ;
        RECT 958.950 49.950 961.050 52.050 ;
        RECT 955.950 43.950 958.050 46.050 ;
        RECT 959.400 27.600 960.450 49.950 ;
        RECT 974.400 40.050 975.450 53.400 ;
        RECT 982.950 52.950 985.050 55.050 ;
        RECT 985.950 52.950 988.050 55.050 ;
        RECT 989.400 53.400 990.600 55.650 ;
        RECT 995.400 53.400 996.600 55.650 ;
        RECT 973.950 37.950 976.050 40.050 ;
        RECT 959.400 25.350 960.600 27.600 ;
        RECT 964.950 26.100 967.050 28.200 ;
        RECT 986.400 27.600 987.450 52.950 ;
        RECT 989.400 37.050 990.450 53.400 ;
        RECT 995.400 46.050 996.450 53.400 ;
        RECT 994.950 43.950 997.050 46.050 ;
        RECT 988.950 34.950 991.050 37.050 ;
        RECT 1010.400 28.200 1011.450 208.950 ;
        RECT 1016.400 115.050 1017.450 235.950 ;
        RECT 1015.950 112.950 1018.050 115.050 ;
        RECT 965.400 25.350 966.600 26.100 ;
        RECT 986.400 25.350 987.600 27.600 ;
        RECT 991.950 26.100 994.050 28.200 ;
        RECT 1009.950 26.100 1012.050 28.200 ;
        RECT 992.400 25.350 993.600 26.100 ;
        RECT 958.950 22.950 961.050 25.050 ;
        RECT 961.950 22.950 964.050 25.050 ;
        RECT 964.950 22.950 967.050 25.050 ;
        RECT 967.950 22.950 970.050 25.050 ;
        RECT 985.950 22.950 988.050 25.050 ;
        RECT 988.950 22.950 991.050 25.050 ;
        RECT 991.950 22.950 994.050 25.050 ;
        RECT 994.950 22.950 997.050 25.050 ;
        RECT 914.400 16.050 915.450 20.400 ;
        RECT 934.950 19.800 937.050 21.900 ;
        RECT 941.400 20.400 946.050 22.050 ;
        RECT 942.000 19.950 946.050 20.400 ;
        RECT 949.950 19.800 952.050 22.050 ;
        RECT 962.400 21.900 963.600 22.650 ;
        RECT 961.950 19.800 964.050 21.900 ;
        RECT 968.400 20.400 969.600 22.650 ;
        RECT 989.400 20.400 990.600 22.650 ;
        RECT 995.400 21.900 996.600 22.650 ;
        RECT 904.950 13.950 907.050 16.050 ;
        RECT 913.950 13.950 916.050 16.050 ;
        RECT 968.400 7.050 969.450 20.400 ;
        RECT 989.400 7.050 990.450 20.400 ;
        RECT 994.950 19.800 997.050 21.900 ;
        RECT 469.950 4.950 472.050 7.050 ;
        RECT 622.950 4.950 625.050 7.050 ;
        RECT 781.950 4.950 784.050 7.050 ;
        RECT 883.950 4.950 886.050 7.050 ;
        RECT 967.950 4.950 970.050 7.050 ;
        RECT 988.950 4.950 991.050 7.050 ;
      LAYER via2 ;
        RECT 67.950 919.950 70.050 922.050 ;
        RECT 142.950 907.950 145.050 910.050 ;
        RECT 67.950 841.950 70.050 844.050 ;
        RECT 130.950 886.950 133.050 889.050 ;
        RECT 91.950 808.950 94.050 811.050 ;
        RECT 247.950 925.950 250.050 928.050 ;
        RECT 295.950 955.800 298.050 957.900 ;
        RECT 346.950 955.950 349.050 958.050 ;
        RECT 259.950 886.950 262.050 889.050 ;
        RECT 268.950 886.950 271.050 889.050 ;
        RECT 247.950 883.950 250.050 886.050 ;
        RECT 118.950 808.950 121.050 811.050 ;
        RECT 319.950 886.950 322.050 889.050 ;
        RECT 475.950 955.800 478.050 957.900 ;
        RECT 190.950 763.950 193.050 766.050 ;
        RECT 52.950 685.950 55.050 688.050 ;
        RECT 88.950 607.950 91.050 610.050 ;
        RECT 64.950 527.100 67.050 529.200 ;
        RECT 259.950 733.800 262.050 735.900 ;
        RECT 139.950 652.950 142.050 655.050 ;
        RECT 103.950 451.950 106.050 454.050 ;
        RECT 337.950 766.950 340.050 769.050 ;
        RECT 484.950 895.950 487.050 898.050 ;
        RECT 487.950 892.950 490.050 895.050 ;
        RECT 328.950 721.950 331.050 724.050 ;
        RECT 295.950 685.950 298.050 688.050 ;
        RECT 163.950 526.950 166.050 529.050 ;
        RECT 151.950 451.950 154.050 454.050 ;
        RECT 55.950 340.950 58.050 343.050 ;
        RECT 46.950 262.950 49.050 265.050 ;
        RECT 208.950 496.950 211.050 499.050 ;
        RECT 169.950 463.950 172.050 466.050 ;
        RECT 172.950 451.950 175.050 454.050 ;
        RECT 121.950 265.950 124.050 268.050 ;
        RECT 283.950 652.950 286.050 655.050 ;
        RECT 352.950 685.950 355.050 688.050 ;
        RECT 370.950 685.950 373.050 688.050 ;
        RECT 343.950 607.950 346.050 610.050 ;
        RECT 349.950 577.950 352.050 580.050 ;
        RECT 205.950 442.950 208.050 445.050 ;
        RECT 226.950 451.950 229.050 454.050 ;
        RECT 478.950 841.950 481.050 844.050 ;
        RECT 400.950 607.950 403.050 610.050 ;
        RECT 463.950 685.950 466.050 688.050 ;
        RECT 463.950 652.950 466.050 655.050 ;
        RECT 430.950 607.950 433.050 610.050 ;
        RECT 454.950 607.950 457.050 610.050 ;
        RECT 334.950 451.950 337.050 454.050 ;
        RECT 163.950 340.950 166.050 343.050 ;
        RECT 124.950 253.800 127.050 255.900 ;
        RECT 85.950 184.950 88.050 187.050 ;
        RECT 37.950 106.950 40.050 109.050 ;
        RECT 67.950 61.950 70.050 64.050 ;
        RECT 298.950 406.950 301.050 409.050 ;
        RECT 250.950 262.950 253.050 265.050 ;
        RECT 244.950 217.950 247.050 220.050 ;
        RECT 169.950 182.100 172.050 184.200 ;
        RECT 223.950 139.950 226.050 142.050 ;
        RECT 196.950 130.800 199.050 132.900 ;
        RECT 373.950 451.950 376.050 454.050 ;
        RECT 523.950 772.950 526.050 775.050 ;
        RECT 670.950 964.950 673.050 967.050 ;
        RECT 691.950 964.950 694.050 967.050 ;
        RECT 733.950 964.950 736.050 967.050 ;
        RECT 580.950 892.950 583.050 895.050 ;
        RECT 763.950 964.950 766.050 967.050 ;
        RECT 808.950 964.950 811.050 967.050 ;
        RECT 622.950 841.950 625.050 844.050 ;
        RECT 601.950 808.950 604.050 811.050 ;
        RECT 598.950 799.800 601.050 801.900 ;
        RECT 529.950 730.950 532.050 733.050 ;
        RECT 496.950 607.950 499.050 610.050 ;
        RECT 430.950 529.950 433.050 532.050 ;
        RECT 457.950 496.950 460.050 499.050 ;
        RECT 556.950 688.950 559.050 691.050 ;
        RECT 391.950 451.950 394.050 454.050 ;
        RECT 373.950 418.950 376.050 421.050 ;
        RECT 394.950 418.950 397.050 421.050 ;
        RECT 274.950 217.950 277.050 220.050 ;
        RECT 112.950 97.800 115.050 99.900 ;
        RECT 184.950 106.950 187.050 109.050 ;
        RECT 214.950 106.950 217.050 109.050 ;
        RECT 130.950 61.950 133.050 64.050 ;
        RECT 100.950 34.950 103.050 37.050 ;
        RECT 61.950 28.950 64.050 31.050 ;
        RECT 91.950 16.950 94.050 19.050 ;
        RECT 232.950 91.950 235.050 94.050 ;
        RECT 310.950 217.950 313.050 220.050 ;
        RECT 544.950 565.800 547.050 567.900 ;
        RECT 550.950 565.950 553.050 568.050 ;
        RECT 589.950 607.950 592.050 610.050 ;
        RECT 883.950 970.950 886.050 973.050 ;
        RECT 892.950 967.950 895.050 970.050 ;
        RECT 844.950 955.950 847.050 958.050 ;
        RECT 868.950 952.950 871.050 955.050 ;
        RECT 757.950 886.950 760.050 889.050 ;
        RECT 781.950 886.950 784.050 889.050 ;
        RECT 613.950 607.950 616.050 610.050 ;
        RECT 700.950 730.950 703.050 733.050 ;
        RECT 541.950 451.950 544.050 454.050 ;
        RECT 481.950 373.950 484.050 376.050 ;
        RECT 475.950 340.950 478.050 343.050 ;
        RECT 391.950 217.950 394.050 220.050 ;
        RECT 226.950 61.950 229.050 64.050 ;
        RECT 226.950 28.950 229.050 31.050 ;
        RECT 109.950 13.950 112.050 16.050 ;
        RECT 394.950 139.950 397.050 142.050 ;
        RECT 541.950 418.950 544.050 421.050 ;
        RECT 598.950 529.800 601.050 531.900 ;
        RECT 556.950 418.950 559.050 421.050 ;
        RECT 523.950 340.950 526.050 343.050 ;
        RECT 487.950 220.950 490.050 223.050 ;
        RECT 685.950 652.950 688.050 655.050 ;
        RECT 880.950 919.950 883.050 922.050 ;
        RECT 925.950 964.950 928.050 967.050 ;
        RECT 934.950 955.800 937.050 957.900 ;
        RECT 790.950 733.950 793.050 736.050 ;
        RECT 676.950 496.950 679.050 499.050 ;
        RECT 787.950 685.950 790.050 688.050 ;
        RECT 757.950 652.950 760.050 655.050 ;
        RECT 784.950 652.950 787.050 655.050 ;
        RECT 697.950 529.950 700.050 532.050 ;
        RECT 700.950 520.800 703.050 522.900 ;
        RECT 868.950 841.950 871.050 844.050 ;
        RECT 838.950 763.950 841.050 766.050 ;
        RECT 859.950 763.950 862.050 766.050 ;
        RECT 868.950 763.950 871.050 766.050 ;
        RECT 862.950 730.950 865.050 733.050 ;
        RECT 727.950 529.950 730.050 532.050 ;
        RECT 604.950 340.950 607.050 343.050 ;
        RECT 535.950 262.950 538.050 265.050 ;
        RECT 403.950 106.950 406.050 109.050 ;
        RECT 346.950 28.950 349.050 31.050 ;
        RECT 607.950 304.800 610.050 306.900 ;
        RECT 610.950 301.950 613.050 304.050 ;
        RECT 625.950 340.950 628.050 343.050 ;
        RECT 631.950 298.950 634.050 301.050 ;
        RECT 562.950 184.950 565.050 187.050 ;
        RECT 604.950 184.950 607.050 187.050 ;
        RECT 568.950 130.800 571.050 132.900 ;
        RECT 481.950 100.950 484.050 103.050 ;
        RECT 460.950 61.950 463.050 64.050 ;
        RECT 463.950 52.800 466.050 54.900 ;
        RECT 835.950 676.800 838.050 678.900 ;
        RECT 946.950 919.950 949.050 922.050 ;
        RECT 952.950 886.950 955.050 889.050 ;
        RECT 865.950 709.950 868.050 712.050 ;
        RECT 769.950 529.950 772.050 532.050 ;
        RECT 835.950 574.950 838.050 577.050 ;
        RECT 682.950 373.950 685.050 376.050 ;
        RECT 670.950 295.950 673.050 298.050 ;
        RECT 943.950 754.800 946.050 756.900 ;
        RECT 949.950 733.950 952.050 736.050 ;
        RECT 871.950 649.950 874.050 652.050 ;
        RECT 859.950 574.950 862.050 577.050 ;
        RECT 847.950 487.950 850.050 490.050 ;
        RECT 682.950 286.950 685.050 289.050 ;
        RECT 697.950 295.800 700.050 297.900 ;
        RECT 655.950 182.100 658.050 184.200 ;
        RECT 655.950 175.800 658.050 177.900 ;
        RECT 727.950 295.800 730.050 297.900 ;
        RECT 874.950 520.950 877.050 523.050 ;
        RECT 934.950 676.800 937.050 678.900 ;
        RECT 895.950 607.950 898.050 610.050 ;
        RECT 964.950 652.950 967.050 655.050 ;
        RECT 892.950 520.800 895.050 522.900 ;
        RECT 709.950 217.950 712.050 220.050 ;
        RECT 580.950 109.950 583.050 112.050 ;
        RECT 562.950 28.950 565.050 31.050 ;
        RECT 535.950 19.800 538.050 21.900 ;
        RECT 580.950 28.950 583.050 31.050 ;
        RECT 661.950 64.950 664.050 67.050 ;
        RECT 787.950 295.950 790.050 298.050 ;
        RECT 850.950 409.800 853.050 411.900 ;
        RECT 802.950 340.950 805.050 343.050 ;
        RECT 997.950 730.950 1000.050 733.050 ;
        RECT 958.950 574.950 961.050 577.050 ;
        RECT 961.950 565.800 964.050 567.900 ;
        RECT 982.950 574.950 985.050 577.050 ;
        RECT 958.950 496.950 961.050 499.050 ;
        RECT 922.950 436.950 925.050 439.050 ;
        RECT 922.950 418.950 925.050 421.050 ;
        RECT 928.950 418.950 931.050 421.050 ;
        RECT 988.950 496.950 991.050 499.050 ;
        RECT 652.950 52.800 655.050 54.900 ;
        RECT 610.950 28.950 613.050 31.050 ;
        RECT 652.950 28.950 655.050 31.050 ;
        RECT 754.950 106.950 757.050 109.050 ;
        RECT 766.950 109.950 769.050 112.050 ;
        RECT 850.950 184.950 853.050 187.050 ;
        RECT 922.950 340.950 925.050 343.050 ;
        RECT 979.950 364.950 982.050 367.050 ;
        RECT 844.950 61.950 847.050 64.050 ;
        RECT 856.950 52.950 859.050 55.050 ;
        RECT 880.950 184.950 883.050 187.050 ;
        RECT 898.950 184.950 901.050 187.050 ;
        RECT 958.950 262.950 961.050 265.050 ;
        RECT 991.950 265.950 994.050 268.050 ;
        RECT 877.950 61.950 880.050 64.050 ;
        RECT 901.950 61.950 904.050 64.050 ;
        RECT 907.950 19.800 910.050 21.900 ;
        RECT 1006.950 217.950 1009.050 220.050 ;
        RECT 988.950 109.950 991.050 112.050 ;
      LAYER metal3 ;
        RECT 79.950 975.600 82.050 976.050 ;
        RECT 190.950 975.600 193.050 976.050 ;
        RECT 349.950 975.600 352.050 976.050 ;
        RECT 79.950 974.400 352.050 975.600 ;
        RECT 79.950 973.950 82.050 974.400 ;
        RECT 190.950 973.950 193.050 974.400 ;
        RECT 349.950 973.950 352.050 974.400 ;
        RECT 553.950 975.600 556.050 976.050 ;
        RECT 595.950 975.600 598.050 976.050 ;
        RECT 553.950 974.400 598.050 975.600 ;
        RECT 553.950 973.950 556.050 974.400 ;
        RECT 595.950 973.950 598.050 974.400 ;
        RECT 835.950 975.600 838.050 976.050 ;
        RECT 919.950 975.600 922.050 976.050 ;
        RECT 835.950 974.400 922.050 975.600 ;
        RECT 835.950 973.950 838.050 974.400 ;
        RECT 919.950 973.950 922.050 974.400 ;
        RECT 403.950 972.600 406.050 973.050 ;
        RECT 427.950 972.600 430.050 973.050 ;
        RECT 403.950 971.400 430.050 972.600 ;
        RECT 403.950 970.950 406.050 971.400 ;
        RECT 427.950 970.950 430.050 971.400 ;
        RECT 433.950 972.600 436.050 973.050 ;
        RECT 478.950 972.600 481.050 973.050 ;
        RECT 433.950 971.400 481.050 972.600 ;
        RECT 433.950 970.950 436.050 971.400 ;
        RECT 478.950 970.950 481.050 971.400 ;
        RECT 514.950 972.600 517.050 973.050 ;
        RECT 526.950 972.600 529.050 973.050 ;
        RECT 622.950 972.600 625.050 973.050 ;
        RECT 733.950 972.600 736.050 973.050 ;
        RECT 514.950 971.400 529.050 972.600 ;
        RECT 514.950 970.950 517.050 971.400 ;
        RECT 526.950 970.950 529.050 971.400 ;
        RECT 530.400 971.400 591.600 972.600 ;
        RECT 25.950 969.600 28.050 970.050 ;
        RECT 85.950 969.600 88.050 970.050 ;
        RECT 208.950 969.600 211.050 970.050 ;
        RECT 220.950 969.600 223.050 970.050 ;
        RECT 25.950 968.400 223.050 969.600 ;
        RECT 25.950 967.950 28.050 968.400 ;
        RECT 85.950 967.950 88.050 968.400 ;
        RECT 208.950 967.950 211.050 968.400 ;
        RECT 220.950 967.950 223.050 968.400 ;
        RECT 226.950 969.600 229.050 970.050 ;
        RECT 259.950 969.600 262.050 970.050 ;
        RECT 226.950 968.400 262.050 969.600 ;
        RECT 226.950 967.950 229.050 968.400 ;
        RECT 259.950 967.950 262.050 968.400 ;
        RECT 409.950 969.600 412.050 970.050 ;
        RECT 490.950 969.600 493.050 970.050 ;
        RECT 530.400 969.600 531.600 971.400 ;
        RECT 409.950 968.400 489.600 969.600 ;
        RECT 409.950 967.950 412.050 968.400 ;
        RECT 488.400 966.600 489.600 968.400 ;
        RECT 490.950 968.400 531.600 969.600 ;
        RECT 590.400 969.600 591.600 971.400 ;
        RECT 622.950 971.400 736.050 972.600 ;
        RECT 622.950 970.950 625.050 971.400 ;
        RECT 733.950 970.950 736.050 971.400 ;
        RECT 739.950 972.600 742.050 973.050 ;
        RECT 781.950 972.600 784.050 973.050 ;
        RECT 739.950 971.400 784.050 972.600 ;
        RECT 739.950 970.950 742.050 971.400 ;
        RECT 781.950 970.950 784.050 971.400 ;
        RECT 856.950 972.600 859.050 973.050 ;
        RECT 883.950 972.600 886.050 973.050 ;
        RECT 856.950 971.400 886.050 972.600 ;
        RECT 856.950 970.950 859.050 971.400 ;
        RECT 883.950 970.950 886.050 971.400 ;
        RECT 991.950 972.600 994.050 973.050 ;
        RECT 1003.950 972.600 1006.050 973.050 ;
        RECT 991.950 971.400 1006.050 972.600 ;
        RECT 991.950 970.950 994.050 971.400 ;
        RECT 1003.950 970.950 1006.050 971.400 ;
        RECT 664.950 969.600 667.050 970.050 ;
        RECT 590.400 968.400 667.050 969.600 ;
        RECT 490.950 967.950 493.050 968.400 ;
        RECT 664.950 967.950 667.050 968.400 ;
        RECT 736.950 969.600 739.050 970.050 ;
        RECT 817.950 969.600 820.050 970.050 ;
        RECT 886.950 969.600 889.050 970.050 ;
        RECT 736.950 968.400 889.050 969.600 ;
        RECT 736.950 967.950 739.050 968.400 ;
        RECT 817.950 967.950 820.050 968.400 ;
        RECT 886.950 967.950 889.050 968.400 ;
        RECT 892.950 969.600 895.050 970.050 ;
        RECT 973.950 969.600 976.050 970.050 ;
        RECT 892.950 968.400 976.050 969.600 ;
        RECT 892.950 967.950 895.050 968.400 ;
        RECT 973.950 967.950 976.050 968.400 ;
        RECT 562.950 966.600 565.050 967.050 ;
        RECT 586.950 966.600 589.050 967.050 ;
        RECT 488.400 965.400 589.050 966.600 ;
        RECT 562.950 964.950 565.050 965.400 ;
        RECT 586.950 964.950 589.050 965.400 ;
        RECT 670.950 966.600 673.050 967.050 ;
        RECT 691.950 966.600 694.050 967.050 ;
        RECT 718.950 966.600 721.050 967.050 ;
        RECT 733.950 966.600 736.050 967.050 ;
        RECT 670.950 965.400 736.050 966.600 ;
        RECT 670.950 964.950 673.050 965.400 ;
        RECT 691.950 964.950 694.050 965.400 ;
        RECT 718.950 964.950 721.050 965.400 ;
        RECT 733.950 964.950 736.050 965.400 ;
        RECT 763.950 966.600 766.050 967.050 ;
        RECT 784.950 966.600 787.050 967.050 ;
        RECT 763.950 965.400 787.050 966.600 ;
        RECT 763.950 964.950 766.050 965.400 ;
        RECT 784.950 964.950 787.050 965.400 ;
        RECT 790.950 966.600 793.050 967.050 ;
        RECT 808.950 966.600 811.050 967.050 ;
        RECT 790.950 965.400 811.050 966.600 ;
        RECT 790.950 964.950 793.050 965.400 ;
        RECT 808.950 964.950 811.050 965.400 ;
        RECT 853.950 966.600 856.050 967.050 ;
        RECT 868.950 966.600 871.050 967.050 ;
        RECT 853.950 965.400 871.050 966.600 ;
        RECT 853.950 964.950 856.050 965.400 ;
        RECT 868.950 964.950 871.050 965.400 ;
        RECT 910.950 966.600 913.050 967.050 ;
        RECT 925.950 966.600 928.050 967.050 ;
        RECT 910.950 965.400 928.050 966.600 ;
        RECT 910.950 964.950 913.050 965.400 ;
        RECT 925.950 964.950 928.050 965.400 ;
        RECT 16.950 963.750 19.050 964.200 ;
        RECT 31.950 963.750 34.050 964.200 ;
        RECT 16.950 962.550 34.050 963.750 ;
        RECT 16.950 962.100 19.050 962.550 ;
        RECT 31.950 962.100 34.050 962.550 ;
        RECT 40.950 963.600 43.050 964.200 ;
        RECT 55.950 963.600 58.050 964.050 ;
        RECT 40.950 962.400 58.050 963.600 ;
        RECT 40.950 962.100 43.050 962.400 ;
        RECT 55.950 961.950 58.050 962.400 ;
        RECT 64.950 963.600 67.050 964.200 ;
        RECT 79.950 963.600 82.050 964.050 ;
        RECT 64.950 962.400 82.050 963.600 ;
        RECT 64.950 962.100 67.050 962.400 ;
        RECT 79.950 961.950 82.050 962.400 ;
        RECT 91.950 963.600 94.050 964.200 ;
        RECT 109.950 963.600 112.050 964.200 ;
        RECT 118.950 963.600 121.050 964.050 ;
        RECT 91.950 962.400 121.050 963.600 ;
        RECT 91.950 962.100 94.050 962.400 ;
        RECT 109.950 962.100 112.050 962.400 ;
        RECT 118.950 961.950 121.050 962.400 ;
        RECT 133.950 963.600 136.050 964.200 ;
        RECT 142.950 963.600 145.050 964.050 ;
        RECT 154.950 963.600 157.050 964.200 ;
        RECT 172.950 963.600 175.050 964.200 ;
        RECT 133.950 962.400 138.600 963.600 ;
        RECT 133.950 962.100 136.050 962.400 ;
        RECT 55.950 957.450 58.050 957.900 ;
        RECT 61.950 957.450 64.050 957.900 ;
        RECT 55.950 956.250 64.050 957.450 ;
        RECT 55.950 955.800 58.050 956.250 ;
        RECT 61.950 955.800 64.050 956.250 ;
        RECT 67.950 957.600 70.050 957.900 ;
        RECT 82.950 957.600 85.050 957.900 ;
        RECT 67.950 956.400 85.050 957.600 ;
        RECT 67.950 955.800 70.050 956.400 ;
        RECT 82.950 955.800 85.050 956.400 ;
        RECT 112.950 957.600 115.050 957.900 ;
        RECT 130.950 957.600 133.050 957.900 ;
        RECT 112.950 956.400 133.050 957.600 ;
        RECT 137.400 957.600 138.600 962.400 ;
        RECT 142.950 962.400 175.050 963.600 ;
        RECT 142.950 961.950 145.050 962.400 ;
        RECT 154.950 962.100 157.050 962.400 ;
        RECT 172.950 962.100 175.050 962.400 ;
        RECT 199.950 963.600 202.050 964.050 ;
        RECT 214.950 963.600 217.050 964.200 ;
        RECT 235.950 963.600 238.050 964.200 ;
        RECT 199.950 962.400 238.050 963.600 ;
        RECT 199.950 961.950 202.050 962.400 ;
        RECT 214.950 962.100 217.050 962.400 ;
        RECT 235.950 962.100 238.050 962.400 ;
        RECT 241.950 963.750 244.050 964.200 ;
        RECT 250.950 963.750 253.050 964.200 ;
        RECT 241.950 962.550 253.050 963.750 ;
        RECT 241.950 962.100 244.050 962.550 ;
        RECT 250.950 962.100 253.050 962.550 ;
        RECT 265.950 963.750 268.050 964.200 ;
        RECT 274.950 963.750 277.050 964.200 ;
        RECT 265.950 963.600 277.050 963.750 ;
        RECT 286.950 963.600 289.050 964.200 ;
        RECT 265.950 962.550 289.050 963.600 ;
        RECT 265.950 962.100 268.050 962.550 ;
        RECT 274.950 962.400 289.050 962.550 ;
        RECT 274.950 962.100 277.050 962.400 ;
        RECT 286.950 962.100 289.050 962.400 ;
        RECT 292.950 963.600 295.050 964.200 ;
        RECT 304.950 963.600 307.050 964.050 ;
        RECT 292.950 962.400 307.050 963.600 ;
        RECT 292.950 962.100 295.050 962.400 ;
        RECT 304.950 961.950 307.050 962.400 ;
        RECT 313.950 962.100 316.050 964.200 ;
        RECT 319.950 963.600 322.050 964.200 ;
        RECT 334.950 963.600 337.050 964.200 ;
        RECT 319.950 962.400 337.050 963.600 ;
        RECT 319.950 962.100 322.050 962.400 ;
        RECT 334.950 962.100 337.050 962.400 ;
        RECT 340.950 963.600 343.050 964.200 ;
        RECT 352.950 963.750 355.050 964.200 ;
        RECT 358.950 963.750 361.050 964.200 ;
        RECT 340.950 962.400 351.600 963.600 ;
        RECT 340.950 962.100 343.050 962.400 ;
        RECT 301.950 960.600 304.050 961.050 ;
        RECT 314.400 960.600 315.600 962.100 ;
        RECT 301.950 959.400 315.600 960.600 ;
        RECT 350.400 960.600 351.600 962.400 ;
        RECT 352.950 962.550 361.050 963.750 ;
        RECT 352.950 962.100 355.050 962.550 ;
        RECT 358.950 962.100 361.050 962.550 ;
        RECT 367.950 963.600 370.050 964.050 ;
        RECT 379.950 963.600 382.050 964.200 ;
        RECT 367.950 962.400 382.050 963.600 ;
        RECT 367.950 961.950 370.050 962.400 ;
        RECT 379.950 962.100 382.050 962.400 ;
        RECT 394.950 963.750 397.050 964.200 ;
        RECT 403.950 963.750 406.050 964.200 ;
        RECT 394.950 962.550 406.050 963.750 ;
        RECT 394.950 962.100 397.050 962.550 ;
        RECT 403.950 962.100 406.050 962.550 ;
        RECT 454.950 963.600 457.050 964.200 ;
        RECT 478.950 963.600 481.050 964.200 ;
        RECT 499.950 963.600 502.050 964.200 ;
        RECT 454.950 962.400 477.600 963.600 ;
        RECT 454.950 962.100 457.050 962.400 ;
        RECT 350.400 959.400 384.600 960.600 ;
        RECT 301.950 958.950 304.050 959.400 ;
        RECT 157.950 957.600 160.050 958.050 ;
        RECT 137.400 956.400 160.050 957.600 ;
        RECT 112.950 955.800 115.050 956.400 ;
        RECT 130.950 955.800 133.050 956.400 ;
        RECT 157.950 955.950 160.050 956.400 ;
        RECT 193.950 957.600 196.050 957.900 ;
        RECT 211.950 957.600 214.050 957.900 ;
        RECT 193.950 956.400 214.050 957.600 ;
        RECT 193.950 955.800 196.050 956.400 ;
        RECT 211.950 955.800 214.050 956.400 ;
        RECT 217.950 957.450 220.050 957.900 ;
        RECT 226.950 957.450 229.050 957.900 ;
        RECT 217.950 956.250 229.050 957.450 ;
        RECT 217.950 955.800 220.050 956.250 ;
        RECT 226.950 955.800 229.050 956.250 ;
        RECT 244.950 957.450 247.050 957.900 ;
        RECT 253.950 957.450 256.050 957.900 ;
        RECT 244.950 956.250 256.050 957.450 ;
        RECT 244.950 955.800 247.050 956.250 ;
        RECT 253.950 955.800 256.050 956.250 ;
        RECT 268.950 957.600 271.050 957.900 ;
        RECT 289.950 957.600 292.050 957.900 ;
        RECT 268.950 957.450 292.050 957.600 ;
        RECT 295.950 957.450 298.050 957.900 ;
        RECT 268.950 956.400 298.050 957.450 ;
        RECT 268.950 955.800 271.050 956.400 ;
        RECT 289.950 956.250 298.050 956.400 ;
        RECT 289.950 955.800 292.050 956.250 ;
        RECT 295.950 955.800 298.050 956.250 ;
        RECT 316.950 957.450 319.050 957.900 ;
        RECT 325.950 957.450 328.050 957.900 ;
        RECT 316.950 956.250 328.050 957.450 ;
        RECT 316.950 955.800 319.050 956.250 ;
        RECT 325.950 955.800 328.050 956.250 ;
        RECT 331.950 957.450 334.050 957.900 ;
        RECT 337.950 957.450 340.050 957.900 ;
        RECT 331.950 956.250 340.050 957.450 ;
        RECT 331.950 955.800 334.050 956.250 ;
        RECT 337.950 955.800 340.050 956.250 ;
        RECT 343.800 955.800 345.900 957.900 ;
        RECT 346.950 957.600 349.050 958.050 ;
        RECT 383.400 957.900 384.600 959.400 ;
        RECT 476.400 957.900 477.600 962.400 ;
        RECT 478.950 962.400 502.050 963.600 ;
        RECT 478.950 962.100 481.050 962.400 ;
        RECT 499.950 962.100 502.050 962.400 ;
        RECT 505.950 963.600 508.050 964.200 ;
        RECT 520.950 963.600 523.050 964.200 ;
        RECT 505.950 962.400 523.050 963.600 ;
        RECT 505.950 962.100 508.050 962.400 ;
        RECT 520.950 962.100 523.050 962.400 ;
        RECT 541.950 963.750 544.050 964.200 ;
        RECT 553.950 963.750 556.050 964.200 ;
        RECT 541.950 962.550 556.050 963.750 ;
        RECT 541.950 962.100 544.050 962.550 ;
        RECT 553.950 962.100 556.050 962.550 ;
        RECT 565.950 963.750 568.050 964.200 ;
        RECT 574.950 963.750 577.050 964.200 ;
        RECT 565.950 962.550 577.050 963.750 ;
        RECT 565.950 962.100 568.050 962.550 ;
        RECT 574.950 962.100 577.050 962.550 ;
        RECT 601.950 962.100 604.050 964.200 ;
        RECT 607.950 963.600 610.050 964.050 ;
        RECT 616.950 963.600 619.050 964.200 ;
        RECT 607.950 962.400 619.050 963.600 ;
        RECT 602.400 960.600 603.600 962.100 ;
        RECT 607.950 961.950 610.050 962.400 ;
        RECT 616.950 962.100 619.050 962.400 ;
        RECT 643.950 963.600 646.050 964.200 ;
        RECT 676.950 963.600 679.050 964.050 ;
        RECT 685.950 963.600 688.050 964.200 ;
        RECT 643.950 962.400 688.050 963.600 ;
        RECT 643.950 962.100 646.050 962.400 ;
        RECT 676.950 961.950 679.050 962.400 ;
        RECT 685.950 962.100 688.050 962.400 ;
        RECT 724.950 963.750 727.050 964.200 ;
        RECT 757.950 963.750 760.050 964.200 ;
        RECT 724.950 962.550 760.050 963.750 ;
        RECT 724.950 962.100 727.050 962.550 ;
        RECT 757.950 962.100 760.050 962.550 ;
        RECT 787.950 962.100 790.050 964.200 ;
        RECT 793.950 963.600 796.050 964.050 ;
        RECT 802.950 963.600 805.050 964.200 ;
        RECT 793.950 962.400 805.050 963.600 ;
        RECT 788.400 960.600 789.600 962.100 ;
        RECT 793.950 961.950 796.050 962.400 ;
        RECT 802.950 962.100 805.050 962.400 ;
        RECT 820.950 963.600 823.050 964.050 ;
        RECT 829.950 963.600 832.050 964.050 ;
        RECT 850.950 963.600 853.050 964.200 ;
        RECT 871.950 963.600 874.050 964.200 ;
        RECT 820.950 962.400 853.050 963.600 ;
        RECT 820.950 961.950 823.050 962.400 ;
        RECT 829.950 961.950 832.050 962.400 ;
        RECT 850.950 962.100 853.050 962.400 ;
        RECT 866.400 962.400 874.050 963.600 ;
        RECT 551.400 959.400 567.600 960.600 ;
        RECT 602.400 959.400 618.600 960.600 ;
        RECT 788.400 959.400 798.600 960.600 ;
        RECT 551.400 957.900 552.600 959.400 ;
        RECT 361.950 957.600 364.050 957.900 ;
        RECT 346.950 956.400 364.050 957.600 ;
        RECT 346.950 955.950 349.050 956.400 ;
        RECT 361.950 955.800 364.050 956.400 ;
        RECT 382.950 957.600 385.050 957.900 ;
        RECT 400.950 957.600 403.050 957.900 ;
        RECT 424.950 957.600 427.050 957.900 ;
        RECT 382.950 956.400 427.050 957.600 ;
        RECT 382.950 955.800 385.050 956.400 ;
        RECT 400.950 955.800 403.050 956.400 ;
        RECT 424.950 955.800 427.050 956.400 ;
        RECT 475.950 955.800 478.050 957.900 ;
        RECT 523.950 957.450 526.050 957.900 ;
        RECT 535.950 957.450 538.050 957.900 ;
        RECT 523.950 956.250 538.050 957.450 ;
        RECT 523.950 955.800 526.050 956.250 ;
        RECT 535.950 955.800 538.050 956.250 ;
        RECT 550.950 955.800 553.050 957.900 ;
        RECT 556.950 957.450 559.050 957.900 ;
        RECT 562.950 957.450 565.050 957.900 ;
        RECT 556.950 956.250 565.050 957.450 ;
        RECT 566.400 957.600 567.600 959.400 ;
        RECT 571.950 957.600 574.050 957.900 ;
        RECT 566.400 956.400 574.050 957.600 ;
        RECT 556.950 955.800 559.050 956.250 ;
        RECT 562.950 955.800 565.050 956.250 ;
        RECT 571.950 955.800 574.050 956.400 ;
        RECT 586.950 957.450 589.050 957.900 ;
        RECT 598.950 957.450 601.050 957.900 ;
        RECT 586.950 956.250 601.050 957.450 ;
        RECT 617.400 957.600 618.600 959.400 ;
        RECT 619.950 957.600 622.050 957.900 ;
        RECT 617.400 956.400 622.050 957.600 ;
        RECT 586.950 955.800 589.050 956.250 ;
        RECT 598.950 955.800 601.050 956.250 ;
        RECT 619.950 955.800 622.050 956.400 ;
        RECT 646.950 957.600 649.050 957.900 ;
        RECT 661.950 957.600 664.050 957.900 ;
        RECT 646.950 956.400 664.050 957.600 ;
        RECT 646.950 955.800 649.050 956.400 ;
        RECT 661.950 955.800 664.050 956.400 ;
        RECT 667.950 957.450 670.050 957.900 ;
        RECT 676.950 957.600 679.050 957.900 ;
        RECT 706.950 957.600 709.050 957.900 ;
        RECT 676.950 957.450 709.050 957.600 ;
        RECT 667.950 956.400 709.050 957.450 ;
        RECT 667.950 956.250 679.050 956.400 ;
        RECT 667.950 955.800 670.050 956.250 ;
        RECT 676.950 955.800 679.050 956.250 ;
        RECT 706.950 955.800 709.050 956.400 ;
        RECT 712.950 957.450 715.050 957.900 ;
        RECT 718.950 957.450 721.050 957.900 ;
        RECT 712.950 956.250 721.050 957.450 ;
        RECT 712.950 955.800 715.050 956.250 ;
        RECT 718.950 955.800 721.050 956.250 ;
        RECT 724.950 957.600 727.050 958.050 ;
        RECT 730.950 957.600 733.050 957.900 ;
        RECT 724.950 956.400 733.050 957.600 ;
        RECT 724.950 955.950 727.050 956.400 ;
        RECT 730.950 955.800 733.050 956.400 ;
        RECT 736.950 957.600 739.050 957.900 ;
        RECT 754.950 957.600 757.050 957.900 ;
        RECT 736.950 956.400 757.050 957.600 ;
        RECT 736.950 955.800 739.050 956.400 ;
        RECT 754.950 955.800 757.050 956.400 ;
        RECT 784.950 957.450 787.050 957.900 ;
        RECT 793.950 957.450 796.050 957.900 ;
        RECT 784.950 956.250 796.050 957.450 ;
        RECT 797.400 957.600 798.600 959.400 ;
        RECT 826.950 957.600 829.050 957.900 ;
        RECT 844.950 957.600 847.050 958.050 ;
        RECT 797.400 956.400 847.050 957.600 ;
        RECT 784.950 955.800 787.050 956.250 ;
        RECT 793.950 955.800 796.050 956.250 ;
        RECT 826.950 955.800 829.050 956.400 ;
        RECT 844.950 955.950 847.050 956.400 ;
        RECT 853.950 957.450 856.050 957.900 ;
        RECT 862.950 957.450 865.050 957.900 ;
        RECT 853.950 956.250 865.050 957.450 ;
        RECT 853.950 955.800 856.050 956.250 ;
        RECT 862.950 955.800 865.050 956.250 ;
        RECT 10.950 954.600 13.050 955.050 ;
        RECT 43.950 954.600 46.050 955.050 ;
        RECT 10.950 953.400 46.050 954.600 ;
        RECT 10.950 952.950 13.050 953.400 ;
        RECT 43.950 952.950 46.050 953.400 ;
        RECT 136.950 954.600 139.050 955.050 ;
        RECT 151.950 954.600 154.050 955.050 ;
        RECT 136.950 953.400 154.050 954.600 ;
        RECT 136.950 952.950 139.050 953.400 ;
        RECT 151.950 952.950 154.050 953.400 ;
        RECT 175.950 954.600 178.050 955.050 ;
        RECT 199.950 954.600 202.050 955.050 ;
        RECT 175.950 953.400 202.050 954.600 ;
        RECT 175.950 952.950 178.050 953.400 ;
        RECT 199.950 952.950 202.050 953.400 ;
        RECT 229.950 954.600 232.050 955.050 ;
        RECT 344.400 954.600 345.600 955.800 ;
        RECT 349.950 954.600 352.050 955.050 ;
        RECT 229.950 953.400 342.600 954.600 ;
        RECT 344.400 953.400 352.050 954.600 ;
        RECT 229.950 952.950 232.050 953.400 ;
        RECT 169.950 951.600 172.050 952.050 ;
        RECT 250.950 951.600 253.050 952.050 ;
        RECT 289.950 951.600 292.050 952.050 ;
        RECT 301.950 951.600 304.050 952.050 ;
        RECT 169.950 950.400 304.050 951.600 ;
        RECT 341.400 951.600 342.600 953.400 ;
        RECT 349.950 952.950 352.050 953.400 ;
        RECT 481.950 954.600 484.050 955.050 ;
        RECT 502.950 954.600 505.050 955.050 ;
        RECT 565.950 954.600 568.050 955.050 ;
        RECT 628.950 954.600 631.050 955.050 ;
        RECT 481.950 953.400 568.050 954.600 ;
        RECT 481.950 952.950 484.050 953.400 ;
        RECT 502.950 952.950 505.050 953.400 ;
        RECT 565.950 952.950 568.050 953.400 ;
        RECT 623.400 953.400 631.050 954.600 ;
        RECT 376.950 951.600 379.050 952.050 ;
        RECT 394.950 951.600 397.050 952.050 ;
        RECT 341.400 950.400 397.050 951.600 ;
        RECT 169.950 949.950 172.050 950.400 ;
        RECT 250.950 949.950 253.050 950.400 ;
        RECT 289.950 949.950 292.050 950.400 ;
        RECT 301.950 949.950 304.050 950.400 ;
        RECT 376.950 949.950 379.050 950.400 ;
        RECT 394.950 949.950 397.050 950.400 ;
        RECT 430.950 951.600 433.050 952.050 ;
        RECT 490.950 951.600 493.050 952.050 ;
        RECT 430.950 950.400 493.050 951.600 ;
        RECT 430.950 949.950 433.050 950.400 ;
        RECT 490.950 949.950 493.050 950.400 ;
        RECT 529.950 951.600 532.050 952.050 ;
        RECT 623.400 951.600 624.600 953.400 ;
        RECT 628.950 952.950 631.050 953.400 ;
        RECT 811.950 954.600 814.050 955.050 ;
        RECT 817.950 954.600 820.050 955.050 ;
        RECT 811.950 953.400 820.050 954.600 ;
        RECT 811.950 952.950 814.050 953.400 ;
        RECT 817.950 952.950 820.050 953.400 ;
        RECT 847.950 954.600 850.050 955.050 ;
        RECT 866.400 954.600 867.600 962.400 ;
        RECT 871.950 962.100 874.050 962.400 ;
        RECT 877.950 963.600 880.050 964.200 ;
        RECT 898.950 963.600 901.050 964.200 ;
        RECT 877.950 962.400 901.050 963.600 ;
        RECT 877.950 962.100 880.050 962.400 ;
        RECT 898.950 962.100 901.050 962.400 ;
        RECT 904.950 963.600 907.050 964.200 ;
        RECT 934.950 963.600 937.050 964.050 ;
        RECT 904.950 962.400 937.050 963.600 ;
        RECT 904.950 962.100 907.050 962.400 ;
        RECT 934.950 961.950 937.050 962.400 ;
        RECT 943.950 963.750 946.050 964.200 ;
        RECT 949.950 963.750 952.050 964.200 ;
        RECT 943.950 962.550 952.050 963.750 ;
        RECT 943.950 962.100 946.050 962.550 ;
        RECT 949.950 962.100 952.050 962.550 ;
        RECT 955.950 963.600 958.050 964.200 ;
        RECT 961.800 963.600 963.900 964.050 ;
        RECT 955.950 962.400 963.900 963.600 ;
        RECT 955.950 962.100 958.050 962.400 ;
        RECT 961.800 961.950 963.900 962.400 ;
        RECT 964.950 963.600 967.050 964.050 ;
        RECT 979.950 963.600 982.050 964.200 ;
        RECT 964.950 962.400 982.050 963.600 ;
        RECT 964.950 961.950 967.050 962.400 ;
        RECT 979.950 962.100 982.050 962.400 ;
        RECT 985.950 963.600 988.050 964.050 ;
        RECT 997.950 963.600 1000.050 964.200 ;
        RECT 985.950 962.400 1000.050 963.600 ;
        RECT 985.950 961.950 988.050 962.400 ;
        RECT 997.950 962.100 1000.050 962.400 ;
        RECT 880.950 957.450 883.050 957.900 ;
        RECT 886.950 957.600 889.050 958.050 ;
        RECT 895.950 957.600 898.050 957.900 ;
        RECT 886.950 957.450 898.050 957.600 ;
        RECT 880.950 956.400 898.050 957.450 ;
        RECT 880.950 956.250 889.050 956.400 ;
        RECT 880.950 955.800 883.050 956.250 ;
        RECT 886.950 955.950 889.050 956.250 ;
        RECT 895.950 955.800 898.050 956.400 ;
        RECT 928.950 957.450 931.050 957.900 ;
        RECT 934.950 957.450 937.050 957.900 ;
        RECT 928.950 956.250 937.050 957.450 ;
        RECT 928.950 955.800 931.050 956.250 ;
        RECT 934.950 955.800 937.050 956.250 ;
        RECT 961.950 957.450 964.050 957.900 ;
        RECT 970.950 957.450 973.050 957.900 ;
        RECT 961.950 956.250 973.050 957.450 ;
        RECT 961.950 955.800 964.050 956.250 ;
        RECT 970.950 955.800 973.050 956.250 ;
        RECT 994.950 957.450 997.050 957.900 ;
        RECT 1000.950 957.450 1003.050 957.900 ;
        RECT 994.950 956.250 1003.050 957.450 ;
        RECT 994.950 955.800 997.050 956.250 ;
        RECT 1000.950 955.800 1003.050 956.250 ;
        RECT 847.950 953.400 867.600 954.600 ;
        RECT 868.950 954.600 871.050 955.050 ;
        RECT 922.950 954.600 925.050 955.050 ;
        RECT 946.950 954.600 949.050 955.050 ;
        RECT 868.950 953.400 949.050 954.600 ;
        RECT 847.950 952.950 850.050 953.400 ;
        RECT 868.950 952.950 871.050 953.400 ;
        RECT 922.950 952.950 925.050 953.400 ;
        RECT 946.950 952.950 949.050 953.400 ;
        RECT 529.950 950.400 624.600 951.600 ;
        RECT 697.950 951.600 700.050 952.050 ;
        RECT 769.950 951.600 772.050 952.050 ;
        RECT 778.950 951.600 781.050 952.050 ;
        RECT 848.400 951.600 849.600 952.950 ;
        RECT 697.950 950.400 849.600 951.600 ;
        RECT 889.950 951.600 892.050 952.050 ;
        RECT 901.950 951.600 904.050 952.050 ;
        RECT 889.950 950.400 904.050 951.600 ;
        RECT 529.950 949.950 532.050 950.400 ;
        RECT 697.950 949.950 700.050 950.400 ;
        RECT 769.950 949.950 772.050 950.400 ;
        RECT 778.950 949.950 781.050 950.400 ;
        RECT 889.950 949.950 892.050 950.400 ;
        RECT 901.950 949.950 904.050 950.400 ;
        RECT 22.950 948.600 25.050 949.050 ;
        RECT 67.950 948.600 70.050 949.050 ;
        RECT 22.950 947.400 70.050 948.600 ;
        RECT 22.950 946.950 25.050 947.400 ;
        RECT 67.950 946.950 70.050 947.400 ;
        RECT 304.950 948.600 307.050 949.050 ;
        RECT 331.950 948.600 334.050 949.050 ;
        RECT 304.950 947.400 334.050 948.600 ;
        RECT 304.950 946.950 307.050 947.400 ;
        RECT 331.950 946.950 334.050 947.400 ;
        RECT 367.950 948.600 370.050 949.050 ;
        RECT 457.950 948.600 460.050 949.050 ;
        RECT 367.950 947.400 460.050 948.600 ;
        RECT 367.950 946.950 370.050 947.400 ;
        RECT 457.950 946.950 460.050 947.400 ;
        RECT 265.950 945.600 268.050 946.050 ;
        RECT 274.950 945.600 277.050 946.050 ;
        RECT 265.950 944.400 277.050 945.600 ;
        RECT 265.950 943.950 268.050 944.400 ;
        RECT 274.950 943.950 277.050 944.400 ;
        RECT 466.950 945.600 469.050 946.050 ;
        RECT 625.950 945.600 628.050 946.050 ;
        RECT 466.950 944.400 628.050 945.600 ;
        RECT 466.950 943.950 469.050 944.400 ;
        RECT 625.950 943.950 628.050 944.400 ;
        RECT 742.950 945.600 745.050 946.050 ;
        RECT 805.950 945.600 808.050 946.050 ;
        RECT 874.950 945.600 877.050 946.050 ;
        RECT 742.950 944.400 877.050 945.600 ;
        RECT 742.950 943.950 745.050 944.400 ;
        RECT 805.950 943.950 808.050 944.400 ;
        RECT 874.950 943.950 877.050 944.400 ;
        RECT 1006.950 945.600 1009.050 946.050 ;
        RECT 1015.950 945.600 1018.050 946.050 ;
        RECT 1006.950 944.400 1018.050 945.600 ;
        RECT 1006.950 943.950 1009.050 944.400 ;
        RECT 1015.950 943.950 1018.050 944.400 ;
        RECT 238.950 942.600 241.050 943.050 ;
        RECT 259.950 942.600 262.050 943.050 ;
        RECT 238.950 941.400 262.050 942.600 ;
        RECT 238.950 940.950 241.050 941.400 ;
        RECT 259.950 940.950 262.050 941.400 ;
        RECT 316.950 942.600 319.050 943.050 ;
        RECT 325.950 942.600 328.050 943.050 ;
        RECT 352.950 942.600 355.050 943.050 ;
        RECT 316.950 941.400 355.050 942.600 ;
        RECT 316.950 940.950 319.050 941.400 ;
        RECT 325.950 940.950 328.050 941.400 ;
        RECT 352.950 940.950 355.050 941.400 ;
        RECT 559.950 942.600 562.050 943.050 ;
        RECT 607.950 942.600 610.050 943.050 ;
        RECT 559.950 941.400 610.050 942.600 ;
        RECT 559.950 940.950 562.050 941.400 ;
        RECT 607.950 940.950 610.050 941.400 ;
        RECT 775.950 942.600 778.050 943.050 ;
        RECT 862.950 942.600 865.050 943.050 ;
        RECT 910.950 942.600 913.050 943.050 ;
        RECT 775.950 941.400 865.050 942.600 ;
        RECT 775.950 940.950 778.050 941.400 ;
        RECT 862.950 940.950 865.050 941.400 ;
        RECT 887.400 941.400 913.050 942.600 ;
        RECT 361.950 939.600 364.050 940.050 ;
        RECT 466.950 939.600 469.050 940.050 ;
        RECT 361.950 938.400 469.050 939.600 ;
        RECT 361.950 937.950 364.050 938.400 ;
        RECT 466.950 937.950 469.050 938.400 ;
        RECT 490.950 939.600 493.050 940.050 ;
        RECT 541.950 939.600 544.050 940.050 ;
        RECT 490.950 938.400 544.050 939.600 ;
        RECT 490.950 937.950 493.050 938.400 ;
        RECT 541.950 937.950 544.050 938.400 ;
        RECT 562.950 939.600 565.050 940.050 ;
        RECT 688.950 939.600 691.050 940.050 ;
        RECT 562.950 938.400 691.050 939.600 ;
        RECT 562.950 937.950 565.050 938.400 ;
        RECT 688.950 937.950 691.050 938.400 ;
        RECT 778.950 939.600 781.050 940.050 ;
        RECT 887.400 939.600 888.600 941.400 ;
        RECT 910.950 940.950 913.050 941.400 ;
        RECT 916.950 942.600 919.050 943.050 ;
        RECT 991.950 942.600 994.050 943.050 ;
        RECT 916.950 941.400 994.050 942.600 ;
        RECT 916.950 940.950 919.050 941.400 ;
        RECT 991.950 940.950 994.050 941.400 ;
        RECT 778.950 938.400 888.600 939.600 ;
        RECT 778.950 937.950 781.050 938.400 ;
        RECT 220.950 936.600 223.050 937.050 ;
        RECT 262.950 936.600 265.050 937.050 ;
        RECT 220.950 935.400 265.050 936.600 ;
        RECT 220.950 934.950 223.050 935.400 ;
        RECT 262.950 934.950 265.050 935.400 ;
        RECT 502.950 936.600 505.050 937.050 ;
        RECT 607.950 936.600 610.050 937.050 ;
        RECT 640.950 936.600 643.050 937.050 ;
        RECT 502.950 935.400 540.600 936.600 ;
        RECT 502.950 934.950 505.050 935.400 ;
        RECT 82.950 933.600 85.050 934.050 ;
        RECT 88.950 933.600 91.050 934.050 ;
        RECT 82.950 932.400 91.050 933.600 ;
        RECT 82.950 931.950 85.050 932.400 ;
        RECT 88.950 931.950 91.050 932.400 ;
        RECT 253.950 933.600 256.050 934.050 ;
        RECT 316.950 933.600 319.050 934.050 ;
        RECT 535.950 933.600 538.050 934.050 ;
        RECT 253.950 932.400 319.050 933.600 ;
        RECT 253.950 931.950 256.050 932.400 ;
        RECT 316.950 931.950 319.050 932.400 ;
        RECT 503.400 932.400 538.050 933.600 ;
        RECT 539.400 933.600 540.600 935.400 ;
        RECT 607.950 935.400 643.050 936.600 ;
        RECT 607.950 934.950 610.050 935.400 ;
        RECT 640.950 934.950 643.050 935.400 ;
        RECT 727.950 936.600 730.050 937.050 ;
        RECT 775.950 936.600 778.050 937.050 ;
        RECT 889.950 936.600 892.050 937.050 ;
        RECT 727.950 935.400 778.050 936.600 ;
        RECT 727.950 934.950 730.050 935.400 ;
        RECT 775.950 934.950 778.050 935.400 ;
        RECT 779.400 935.400 892.050 936.600 ;
        RECT 562.950 933.600 565.050 934.050 ;
        RECT 539.400 932.400 565.050 933.600 ;
        RECT 157.950 930.600 160.050 931.050 ;
        RECT 184.950 930.600 187.050 931.050 ;
        RECT 157.950 929.400 187.050 930.600 ;
        RECT 157.950 928.950 160.050 929.400 ;
        RECT 184.950 928.950 187.050 929.400 ;
        RECT 193.950 930.600 196.050 931.050 ;
        RECT 235.950 930.600 238.050 931.050 ;
        RECT 193.950 929.400 238.050 930.600 ;
        RECT 193.950 928.950 196.050 929.400 ;
        RECT 235.950 928.950 238.050 929.400 ;
        RECT 250.950 930.600 253.050 931.050 ;
        RECT 319.950 930.600 322.050 931.050 ;
        RECT 250.950 929.400 322.050 930.600 ;
        RECT 250.950 928.950 253.050 929.400 ;
        RECT 319.950 928.950 322.050 929.400 ;
        RECT 376.950 930.600 379.050 931.050 ;
        RECT 406.950 930.600 409.050 931.050 ;
        RECT 451.950 930.600 454.050 931.050 ;
        RECT 503.400 930.600 504.600 932.400 ;
        RECT 535.950 931.950 538.050 932.400 ;
        RECT 562.950 931.950 565.050 932.400 ;
        RECT 733.950 933.600 736.050 934.050 ;
        RECT 779.400 933.600 780.600 935.400 ;
        RECT 889.950 934.950 892.050 935.400 ;
        RECT 733.950 932.400 780.600 933.600 ;
        RECT 943.950 933.600 946.050 934.050 ;
        RECT 994.950 933.600 997.050 934.050 ;
        RECT 943.950 932.400 997.050 933.600 ;
        RECT 733.950 931.950 736.050 932.400 ;
        RECT 943.950 931.950 946.050 932.400 ;
        RECT 994.950 931.950 997.050 932.400 ;
        RECT 376.950 929.400 504.600 930.600 ;
        RECT 532.950 930.600 535.050 931.050 ;
        RECT 646.950 930.600 649.050 931.050 ;
        RECT 532.950 929.400 649.050 930.600 ;
        RECT 376.950 928.950 379.050 929.400 ;
        RECT 406.950 928.950 409.050 929.400 ;
        RECT 451.950 928.950 454.050 929.400 ;
        RECT 532.950 928.950 535.050 929.400 ;
        RECT 646.950 928.950 649.050 929.400 ;
        RECT 673.950 930.600 676.050 931.050 ;
        RECT 781.950 930.600 784.050 931.050 ;
        RECT 673.950 929.400 784.050 930.600 ;
        RECT 673.950 928.950 676.050 929.400 ;
        RECT 781.950 928.950 784.050 929.400 ;
        RECT 805.950 930.600 808.050 931.050 ;
        RECT 835.950 930.600 838.050 931.050 ;
        RECT 805.950 929.400 838.050 930.600 ;
        RECT 805.950 928.950 808.050 929.400 ;
        RECT 835.950 928.950 838.050 929.400 ;
        RECT 88.950 927.600 91.050 928.050 ;
        RECT 121.950 927.600 124.050 928.050 ;
        RECT 139.950 927.600 142.050 928.050 ;
        RECT 88.950 926.400 142.050 927.600 ;
        RECT 88.950 925.950 91.050 926.400 ;
        RECT 121.950 925.950 124.050 926.400 ;
        RECT 139.950 925.950 142.050 926.400 ;
        RECT 178.950 927.600 181.050 928.050 ;
        RECT 238.950 927.600 241.050 928.050 ;
        RECT 178.950 926.400 241.050 927.600 ;
        RECT 178.950 925.950 181.050 926.400 ;
        RECT 238.950 925.950 241.050 926.400 ;
        RECT 247.950 927.600 250.050 928.050 ;
        RECT 331.950 927.600 334.050 928.050 ;
        RECT 247.950 926.400 334.050 927.600 ;
        RECT 247.950 925.950 250.050 926.400 ;
        RECT 331.950 925.950 334.050 926.400 ;
        RECT 412.950 927.600 415.050 928.050 ;
        RECT 448.950 927.600 451.050 928.050 ;
        RECT 412.950 926.400 451.050 927.600 ;
        RECT 412.950 925.950 415.050 926.400 ;
        RECT 448.950 925.950 451.050 926.400 ;
        RECT 457.950 927.600 460.050 928.050 ;
        RECT 496.950 927.600 499.050 928.050 ;
        RECT 457.950 926.400 499.050 927.600 ;
        RECT 457.950 925.950 460.050 926.400 ;
        RECT 496.950 925.950 499.050 926.400 ;
        RECT 688.950 927.600 691.050 928.050 ;
        RECT 700.950 927.600 703.050 928.050 ;
        RECT 688.950 926.400 703.050 927.600 ;
        RECT 688.950 925.950 691.050 926.400 ;
        RECT 700.950 925.950 703.050 926.400 ;
        RECT 748.950 927.600 751.050 928.050 ;
        RECT 778.950 927.600 781.050 928.050 ;
        RECT 748.950 926.400 781.050 927.600 ;
        RECT 748.950 925.950 751.050 926.400 ;
        RECT 778.950 925.950 781.050 926.400 ;
        RECT 865.950 927.600 868.050 928.050 ;
        RECT 898.950 927.600 901.050 928.050 ;
        RECT 865.950 926.400 901.050 927.600 ;
        RECT 865.950 925.950 868.050 926.400 ;
        RECT 898.950 925.950 901.050 926.400 ;
        RECT 913.950 927.600 916.050 928.050 ;
        RECT 964.950 927.600 967.050 928.050 ;
        RECT 913.950 926.400 967.050 927.600 ;
        RECT 913.950 925.950 916.050 926.400 ;
        RECT 964.950 925.950 967.050 926.400 ;
        RECT 43.950 924.600 46.050 925.050 ;
        RECT 109.950 924.600 112.050 925.050 ;
        RECT 127.950 924.600 130.050 925.050 ;
        RECT 142.950 924.600 145.050 925.050 ;
        RECT 43.950 923.400 69.600 924.600 ;
        RECT 43.950 922.950 46.050 923.400 ;
        RECT 68.400 922.050 69.600 923.400 ;
        RECT 109.950 923.400 145.050 924.600 ;
        RECT 109.950 922.950 112.050 923.400 ;
        RECT 127.950 922.950 130.050 923.400 ;
        RECT 142.950 922.950 145.050 923.400 ;
        RECT 205.950 924.600 208.050 925.050 ;
        RECT 229.950 924.600 232.050 925.050 ;
        RECT 241.950 924.600 244.050 924.900 ;
        RECT 205.950 923.400 244.050 924.600 ;
        RECT 205.950 922.950 208.050 923.400 ;
        RECT 229.950 922.950 232.050 923.400 ;
        RECT 241.950 922.800 244.050 923.400 ;
        RECT 259.950 924.600 262.050 925.050 ;
        RECT 310.950 924.600 313.050 925.050 ;
        RECT 259.950 923.400 313.050 924.600 ;
        RECT 259.950 922.950 262.050 923.400 ;
        RECT 310.950 922.950 313.050 923.400 ;
        RECT 430.950 924.600 433.050 925.050 ;
        RECT 436.950 924.600 439.050 925.050 ;
        RECT 472.950 924.600 475.050 925.050 ;
        RECT 430.950 923.400 475.050 924.600 ;
        RECT 430.950 922.950 433.050 923.400 ;
        RECT 436.950 922.950 439.050 923.400 ;
        RECT 472.950 922.950 475.050 923.400 ;
        RECT 511.950 924.600 514.050 925.050 ;
        RECT 523.950 924.600 526.050 925.050 ;
        RECT 544.950 924.600 547.050 925.050 ;
        RECT 511.950 923.400 547.050 924.600 ;
        RECT 511.950 922.950 514.050 923.400 ;
        RECT 523.950 922.950 526.050 923.400 ;
        RECT 544.950 922.950 547.050 923.400 ;
        RECT 550.950 924.600 553.050 925.050 ;
        RECT 613.950 924.600 616.050 925.050 ;
        RECT 550.950 923.400 616.050 924.600 ;
        RECT 550.950 922.950 553.050 923.400 ;
        RECT 613.950 922.950 616.050 923.400 ;
        RECT 640.950 924.600 643.050 925.050 ;
        RECT 736.950 924.600 739.050 925.050 ;
        RECT 640.950 923.400 739.050 924.600 ;
        RECT 640.950 922.950 643.050 923.400 ;
        RECT 736.950 922.950 739.050 923.400 ;
        RECT 781.950 924.600 784.050 925.050 ;
        RECT 820.950 924.600 823.050 925.050 ;
        RECT 781.950 923.400 823.050 924.600 ;
        RECT 781.950 922.950 784.050 923.400 ;
        RECT 820.950 922.950 823.050 923.400 ;
        RECT 850.950 924.600 853.050 925.050 ;
        RECT 868.950 924.600 871.050 925.050 ;
        RECT 850.950 923.400 871.050 924.600 ;
        RECT 850.950 922.950 853.050 923.400 ;
        RECT 868.950 922.950 871.050 923.400 ;
        RECT 967.950 924.600 970.050 925.050 ;
        RECT 985.950 924.600 988.050 925.050 ;
        RECT 967.950 923.400 988.050 924.600 ;
        RECT 967.950 922.950 970.050 923.400 ;
        RECT 985.950 922.950 988.050 923.400 ;
        RECT 67.950 921.600 70.050 922.050 ;
        RECT 97.950 921.600 100.050 922.050 ;
        RECT 67.950 920.400 100.050 921.600 ;
        RECT 67.950 919.950 70.050 920.400 ;
        RECT 97.950 919.950 100.050 920.400 ;
        RECT 19.950 918.750 22.050 919.200 ;
        RECT 31.950 918.750 34.050 919.200 ;
        RECT 19.950 918.600 34.050 918.750 ;
        RECT 37.950 918.600 40.050 919.050 ;
        RECT 19.950 917.550 40.050 918.600 ;
        RECT 19.950 917.100 22.050 917.550 ;
        RECT 31.950 917.400 40.050 917.550 ;
        RECT 31.950 917.100 34.050 917.400 ;
        RECT 37.950 916.950 40.050 917.400 ;
        RECT 49.950 917.100 52.050 919.200 ;
        RECT 115.950 918.600 118.050 919.200 ;
        RECT 133.950 918.600 136.050 919.200 ;
        RECT 115.950 917.400 136.050 918.600 ;
        RECT 115.950 917.100 118.050 917.400 ;
        RECT 133.950 917.100 136.050 917.400 ;
        RECT 151.950 918.750 154.050 919.200 ;
        RECT 163.950 918.750 166.050 919.200 ;
        RECT 151.950 917.550 166.050 918.750 ;
        RECT 151.950 917.100 154.050 917.550 ;
        RECT 163.950 917.100 166.050 917.550 ;
        RECT 211.950 918.750 214.050 919.200 ;
        RECT 217.950 918.750 220.050 919.200 ;
        RECT 211.950 917.550 220.050 918.750 ;
        RECT 211.950 917.100 214.050 917.550 ;
        RECT 217.950 917.100 220.050 917.550 ;
        RECT 235.950 918.600 238.050 919.200 ;
        RECT 250.950 918.600 253.050 919.200 ;
        RECT 262.950 918.600 265.050 919.050 ;
        RECT 235.950 917.400 265.050 918.600 ;
        RECT 235.950 917.100 238.050 917.400 ;
        RECT 250.950 917.100 253.050 917.400 ;
        RECT 50.400 915.600 51.600 917.100 ;
        RECT 262.950 916.950 265.050 917.400 ;
        RECT 274.950 917.100 277.050 919.200 ;
        RECT 287.400 917.400 294.600 918.600 ;
        RECT 79.950 915.600 82.050 916.050 ;
        RECT 50.400 914.400 82.050 915.600 ;
        RECT 275.400 915.600 276.600 917.100 ;
        RECT 287.400 915.600 288.600 917.400 ;
        RECT 275.400 914.400 288.600 915.600 ;
        RECT 293.400 915.600 294.600 917.400 ;
        RECT 298.950 917.100 301.050 919.200 ;
        RECT 325.950 918.600 328.050 919.200 ;
        RECT 343.950 918.600 346.050 919.200 ;
        RECT 325.950 917.400 346.050 918.600 ;
        RECT 325.950 917.100 328.050 917.400 ;
        RECT 343.950 917.100 346.050 917.400 ;
        RECT 385.950 917.100 388.050 919.200 ;
        RECT 391.950 918.750 394.050 919.200 ;
        RECT 421.950 918.750 424.050 919.200 ;
        RECT 391.950 917.550 424.050 918.750 ;
        RECT 391.950 917.100 394.050 917.550 ;
        RECT 421.950 917.100 424.050 917.550 ;
        RECT 451.950 918.600 454.050 919.200 ;
        RECT 466.950 918.600 469.050 919.050 ;
        RECT 451.950 917.400 469.050 918.600 ;
        RECT 475.950 918.600 478.050 922.050 ;
        RECT 610.950 921.600 613.050 922.050 ;
        RECT 730.950 921.600 733.050 922.050 ;
        RECT 581.400 920.400 733.050 921.600 ;
        RECT 581.400 919.200 582.600 920.400 ;
        RECT 610.950 919.950 613.050 920.400 ;
        RECT 478.950 918.600 481.050 919.200 ;
        RECT 475.950 918.000 481.050 918.600 ;
        RECT 476.400 917.400 481.050 918.000 ;
        RECT 451.950 917.100 454.050 917.400 ;
        RECT 299.400 915.600 300.600 917.100 ;
        RECT 313.950 915.600 316.050 916.050 ;
        RECT 293.400 914.400 316.050 915.600 ;
        RECT 79.950 913.950 82.050 914.400 ;
        RECT 313.950 913.950 316.050 914.400 ;
        RECT 386.400 913.050 387.600 917.100 ;
        RECT 466.950 916.950 469.050 917.400 ;
        RECT 478.950 917.100 481.050 917.400 ;
        RECT 574.950 918.750 577.050 919.200 ;
        RECT 580.950 918.750 583.050 919.200 ;
        RECT 574.950 917.550 583.050 918.750 ;
        RECT 574.950 917.100 577.050 917.550 ;
        RECT 580.950 917.100 583.050 917.550 ;
        RECT 592.950 917.100 595.050 919.200 ;
        RECT 598.950 918.750 601.050 919.200 ;
        RECT 604.950 918.750 607.050 919.200 ;
        RECT 598.950 917.550 607.050 918.750 ;
        RECT 598.950 917.100 601.050 917.550 ;
        RECT 604.950 917.100 607.050 917.550 ;
        RECT 625.950 918.750 628.050 919.200 ;
        RECT 640.950 918.750 643.050 919.200 ;
        RECT 625.950 917.550 643.050 918.750 ;
        RECT 625.950 917.100 628.050 917.550 ;
        RECT 640.950 917.100 643.050 917.550 ;
        RECT 562.950 915.600 565.050 916.050 ;
        RECT 562.950 914.400 570.600 915.600 ;
        RECT 562.950 913.950 565.050 914.400 ;
        RECT 22.950 912.600 25.050 912.900 ;
        RECT 46.950 912.600 49.050 912.900 ;
        RECT 22.950 911.400 49.050 912.600 ;
        RECT 22.950 910.800 25.050 911.400 ;
        RECT 46.950 910.800 49.050 911.400 ;
        RECT 70.950 912.600 73.050 912.900 ;
        RECT 82.950 912.600 85.050 913.050 ;
        RECT 91.950 912.600 94.050 912.900 ;
        RECT 112.950 912.600 115.050 912.900 ;
        RECT 70.950 911.400 85.050 912.600 ;
        RECT 70.950 910.800 73.050 911.400 ;
        RECT 82.950 910.950 85.050 911.400 ;
        RECT 89.400 911.400 115.050 912.600 ;
        RECT 52.950 909.600 55.050 910.050 ;
        RECT 89.400 909.600 90.600 911.400 ;
        RECT 91.950 910.800 94.050 911.400 ;
        RECT 112.950 910.800 115.050 911.400 ;
        RECT 127.950 912.450 130.050 912.900 ;
        RECT 136.950 912.450 139.050 912.900 ;
        RECT 127.950 911.250 139.050 912.450 ;
        RECT 127.950 910.800 130.050 911.250 ;
        RECT 136.950 910.800 139.050 911.250 ;
        RECT 208.950 912.600 211.050 912.900 ;
        RECT 220.950 912.600 223.050 913.050 ;
        RECT 208.950 911.400 223.050 912.600 ;
        RECT 208.950 910.800 211.050 911.400 ;
        RECT 220.950 910.950 223.050 911.400 ;
        RECT 232.950 912.600 235.050 912.900 ;
        RECT 259.950 912.600 262.050 913.050 ;
        RECT 232.950 911.400 262.050 912.600 ;
        RECT 232.950 910.800 235.050 911.400 ;
        RECT 259.950 910.950 262.050 911.400 ;
        RECT 265.950 912.600 268.050 913.050 ;
        RECT 271.950 912.600 274.050 912.900 ;
        RECT 265.950 911.400 274.050 912.600 ;
        RECT 265.950 910.950 268.050 911.400 ;
        RECT 271.950 910.800 274.050 911.400 ;
        RECT 289.950 912.600 292.050 913.050 ;
        RECT 295.950 912.600 298.050 912.900 ;
        RECT 289.950 911.400 298.050 912.600 ;
        RECT 289.950 910.950 292.050 911.400 ;
        RECT 295.950 910.800 298.050 911.400 ;
        RECT 331.950 912.600 334.050 913.050 ;
        RECT 346.950 912.600 349.050 912.900 ;
        RECT 364.950 912.600 367.050 912.900 ;
        RECT 331.950 911.400 367.050 912.600 ;
        RECT 331.950 910.950 334.050 911.400 ;
        RECT 346.950 910.800 349.050 911.400 ;
        RECT 364.950 910.800 367.050 911.400 ;
        RECT 382.950 911.400 387.600 913.050 ;
        RECT 436.950 912.450 439.050 912.900 ;
        RECT 448.950 912.450 451.050 912.900 ;
        RECT 382.950 910.950 387.000 911.400 ;
        RECT 436.950 911.250 451.050 912.450 ;
        RECT 436.950 910.800 439.050 911.250 ;
        RECT 448.950 910.800 451.050 911.250 ;
        RECT 466.950 912.450 469.050 912.900 ;
        RECT 475.950 912.450 478.050 912.900 ;
        RECT 466.950 911.250 478.050 912.450 ;
        RECT 466.950 910.800 469.050 911.250 ;
        RECT 475.950 910.800 478.050 911.250 ;
        RECT 490.950 912.600 493.050 913.050 ;
        RECT 499.950 912.600 502.050 912.900 ;
        RECT 490.950 911.400 502.050 912.600 ;
        RECT 490.950 910.950 493.050 911.400 ;
        RECT 499.950 910.800 502.050 911.400 ;
        RECT 505.950 912.450 508.050 912.900 ;
        RECT 511.950 912.450 514.050 912.900 ;
        RECT 505.950 911.250 514.050 912.450 ;
        RECT 505.950 910.800 508.050 911.250 ;
        RECT 511.950 910.800 514.050 911.250 ;
        RECT 526.950 912.600 529.050 912.900 ;
        RECT 532.950 912.600 535.050 913.050 ;
        RECT 526.950 911.400 535.050 912.600 ;
        RECT 569.400 912.600 570.600 914.400 ;
        RECT 571.950 912.600 574.050 912.900 ;
        RECT 569.400 911.400 574.050 912.600 ;
        RECT 526.950 910.800 529.050 911.400 ;
        RECT 532.950 910.950 535.050 911.400 ;
        RECT 571.950 910.800 574.050 911.400 ;
        RECT 580.950 912.600 583.050 913.050 ;
        RECT 589.950 912.600 592.050 912.900 ;
        RECT 580.950 911.400 592.050 912.600 ;
        RECT 580.950 910.950 583.050 911.400 ;
        RECT 589.950 910.800 592.050 911.400 ;
        RECT 141.000 909.600 145.050 910.050 ;
        RECT 151.950 909.600 154.050 910.050 ;
        RECT 181.950 909.600 184.050 910.050 ;
        RECT 52.950 908.400 90.600 909.600 ;
        RECT 140.400 908.400 184.050 909.600 ;
        RECT 52.950 907.950 55.050 908.400 ;
        RECT 141.000 907.950 145.050 908.400 ;
        RECT 151.950 907.950 154.050 908.400 ;
        RECT 181.950 907.950 184.050 908.400 ;
        RECT 262.950 909.600 265.050 910.050 ;
        RECT 277.950 909.600 280.050 910.050 ;
        RECT 262.950 908.400 280.050 909.600 ;
        RECT 262.950 907.950 265.050 908.400 ;
        RECT 277.950 907.950 280.050 908.400 ;
        RECT 394.950 909.600 397.050 910.050 ;
        RECT 409.950 909.600 412.050 910.050 ;
        RECT 448.950 909.600 451.050 909.750 ;
        RECT 394.950 908.400 451.050 909.600 ;
        RECT 593.400 909.600 594.600 917.100 ;
        RECT 644.400 912.900 645.600 920.400 ;
        RECT 730.950 919.950 733.050 920.400 ;
        RECT 880.950 921.600 883.050 922.050 ;
        RECT 910.950 921.600 913.050 922.050 ;
        RECT 946.950 921.600 949.050 922.050 ;
        RECT 880.950 920.400 949.050 921.600 ;
        RECT 880.950 919.950 883.050 920.400 ;
        RECT 910.950 919.950 913.050 920.400 ;
        RECT 946.950 919.950 949.050 920.400 ;
        RECT 979.950 919.950 982.050 922.050 ;
        RECT 646.950 918.750 649.050 919.200 ;
        RECT 655.950 918.750 658.050 919.200 ;
        RECT 646.950 917.550 658.050 918.750 ;
        RECT 646.950 917.100 649.050 917.550 ;
        RECT 655.950 917.100 658.050 917.550 ;
        RECT 667.950 918.600 670.050 919.200 ;
        RECT 691.950 918.600 694.050 919.200 ;
        RECT 696.000 918.600 700.050 919.050 ;
        RECT 667.950 917.400 694.050 918.600 ;
        RECT 667.950 917.100 670.050 917.400 ;
        RECT 691.950 917.100 694.050 917.400 ;
        RECT 695.400 916.950 700.050 918.600 ;
        RECT 703.950 918.750 706.050 919.200 ;
        RECT 712.950 918.750 715.050 919.200 ;
        RECT 703.950 918.600 715.050 918.750 ;
        RECT 736.950 918.600 739.050 919.200 ;
        RECT 703.950 917.550 739.050 918.600 ;
        RECT 703.950 917.100 706.050 917.550 ;
        RECT 712.950 917.400 739.050 917.550 ;
        RECT 712.950 917.100 715.050 917.400 ;
        RECT 736.950 917.100 739.050 917.400 ;
        RECT 757.950 918.600 760.050 919.200 ;
        RECT 766.950 918.600 769.050 919.050 ;
        RECT 757.950 917.400 769.050 918.600 ;
        RECT 757.950 917.100 760.050 917.400 ;
        RECT 766.950 916.950 769.050 917.400 ;
        RECT 811.950 918.750 814.050 919.200 ;
        RECT 817.950 918.750 820.050 919.200 ;
        RECT 811.950 917.550 820.050 918.750 ;
        RECT 811.950 917.100 814.050 917.550 ;
        RECT 817.950 917.100 820.050 917.550 ;
        RECT 835.950 918.750 838.050 919.200 ;
        RECT 841.950 918.750 844.050 919.200 ;
        RECT 835.950 918.600 844.050 918.750 ;
        RECT 856.950 918.600 859.050 919.200 ;
        RECT 835.950 917.550 859.050 918.600 ;
        RECT 835.950 917.100 838.050 917.550 ;
        RECT 841.950 917.400 859.050 917.550 ;
        RECT 841.950 917.100 844.050 917.400 ;
        RECT 856.950 917.100 859.050 917.400 ;
        RECT 868.950 918.600 871.050 919.050 ;
        RECT 922.950 918.600 925.050 919.050 ;
        RECT 937.950 918.600 940.050 919.050 ;
        RECT 868.950 917.400 940.050 918.600 ;
        RECT 868.950 916.950 871.050 917.400 ;
        RECT 922.950 916.950 925.050 917.400 ;
        RECT 937.950 916.950 940.050 917.400 ;
        RECT 976.950 917.100 979.050 919.200 ;
        RECT 695.400 912.900 696.600 916.950 ;
        RECT 610.950 912.450 613.050 912.900 ;
        RECT 616.950 912.450 619.050 912.900 ;
        RECT 610.950 911.250 619.050 912.450 ;
        RECT 610.950 910.800 613.050 911.250 ;
        RECT 616.950 910.800 619.050 911.250 ;
        RECT 643.950 910.800 646.050 912.900 ;
        RECT 694.950 910.800 697.050 912.900 ;
        RECT 700.950 912.450 703.050 912.900 ;
        RECT 709.950 912.600 712.050 912.900 ;
        RECT 733.950 912.600 736.050 912.900 ;
        RECT 709.950 912.450 736.050 912.600 ;
        RECT 700.950 911.400 736.050 912.450 ;
        RECT 700.950 911.250 712.050 911.400 ;
        RECT 700.950 910.800 703.050 911.250 ;
        RECT 709.950 910.800 712.050 911.250 ;
        RECT 733.950 910.800 736.050 911.400 ;
        RECT 769.950 912.450 772.050 912.900 ;
        RECT 778.950 912.450 781.050 912.900 ;
        RECT 769.950 911.250 781.050 912.450 ;
        RECT 769.950 910.800 772.050 911.250 ;
        RECT 778.950 910.800 781.050 911.250 ;
        RECT 784.950 912.600 787.050 912.900 ;
        RECT 802.950 912.600 805.050 912.900 ;
        RECT 784.950 911.400 805.050 912.600 ;
        RECT 784.950 910.800 787.050 911.400 ;
        RECT 802.950 910.800 805.050 911.400 ;
        RECT 820.950 912.600 823.050 913.050 ;
        RECT 832.950 912.600 835.050 912.900 ;
        RECT 820.950 911.400 835.050 912.600 ;
        RECT 820.950 910.950 823.050 911.400 ;
        RECT 832.950 910.800 835.050 911.400 ;
        RECT 877.950 912.600 880.050 912.900 ;
        RECT 886.800 912.600 888.900 913.050 ;
        RECT 877.950 911.400 888.900 912.600 ;
        RECT 877.950 910.800 880.050 911.400 ;
        RECT 886.800 910.950 888.900 911.400 ;
        RECT 889.950 912.600 892.050 913.050 ;
        RECT 895.950 912.600 898.050 912.900 ;
        RECT 889.950 911.400 898.050 912.600 ;
        RECT 889.950 910.950 892.050 911.400 ;
        RECT 895.950 910.800 898.050 911.400 ;
        RECT 901.950 912.600 904.050 912.900 ;
        RECT 934.950 912.600 937.050 913.050 ;
        RECT 952.950 912.600 955.050 912.900 ;
        RECT 901.950 911.400 955.050 912.600 ;
        RECT 901.950 910.800 904.050 911.400 ;
        RECT 934.950 910.950 937.050 911.400 ;
        RECT 952.950 910.800 955.050 911.400 ;
        RECT 598.950 909.600 601.050 910.050 ;
        RECT 593.400 908.400 601.050 909.600 ;
        RECT 394.950 907.950 397.050 908.400 ;
        RECT 409.950 907.950 412.050 908.400 ;
        RECT 448.950 907.650 451.050 908.400 ;
        RECT 598.950 907.950 601.050 908.400 ;
        RECT 625.950 909.600 628.050 910.050 ;
        RECT 640.950 909.600 643.050 910.050 ;
        RECT 625.950 908.400 643.050 909.600 ;
        RECT 625.950 907.950 628.050 908.400 ;
        RECT 640.950 907.950 643.050 908.400 ;
        RECT 742.950 909.600 745.050 910.050 ;
        RECT 760.950 909.600 763.050 910.050 ;
        RECT 742.950 908.400 763.050 909.600 ;
        RECT 742.950 907.950 745.050 908.400 ;
        RECT 760.950 907.950 763.050 908.400 ;
        RECT 847.950 909.600 850.050 910.050 ;
        RECT 853.950 909.600 856.050 910.050 ;
        RECT 862.950 909.600 865.050 910.050 ;
        RECT 847.950 908.400 865.050 909.600 ;
        RECT 847.950 907.950 850.050 908.400 ;
        RECT 853.950 907.950 856.050 908.400 ;
        RECT 862.950 907.950 865.050 908.400 ;
        RECT 961.950 909.600 964.050 910.050 ;
        RECT 967.950 909.600 970.050 910.050 ;
        RECT 961.950 908.400 970.050 909.600 ;
        RECT 961.950 907.950 964.050 908.400 ;
        RECT 967.950 907.950 970.050 908.400 ;
        RECT 977.400 907.050 978.600 917.100 ;
        RECT 980.400 912.900 981.600 919.950 ;
        RECT 994.950 918.750 997.050 919.200 ;
        RECT 1000.950 918.750 1003.050 919.200 ;
        RECT 994.950 917.550 1003.050 918.750 ;
        RECT 994.950 917.100 997.050 917.550 ;
        RECT 1000.950 917.100 1003.050 917.550 ;
        RECT 979.950 910.800 982.050 912.900 ;
        RECT 994.950 909.600 997.050 910.050 ;
        RECT 1009.950 909.600 1012.050 910.050 ;
        RECT 994.950 908.400 1012.050 909.600 ;
        RECT 994.950 907.950 997.050 908.400 ;
        RECT 1009.950 907.950 1012.050 908.400 ;
        RECT 160.950 906.600 163.050 907.050 ;
        RECT 193.950 906.600 196.050 907.050 ;
        RECT 160.950 905.400 196.050 906.600 ;
        RECT 160.950 904.950 163.050 905.400 ;
        RECT 193.950 904.950 196.050 905.400 ;
        RECT 322.950 906.600 325.050 907.050 ;
        RECT 379.950 906.600 382.050 907.050 ;
        RECT 322.950 905.400 382.050 906.600 ;
        RECT 322.950 904.950 325.050 905.400 ;
        RECT 379.950 904.950 382.050 905.400 ;
        RECT 421.950 906.600 424.050 907.050 ;
        RECT 427.950 906.600 430.050 907.050 ;
        RECT 457.950 906.600 460.050 907.050 ;
        RECT 421.950 905.400 460.050 906.600 ;
        RECT 421.950 904.950 424.050 905.400 ;
        RECT 427.950 904.950 430.050 905.400 ;
        RECT 457.950 904.950 460.050 905.400 ;
        RECT 553.950 906.600 556.050 907.050 ;
        RECT 595.950 906.600 598.050 907.050 ;
        RECT 553.950 905.400 598.050 906.600 ;
        RECT 553.950 904.950 556.050 905.400 ;
        RECT 595.950 904.950 598.050 905.400 ;
        RECT 628.950 906.600 631.050 907.050 ;
        RECT 664.950 906.600 667.050 907.050 ;
        RECT 628.950 905.400 667.050 906.600 ;
        RECT 628.950 904.950 631.050 905.400 ;
        RECT 664.950 904.950 667.050 905.400 ;
        RECT 670.950 906.600 673.050 907.050 ;
        RECT 715.950 906.600 718.050 907.050 ;
        RECT 727.950 906.600 730.050 907.050 ;
        RECT 670.950 905.400 730.050 906.600 ;
        RECT 670.950 904.950 673.050 905.400 ;
        RECT 715.950 904.950 718.050 905.400 ;
        RECT 727.950 904.950 730.050 905.400 ;
        RECT 739.950 906.600 742.050 907.050 ;
        RECT 748.950 906.600 751.050 907.050 ;
        RECT 739.950 905.400 751.050 906.600 ;
        RECT 739.950 904.950 742.050 905.400 ;
        RECT 748.950 904.950 751.050 905.400 ;
        RECT 838.950 906.600 841.050 907.050 ;
        RECT 922.950 906.600 925.050 907.050 ;
        RECT 928.950 906.600 931.050 907.050 ;
        RECT 838.950 905.400 931.050 906.600 ;
        RECT 838.950 904.950 841.050 905.400 ;
        RECT 922.950 904.950 925.050 905.400 ;
        RECT 928.950 904.950 931.050 905.400 ;
        RECT 967.950 906.600 970.050 906.900 ;
        RECT 973.950 906.600 976.050 907.050 ;
        RECT 967.950 905.400 976.050 906.600 ;
        RECT 977.400 905.400 982.050 907.050 ;
        RECT 967.950 904.800 970.050 905.400 ;
        RECT 973.950 904.950 976.050 905.400 ;
        RECT 978.000 904.950 982.050 905.400 ;
        RECT 10.950 903.600 13.050 904.050 ;
        RECT 16.950 903.600 19.050 904.050 ;
        RECT 52.950 903.600 55.050 904.050 ;
        RECT 10.950 902.400 55.050 903.600 ;
        RECT 10.950 901.950 13.050 902.400 ;
        RECT 16.950 901.950 19.050 902.400 ;
        RECT 52.950 901.950 55.050 902.400 ;
        RECT 382.950 903.600 385.050 904.050 ;
        RECT 538.950 903.600 541.050 904.050 ;
        RECT 610.950 903.600 613.050 904.050 ;
        RECT 382.950 902.400 411.600 903.600 ;
        RECT 382.950 901.950 385.050 902.400 ;
        RECT 410.400 901.050 411.600 902.400 ;
        RECT 538.950 902.400 613.050 903.600 ;
        RECT 538.950 901.950 541.050 902.400 ;
        RECT 610.950 901.950 613.050 902.400 ;
        RECT 655.950 903.600 658.050 904.050 ;
        RECT 751.950 903.600 754.050 904.050 ;
        RECT 913.950 903.600 916.050 904.050 ;
        RECT 655.950 902.400 754.050 903.600 ;
        RECT 655.950 901.950 658.050 902.400 ;
        RECT 751.950 901.950 754.050 902.400 ;
        RECT 842.400 902.400 916.050 903.600 ;
        RECT 202.950 900.600 205.050 901.050 ;
        RECT 226.950 900.600 229.050 901.050 ;
        RECT 202.950 899.400 229.050 900.600 ;
        RECT 202.950 898.950 205.050 899.400 ;
        RECT 226.950 898.950 229.050 899.400 ;
        RECT 286.950 900.600 289.050 901.050 ;
        RECT 301.950 900.600 304.050 901.050 ;
        RECT 346.950 900.600 349.050 901.050 ;
        RECT 286.950 899.400 349.050 900.600 ;
        RECT 286.950 898.950 289.050 899.400 ;
        RECT 301.950 898.950 304.050 899.400 ;
        RECT 346.950 898.950 349.050 899.400 ;
        RECT 409.950 900.600 412.050 901.050 ;
        RECT 439.950 900.600 442.050 901.050 ;
        RECT 460.950 900.600 463.050 901.050 ;
        RECT 409.950 899.400 463.050 900.600 ;
        RECT 409.950 898.950 412.050 899.400 ;
        RECT 439.950 898.950 442.050 899.400 ;
        RECT 460.950 898.950 463.050 899.400 ;
        RECT 547.950 900.600 550.050 901.050 ;
        RECT 586.950 900.600 589.050 901.050 ;
        RECT 607.950 900.600 610.050 901.050 ;
        RECT 547.950 899.400 610.050 900.600 ;
        RECT 547.950 898.950 550.050 899.400 ;
        RECT 586.950 898.950 589.050 899.400 ;
        RECT 607.950 898.950 610.050 899.400 ;
        RECT 649.950 900.600 652.050 901.050 ;
        RECT 703.950 900.600 706.050 901.050 ;
        RECT 649.950 899.400 706.050 900.600 ;
        RECT 649.950 898.950 652.050 899.400 ;
        RECT 703.950 898.950 706.050 899.400 ;
        RECT 772.950 900.600 775.050 901.050 ;
        RECT 842.400 900.600 843.600 902.400 ;
        RECT 913.950 901.950 916.050 902.400 ;
        RECT 985.950 903.600 988.050 904.050 ;
        RECT 991.950 903.600 994.050 904.050 ;
        RECT 1003.950 903.600 1006.050 904.050 ;
        RECT 985.950 902.400 1006.050 903.600 ;
        RECT 985.950 901.950 988.050 902.400 ;
        RECT 991.950 901.950 994.050 902.400 ;
        RECT 1003.950 901.950 1006.050 902.400 ;
        RECT 772.950 899.400 843.600 900.600 ;
        RECT 862.950 900.600 865.050 901.050 ;
        RECT 871.950 900.600 874.050 901.050 ;
        RECT 862.950 899.400 874.050 900.600 ;
        RECT 772.950 898.950 775.050 899.400 ;
        RECT 862.950 898.950 865.050 899.400 ;
        RECT 871.950 898.950 874.050 899.400 ;
        RECT 79.950 897.600 82.050 898.050 ;
        RECT 85.950 897.600 88.050 898.050 ;
        RECT 79.950 896.400 88.050 897.600 ;
        RECT 79.950 895.950 82.050 896.400 ;
        RECT 85.950 895.950 88.050 896.400 ;
        RECT 241.950 897.600 244.050 898.050 ;
        RECT 286.950 897.600 289.050 897.900 ;
        RECT 241.950 896.400 289.050 897.600 ;
        RECT 241.950 895.950 244.050 896.400 ;
        RECT 286.950 895.800 289.050 896.400 ;
        RECT 352.950 897.600 355.050 898.050 ;
        RECT 388.950 897.600 391.050 898.050 ;
        RECT 352.950 896.400 391.050 897.600 ;
        RECT 352.950 895.950 355.050 896.400 ;
        RECT 388.950 895.950 391.050 896.400 ;
        RECT 484.950 897.600 487.050 898.050 ;
        RECT 538.950 897.600 541.050 898.050 ;
        RECT 484.950 896.400 541.050 897.600 ;
        RECT 484.950 895.950 487.050 896.400 ;
        RECT 538.950 895.950 541.050 896.400 ;
        RECT 604.950 897.600 607.050 898.050 ;
        RECT 664.950 897.600 667.050 898.050 ;
        RECT 604.950 896.400 667.050 897.600 ;
        RECT 604.950 895.950 607.050 896.400 ;
        RECT 664.950 895.950 667.050 896.400 ;
        RECT 892.950 897.600 895.050 898.050 ;
        RECT 943.950 897.600 946.050 898.050 ;
        RECT 892.950 896.400 946.050 897.600 ;
        RECT 892.950 895.950 895.050 896.400 ;
        RECT 943.950 895.950 946.050 896.400 ;
        RECT 97.950 894.600 100.050 895.050 ;
        RECT 124.950 894.600 127.050 895.050 ;
        RECT 97.950 893.400 127.050 894.600 ;
        RECT 97.950 892.950 100.050 893.400 ;
        RECT 124.950 892.950 127.050 893.400 ;
        RECT 253.950 894.600 256.050 895.050 ;
        RECT 310.950 894.600 313.050 895.050 ;
        RECT 358.950 894.600 361.050 895.050 ;
        RECT 253.950 893.400 361.050 894.600 ;
        RECT 253.950 892.950 256.050 893.400 ;
        RECT 310.950 892.950 313.050 893.400 ;
        RECT 358.950 892.950 361.050 893.400 ;
        RECT 457.950 894.600 460.050 895.050 ;
        RECT 481.950 894.600 484.050 895.050 ;
        RECT 457.950 893.400 484.050 894.600 ;
        RECT 457.950 892.950 460.050 893.400 ;
        RECT 481.950 892.950 484.050 893.400 ;
        RECT 487.950 894.600 490.050 895.050 ;
        RECT 532.950 894.600 535.050 895.050 ;
        RECT 547.950 894.600 550.050 895.050 ;
        RECT 487.950 893.400 550.050 894.600 ;
        RECT 487.950 892.950 490.050 893.400 ;
        RECT 532.950 892.950 535.050 893.400 ;
        RECT 547.950 892.950 550.050 893.400 ;
        RECT 571.950 894.600 574.050 895.050 ;
        RECT 580.950 894.600 583.050 895.050 ;
        RECT 571.950 893.400 583.050 894.600 ;
        RECT 571.950 892.950 574.050 893.400 ;
        RECT 580.950 892.950 583.050 893.400 ;
        RECT 727.950 894.600 730.050 895.050 ;
        RECT 808.950 894.600 811.050 895.050 ;
        RECT 727.950 893.400 811.050 894.600 ;
        RECT 727.950 892.950 730.050 893.400 ;
        RECT 808.950 892.950 811.050 893.400 ;
        RECT 64.950 891.600 67.050 892.050 ;
        RECT 76.950 891.600 79.050 892.050 ;
        RECT 106.950 891.600 109.050 892.050 ;
        RECT 64.950 890.400 109.050 891.600 ;
        RECT 64.950 889.950 67.050 890.400 ;
        RECT 76.950 889.950 79.050 890.400 ;
        RECT 106.950 889.950 109.050 890.400 ;
        RECT 157.950 891.600 160.050 892.050 ;
        RECT 184.950 891.600 187.050 892.050 ;
        RECT 211.950 891.600 214.050 892.050 ;
        RECT 157.950 890.400 214.050 891.600 ;
        RECT 157.950 889.950 160.050 890.400 ;
        RECT 184.950 889.950 187.050 890.400 ;
        RECT 211.950 889.950 214.050 890.400 ;
        RECT 217.950 891.600 220.050 892.050 ;
        RECT 254.400 891.600 255.600 892.950 ;
        RECT 217.950 890.400 255.600 891.600 ;
        RECT 454.950 891.600 457.050 892.050 ;
        RECT 583.950 891.600 586.050 892.050 ;
        RECT 454.950 890.400 586.050 891.600 ;
        RECT 217.950 889.950 220.050 890.400 ;
        RECT 454.950 889.950 457.050 890.400 ;
        RECT 583.950 889.950 586.050 890.400 ;
        RECT 589.950 891.600 592.050 892.050 ;
        RECT 634.950 891.600 637.050 892.050 ;
        RECT 589.950 890.400 637.050 891.600 ;
        RECT 589.950 889.950 592.050 890.400 ;
        RECT 634.950 889.950 637.050 890.400 ;
        RECT 664.950 891.600 667.050 892.050 ;
        RECT 712.950 891.600 715.050 892.050 ;
        RECT 664.950 890.400 715.050 891.600 ;
        RECT 664.950 889.950 667.050 890.400 ;
        RECT 712.950 889.950 715.050 890.400 ;
        RECT 856.950 891.600 859.050 892.050 ;
        RECT 889.950 891.600 892.050 892.050 ;
        RECT 856.950 890.400 912.600 891.600 ;
        RECT 856.950 889.950 859.050 890.400 ;
        RECT 889.950 889.950 892.050 890.400 ;
        RECT 118.950 888.600 121.050 889.050 ;
        RECT 130.950 888.600 133.050 889.050 ;
        RECT 118.950 887.400 133.050 888.600 ;
        RECT 118.950 886.950 121.050 887.400 ;
        RECT 130.950 886.950 133.050 887.400 ;
        RECT 220.950 888.600 223.050 889.050 ;
        RECT 229.950 888.600 234.000 889.050 ;
        RECT 259.950 888.600 262.050 889.050 ;
        RECT 268.950 888.600 271.050 889.050 ;
        RECT 220.950 887.400 234.600 888.600 ;
        RECT 259.950 887.400 271.050 888.600 ;
        RECT 220.950 886.950 223.050 887.400 ;
        RECT 229.950 886.950 234.000 887.400 ;
        RECT 259.950 886.950 262.050 887.400 ;
        RECT 268.950 886.950 271.050 887.400 ;
        RECT 301.950 888.600 304.050 889.050 ;
        RECT 319.950 888.600 322.050 889.050 ;
        RECT 355.950 888.600 358.050 889.050 ;
        RECT 301.950 887.400 358.050 888.600 ;
        RECT 301.950 886.950 304.050 887.400 ;
        RECT 319.950 886.950 322.050 887.400 ;
        RECT 355.950 886.950 358.050 887.400 ;
        RECT 757.950 888.600 760.050 889.050 ;
        RECT 766.950 888.600 769.050 889.050 ;
        RECT 781.950 888.600 784.050 889.050 ;
        RECT 757.950 887.400 784.050 888.600 ;
        RECT 911.400 888.600 912.600 890.400 ;
        RECT 952.950 888.600 955.050 889.050 ;
        RECT 911.400 887.400 955.050 888.600 ;
        RECT 757.950 886.950 760.050 887.400 ;
        RECT 766.950 886.950 769.050 887.400 ;
        RECT 781.950 886.950 784.050 887.400 ;
        RECT 952.950 886.950 955.050 887.400 ;
        RECT 22.950 885.750 25.050 886.200 ;
        RECT 34.950 885.750 37.050 886.200 ;
        RECT 22.950 884.550 37.050 885.750 ;
        RECT 22.950 884.100 25.050 884.550 ;
        RECT 34.950 884.100 37.050 884.550 ;
        RECT 43.950 885.600 46.050 886.200 ;
        RECT 55.950 885.600 58.050 886.050 ;
        RECT 43.950 884.400 58.050 885.600 ;
        RECT 43.950 884.100 46.050 884.400 ;
        RECT 55.950 883.950 58.050 884.400 ;
        RECT 91.950 885.750 94.050 886.200 ;
        RECT 163.950 885.750 166.050 886.200 ;
        RECT 91.950 884.550 166.050 885.750 ;
        RECT 91.950 884.100 94.050 884.550 ;
        RECT 163.950 884.100 166.050 884.550 ;
        RECT 172.950 885.750 175.050 886.200 ;
        RECT 178.950 885.750 181.050 886.200 ;
        RECT 172.950 884.550 181.050 885.750 ;
        RECT 172.950 884.100 175.050 884.550 ;
        RECT 178.950 884.100 181.050 884.550 ;
        RECT 193.950 885.600 196.050 886.050 ;
        RECT 202.950 885.600 205.050 886.200 ;
        RECT 193.950 884.400 205.050 885.600 ;
        RECT 193.950 883.950 196.050 884.400 ;
        RECT 202.950 884.100 205.050 884.400 ;
        RECT 220.950 885.750 223.050 885.900 ;
        RECT 235.950 885.750 238.050 886.200 ;
        RECT 220.950 884.550 238.050 885.750 ;
        RECT 220.950 883.800 223.050 884.550 ;
        RECT 235.950 884.100 238.050 884.550 ;
        RECT 247.950 885.600 250.050 886.050 ;
        RECT 262.950 885.600 265.050 886.200 ;
        RECT 247.950 884.400 265.050 885.600 ;
        RECT 247.950 883.950 250.050 884.400 ;
        RECT 262.950 884.100 265.050 884.400 ;
        RECT 280.950 885.750 283.050 886.200 ;
        RECT 292.950 885.750 295.050 886.200 ;
        RECT 280.950 884.550 295.050 885.750 ;
        RECT 280.950 884.100 283.050 884.550 ;
        RECT 292.950 884.100 295.050 884.550 ;
        RECT 334.950 885.750 337.050 886.200 ;
        RECT 340.950 885.750 343.050 886.200 ;
        RECT 334.950 884.550 343.050 885.750 ;
        RECT 367.950 885.600 370.050 886.200 ;
        RECT 388.950 885.600 391.050 886.200 ;
        RECT 457.950 885.600 460.050 886.200 ;
        RECT 334.950 884.100 337.050 884.550 ;
        RECT 340.950 884.100 343.050 884.550 ;
        RECT 350.400 884.400 391.050 885.600 ;
        RECT 263.400 882.600 264.600 884.100 ;
        RECT 350.400 882.600 351.600 884.400 ;
        RECT 367.950 884.100 370.050 884.400 ;
        RECT 388.950 884.100 391.050 884.400 ;
        RECT 440.400 884.400 460.050 885.600 ;
        RECT 263.400 881.400 351.600 882.600 ;
        RECT 25.950 879.600 28.050 879.900 ;
        RECT 46.950 879.600 49.050 879.900 ;
        RECT 25.950 878.400 49.050 879.600 ;
        RECT 25.950 877.800 28.050 878.400 ;
        RECT 46.950 877.800 49.050 878.400 ;
        RECT 55.950 879.450 58.050 879.900 ;
        RECT 61.950 879.450 64.050 879.900 ;
        RECT 55.950 878.250 64.050 879.450 ;
        RECT 55.950 877.800 58.050 878.250 ;
        RECT 61.950 877.800 64.050 878.250 ;
        RECT 76.950 879.450 79.050 879.900 ;
        RECT 82.950 879.450 85.050 879.900 ;
        RECT 76.950 878.250 85.050 879.450 ;
        RECT 76.950 877.800 79.050 878.250 ;
        RECT 82.950 877.800 85.050 878.250 ;
        RECT 109.950 879.600 112.050 879.900 ;
        RECT 118.950 879.600 121.050 880.050 ;
        RECT 109.950 878.400 121.050 879.600 ;
        RECT 109.950 877.800 112.050 878.400 ;
        RECT 118.950 877.950 121.050 878.400 ;
        RECT 127.950 879.600 130.050 879.900 ;
        RECT 151.950 879.600 154.050 879.900 ;
        RECT 127.950 878.400 154.050 879.600 ;
        RECT 127.950 877.800 130.050 878.400 ;
        RECT 151.950 877.800 154.050 878.400 ;
        RECT 163.950 879.600 166.050 880.050 ;
        RECT 181.950 879.600 184.050 879.900 ;
        RECT 163.950 878.400 184.050 879.600 ;
        RECT 163.950 877.950 166.050 878.400 ;
        RECT 181.950 877.800 184.050 878.400 ;
        RECT 205.950 879.600 208.050 879.900 ;
        RECT 226.950 879.600 229.050 880.050 ;
        RECT 350.400 879.900 351.600 881.400 ;
        RECT 229.950 879.600 232.050 879.900 ;
        RECT 205.950 878.400 232.050 879.600 ;
        RECT 205.950 877.800 208.050 878.400 ;
        RECT 226.950 877.950 229.050 878.400 ;
        RECT 229.950 877.800 232.050 878.400 ;
        RECT 295.950 879.600 298.050 879.900 ;
        RECT 316.950 879.600 319.050 879.900 ;
        RECT 295.950 878.400 319.050 879.600 ;
        RECT 295.950 877.800 298.050 878.400 ;
        RECT 316.950 877.800 319.050 878.400 ;
        RECT 325.950 879.450 328.050 879.900 ;
        RECT 343.950 879.450 346.050 879.900 ;
        RECT 325.950 878.250 346.050 879.450 ;
        RECT 325.950 877.800 328.050 878.250 ;
        RECT 343.950 877.800 346.050 878.250 ;
        RECT 349.950 877.800 352.050 879.900 ;
        RECT 355.950 879.600 358.050 880.050 ;
        RECT 364.950 879.600 367.050 879.900 ;
        RECT 355.950 878.400 367.050 879.600 ;
        RECT 355.950 877.950 358.050 878.400 ;
        RECT 364.950 877.800 367.050 878.400 ;
        RECT 418.950 879.450 421.050 879.900 ;
        RECT 430.950 879.450 433.050 879.900 ;
        RECT 418.950 878.250 433.050 879.450 ;
        RECT 418.950 877.800 421.050 878.250 ;
        RECT 430.950 877.800 433.050 878.250 ;
        RECT 436.950 879.600 439.050 879.900 ;
        RECT 440.400 879.600 441.600 884.400 ;
        RECT 457.950 884.100 460.050 884.400 ;
        RECT 463.950 885.600 466.050 886.050 ;
        RECT 478.950 885.600 481.050 886.050 ;
        RECT 463.950 884.400 481.050 885.600 ;
        RECT 463.950 883.950 466.050 884.400 ;
        RECT 478.950 883.950 481.050 884.400 ;
        RECT 487.950 884.100 490.050 886.200 ;
        RECT 577.950 885.600 580.050 886.200 ;
        RECT 592.950 885.600 595.050 886.200 ;
        RECT 577.950 884.400 595.050 885.600 ;
        RECT 577.950 884.100 580.050 884.400 ;
        RECT 592.950 884.100 595.050 884.400 ;
        RECT 607.950 885.750 610.050 886.200 ;
        RECT 619.950 885.750 622.050 886.200 ;
        RECT 607.950 884.550 622.050 885.750 ;
        RECT 607.950 884.100 610.050 884.550 ;
        RECT 619.950 884.100 622.050 884.550 ;
        RECT 625.950 885.600 628.050 886.200 ;
        RECT 646.950 885.600 649.050 886.200 ;
        RECT 625.950 884.400 649.050 885.600 ;
        RECT 625.950 884.100 628.050 884.400 ;
        RECT 646.950 884.100 649.050 884.400 ;
        RECT 700.950 885.750 703.050 886.200 ;
        RECT 718.950 885.750 721.050 886.200 ;
        RECT 700.950 885.600 721.050 885.750 ;
        RECT 733.950 885.600 736.050 886.200 ;
        RECT 700.950 884.550 736.050 885.600 ;
        RECT 700.950 884.100 703.050 884.550 ;
        RECT 718.950 884.400 736.050 884.550 ;
        RECT 718.950 884.100 721.050 884.400 ;
        RECT 733.950 884.100 736.050 884.400 ;
        RECT 787.950 885.600 790.050 886.200 ;
        RECT 796.950 885.600 799.050 886.050 ;
        RECT 787.950 884.400 799.050 885.600 ;
        RECT 787.950 884.100 790.050 884.400 ;
        RECT 488.400 882.600 489.600 884.100 ;
        RECT 578.400 882.600 579.600 884.100 ;
        RECT 796.950 883.950 799.050 884.400 ;
        RECT 805.950 884.100 808.050 886.200 ;
        RECT 811.950 885.600 814.050 886.200 ;
        RECT 823.950 885.600 826.050 886.050 ;
        RECT 832.950 885.600 835.050 886.200 ;
        RECT 811.950 884.400 835.050 885.600 ;
        RECT 811.950 884.100 814.050 884.400 ;
        RECT 479.400 881.400 489.600 882.600 ;
        RECT 572.400 881.400 579.600 882.600 ;
        RECT 436.950 878.400 441.600 879.600 ;
        RECT 448.950 879.450 451.050 879.900 ;
        RECT 466.950 879.600 469.050 879.900 ;
        RECT 479.400 879.600 480.600 881.400 ;
        RECT 466.950 879.450 480.600 879.600 ;
        RECT 448.950 878.400 480.600 879.450 ;
        RECT 481.950 879.450 484.050 879.900 ;
        RECT 493.950 879.450 496.050 879.900 ;
        RECT 436.950 877.800 439.050 878.400 ;
        RECT 448.950 878.250 469.050 878.400 ;
        RECT 448.950 877.800 451.050 878.250 ;
        RECT 466.950 877.800 469.050 878.250 ;
        RECT 481.950 878.250 496.050 879.450 ;
        RECT 481.950 877.800 484.050 878.250 ;
        RECT 493.950 877.800 496.050 878.250 ;
        RECT 550.950 879.600 553.050 879.900 ;
        RECT 562.950 879.600 565.050 879.900 ;
        RECT 550.950 879.450 565.050 879.600 ;
        RECT 568.950 879.450 571.050 879.900 ;
        RECT 550.950 878.400 571.050 879.450 ;
        RECT 550.950 877.800 553.050 878.400 ;
        RECT 562.950 878.250 571.050 878.400 ;
        RECT 562.950 877.800 565.050 878.250 ;
        RECT 568.950 877.800 571.050 878.250 ;
        RECT 124.950 876.600 127.050 877.050 ;
        RECT 133.950 876.600 136.050 877.050 ;
        RECT 142.950 876.600 145.050 877.050 ;
        RECT 193.950 876.600 196.050 877.050 ;
        RECT 124.950 875.400 196.050 876.600 ;
        RECT 124.950 874.950 127.050 875.400 ;
        RECT 133.950 874.950 136.050 875.400 ;
        RECT 142.950 874.950 145.050 875.400 ;
        RECT 193.950 874.950 196.050 875.400 ;
        RECT 502.950 876.600 505.050 877.050 ;
        RECT 572.400 876.600 573.600 881.400 ;
        RECT 574.950 879.450 577.050 879.900 ;
        RECT 583.950 879.600 586.050 879.900 ;
        RECT 595.950 879.600 598.050 879.900 ;
        RECT 583.950 879.450 598.050 879.600 ;
        RECT 574.950 878.400 598.050 879.450 ;
        RECT 574.950 878.250 586.050 878.400 ;
        RECT 574.950 877.800 577.050 878.250 ;
        RECT 583.950 877.800 586.050 878.250 ;
        RECT 595.950 877.800 598.050 878.400 ;
        RECT 610.950 879.450 613.050 879.900 ;
        RECT 616.950 879.450 619.050 879.900 ;
        RECT 610.950 878.250 619.050 879.450 ;
        RECT 610.950 877.800 613.050 878.250 ;
        RECT 616.950 877.800 619.050 878.250 ;
        RECT 649.950 879.600 652.050 879.900 ;
        RECT 667.950 879.600 670.050 879.900 ;
        RECT 754.950 879.600 757.050 879.900 ;
        RECT 784.950 879.600 787.050 879.900 ;
        RECT 649.950 878.400 670.050 879.600 ;
        RECT 649.950 877.800 652.050 878.400 ;
        RECT 667.950 877.800 670.050 878.400 ;
        RECT 752.400 878.400 787.050 879.600 ;
        RECT 806.400 879.600 807.600 884.100 ;
        RECT 823.950 883.950 826.050 884.400 ;
        RECT 832.950 884.100 835.050 884.400 ;
        RECT 862.950 884.100 865.050 886.200 ;
        RECT 871.950 885.750 874.050 886.200 ;
        RECT 877.950 885.750 880.050 886.200 ;
        RECT 871.950 884.550 880.050 885.750 ;
        RECT 871.950 884.100 874.050 884.550 ;
        RECT 877.950 884.100 880.050 884.550 ;
        RECT 883.950 884.100 886.050 886.200 ;
        RECT 910.950 885.750 913.050 886.200 ;
        RECT 928.950 885.750 931.050 886.200 ;
        RECT 910.950 884.550 931.050 885.750 ;
        RECT 933.000 885.600 937.050 886.050 ;
        RECT 910.950 884.100 913.050 884.550 ;
        RECT 928.950 884.100 931.050 884.550 ;
        RECT 863.400 880.050 864.600 884.100 ;
        RECT 884.400 882.600 885.600 884.100 ;
        RECT 932.400 883.950 937.050 885.600 ;
        RECT 940.950 885.600 943.050 886.050 ;
        RECT 946.950 885.600 949.050 886.200 ;
        RECT 957.000 885.600 961.050 886.050 ;
        RECT 940.950 884.400 949.050 885.600 ;
        RECT 940.950 883.950 943.050 884.400 ;
        RECT 946.950 884.100 949.050 884.400 ;
        RECT 956.400 883.950 961.050 885.600 ;
        RECT 967.950 883.950 970.050 886.050 ;
        RECT 973.950 885.600 976.050 886.200 ;
        RECT 997.950 885.600 1000.050 886.200 ;
        RECT 973.950 884.400 1000.050 885.600 ;
        RECT 973.950 884.100 976.050 884.400 ;
        RECT 997.950 884.100 1000.050 884.400 ;
        RECT 1006.950 883.950 1009.050 886.050 ;
        RECT 1014.000 885.600 1018.050 886.050 ;
        RECT 1013.400 883.950 1018.050 885.600 ;
        RECT 884.400 881.400 894.600 882.600 ;
        RECT 814.950 879.600 817.050 880.050 ;
        RECT 806.400 878.400 817.050 879.600 ;
        RECT 863.400 878.400 867.900 880.050 ;
        RECT 502.950 875.400 573.600 876.600 ;
        RECT 622.950 876.600 625.050 877.050 ;
        RECT 637.950 876.600 640.050 877.050 ;
        RECT 622.950 875.400 640.050 876.600 ;
        RECT 502.950 874.950 505.050 875.400 ;
        RECT 622.950 874.950 625.050 875.400 ;
        RECT 637.950 874.950 640.050 875.400 ;
        RECT 679.950 876.600 682.050 877.050 ;
        RECT 709.950 876.600 712.050 877.050 ;
        RECT 679.950 875.400 712.050 876.600 ;
        RECT 679.950 874.950 682.050 875.400 ;
        RECT 709.950 874.950 712.050 875.400 ;
        RECT 736.950 876.600 739.050 877.050 ;
        RECT 752.400 876.600 753.600 878.400 ;
        RECT 754.950 877.800 757.050 878.400 ;
        RECT 784.950 877.800 787.050 878.400 ;
        RECT 814.950 877.950 817.050 878.400 ;
        RECT 864.000 877.950 867.900 878.400 ;
        RECT 868.950 879.600 871.050 880.050 ;
        RECT 880.950 879.600 883.050 879.900 ;
        RECT 868.950 878.400 883.050 879.600 ;
        RECT 893.400 879.600 894.600 881.400 ;
        RECT 932.400 879.900 933.600 883.950 ;
        RECT 956.400 879.900 957.600 883.950 ;
        RECT 968.400 880.050 969.600 883.950 ;
        RECT 904.950 879.600 907.050 879.900 ;
        RECT 893.400 878.400 907.050 879.600 ;
        RECT 868.950 877.950 871.050 878.400 ;
        RECT 736.950 875.400 753.600 876.600 ;
        RECT 847.950 876.600 850.050 877.050 ;
        RECT 853.950 876.600 856.050 877.050 ;
        RECT 847.950 875.400 856.050 876.600 ;
        RECT 736.950 874.950 739.050 875.400 ;
        RECT 847.950 874.950 850.050 875.400 ;
        RECT 853.950 874.950 856.050 875.400 ;
        RECT 859.950 876.600 862.050 877.050 ;
        RECT 869.400 876.600 870.600 877.950 ;
        RECT 880.950 877.800 883.050 878.400 ;
        RECT 904.950 877.800 907.050 878.400 ;
        RECT 931.950 877.800 934.050 879.900 ;
        RECT 943.950 879.450 946.050 879.900 ;
        RECT 949.950 879.450 952.050 879.900 ;
        RECT 943.950 878.250 952.050 879.450 ;
        RECT 943.950 877.800 946.050 878.250 ;
        RECT 949.950 877.800 952.050 878.250 ;
        RECT 955.950 877.800 958.050 879.900 ;
        RECT 967.950 877.950 970.050 880.050 ;
        RECT 982.950 879.600 985.050 880.050 ;
        RECT 1007.400 879.600 1008.600 883.950 ;
        RECT 982.950 878.400 1008.600 879.600 ;
        RECT 982.950 877.950 985.050 878.400 ;
        RECT 1013.400 877.050 1014.600 883.950 ;
        RECT 859.950 875.400 870.600 876.600 ;
        RECT 1009.950 875.400 1014.600 877.050 ;
        RECT 859.950 874.950 862.050 875.400 ;
        RECT 1009.950 874.950 1014.000 875.400 ;
        RECT 16.950 873.600 19.050 874.050 ;
        RECT 67.950 873.600 70.050 874.050 ;
        RECT 16.950 872.400 70.050 873.600 ;
        RECT 16.950 871.950 19.050 872.400 ;
        RECT 67.950 871.950 70.050 872.400 ;
        RECT 88.950 873.600 91.050 874.050 ;
        RECT 115.950 873.600 118.050 874.050 ;
        RECT 88.950 872.400 118.050 873.600 ;
        RECT 88.950 871.950 91.050 872.400 ;
        RECT 115.950 871.950 118.050 872.400 ;
        RECT 271.950 873.600 274.050 874.050 ;
        RECT 295.950 873.600 298.050 874.050 ;
        RECT 271.950 872.400 298.050 873.600 ;
        RECT 271.950 871.950 274.050 872.400 ;
        RECT 295.950 871.950 298.050 872.400 ;
        RECT 385.950 873.600 388.050 874.050 ;
        RECT 442.950 873.600 445.050 874.050 ;
        RECT 385.950 872.400 445.050 873.600 ;
        RECT 385.950 871.950 388.050 872.400 ;
        RECT 442.950 871.950 445.050 872.400 ;
        RECT 460.950 873.600 463.050 874.050 ;
        RECT 472.950 873.600 475.050 874.050 ;
        RECT 460.950 872.400 475.050 873.600 ;
        RECT 460.950 871.950 463.050 872.400 ;
        RECT 472.950 871.950 475.050 872.400 ;
        RECT 532.950 873.600 535.050 874.050 ;
        RECT 607.950 873.600 610.050 874.050 ;
        RECT 532.950 872.400 610.050 873.600 ;
        RECT 532.950 871.950 535.050 872.400 ;
        RECT 607.950 871.950 610.050 872.400 ;
        RECT 634.950 873.600 637.050 874.050 ;
        RECT 643.950 873.600 646.050 874.050 ;
        RECT 634.950 872.400 646.050 873.600 ;
        RECT 634.950 871.950 637.050 872.400 ;
        RECT 643.950 871.950 646.050 872.400 ;
        RECT 919.950 873.600 922.050 874.050 ;
        RECT 937.950 873.600 940.050 874.050 ;
        RECT 919.950 872.400 940.050 873.600 ;
        RECT 919.950 871.950 922.050 872.400 ;
        RECT 937.950 871.950 940.050 872.400 ;
        RECT 160.950 870.600 163.050 871.050 ;
        RECT 172.950 870.600 175.050 871.050 ;
        RECT 199.950 870.600 202.050 871.050 ;
        RECT 160.950 869.400 202.050 870.600 ;
        RECT 160.950 868.950 163.050 869.400 ;
        RECT 172.950 868.950 175.050 869.400 ;
        RECT 199.950 868.950 202.050 869.400 ;
        RECT 220.950 870.600 223.050 871.050 ;
        RECT 325.950 870.600 328.050 871.050 ;
        RECT 220.950 869.400 328.050 870.600 ;
        RECT 220.950 868.950 223.050 869.400 ;
        RECT 325.950 868.950 328.050 869.400 ;
        RECT 589.950 870.600 592.050 871.050 ;
        RECT 655.950 870.600 658.050 871.050 ;
        RECT 589.950 869.400 658.050 870.600 ;
        RECT 589.950 868.950 592.050 869.400 ;
        RECT 655.950 868.950 658.050 869.400 ;
        RECT 709.950 870.600 712.050 871.050 ;
        RECT 760.950 870.600 763.050 871.050 ;
        RECT 778.950 870.600 781.050 871.050 ;
        RECT 709.950 869.400 781.050 870.600 ;
        RECT 709.950 868.950 712.050 869.400 ;
        RECT 760.950 868.950 763.050 869.400 ;
        RECT 778.950 868.950 781.050 869.400 ;
        RECT 964.950 870.600 967.050 871.050 ;
        RECT 976.950 870.600 979.050 871.050 ;
        RECT 994.950 870.600 997.050 871.050 ;
        RECT 964.950 869.400 997.050 870.600 ;
        RECT 964.950 868.950 967.050 869.400 ;
        RECT 976.950 868.950 979.050 869.400 ;
        RECT 994.950 868.950 997.050 869.400 ;
        RECT 265.950 867.600 268.050 868.050 ;
        RECT 280.950 867.600 283.050 868.050 ;
        RECT 322.950 867.600 325.050 868.050 ;
        RECT 265.950 866.400 325.050 867.600 ;
        RECT 265.950 865.950 268.050 866.400 ;
        RECT 280.950 865.950 283.050 866.400 ;
        RECT 322.950 865.950 325.050 866.400 ;
        RECT 337.950 867.600 340.050 868.050 ;
        RECT 469.950 867.600 472.050 868.050 ;
        RECT 337.950 866.400 472.050 867.600 ;
        RECT 337.950 865.950 340.050 866.400 ;
        RECT 469.950 865.950 472.050 866.400 ;
        RECT 514.950 867.600 517.050 868.050 ;
        RECT 541.950 867.600 544.050 868.050 ;
        RECT 514.950 866.400 544.050 867.600 ;
        RECT 514.950 865.950 517.050 866.400 ;
        RECT 541.950 865.950 544.050 866.400 ;
        RECT 769.950 867.600 772.050 868.050 ;
        RECT 802.950 867.600 805.050 868.050 ;
        RECT 841.950 867.600 844.050 868.050 ;
        RECT 769.950 866.400 844.050 867.600 ;
        RECT 769.950 865.950 772.050 866.400 ;
        RECT 802.950 865.950 805.050 866.400 ;
        RECT 841.950 865.950 844.050 866.400 ;
        RECT 889.950 867.600 892.050 868.050 ;
        RECT 970.950 867.600 973.050 868.050 ;
        RECT 1000.950 867.600 1003.050 868.050 ;
        RECT 889.950 866.400 1003.050 867.600 ;
        RECT 889.950 865.950 892.050 866.400 ;
        RECT 970.950 865.950 973.050 866.400 ;
        RECT 1000.950 865.950 1003.050 866.400 ;
        RECT 301.950 864.600 304.050 865.050 ;
        RECT 307.950 864.600 310.050 865.050 ;
        RECT 301.950 863.400 310.050 864.600 ;
        RECT 301.950 862.950 304.050 863.400 ;
        RECT 307.950 862.950 310.050 863.400 ;
        RECT 412.950 864.600 415.050 865.050 ;
        RECT 682.950 864.600 685.050 865.050 ;
        RECT 412.950 863.400 685.050 864.600 ;
        RECT 412.950 862.950 415.050 863.400 ;
        RECT 682.950 862.950 685.050 863.400 ;
        RECT 880.950 864.600 883.050 865.050 ;
        RECT 892.950 864.600 895.050 865.050 ;
        RECT 880.950 863.400 895.050 864.600 ;
        RECT 880.950 862.950 883.050 863.400 ;
        RECT 892.950 862.950 895.050 863.400 ;
        RECT 970.950 864.600 973.050 864.900 ;
        RECT 982.800 864.600 984.900 865.050 ;
        RECT 970.950 863.400 984.900 864.600 ;
        RECT 970.950 862.800 973.050 863.400 ;
        RECT 982.800 862.950 984.900 863.400 ;
        RECT 985.950 864.600 988.050 865.050 ;
        RECT 997.950 864.600 1000.050 865.050 ;
        RECT 985.950 863.400 1000.050 864.600 ;
        RECT 985.950 862.950 988.050 863.400 ;
        RECT 997.950 862.950 1000.050 863.400 ;
        RECT 256.950 861.600 259.050 862.050 ;
        RECT 268.950 861.600 271.050 862.050 ;
        RECT 334.950 861.600 337.050 862.050 ;
        RECT 256.950 860.400 337.050 861.600 ;
        RECT 256.950 859.950 259.050 860.400 ;
        RECT 268.950 859.950 271.050 860.400 ;
        RECT 334.950 859.950 337.050 860.400 ;
        RECT 358.950 861.600 361.050 862.050 ;
        RECT 370.950 861.600 373.050 862.050 ;
        RECT 412.950 861.600 415.050 861.900 ;
        RECT 358.950 860.400 415.050 861.600 ;
        RECT 358.950 859.950 361.050 860.400 ;
        RECT 370.950 859.950 373.050 860.400 ;
        RECT 412.950 859.800 415.050 860.400 ;
        RECT 52.950 858.600 55.050 859.050 ;
        RECT 229.950 858.600 232.050 859.050 ;
        RECT 301.950 858.600 304.050 859.050 ;
        RECT 52.950 857.400 304.050 858.600 ;
        RECT 52.950 856.950 55.050 857.400 ;
        RECT 229.950 856.950 232.050 857.400 ;
        RECT 301.950 856.950 304.050 857.400 ;
        RECT 307.950 858.600 310.050 859.050 ;
        RECT 337.950 858.600 340.050 859.050 ;
        RECT 307.950 857.400 340.050 858.600 ;
        RECT 307.950 856.950 310.050 857.400 ;
        RECT 337.950 856.950 340.050 857.400 ;
        RECT 451.950 858.600 454.050 859.050 ;
        RECT 505.950 858.600 508.050 859.050 ;
        RECT 451.950 857.400 508.050 858.600 ;
        RECT 451.950 856.950 454.050 857.400 ;
        RECT 505.950 856.950 508.050 857.400 ;
        RECT 514.950 858.600 517.050 859.050 ;
        RECT 604.950 858.600 607.050 859.050 ;
        RECT 514.950 857.400 607.050 858.600 ;
        RECT 514.950 856.950 517.050 857.400 ;
        RECT 604.950 856.950 607.050 857.400 ;
        RECT 622.950 858.600 625.050 859.050 ;
        RECT 685.950 858.600 688.050 859.050 ;
        RECT 691.950 858.600 694.050 859.050 ;
        RECT 622.950 857.400 694.050 858.600 ;
        RECT 622.950 856.950 625.050 857.400 ;
        RECT 685.950 856.950 688.050 857.400 ;
        RECT 691.950 856.950 694.050 857.400 ;
        RECT 817.950 858.600 820.050 859.050 ;
        RECT 988.950 858.600 991.050 859.050 ;
        RECT 817.950 857.400 991.050 858.600 ;
        RECT 817.950 856.950 820.050 857.400 ;
        RECT 988.950 856.950 991.050 857.400 ;
        RECT 40.950 855.600 43.050 856.050 ;
        RECT 46.950 855.600 49.050 856.050 ;
        RECT 406.950 855.600 409.050 856.050 ;
        RECT 40.950 854.400 49.050 855.600 ;
        RECT 40.950 853.950 43.050 854.400 ;
        RECT 46.950 853.950 49.050 854.400 ;
        RECT 305.400 854.400 409.050 855.600 ;
        RECT 305.400 853.050 306.600 854.400 ;
        RECT 406.950 853.950 409.050 854.400 ;
        RECT 508.950 855.600 511.050 856.050 ;
        RECT 580.950 855.600 583.050 856.050 ;
        RECT 508.950 854.400 583.050 855.600 ;
        RECT 508.950 853.950 511.050 854.400 ;
        RECT 580.950 853.950 583.050 854.400 ;
        RECT 709.950 855.600 712.050 856.050 ;
        RECT 721.950 855.600 724.050 856.050 ;
        RECT 772.950 855.600 775.050 856.050 ;
        RECT 709.950 854.400 775.050 855.600 ;
        RECT 709.950 853.950 712.050 854.400 ;
        RECT 721.950 853.950 724.050 854.400 ;
        RECT 772.950 853.950 775.050 854.400 ;
        RECT 853.950 855.600 856.050 856.050 ;
        RECT 919.950 855.600 922.050 856.050 ;
        RECT 853.950 854.400 922.050 855.600 ;
        RECT 853.950 853.950 856.050 854.400 ;
        RECT 919.950 853.950 922.050 854.400 ;
        RECT 169.950 852.600 172.050 853.050 ;
        RECT 184.950 852.600 187.050 853.050 ;
        RECT 169.950 851.400 187.050 852.600 ;
        RECT 169.950 850.950 172.050 851.400 ;
        RECT 184.950 850.950 187.050 851.400 ;
        RECT 244.950 852.600 247.050 853.050 ;
        RECT 283.800 852.600 285.900 853.050 ;
        RECT 244.950 851.400 285.900 852.600 ;
        RECT 244.950 850.950 247.050 851.400 ;
        RECT 283.800 850.950 285.900 851.400 ;
        RECT 286.950 852.600 289.050 853.050 ;
        RECT 304.800 852.600 306.900 853.050 ;
        RECT 286.950 851.400 306.900 852.600 ;
        RECT 286.950 850.950 289.050 851.400 ;
        RECT 304.800 850.950 306.900 851.400 ;
        RECT 307.950 852.600 310.050 853.050 ;
        RECT 355.950 852.600 358.050 853.050 ;
        RECT 307.950 851.400 358.050 852.600 ;
        RECT 307.950 850.950 310.050 851.400 ;
        RECT 355.950 850.950 358.050 851.400 ;
        RECT 418.950 852.600 421.050 853.050 ;
        RECT 442.950 852.600 445.050 853.050 ;
        RECT 472.950 852.600 475.050 853.050 ;
        RECT 418.950 851.400 475.050 852.600 ;
        RECT 418.950 850.950 421.050 851.400 ;
        RECT 442.950 850.950 445.050 851.400 ;
        RECT 472.950 850.950 475.050 851.400 ;
        RECT 715.950 852.600 718.050 853.050 ;
        RECT 742.950 852.600 745.050 853.050 ;
        RECT 715.950 851.400 745.050 852.600 ;
        RECT 715.950 850.950 718.050 851.400 ;
        RECT 742.950 850.950 745.050 851.400 ;
        RECT 994.950 852.600 997.050 853.050 ;
        RECT 1003.950 852.600 1006.050 853.050 ;
        RECT 994.950 851.400 1006.050 852.600 ;
        RECT 994.950 850.950 997.050 851.400 ;
        RECT 1003.950 850.950 1006.050 851.400 ;
        RECT 61.950 849.600 64.050 850.050 ;
        RECT 67.950 849.600 70.050 850.050 ;
        RECT 91.950 849.600 94.050 850.050 ;
        RECT 61.950 848.400 94.050 849.600 ;
        RECT 61.950 847.950 64.050 848.400 ;
        RECT 67.950 847.950 70.050 848.400 ;
        RECT 91.950 847.950 94.050 848.400 ;
        RECT 187.950 849.600 190.050 850.050 ;
        RECT 403.950 849.600 406.050 850.050 ;
        RECT 484.950 849.600 487.050 850.050 ;
        RECT 499.950 849.600 502.050 850.050 ;
        RECT 187.950 848.400 406.050 849.600 ;
        RECT 187.950 847.950 190.050 848.400 ;
        RECT 403.950 847.950 406.050 848.400 ;
        RECT 434.400 848.400 502.050 849.600 ;
        RECT 211.950 846.600 214.050 847.050 ;
        RECT 220.950 846.600 223.050 847.050 ;
        RECT 364.950 846.600 367.050 847.050 ;
        RECT 211.950 845.400 367.050 846.600 ;
        RECT 211.950 844.950 214.050 845.400 ;
        RECT 220.950 844.950 223.050 845.400 ;
        RECT 364.950 844.950 367.050 845.400 ;
        RECT 382.950 846.600 385.050 847.050 ;
        RECT 434.400 846.600 435.600 848.400 ;
        RECT 484.950 847.950 487.050 848.400 ;
        RECT 499.950 847.950 502.050 848.400 ;
        RECT 535.950 849.600 538.050 850.050 ;
        RECT 559.950 849.600 562.050 850.050 ;
        RECT 535.950 848.400 562.050 849.600 ;
        RECT 535.950 847.950 538.050 848.400 ;
        RECT 559.950 847.950 562.050 848.400 ;
        RECT 640.950 849.600 643.050 850.050 ;
        RECT 694.950 849.600 697.050 850.050 ;
        RECT 640.950 848.400 697.050 849.600 ;
        RECT 640.950 847.950 643.050 848.400 ;
        RECT 694.950 847.950 697.050 848.400 ;
        RECT 775.950 849.600 778.050 850.050 ;
        RECT 814.950 849.600 817.050 850.050 ;
        RECT 847.950 849.600 850.050 850.050 ;
        RECT 775.950 848.400 850.050 849.600 ;
        RECT 775.950 847.950 778.050 848.400 ;
        RECT 814.950 847.950 817.050 848.400 ;
        RECT 847.950 847.950 850.050 848.400 ;
        RECT 955.950 849.600 958.050 850.050 ;
        RECT 973.950 849.600 976.050 850.050 ;
        RECT 955.950 848.400 976.050 849.600 ;
        RECT 955.950 847.950 958.050 848.400 ;
        RECT 973.950 847.950 976.050 848.400 ;
        RECT 382.950 845.400 435.600 846.600 ;
        RECT 523.950 846.600 526.050 847.050 ;
        RECT 550.950 846.600 553.050 847.050 ;
        RECT 523.950 845.400 553.050 846.600 ;
        RECT 382.950 844.950 385.050 845.400 ;
        RECT 523.950 844.950 526.050 845.400 ;
        RECT 550.950 844.950 553.050 845.400 ;
        RECT 568.950 846.600 571.050 846.900 ;
        RECT 586.950 846.600 589.050 847.050 ;
        RECT 568.950 845.400 589.050 846.600 ;
        RECT 568.950 844.800 571.050 845.400 ;
        RECT 586.950 844.950 589.050 845.400 ;
        RECT 682.950 846.600 685.050 847.050 ;
        RECT 700.950 846.600 703.050 847.050 ;
        RECT 760.950 846.600 763.050 847.050 ;
        RECT 766.950 846.600 769.050 847.050 ;
        RECT 682.950 845.400 693.600 846.600 ;
        RECT 682.950 844.950 685.050 845.400 ;
        RECT 33.000 843.600 37.050 844.050 ;
        RECT 32.400 841.950 37.050 843.600 ;
        RECT 67.950 843.600 70.050 844.050 ;
        RECT 97.950 843.600 100.050 844.050 ;
        RECT 67.950 842.400 100.050 843.600 ;
        RECT 67.950 841.950 70.050 842.400 ;
        RECT 97.950 841.950 100.050 842.400 ;
        RECT 283.950 843.600 286.050 844.050 ;
        RECT 307.950 843.600 310.050 844.050 ;
        RECT 283.950 842.400 310.050 843.600 ;
        RECT 283.950 841.950 286.050 842.400 ;
        RECT 307.950 841.950 310.050 842.400 ;
        RECT 478.950 843.600 481.050 844.050 ;
        RECT 496.950 843.600 499.050 844.050 ;
        RECT 478.950 842.400 499.050 843.600 ;
        RECT 478.950 841.950 481.050 842.400 ;
        RECT 496.950 841.950 499.050 842.400 ;
        RECT 505.950 843.600 508.050 844.050 ;
        RECT 622.950 843.600 625.050 844.050 ;
        RECT 505.950 842.400 625.050 843.600 ;
        RECT 505.950 841.950 508.050 842.400 ;
        RECT 622.950 841.950 625.050 842.400 ;
        RECT 32.400 837.600 33.600 841.950 ;
        RECT 46.950 840.600 49.050 841.200 ;
        RECT 29.400 836.400 33.600 837.600 ;
        RECT 35.400 839.400 49.050 840.600 ;
        RECT 7.950 834.450 10.050 834.900 ;
        RECT 16.950 834.450 19.050 834.900 ;
        RECT 7.950 833.250 19.050 834.450 ;
        RECT 7.950 832.800 10.050 833.250 ;
        RECT 16.950 832.800 19.050 833.250 ;
        RECT 29.400 831.600 30.600 836.400 ;
        RECT 35.400 832.050 36.600 839.400 ;
        RECT 46.950 839.100 49.050 839.400 ;
        RECT 73.950 840.750 76.050 841.200 ;
        RECT 82.950 840.750 85.050 841.200 ;
        RECT 73.950 839.550 85.050 840.750 ;
        RECT 73.950 839.100 76.050 839.550 ;
        RECT 82.950 839.100 85.050 839.550 ;
        RECT 109.950 840.600 112.050 841.050 ;
        RECT 115.950 840.600 118.050 841.200 ;
        RECT 109.950 839.400 118.050 840.600 ;
        RECT 109.950 838.950 112.050 839.400 ;
        RECT 115.950 839.100 118.050 839.400 ;
        RECT 136.950 840.600 139.050 841.200 ;
        RECT 160.950 840.600 163.050 841.200 ;
        RECT 136.950 839.400 163.050 840.600 ;
        RECT 136.950 839.100 139.050 839.400 ;
        RECT 160.950 839.100 163.050 839.400 ;
        RECT 178.950 839.100 181.050 841.200 ;
        RECT 232.950 840.750 235.050 841.200 ;
        RECT 238.950 840.750 241.050 841.200 ;
        RECT 232.950 839.550 241.050 840.750 ;
        RECT 232.950 839.100 235.050 839.550 ;
        RECT 238.950 839.100 241.050 839.550 ;
        RECT 280.950 839.100 283.050 841.200 ;
        RECT 349.950 840.750 352.050 841.200 ;
        RECT 358.950 840.750 361.050 841.200 ;
        RECT 349.950 839.550 361.050 840.750 ;
        RECT 349.950 839.100 352.050 839.550 ;
        RECT 358.950 839.100 361.050 839.550 ;
        RECT 391.950 839.100 394.050 841.200 ;
        RECT 397.950 840.600 400.050 841.200 ;
        RECT 421.950 840.600 424.050 841.200 ;
        RECT 397.950 839.400 424.050 840.600 ;
        RECT 397.950 839.100 400.050 839.400 ;
        RECT 421.950 839.100 424.050 839.400 ;
        RECT 469.950 840.750 472.050 841.200 ;
        RECT 478.950 840.750 481.050 841.200 ;
        RECT 469.950 839.550 481.050 840.750 ;
        RECT 469.950 839.100 472.050 839.550 ;
        RECT 478.950 839.100 481.050 839.550 ;
        RECT 490.950 840.600 493.050 841.050 ;
        RECT 517.950 840.750 520.050 841.200 ;
        RECT 523.950 840.750 526.050 841.200 ;
        RECT 490.950 839.400 513.600 840.600 ;
        RECT 179.400 837.600 180.600 839.100 ;
        RECT 176.400 836.400 180.600 837.600 ;
        RECT 281.400 837.600 282.600 839.100 ;
        RECT 298.950 837.600 301.050 838.050 ;
        RECT 281.400 836.400 301.050 837.600 ;
        RECT 392.400 837.600 393.600 839.100 ;
        RECT 490.950 838.950 493.050 839.400 ;
        RECT 406.950 837.600 409.050 838.050 ;
        RECT 392.400 836.400 409.050 837.600 ;
        RECT 512.400 837.600 513.600 839.400 ;
        RECT 517.950 839.550 526.050 840.750 ;
        RECT 517.950 839.100 520.050 839.550 ;
        RECT 523.950 839.100 526.050 839.550 ;
        RECT 529.950 840.750 532.050 841.200 ;
        RECT 538.950 840.750 541.050 841.200 ;
        RECT 529.950 839.550 541.050 840.750 ;
        RECT 529.950 839.100 532.050 839.550 ;
        RECT 538.950 839.100 541.050 839.550 ;
        RECT 556.950 840.600 559.050 841.200 ;
        RECT 565.950 840.750 568.050 841.200 ;
        RECT 574.950 840.750 577.050 841.200 ;
        RECT 565.950 840.600 577.050 840.750 ;
        RECT 556.950 839.550 577.050 840.600 ;
        RECT 556.950 839.400 568.050 839.550 ;
        RECT 556.950 839.100 559.050 839.400 ;
        RECT 565.950 839.100 568.050 839.400 ;
        RECT 574.950 839.100 577.050 839.550 ;
        RECT 592.950 840.750 595.050 841.200 ;
        RECT 598.950 840.750 601.050 841.200 ;
        RECT 592.950 839.550 601.050 840.750 ;
        RECT 592.950 839.100 595.050 839.550 ;
        RECT 598.950 839.100 601.050 839.550 ;
        RECT 649.950 840.600 652.050 841.200 ;
        RECT 664.950 840.600 667.050 841.200 ;
        RECT 649.950 839.400 667.050 840.600 ;
        RECT 649.950 839.100 652.050 839.400 ;
        RECT 664.950 839.100 667.050 839.400 ;
        RECT 670.950 839.100 673.050 841.200 ;
        RECT 676.950 840.750 679.050 841.200 ;
        RECT 688.950 840.750 691.050 841.200 ;
        RECT 676.950 839.550 691.050 840.750 ;
        RECT 676.950 839.100 679.050 839.550 ;
        RECT 688.950 839.100 691.050 839.550 ;
        RECT 692.400 840.600 693.600 845.400 ;
        RECT 700.950 845.400 769.050 846.600 ;
        RECT 700.950 844.950 703.050 845.400 ;
        RECT 760.950 844.950 763.050 845.400 ;
        RECT 766.950 844.950 769.050 845.400 ;
        RECT 796.950 846.600 799.050 847.050 ;
        RECT 805.950 846.600 808.050 847.050 ;
        RECT 796.950 845.400 808.050 846.600 ;
        RECT 796.950 844.950 799.050 845.400 ;
        RECT 805.950 844.950 808.050 845.400 ;
        RECT 871.950 846.600 874.050 847.050 ;
        RECT 886.950 846.600 889.050 847.050 ;
        RECT 898.950 846.600 901.050 847.050 ;
        RECT 871.950 845.400 901.050 846.600 ;
        RECT 871.950 844.950 874.050 845.400 ;
        RECT 886.950 844.950 889.050 845.400 ;
        RECT 898.950 844.950 901.050 845.400 ;
        RECT 916.950 846.600 919.050 847.050 ;
        RECT 946.950 846.600 949.050 847.050 ;
        RECT 916.950 845.400 949.050 846.600 ;
        RECT 916.950 844.950 919.050 845.400 ;
        RECT 946.950 844.950 949.050 845.400 ;
        RECT 859.950 843.600 862.050 844.050 ;
        RECT 868.950 843.600 871.050 844.050 ;
        RECT 948.000 843.600 952.050 844.050 ;
        RECT 859.950 842.400 871.050 843.600 ;
        RECT 859.950 841.950 862.050 842.400 ;
        RECT 868.950 841.950 871.050 842.400 ;
        RECT 947.400 841.950 952.050 843.600 ;
        RECT 961.950 843.600 964.050 844.050 ;
        RECT 976.950 843.600 979.050 844.200 ;
        RECT 961.950 842.400 979.050 843.600 ;
        RECT 961.950 841.950 964.050 842.400 ;
        RECT 976.950 842.100 979.050 842.400 ;
        RECT 694.950 840.600 697.050 841.050 ;
        RECT 692.400 839.400 697.050 840.600 ;
        RECT 512.400 836.400 606.600 837.600 ;
        RECT 40.950 834.600 43.050 835.050 ;
        RECT 49.950 834.600 52.050 834.900 ;
        RECT 40.950 833.400 52.050 834.600 ;
        RECT 40.950 832.950 43.050 833.400 ;
        RECT 49.950 832.800 52.050 833.400 ;
        RECT 61.950 834.450 64.050 834.900 ;
        RECT 70.950 834.450 73.050 834.900 ;
        RECT 61.950 833.250 73.050 834.450 ;
        RECT 61.950 832.800 64.050 833.250 ;
        RECT 70.950 832.800 73.050 833.250 ;
        RECT 166.950 834.600 169.050 835.050 ;
        RECT 176.400 834.600 177.600 836.400 ;
        RECT 298.950 835.950 301.050 836.400 ;
        RECT 406.950 835.950 409.050 836.400 ;
        RECT 166.950 833.400 177.600 834.600 ;
        RECT 196.950 834.600 199.050 834.900 ;
        RECT 217.950 834.600 220.050 834.900 ;
        RECT 232.950 834.600 235.050 835.050 ;
        RECT 196.950 833.400 235.050 834.600 ;
        RECT 166.950 832.950 169.050 833.400 ;
        RECT 196.950 832.800 199.050 833.400 ;
        RECT 217.950 832.800 220.050 833.400 ;
        RECT 232.950 832.950 235.050 833.400 ;
        RECT 256.950 834.450 259.050 834.900 ;
        RECT 262.950 834.450 265.050 834.900 ;
        RECT 256.950 833.250 265.050 834.450 ;
        RECT 256.950 832.800 259.050 833.250 ;
        RECT 262.950 832.800 265.050 833.250 ;
        RECT 283.950 834.600 286.050 834.900 ;
        RECT 295.950 834.600 298.050 835.050 ;
        RECT 283.950 833.400 298.050 834.600 ;
        RECT 283.950 832.800 286.050 833.400 ;
        RECT 295.950 832.950 298.050 833.400 ;
        RECT 307.950 834.600 310.050 834.900 ;
        RECT 322.950 834.600 325.050 834.900 ;
        RECT 307.950 833.400 325.050 834.600 ;
        RECT 307.950 832.800 310.050 833.400 ;
        RECT 322.950 832.800 325.050 833.400 ;
        RECT 328.950 834.600 331.050 834.900 ;
        RECT 346.950 834.600 349.050 834.900 ;
        RECT 328.950 833.400 349.050 834.600 ;
        RECT 328.950 832.800 331.050 833.400 ;
        RECT 346.950 832.800 349.050 833.400 ;
        RECT 367.950 834.600 370.050 834.900 ;
        RECT 382.950 834.600 385.050 835.050 ;
        RECT 367.950 833.400 385.050 834.600 ;
        RECT 367.950 832.800 370.050 833.400 ;
        RECT 382.950 832.950 385.050 833.400 ;
        RECT 439.950 834.600 442.050 834.900 ;
        RECT 457.950 834.600 460.050 834.900 ;
        RECT 439.950 833.400 460.050 834.600 ;
        RECT 439.950 832.800 442.050 833.400 ;
        RECT 457.950 832.800 460.050 833.400 ;
        RECT 463.950 834.450 466.050 834.900 ;
        RECT 490.950 834.450 493.050 834.900 ;
        RECT 463.950 833.250 493.050 834.450 ;
        RECT 463.950 832.800 466.050 833.250 ;
        RECT 490.950 832.800 493.050 833.250 ;
        RECT 496.950 834.450 499.050 834.900 ;
        RECT 505.950 834.450 508.050 834.900 ;
        RECT 496.950 833.250 508.050 834.450 ;
        RECT 496.950 832.800 499.050 833.250 ;
        RECT 505.950 832.800 508.050 833.250 ;
        RECT 514.950 834.600 517.050 835.050 ;
        RECT 526.950 834.600 529.050 834.900 ;
        RECT 514.950 833.400 529.050 834.600 ;
        RECT 514.950 832.950 517.050 833.400 ;
        RECT 526.950 832.800 529.050 833.400 ;
        RECT 547.950 834.600 550.050 834.900 ;
        RECT 568.950 834.600 571.050 835.050 ;
        RECT 547.950 833.400 571.050 834.600 ;
        RECT 547.950 832.800 550.050 833.400 ;
        RECT 568.950 832.950 571.050 833.400 ;
        RECT 589.950 834.600 592.050 835.050 ;
        RECT 601.950 834.600 604.050 834.900 ;
        RECT 589.950 833.400 604.050 834.600 ;
        RECT 605.400 834.600 606.600 836.400 ;
        RECT 671.400 835.050 672.600 839.100 ;
        RECT 694.950 838.950 697.050 839.400 ;
        RECT 715.950 840.750 718.050 841.200 ;
        RECT 727.950 840.750 730.050 841.200 ;
        RECT 715.950 839.550 730.050 840.750 ;
        RECT 715.950 839.100 718.050 839.550 ;
        RECT 727.950 839.100 730.050 839.550 ;
        RECT 733.950 840.600 736.050 841.200 ;
        RECT 754.950 840.600 757.050 841.200 ;
        RECT 772.950 840.600 775.050 841.050 ;
        RECT 733.950 839.400 775.050 840.600 ;
        RECT 733.950 839.100 736.050 839.400 ;
        RECT 754.950 839.100 757.050 839.400 ;
        RECT 772.950 838.950 775.050 839.400 ;
        RECT 787.950 839.100 790.050 841.200 ;
        RECT 796.950 840.600 799.050 841.200 ;
        RECT 808.950 840.600 811.050 841.050 ;
        RECT 817.950 840.600 820.050 841.200 ;
        RECT 796.950 839.400 820.050 840.600 ;
        RECT 796.950 839.100 799.050 839.400 ;
        RECT 788.400 837.600 789.600 839.100 ;
        RECT 808.950 838.950 811.050 839.400 ;
        RECT 817.950 839.100 820.050 839.400 ;
        RECT 823.950 840.750 826.050 841.200 ;
        RECT 835.950 840.750 838.050 841.200 ;
        RECT 823.950 839.550 838.050 840.750 ;
        RECT 823.950 839.100 826.050 839.550 ;
        RECT 835.950 839.100 838.050 839.550 ;
        RECT 853.950 838.950 856.050 841.050 ;
        RECT 862.950 838.950 865.050 841.050 ;
        RECT 874.950 840.600 877.050 841.200 ;
        RECT 883.950 840.750 886.050 841.200 ;
        RECT 889.950 840.750 892.050 841.200 ;
        RECT 883.950 840.600 892.050 840.750 ;
        RECT 909.000 840.600 913.050 841.050 ;
        RECT 874.950 839.550 892.050 840.600 ;
        RECT 874.950 839.400 886.050 839.550 ;
        RECT 874.950 839.100 877.050 839.400 ;
        RECT 883.950 839.100 886.050 839.400 ;
        RECT 889.950 839.100 892.050 839.550 ;
        RECT 908.400 838.950 913.050 840.600 ;
        RECT 916.950 839.100 919.050 841.200 ;
        RECT 922.950 840.750 925.050 841.200 ;
        RECT 928.950 840.750 931.050 841.200 ;
        RECT 922.950 840.600 931.050 840.750 ;
        RECT 943.950 840.600 946.050 841.050 ;
        RECT 922.950 839.550 946.050 840.600 ;
        RECT 922.950 839.100 925.050 839.550 ;
        RECT 928.950 839.400 946.050 839.550 ;
        RECT 928.950 839.100 931.050 839.400 ;
        RECT 755.400 836.400 789.600 837.600 ;
        RECT 625.950 834.600 628.050 834.900 ;
        RECT 640.950 834.600 643.050 835.050 ;
        RECT 605.400 833.400 643.050 834.600 ;
        RECT 671.400 833.400 676.050 835.050 ;
        RECT 589.950 832.950 592.050 833.400 ;
        RECT 601.950 832.800 604.050 833.400 ;
        RECT 625.950 832.800 628.050 833.400 ;
        RECT 640.950 832.950 643.050 833.400 ;
        RECT 672.000 832.950 676.050 833.400 ;
        RECT 751.950 834.600 754.050 834.900 ;
        RECT 755.400 834.600 756.600 836.400 ;
        RECT 751.950 833.400 756.600 834.600 ;
        RECT 757.950 834.600 760.050 834.900 ;
        RECT 775.950 834.600 778.050 835.050 ;
        RECT 757.950 833.400 778.050 834.600 ;
        RECT 751.950 832.800 754.050 833.400 ;
        RECT 757.950 832.800 760.050 833.400 ;
        RECT 775.950 832.950 778.050 833.400 ;
        RECT 805.950 834.450 808.050 834.900 ;
        RECT 814.950 834.450 817.050 834.900 ;
        RECT 805.950 833.250 817.050 834.450 ;
        RECT 805.950 832.800 808.050 833.250 ;
        RECT 814.950 832.800 817.050 833.250 ;
        RECT 820.950 834.600 823.050 834.900 ;
        RECT 832.950 834.600 835.050 835.050 ;
        RECT 820.950 833.400 835.050 834.600 ;
        RECT 820.950 832.800 823.050 833.400 ;
        RECT 832.950 832.950 835.050 833.400 ;
        RECT 838.950 834.600 841.050 835.050 ;
        RECT 854.400 834.600 855.600 838.950 ;
        RECT 838.950 833.400 855.600 834.600 ;
        RECT 863.400 834.600 864.600 838.950 ;
        RECT 865.950 834.600 868.050 834.900 ;
        RECT 863.400 833.400 868.050 834.600 ;
        RECT 838.950 832.950 841.050 833.400 ;
        RECT 865.950 832.800 868.050 833.400 ;
        RECT 871.950 834.600 874.050 834.900 ;
        RECT 892.950 834.600 895.050 834.900 ;
        RECT 871.950 833.400 895.050 834.600 ;
        RECT 871.950 832.800 874.050 833.400 ;
        RECT 892.950 832.800 895.050 833.400 ;
        RECT 898.950 834.600 901.050 834.900 ;
        RECT 908.400 834.600 909.600 838.950 ;
        RECT 898.950 833.400 909.600 834.600 ;
        RECT 910.950 834.600 913.050 835.050 ;
        RECT 917.400 834.600 918.600 839.100 ;
        RECT 943.950 838.950 946.050 839.400 ;
        RECT 910.950 833.400 918.600 834.600 ;
        RECT 898.950 832.800 901.050 833.400 ;
        RECT 910.950 832.950 913.050 833.400 ;
        RECT 947.400 832.050 948.600 841.950 ;
        RECT 973.950 840.600 976.050 841.050 ;
        RECT 979.950 840.600 982.050 841.050 ;
        RECT 973.950 839.400 982.050 840.600 ;
        RECT 973.950 838.950 976.050 839.400 ;
        RECT 979.950 838.950 982.050 839.400 ;
        RECT 1009.950 838.950 1012.050 841.050 ;
        RECT 1010.400 835.050 1011.600 838.950 ;
        RECT 958.950 834.600 961.050 834.900 ;
        RECT 991.950 834.600 994.050 835.050 ;
        RECT 958.950 833.400 994.050 834.600 ;
        RECT 958.950 832.800 961.050 833.400 ;
        RECT 991.950 832.950 994.050 833.400 ;
        RECT 1009.950 832.950 1012.050 835.050 ;
        RECT 23.400 831.000 30.600 831.600 ;
        RECT 22.950 830.400 30.600 831.000 ;
        RECT 31.950 830.400 36.600 832.050 ;
        RECT 76.950 831.600 79.050 832.050 ;
        RECT 133.950 831.600 136.050 832.050 ;
        RECT 76.950 830.400 136.050 831.600 ;
        RECT 22.950 826.950 25.050 830.400 ;
        RECT 31.950 829.950 36.000 830.400 ;
        RECT 76.950 829.950 79.050 830.400 ;
        RECT 133.950 829.950 136.050 830.400 ;
        RECT 178.950 831.600 181.050 832.050 ;
        RECT 184.950 831.600 187.050 832.050 ;
        RECT 178.950 830.400 187.050 831.600 ;
        RECT 178.950 829.950 181.050 830.400 ;
        RECT 184.950 829.950 187.050 830.400 ;
        RECT 229.950 831.600 232.050 832.050 ;
        RECT 241.950 831.600 244.050 832.050 ;
        RECT 229.950 830.400 244.050 831.600 ;
        RECT 229.950 829.950 232.050 830.400 ;
        RECT 241.950 829.950 244.050 830.400 ;
        RECT 613.950 831.600 616.050 832.050 ;
        RECT 688.950 831.600 691.050 832.050 ;
        RECT 613.950 830.400 691.050 831.600 ;
        RECT 613.950 829.950 616.050 830.400 ;
        RECT 688.950 829.950 691.050 830.400 ;
        RECT 703.950 831.600 706.050 832.050 ;
        RECT 736.950 831.600 739.050 832.050 ;
        RECT 703.950 830.400 739.050 831.600 ;
        RECT 703.950 829.950 706.050 830.400 ;
        RECT 736.950 829.950 739.050 830.400 ;
        RECT 832.950 831.600 835.050 831.900 ;
        RECT 850.950 831.600 853.050 832.050 ;
        RECT 832.950 830.400 853.050 831.600 ;
        RECT 832.950 829.800 835.050 830.400 ;
        RECT 850.950 829.950 853.050 830.400 ;
        RECT 874.950 831.600 877.050 832.050 ;
        RECT 880.950 831.600 883.050 832.050 ;
        RECT 874.950 830.400 883.050 831.600 ;
        RECT 874.950 829.950 877.050 830.400 ;
        RECT 880.950 829.950 883.050 830.400 ;
        RECT 934.950 831.600 937.050 832.050 ;
        RECT 940.950 831.600 943.050 832.050 ;
        RECT 934.950 830.400 943.050 831.600 ;
        RECT 934.950 829.950 937.050 830.400 ;
        RECT 940.950 829.950 943.050 830.400 ;
        RECT 946.950 829.950 949.050 832.050 ;
        RECT 148.950 828.600 151.050 829.050 ;
        RECT 247.950 828.600 250.050 829.050 ;
        RECT 325.950 828.600 328.050 829.050 ;
        RECT 148.950 827.400 328.050 828.600 ;
        RECT 148.950 826.950 151.050 827.400 ;
        RECT 247.950 826.950 250.050 827.400 ;
        RECT 325.950 826.950 328.050 827.400 ;
        RECT 331.950 828.600 334.050 829.050 ;
        RECT 349.950 828.600 352.050 829.050 ;
        RECT 331.950 827.400 352.050 828.600 ;
        RECT 331.950 826.950 334.050 827.400 ;
        RECT 349.950 826.950 352.050 827.400 ;
        RECT 355.950 828.600 358.050 829.050 ;
        RECT 388.950 828.600 391.050 829.050 ;
        RECT 355.950 827.400 391.050 828.600 ;
        RECT 355.950 826.950 358.050 827.400 ;
        RECT 388.950 826.950 391.050 827.400 ;
        RECT 394.950 828.600 397.050 829.050 ;
        RECT 415.950 828.600 418.050 829.050 ;
        RECT 505.950 828.600 508.050 829.050 ;
        RECT 394.950 827.400 508.050 828.600 ;
        RECT 394.950 826.950 397.050 827.400 ;
        RECT 415.950 826.950 418.050 827.400 ;
        RECT 505.950 826.950 508.050 827.400 ;
        RECT 625.950 828.600 628.050 829.050 ;
        RECT 640.950 828.600 643.050 829.050 ;
        RECT 646.950 828.600 649.050 829.050 ;
        RECT 625.950 827.400 649.050 828.600 ;
        RECT 625.950 826.950 628.050 827.400 ;
        RECT 640.950 826.950 643.050 827.400 ;
        RECT 646.950 826.950 649.050 827.400 ;
        RECT 664.950 828.600 667.050 829.050 ;
        RECT 676.800 828.600 678.900 829.050 ;
        RECT 664.950 827.400 678.900 828.600 ;
        RECT 664.950 826.950 667.050 827.400 ;
        RECT 676.800 826.950 678.900 827.400 ;
        RECT 679.950 828.600 682.050 829.050 ;
        RECT 691.950 828.600 694.050 829.050 ;
        RECT 679.950 827.400 694.050 828.600 ;
        RECT 679.950 826.950 682.050 827.400 ;
        RECT 691.950 826.950 694.050 827.400 ;
        RECT 823.950 828.600 826.050 829.050 ;
        RECT 829.950 828.600 832.050 829.050 ;
        RECT 823.950 827.400 832.050 828.600 ;
        RECT 823.950 826.950 826.050 827.400 ;
        RECT 829.950 826.950 832.050 827.400 ;
        RECT 955.950 828.600 958.050 829.050 ;
        RECT 961.950 828.600 964.050 829.050 ;
        RECT 955.950 827.400 964.050 828.600 ;
        RECT 955.950 826.950 958.050 827.400 ;
        RECT 961.950 826.950 964.050 827.400 ;
        RECT 970.950 828.600 973.050 829.050 ;
        RECT 985.950 828.600 988.050 829.050 ;
        RECT 970.950 827.400 988.050 828.600 ;
        RECT 970.950 826.950 973.050 827.400 ;
        RECT 985.950 826.950 988.050 827.400 ;
        RECT 991.950 828.600 994.050 829.050 ;
        RECT 1006.950 828.600 1009.050 829.050 ;
        RECT 991.950 827.400 1009.050 828.600 ;
        RECT 991.950 826.950 994.050 827.400 ;
        RECT 1006.950 826.950 1009.050 827.400 ;
        RECT 34.950 825.600 37.050 826.050 ;
        RECT 58.950 825.600 61.050 826.050 ;
        RECT 395.400 825.600 396.600 826.950 ;
        RECT 34.950 824.400 396.600 825.600 ;
        RECT 448.950 825.600 451.050 826.050 ;
        RECT 460.950 825.600 463.050 826.050 ;
        RECT 448.950 824.400 463.050 825.600 ;
        RECT 34.950 823.950 37.050 824.400 ;
        RECT 58.950 823.950 61.050 824.400 ;
        RECT 448.950 823.950 451.050 824.400 ;
        RECT 460.950 823.950 463.050 824.400 ;
        RECT 481.950 825.600 484.050 826.050 ;
        RECT 517.950 825.600 520.050 826.050 ;
        RECT 481.950 824.400 520.050 825.600 ;
        RECT 481.950 823.950 484.050 824.400 ;
        RECT 517.950 823.950 520.050 824.400 ;
        RECT 565.950 825.600 568.050 826.050 ;
        RECT 580.950 825.600 583.050 826.050 ;
        RECT 565.950 824.400 583.050 825.600 ;
        RECT 565.950 823.950 568.050 824.400 ;
        RECT 580.950 823.950 583.050 824.400 ;
        RECT 655.950 825.600 658.050 826.050 ;
        RECT 703.950 825.600 706.050 826.050 ;
        RECT 655.950 824.400 706.050 825.600 ;
        RECT 655.950 823.950 658.050 824.400 ;
        RECT 703.950 823.950 706.050 824.400 ;
        RECT 733.950 825.600 736.050 826.050 ;
        RECT 742.950 825.600 745.050 826.050 ;
        RECT 751.950 825.600 754.050 826.050 ;
        RECT 733.950 824.400 754.050 825.600 ;
        RECT 733.950 823.950 736.050 824.400 ;
        RECT 742.950 823.950 745.050 824.400 ;
        RECT 751.950 823.950 754.050 824.400 ;
        RECT 781.950 825.600 784.050 825.900 ;
        RECT 835.950 825.600 838.050 826.050 ;
        RECT 844.950 825.600 847.050 826.050 ;
        RECT 781.950 824.400 847.050 825.600 ;
        RECT 781.950 823.800 784.050 824.400 ;
        RECT 835.950 823.950 838.050 824.400 ;
        RECT 844.950 823.950 847.050 824.400 ;
        RECT 859.950 825.600 862.050 826.050 ;
        RECT 871.950 825.600 874.050 826.050 ;
        RECT 859.950 824.400 874.050 825.600 ;
        RECT 859.950 823.950 862.050 824.400 ;
        RECT 871.950 823.950 874.050 824.400 ;
        RECT 895.950 825.600 898.050 826.050 ;
        RECT 904.950 825.600 907.050 826.050 ;
        RECT 895.950 824.400 907.050 825.600 ;
        RECT 895.950 823.950 898.050 824.400 ;
        RECT 904.950 823.950 907.050 824.400 ;
        RECT 928.950 825.600 931.050 826.050 ;
        RECT 940.950 825.600 943.050 826.050 ;
        RECT 949.950 825.600 952.050 826.050 ;
        RECT 928.950 824.400 952.050 825.600 ;
        RECT 928.950 823.950 931.050 824.400 ;
        RECT 940.950 823.950 943.050 824.400 ;
        RECT 949.950 823.950 952.050 824.400 ;
        RECT 79.950 822.600 82.050 823.050 ;
        RECT 94.950 822.600 97.050 823.050 ;
        RECT 79.950 821.400 97.050 822.600 ;
        RECT 79.950 820.950 82.050 821.400 ;
        RECT 94.950 820.950 97.050 821.400 ;
        RECT 196.950 822.600 199.050 823.050 ;
        RECT 319.800 822.600 321.900 823.050 ;
        RECT 196.950 821.400 321.900 822.600 ;
        RECT 196.950 820.950 199.050 821.400 ;
        RECT 319.800 820.950 321.900 821.400 ;
        RECT 322.950 822.600 325.050 823.050 ;
        RECT 391.950 822.600 394.050 823.050 ;
        RECT 322.950 821.400 394.050 822.600 ;
        RECT 322.950 820.950 325.050 821.400 ;
        RECT 391.950 820.950 394.050 821.400 ;
        RECT 397.950 822.600 400.050 823.050 ;
        RECT 439.950 822.600 442.050 823.050 ;
        RECT 397.950 821.400 442.050 822.600 ;
        RECT 397.950 820.950 400.050 821.400 ;
        RECT 439.950 820.950 442.050 821.400 ;
        RECT 694.950 822.600 697.050 823.050 ;
        RECT 700.950 822.600 703.050 823.050 ;
        RECT 694.950 821.400 703.050 822.600 ;
        RECT 694.950 820.950 697.050 821.400 ;
        RECT 700.950 820.950 703.050 821.400 ;
        RECT 706.950 822.600 709.050 823.050 ;
        RECT 721.950 822.600 724.050 823.050 ;
        RECT 706.950 821.400 724.050 822.600 ;
        RECT 706.950 820.950 709.050 821.400 ;
        RECT 721.950 820.950 724.050 821.400 ;
        RECT 919.950 822.600 922.050 823.050 ;
        RECT 982.950 822.600 985.050 823.050 ;
        RECT 1009.950 822.600 1012.050 823.050 ;
        RECT 919.950 821.400 1012.050 822.600 ;
        RECT 919.950 820.950 922.050 821.400 ;
        RECT 982.950 820.950 985.050 821.400 ;
        RECT 1009.950 820.950 1012.050 821.400 ;
        RECT 118.950 819.600 121.050 820.050 ;
        RECT 163.950 819.600 166.050 820.050 ;
        RECT 118.950 818.400 166.050 819.600 ;
        RECT 118.950 817.950 121.050 818.400 ;
        RECT 163.950 817.950 166.050 818.400 ;
        RECT 202.950 819.600 205.050 820.050 ;
        RECT 280.950 819.600 283.050 820.050 ;
        RECT 202.950 818.400 283.050 819.600 ;
        RECT 202.950 817.950 205.050 818.400 ;
        RECT 280.950 817.950 283.050 818.400 ;
        RECT 349.950 819.600 352.050 820.050 ;
        RECT 376.950 819.600 379.050 820.050 ;
        RECT 349.950 818.400 379.050 819.600 ;
        RECT 349.950 817.950 352.050 818.400 ;
        RECT 376.950 817.950 379.050 818.400 ;
        RECT 529.950 819.600 532.050 820.050 ;
        RECT 535.950 819.600 538.050 820.050 ;
        RECT 529.950 818.400 538.050 819.600 ;
        RECT 529.950 817.950 532.050 818.400 ;
        RECT 535.950 817.950 538.050 818.400 ;
        RECT 553.950 819.600 556.050 820.050 ;
        RECT 577.950 819.600 580.050 820.050 ;
        RECT 655.950 819.600 658.050 820.050 ;
        RECT 553.950 818.400 658.050 819.600 ;
        RECT 553.950 817.950 556.050 818.400 ;
        RECT 577.950 817.950 580.050 818.400 ;
        RECT 655.950 817.950 658.050 818.400 ;
        RECT 667.950 819.600 670.050 820.050 ;
        RECT 844.950 819.600 847.050 820.050 ;
        RECT 883.950 819.600 886.050 820.050 ;
        RECT 667.950 818.400 886.050 819.600 ;
        RECT 667.950 817.950 670.050 818.400 ;
        RECT 844.950 817.950 847.050 818.400 ;
        RECT 883.950 817.950 886.050 818.400 ;
        RECT 892.950 819.600 895.050 820.050 ;
        RECT 901.950 819.600 904.050 820.050 ;
        RECT 892.950 818.400 904.050 819.600 ;
        RECT 892.950 817.950 895.050 818.400 ;
        RECT 901.950 817.950 904.050 818.400 ;
        RECT 373.950 816.600 376.050 817.050 ;
        RECT 406.950 816.600 409.050 817.050 ;
        RECT 445.950 816.600 448.050 817.050 ;
        RECT 373.950 815.400 448.050 816.600 ;
        RECT 373.950 814.950 376.050 815.400 ;
        RECT 406.950 814.950 409.050 815.400 ;
        RECT 445.950 814.950 448.050 815.400 ;
        RECT 688.950 816.600 691.050 817.050 ;
        RECT 712.950 816.600 715.050 817.050 ;
        RECT 688.950 815.400 715.050 816.600 ;
        RECT 688.950 814.950 691.050 815.400 ;
        RECT 712.950 814.950 715.050 815.400 ;
        RECT 742.950 816.600 745.050 817.050 ;
        RECT 787.950 816.600 790.050 817.050 ;
        RECT 742.950 815.400 790.050 816.600 ;
        RECT 742.950 814.950 745.050 815.400 ;
        RECT 787.950 814.950 790.050 815.400 ;
        RECT 913.950 816.600 916.050 817.050 ;
        RECT 934.950 816.600 937.050 817.050 ;
        RECT 913.950 815.400 937.050 816.600 ;
        RECT 913.950 814.950 916.050 815.400 ;
        RECT 934.950 814.950 937.050 815.400 ;
        RECT 973.950 816.600 976.050 817.050 ;
        RECT 997.950 816.600 1000.050 817.050 ;
        RECT 973.950 815.400 1000.050 816.600 ;
        RECT 973.950 814.950 976.050 815.400 ;
        RECT 997.950 814.950 1000.050 815.400 ;
        RECT 169.950 813.600 172.050 814.050 ;
        RECT 211.950 813.600 214.050 814.050 ;
        RECT 169.950 812.400 214.050 813.600 ;
        RECT 169.950 811.950 172.050 812.400 ;
        RECT 211.950 811.950 214.050 812.400 ;
        RECT 313.950 811.950 316.050 814.050 ;
        RECT 328.950 813.600 331.050 814.050 ;
        RECT 334.950 813.600 337.050 814.050 ;
        RECT 328.950 812.400 337.050 813.600 ;
        RECT 328.950 811.950 331.050 812.400 ;
        RECT 334.950 811.950 337.050 812.400 ;
        RECT 397.950 813.600 400.050 814.050 ;
        RECT 409.950 813.600 412.050 814.050 ;
        RECT 397.950 812.400 412.050 813.600 ;
        RECT 397.950 811.950 400.050 812.400 ;
        RECT 409.950 811.950 412.050 812.400 ;
        RECT 523.950 813.600 526.050 814.050 ;
        RECT 532.950 813.600 535.050 814.050 ;
        RECT 547.950 813.600 550.050 814.050 ;
        RECT 523.950 812.400 550.050 813.600 ;
        RECT 523.950 811.950 526.050 812.400 ;
        RECT 532.950 811.950 535.050 812.400 ;
        RECT 547.950 811.950 550.050 812.400 ;
        RECT 808.950 813.600 811.050 814.050 ;
        RECT 820.950 813.600 823.050 814.050 ;
        RECT 808.950 812.400 823.050 813.600 ;
        RECT 808.950 811.950 811.050 812.400 ;
        RECT 820.950 811.950 823.050 812.400 ;
        RECT 850.950 813.600 853.050 814.050 ;
        RECT 859.950 813.600 862.050 814.050 ;
        RECT 877.950 813.600 880.050 814.050 ;
        RECT 850.950 812.400 880.050 813.600 ;
        RECT 850.950 811.950 853.050 812.400 ;
        RECT 859.950 811.950 862.050 812.400 ;
        RECT 877.950 811.950 880.050 812.400 ;
        RECT 943.950 813.600 946.050 814.050 ;
        RECT 967.950 813.600 970.050 814.050 ;
        RECT 943.950 812.400 970.050 813.600 ;
        RECT 943.950 811.950 946.050 812.400 ;
        RECT 967.950 811.950 970.050 812.400 ;
        RECT 988.950 813.600 991.050 814.050 ;
        RECT 994.950 813.600 997.050 814.050 ;
        RECT 988.950 812.400 997.050 813.600 ;
        RECT 988.950 811.950 991.050 812.400 ;
        RECT 994.950 811.950 997.050 812.400 ;
        RECT 91.950 810.600 94.050 811.050 ;
        RECT 100.950 810.600 103.050 811.050 ;
        RECT 118.950 810.600 121.050 811.050 ;
        RECT 91.950 809.400 121.050 810.600 ;
        RECT 91.950 808.950 94.050 809.400 ;
        RECT 100.950 808.950 103.050 809.400 ;
        RECT 118.950 808.950 121.050 809.400 ;
        RECT 133.950 810.600 136.050 811.050 ;
        RECT 139.950 810.600 142.050 811.050 ;
        RECT 133.950 809.400 142.050 810.600 ;
        RECT 133.950 808.950 136.050 809.400 ;
        RECT 139.950 808.950 142.050 809.400 ;
        RECT 16.950 807.600 19.050 808.200 ;
        RECT 22.950 807.600 25.050 808.200 ;
        RECT 31.950 807.600 34.050 808.050 ;
        RECT 16.950 806.400 34.050 807.600 ;
        RECT 16.950 806.100 19.050 806.400 ;
        RECT 22.950 806.100 25.050 806.400 ;
        RECT 31.950 805.950 34.050 806.400 ;
        RECT 124.950 807.600 127.050 808.200 ;
        RECT 142.950 807.600 145.050 808.200 ;
        RECT 151.950 807.600 154.050 808.050 ;
        RECT 124.950 806.400 141.600 807.600 ;
        RECT 124.950 806.100 127.050 806.400 ;
        RECT 140.400 804.600 141.600 806.400 ;
        RECT 142.950 806.400 154.050 807.600 ;
        RECT 142.950 806.100 145.050 806.400 ;
        RECT 151.950 805.950 154.050 806.400 ;
        RECT 190.950 807.600 193.050 808.200 ;
        RECT 217.950 807.600 220.050 808.050 ;
        RECT 190.950 806.400 220.050 807.600 ;
        RECT 190.950 806.100 193.050 806.400 ;
        RECT 217.950 805.950 220.050 806.400 ;
        RECT 229.950 807.750 232.050 808.200 ;
        RECT 235.950 807.750 238.050 808.200 ;
        RECT 229.950 806.550 238.050 807.750 ;
        RECT 229.950 806.100 232.050 806.550 ;
        RECT 235.950 806.100 238.050 806.550 ;
        RECT 241.950 807.600 244.050 808.050 ;
        RECT 253.950 807.600 256.050 808.200 ;
        RECT 241.950 806.400 256.050 807.600 ;
        RECT 314.400 807.600 315.600 811.950 ;
        RECT 526.950 810.600 529.050 811.050 ;
        RECT 541.950 810.600 544.050 811.050 ;
        RECT 526.950 809.400 544.050 810.600 ;
        RECT 526.950 808.950 529.050 809.400 ;
        RECT 541.950 808.950 544.050 809.400 ;
        RECT 601.950 810.600 604.050 811.050 ;
        RECT 607.950 810.600 610.050 811.050 ;
        RECT 601.950 809.400 610.050 810.600 ;
        RECT 601.950 808.950 604.050 809.400 ;
        RECT 607.950 808.950 610.050 809.400 ;
        RECT 847.950 810.600 850.050 811.050 ;
        RECT 856.950 810.600 859.050 811.050 ;
        RECT 975.000 810.600 979.050 811.050 ;
        RECT 847.950 809.400 859.050 810.600 ;
        RECT 847.950 808.950 850.050 809.400 ;
        RECT 856.950 808.950 859.050 809.400 ;
        RECT 974.400 808.950 979.050 810.600 ;
        RECT 319.950 807.750 322.050 808.200 ;
        RECT 325.950 807.750 328.050 808.200 ;
        RECT 314.400 806.400 318.600 807.600 ;
        RECT 241.950 805.950 244.050 806.400 ;
        RECT 253.950 806.100 256.050 806.400 ;
        RECT 154.950 804.600 157.050 805.050 ;
        RECT 140.400 803.400 157.050 804.600 ;
        RECT 317.400 804.600 318.600 806.400 ;
        RECT 319.950 806.550 328.050 807.750 ;
        RECT 319.950 806.100 322.050 806.550 ;
        RECT 325.950 806.100 328.050 806.550 ;
        RECT 355.950 807.600 358.050 808.050 ;
        RECT 367.950 807.600 370.050 808.200 ;
        RECT 355.950 806.400 370.050 807.600 ;
        RECT 355.950 805.950 358.050 806.400 ;
        RECT 367.950 806.100 370.050 806.400 ;
        RECT 391.950 807.750 394.050 808.200 ;
        RECT 403.950 807.750 406.050 808.200 ;
        RECT 391.950 806.550 406.050 807.750 ;
        RECT 391.950 806.100 394.050 806.550 ;
        RECT 403.950 806.100 406.050 806.550 ;
        RECT 415.950 807.600 418.050 808.200 ;
        RECT 421.950 807.600 424.050 808.050 ;
        RECT 415.950 806.400 424.050 807.600 ;
        RECT 415.950 806.100 418.050 806.400 ;
        RECT 421.950 805.950 424.050 806.400 ;
        RECT 439.950 806.100 442.050 808.200 ;
        RECT 556.950 807.600 559.050 808.200 ;
        RECT 571.950 807.600 574.050 808.050 ;
        RECT 631.950 807.600 634.050 808.200 ;
        RECT 556.950 806.400 634.050 807.600 ;
        RECT 556.950 806.100 559.050 806.400 ;
        RECT 322.950 804.600 325.050 805.050 ;
        RECT 317.400 803.400 325.050 804.600 ;
        RECT 154.950 802.950 157.050 803.400 ;
        RECT 322.950 802.950 325.050 803.400 ;
        RECT 7.950 801.600 10.050 802.050 ;
        RECT 13.950 801.600 16.050 801.900 ;
        RECT 7.950 800.400 16.050 801.600 ;
        RECT 7.950 799.950 10.050 800.400 ;
        RECT 13.950 799.800 16.050 800.400 ;
        RECT 31.950 801.450 34.050 801.900 ;
        RECT 40.950 801.450 43.050 801.900 ;
        RECT 31.950 800.250 43.050 801.450 ;
        RECT 31.950 799.800 34.050 800.250 ;
        RECT 40.950 799.800 43.050 800.250 ;
        RECT 88.950 801.600 91.050 801.900 ;
        RECT 109.950 801.600 112.050 801.900 ;
        RECT 88.950 801.450 112.050 801.600 ;
        RECT 115.950 801.450 118.050 801.900 ;
        RECT 88.950 800.400 118.050 801.450 ;
        RECT 88.950 799.800 91.050 800.400 ;
        RECT 109.950 800.250 118.050 800.400 ;
        RECT 109.950 799.800 112.050 800.250 ;
        RECT 115.950 799.800 118.050 800.250 ;
        RECT 121.950 801.450 124.050 801.900 ;
        RECT 130.800 801.450 132.900 801.900 ;
        RECT 121.950 800.250 132.900 801.450 ;
        RECT 121.950 799.800 124.050 800.250 ;
        RECT 130.800 799.800 132.900 800.250 ;
        RECT 133.950 801.450 136.050 801.900 ;
        RECT 139.950 801.450 142.050 801.900 ;
        RECT 133.950 800.250 142.050 801.450 ;
        RECT 133.950 799.800 136.050 800.250 ;
        RECT 139.950 799.800 142.050 800.250 ;
        RECT 166.950 801.600 169.050 801.900 ;
        RECT 193.950 801.600 196.050 801.900 ;
        RECT 166.950 800.400 196.050 801.600 ;
        RECT 166.950 799.800 169.050 800.400 ;
        RECT 193.950 799.800 196.050 800.400 ;
        RECT 211.950 801.450 214.050 801.900 ;
        RECT 217.950 801.450 220.050 801.900 ;
        RECT 211.950 800.250 220.050 801.450 ;
        RECT 211.950 799.800 214.050 800.250 ;
        RECT 217.950 799.800 220.050 800.250 ;
        RECT 262.950 801.450 265.050 801.900 ;
        RECT 271.950 801.450 274.050 801.900 ;
        RECT 262.950 800.250 274.050 801.450 ;
        RECT 262.950 799.800 265.050 800.250 ;
        RECT 271.950 799.800 274.050 800.250 ;
        RECT 328.950 801.600 331.050 802.050 ;
        RECT 340.950 801.600 343.050 801.900 ;
        RECT 328.950 800.400 343.050 801.600 ;
        RECT 328.950 799.950 331.050 800.400 ;
        RECT 340.950 799.800 343.050 800.400 ;
        RECT 370.950 801.600 373.050 801.900 ;
        RECT 388.950 801.600 391.050 801.900 ;
        RECT 370.950 800.400 391.050 801.600 ;
        RECT 370.950 799.800 373.050 800.400 ;
        RECT 388.950 799.800 391.050 800.400 ;
        RECT 400.950 801.450 403.050 801.900 ;
        RECT 406.950 801.600 409.050 801.900 ;
        RECT 440.400 801.600 441.600 806.100 ;
        RECT 571.950 805.950 574.050 806.400 ;
        RECT 631.950 806.100 634.050 806.400 ;
        RECT 649.950 807.750 652.050 808.200 ;
        RECT 661.950 807.750 664.050 808.200 ;
        RECT 649.950 806.550 664.050 807.750 ;
        RECT 649.950 806.100 652.050 806.550 ;
        RECT 661.950 806.100 664.050 806.550 ;
        RECT 742.950 807.600 745.050 808.200 ;
        RECT 742.950 806.400 750.600 807.600 ;
        RECT 742.950 806.100 745.050 806.400 ;
        RECT 406.950 801.450 441.600 801.600 ;
        RECT 400.950 800.400 441.600 801.450 ;
        RECT 445.950 801.600 448.050 802.050 ;
        RECT 487.950 801.600 490.050 801.900 ;
        RECT 445.950 800.400 490.050 801.600 ;
        RECT 400.950 800.250 409.050 800.400 ;
        RECT 400.950 799.800 403.050 800.250 ;
        RECT 406.950 799.800 409.050 800.250 ;
        RECT 445.950 799.950 448.050 800.400 ;
        RECT 487.950 799.800 490.050 800.400 ;
        RECT 493.950 801.600 496.050 801.900 ;
        RECT 517.950 801.600 520.050 801.900 ;
        RECT 493.950 800.400 520.050 801.600 ;
        RECT 493.950 799.800 496.050 800.400 ;
        RECT 517.950 799.800 520.050 800.400 ;
        RECT 547.950 801.600 550.050 802.050 ;
        RECT 559.950 801.600 562.050 801.900 ;
        RECT 547.950 800.400 562.050 801.600 ;
        RECT 547.950 799.950 550.050 800.400 ;
        RECT 559.950 799.800 562.050 800.400 ;
        RECT 571.950 801.450 574.050 801.900 ;
        RECT 577.950 801.450 580.050 801.900 ;
        RECT 571.950 800.250 580.050 801.450 ;
        RECT 571.950 799.800 574.050 800.250 ;
        RECT 577.950 799.800 580.050 800.250 ;
        RECT 583.950 801.600 586.050 801.900 ;
        RECT 598.950 801.600 601.050 801.900 ;
        RECT 583.950 800.400 601.050 801.600 ;
        RECT 583.950 799.800 586.050 800.400 ;
        RECT 598.950 799.800 601.050 800.400 ;
        RECT 604.950 801.450 607.050 801.900 ;
        RECT 616.950 801.450 619.050 801.900 ;
        RECT 604.950 800.250 619.050 801.450 ;
        RECT 604.950 799.800 607.050 800.250 ;
        RECT 616.950 799.800 619.050 800.250 ;
        RECT 640.950 801.450 643.050 801.900 ;
        RECT 646.950 801.450 649.050 801.900 ;
        RECT 640.950 800.250 649.050 801.450 ;
        RECT 640.950 799.800 643.050 800.250 ;
        RECT 646.950 799.800 649.050 800.250 ;
        RECT 652.950 801.600 655.050 801.900 ;
        RECT 670.950 801.600 673.050 801.900 ;
        RECT 652.950 800.400 673.050 801.600 ;
        RECT 749.400 801.600 750.600 806.400 ;
        RECT 763.950 806.100 766.050 808.200 ;
        RECT 769.950 807.750 772.050 808.200 ;
        RECT 778.950 807.750 781.050 808.200 ;
        RECT 769.950 806.550 781.050 807.750 ;
        RECT 769.950 806.100 772.050 806.550 ;
        RECT 778.950 806.100 781.050 806.550 ;
        RECT 808.950 807.600 811.050 808.200 ;
        RECT 868.950 807.750 871.050 808.200 ;
        RECT 880.950 807.750 883.050 808.200 ;
        RECT 808.950 806.400 837.600 807.600 ;
        RECT 808.950 806.100 811.050 806.400 ;
        RECT 754.950 804.600 757.050 805.050 ;
        RECT 764.400 804.600 765.600 806.100 ;
        RECT 781.950 804.600 784.050 805.050 ;
        RECT 754.950 803.400 765.600 804.600 ;
        RECT 776.400 803.400 784.050 804.600 ;
        RECT 754.950 802.950 757.050 803.400 ;
        RECT 766.950 801.600 769.050 801.900 ;
        RECT 776.400 801.600 777.600 803.400 ;
        RECT 781.950 802.950 784.050 803.400 ;
        RECT 749.400 800.400 753.600 801.600 ;
        RECT 652.950 799.800 655.050 800.400 ;
        RECT 670.950 799.800 673.050 800.400 ;
        RECT 598.950 798.600 601.050 799.050 ;
        RECT 634.950 798.600 637.050 799.050 ;
        RECT 598.950 797.400 637.050 798.600 ;
        RECT 752.400 798.600 753.600 800.400 ;
        RECT 766.950 800.400 777.600 801.600 ;
        RECT 778.950 801.600 781.050 802.050 ;
        RECT 790.950 801.600 793.050 801.900 ;
        RECT 778.950 800.400 793.050 801.600 ;
        RECT 766.950 799.800 769.050 800.400 ;
        RECT 778.950 799.950 781.050 800.400 ;
        RECT 790.950 799.800 793.050 800.400 ;
        RECT 799.950 801.600 802.050 802.050 ;
        RECT 836.400 801.900 837.600 806.400 ;
        RECT 868.950 806.550 883.050 807.750 ;
        RECT 868.950 806.100 871.050 806.550 ;
        RECT 880.950 806.100 883.050 806.550 ;
        RECT 886.950 807.600 889.050 808.200 ;
        RECT 904.950 807.600 907.050 808.200 ;
        RECT 886.950 806.400 907.050 807.600 ;
        RECT 886.950 806.100 889.050 806.400 ;
        RECT 904.950 806.100 907.050 806.400 ;
        RECT 910.950 807.600 913.050 808.200 ;
        RECT 916.800 807.600 918.900 808.050 ;
        RECT 910.950 806.400 918.900 807.600 ;
        RECT 910.950 806.100 913.050 806.400 ;
        RECT 916.800 805.950 918.900 806.400 ;
        RECT 919.950 807.600 922.050 808.050 ;
        RECT 928.950 807.600 931.050 808.200 ;
        RECT 919.950 806.400 931.050 807.600 ;
        RECT 919.950 805.950 922.050 806.400 ;
        RECT 928.950 806.100 931.050 806.400 ;
        RECT 949.950 807.750 952.050 808.200 ;
        RECT 955.950 807.750 958.050 808.200 ;
        RECT 949.950 806.550 958.050 807.750 ;
        RECT 949.950 806.100 952.050 806.550 ;
        RECT 955.950 806.100 958.050 806.550 ;
        RECT 863.400 803.400 879.600 804.600 ;
        RECT 863.400 801.900 864.600 803.400 ;
        RECT 878.400 801.900 879.600 803.400 ;
        RECT 805.950 801.600 808.050 801.900 ;
        RECT 799.950 800.400 808.050 801.600 ;
        RECT 799.950 799.950 802.050 800.400 ;
        RECT 805.950 799.800 808.050 800.400 ;
        RECT 811.950 801.450 814.050 801.900 ;
        RECT 820.950 801.450 823.050 801.900 ;
        RECT 811.950 800.250 823.050 801.450 ;
        RECT 811.950 799.800 814.050 800.250 ;
        RECT 820.950 799.800 823.050 800.250 ;
        RECT 835.950 799.800 838.050 801.900 ;
        RECT 844.950 801.450 847.050 801.900 ;
        RECT 862.950 801.450 865.050 801.900 ;
        RECT 844.950 800.250 865.050 801.450 ;
        RECT 844.950 799.800 847.050 800.250 ;
        RECT 862.950 799.800 865.050 800.250 ;
        RECT 877.950 799.800 880.050 801.900 ;
        RECT 883.950 801.600 886.050 801.900 ;
        RECT 892.950 801.600 895.050 802.050 ;
        RECT 883.950 800.400 895.050 801.600 ;
        RECT 883.950 799.800 886.050 800.400 ;
        RECT 892.950 799.950 895.050 800.400 ;
        RECT 916.950 801.450 919.050 801.900 ;
        RECT 931.950 801.450 934.050 801.900 ;
        RECT 916.950 800.250 934.050 801.450 ;
        RECT 916.950 799.800 919.050 800.250 ;
        RECT 931.950 799.800 934.050 800.250 ;
        RECT 943.950 801.600 946.050 802.050 ;
        RECT 952.950 801.600 955.050 801.900 ;
        RECT 970.950 801.600 973.050 801.900 ;
        RECT 943.950 800.400 973.050 801.600 ;
        RECT 943.950 799.950 946.050 800.400 ;
        RECT 952.950 799.800 955.050 800.400 ;
        RECT 970.950 799.800 973.050 800.400 ;
        RECT 974.400 799.050 975.600 808.950 ;
        RECT 994.950 807.600 997.050 808.200 ;
        RECT 992.400 806.400 997.050 807.600 ;
        RECT 992.400 802.050 993.600 806.400 ;
        RECT 994.950 806.100 997.050 806.400 ;
        RECT 1006.950 805.950 1009.050 808.050 ;
        RECT 1007.400 802.050 1008.600 805.950 ;
        RECT 976.950 801.600 979.050 801.900 ;
        RECT 976.950 800.400 981.600 801.600 ;
        RECT 976.950 799.800 979.050 800.400 ;
        RECT 763.950 798.600 766.050 799.050 ;
        RECT 752.400 797.400 766.050 798.600 ;
        RECT 598.950 796.950 601.050 797.400 ;
        RECT 634.950 796.950 637.050 797.400 ;
        RECT 763.950 796.950 766.050 797.400 ;
        RECT 934.950 798.600 937.050 799.050 ;
        RECT 940.950 798.600 943.050 799.050 ;
        RECT 934.950 797.400 943.050 798.600 ;
        RECT 934.950 796.950 937.050 797.400 ;
        RECT 940.950 796.950 943.050 797.400 ;
        RECT 973.950 796.950 976.050 799.050 ;
        RECT 980.400 798.600 981.600 800.400 ;
        RECT 991.950 799.950 994.050 802.050 ;
        RECT 1006.950 799.950 1009.050 802.050 ;
        RECT 1003.950 798.600 1006.050 799.050 ;
        RECT 1009.950 798.600 1012.050 799.050 ;
        RECT 980.400 797.400 1012.050 798.600 ;
        RECT 1003.950 796.950 1006.050 797.400 ;
        RECT 1009.950 796.950 1012.050 797.400 ;
        RECT 103.950 795.600 106.050 796.050 ;
        RECT 145.950 795.600 148.050 796.050 ;
        RECT 103.950 794.400 148.050 795.600 ;
        RECT 103.950 793.950 106.050 794.400 ;
        RECT 145.950 793.950 148.050 794.400 ;
        RECT 379.950 795.600 382.050 796.050 ;
        RECT 412.950 795.600 415.050 796.050 ;
        RECT 433.950 795.600 436.050 796.050 ;
        RECT 379.950 794.400 436.050 795.600 ;
        RECT 379.950 793.950 382.050 794.400 ;
        RECT 412.950 793.950 415.050 794.400 ;
        RECT 433.950 793.950 436.050 794.400 ;
        RECT 502.950 795.600 505.050 796.050 ;
        RECT 706.950 795.600 709.050 796.050 ;
        RECT 502.950 794.400 709.050 795.600 ;
        RECT 502.950 793.950 505.050 794.400 ;
        RECT 706.950 793.950 709.050 794.400 ;
        RECT 715.950 795.600 718.050 796.050 ;
        RECT 757.950 795.600 760.050 796.050 ;
        RECT 715.950 794.400 760.050 795.600 ;
        RECT 715.950 793.950 718.050 794.400 ;
        RECT 757.950 793.950 760.050 794.400 ;
        RECT 823.950 795.600 826.050 796.050 ;
        RECT 829.950 795.600 832.050 796.050 ;
        RECT 823.950 794.400 832.050 795.600 ;
        RECT 823.950 793.950 826.050 794.400 ;
        RECT 829.950 793.950 832.050 794.400 ;
        RECT 853.950 795.600 856.050 796.050 ;
        RECT 868.950 795.600 871.050 796.050 ;
        RECT 853.950 794.400 871.050 795.600 ;
        RECT 853.950 793.950 856.050 794.400 ;
        RECT 868.950 793.950 871.050 794.400 ;
        RECT 877.950 795.600 880.050 796.050 ;
        RECT 895.950 795.600 898.050 796.050 ;
        RECT 961.950 795.600 964.050 796.050 ;
        RECT 877.950 794.400 898.050 795.600 ;
        RECT 877.950 793.950 880.050 794.400 ;
        RECT 895.950 793.950 898.050 794.400 ;
        RECT 953.400 794.400 964.050 795.600 ;
        RECT 151.950 792.600 154.050 793.050 ;
        RECT 250.950 792.600 253.050 793.050 ;
        RECT 301.950 792.600 304.050 793.050 ;
        RECT 151.950 791.400 304.050 792.600 ;
        RECT 151.950 790.950 154.050 791.400 ;
        RECT 250.950 790.950 253.050 791.400 ;
        RECT 301.950 790.950 304.050 791.400 ;
        RECT 346.950 792.600 349.050 793.050 ;
        RECT 358.950 792.600 361.050 792.900 ;
        RECT 475.950 792.600 478.050 793.050 ;
        RECT 346.950 791.400 478.050 792.600 ;
        RECT 346.950 790.950 349.050 791.400 ;
        RECT 358.950 790.800 361.050 791.400 ;
        RECT 475.950 790.950 478.050 791.400 ;
        RECT 535.950 792.600 538.050 793.050 ;
        RECT 604.950 792.600 607.050 793.050 ;
        RECT 535.950 791.400 607.050 792.600 ;
        RECT 535.950 790.950 538.050 791.400 ;
        RECT 604.950 790.950 607.050 791.400 ;
        RECT 610.950 792.600 613.050 793.050 ;
        RECT 700.950 792.600 703.050 793.050 ;
        RECT 610.950 791.400 703.050 792.600 ;
        RECT 610.950 790.950 613.050 791.400 ;
        RECT 700.950 790.950 703.050 791.400 ;
        RECT 706.950 792.600 709.050 792.900 ;
        RECT 760.950 792.600 763.050 793.050 ;
        RECT 706.950 791.400 763.050 792.600 ;
        RECT 706.950 790.800 709.050 791.400 ;
        RECT 760.950 790.950 763.050 791.400 ;
        RECT 925.950 792.600 928.050 793.050 ;
        RECT 953.400 792.600 954.600 794.400 ;
        RECT 961.950 793.950 964.050 794.400 ;
        RECT 925.950 791.400 954.600 792.600 ;
        RECT 955.950 792.600 958.050 793.050 ;
        RECT 997.950 792.600 1000.050 793.050 ;
        RECT 955.950 791.400 1000.050 792.600 ;
        RECT 925.950 790.950 928.050 791.400 ;
        RECT 955.950 790.950 958.050 791.400 ;
        RECT 997.950 790.950 1000.050 791.400 ;
        RECT 34.950 789.600 37.050 790.050 ;
        RECT 43.950 789.600 46.050 790.050 ;
        RECT 34.950 788.400 46.050 789.600 ;
        RECT 34.950 787.950 37.050 788.400 ;
        RECT 43.950 787.950 46.050 788.400 ;
        RECT 307.950 789.600 310.050 790.050 ;
        RECT 325.950 789.600 328.050 790.050 ;
        RECT 307.950 788.400 328.050 789.600 ;
        RECT 307.950 787.950 310.050 788.400 ;
        RECT 325.950 787.950 328.050 788.400 ;
        RECT 376.950 789.600 379.050 790.050 ;
        RECT 523.950 789.600 526.050 790.050 ;
        RECT 376.950 788.400 526.050 789.600 ;
        RECT 376.950 787.950 379.050 788.400 ;
        RECT 523.950 787.950 526.050 788.400 ;
        RECT 559.950 789.600 562.050 790.050 ;
        RECT 565.950 789.600 568.050 790.050 ;
        RECT 559.950 788.400 568.050 789.600 ;
        RECT 559.950 787.950 562.050 788.400 ;
        RECT 565.950 787.950 568.050 788.400 ;
        RECT 628.950 789.600 631.050 790.050 ;
        RECT 637.950 789.600 640.050 790.050 ;
        RECT 628.950 788.400 640.050 789.600 ;
        RECT 628.950 787.950 631.050 788.400 ;
        RECT 637.950 787.950 640.050 788.400 ;
        RECT 661.950 789.600 664.050 790.050 ;
        RECT 676.950 789.600 679.050 790.050 ;
        RECT 661.950 788.400 679.050 789.600 ;
        RECT 661.950 787.950 664.050 788.400 ;
        RECT 676.950 787.950 679.050 788.400 ;
        RECT 691.950 789.600 694.050 790.050 ;
        RECT 697.950 789.600 700.050 790.050 ;
        RECT 691.950 788.400 700.050 789.600 ;
        RECT 691.950 787.950 694.050 788.400 ;
        RECT 697.950 787.950 700.050 788.400 ;
        RECT 703.950 789.600 706.050 790.050 ;
        RECT 853.950 789.600 856.050 790.050 ;
        RECT 703.950 788.400 856.050 789.600 ;
        RECT 703.950 787.950 706.050 788.400 ;
        RECT 853.950 787.950 856.050 788.400 ;
        RECT 49.950 786.600 52.050 787.050 ;
        RECT 178.950 786.600 181.050 787.050 ;
        RECT 202.950 786.600 205.050 787.050 ;
        RECT 49.950 785.400 205.050 786.600 ;
        RECT 49.950 784.950 52.050 785.400 ;
        RECT 178.950 784.950 181.050 785.400 ;
        RECT 202.950 784.950 205.050 785.400 ;
        RECT 328.950 786.600 331.050 787.050 ;
        RECT 349.950 786.600 352.050 787.050 ;
        RECT 328.950 785.400 352.050 786.600 ;
        RECT 328.950 784.950 331.050 785.400 ;
        RECT 349.950 784.950 352.050 785.400 ;
        RECT 682.950 786.600 685.050 787.050 ;
        RECT 724.950 786.600 727.050 787.050 ;
        RECT 739.950 786.600 742.050 787.050 ;
        RECT 682.950 785.400 742.050 786.600 ;
        RECT 682.950 784.950 685.050 785.400 ;
        RECT 724.950 784.950 727.050 785.400 ;
        RECT 739.950 784.950 742.050 785.400 ;
        RECT 757.950 786.600 760.050 787.050 ;
        RECT 772.950 786.600 775.050 787.050 ;
        RECT 808.950 786.600 811.050 787.050 ;
        RECT 757.950 785.400 811.050 786.600 ;
        RECT 757.950 784.950 760.050 785.400 ;
        RECT 772.950 784.950 775.050 785.400 ;
        RECT 808.950 784.950 811.050 785.400 ;
        RECT 256.950 783.600 259.050 784.050 ;
        RECT 355.950 783.600 358.050 784.050 ;
        RECT 256.950 782.400 358.050 783.600 ;
        RECT 256.950 781.950 259.050 782.400 ;
        RECT 355.950 781.950 358.050 782.400 ;
        RECT 400.950 783.600 403.050 784.050 ;
        RECT 571.950 783.600 574.050 784.050 ;
        RECT 610.950 783.600 613.050 784.050 ;
        RECT 400.950 782.400 574.050 783.600 ;
        RECT 400.950 781.950 403.050 782.400 ;
        RECT 571.950 781.950 574.050 782.400 ;
        RECT 581.400 782.400 613.050 783.600 ;
        RECT 34.950 780.600 37.050 781.050 ;
        RECT 160.950 780.600 163.050 781.050 ;
        RECT 34.950 779.400 163.050 780.600 ;
        RECT 34.950 778.950 37.050 779.400 ;
        RECT 160.950 778.950 163.050 779.400 ;
        RECT 322.950 780.600 325.050 781.050 ;
        RECT 364.950 780.600 367.050 781.050 ;
        RECT 394.950 780.600 397.050 781.050 ;
        RECT 322.950 779.400 397.050 780.600 ;
        RECT 322.950 778.950 325.050 779.400 ;
        RECT 364.950 778.950 367.050 779.400 ;
        RECT 394.950 778.950 397.050 779.400 ;
        RECT 412.950 780.600 415.050 781.050 ;
        RECT 463.950 780.600 466.050 781.050 ;
        RECT 581.400 780.600 582.600 782.400 ;
        RECT 610.950 781.950 613.050 782.400 ;
        RECT 619.950 783.600 622.050 784.050 ;
        RECT 649.950 783.600 652.050 784.050 ;
        RECT 619.950 782.400 652.050 783.600 ;
        RECT 619.950 781.950 622.050 782.400 ;
        RECT 649.950 781.950 652.050 782.400 ;
        RECT 412.950 779.400 582.600 780.600 ;
        RECT 583.950 780.600 586.050 781.050 ;
        RECT 652.950 780.600 655.050 781.050 ;
        RECT 583.950 779.400 655.050 780.600 ;
        RECT 412.950 778.950 415.050 779.400 ;
        RECT 463.950 778.950 466.050 779.400 ;
        RECT 583.950 778.950 586.050 779.400 ;
        RECT 652.950 778.950 655.050 779.400 ;
        RECT 847.950 780.600 850.050 781.050 ;
        RECT 907.950 780.600 910.050 781.050 ;
        RECT 847.950 779.400 910.050 780.600 ;
        RECT 847.950 778.950 850.050 779.400 ;
        RECT 907.950 778.950 910.050 779.400 ;
        RECT 289.950 777.600 292.050 778.050 ;
        RECT 304.950 777.600 307.050 778.050 ;
        RECT 349.950 777.600 352.050 778.050 ;
        RECT 289.950 776.400 352.050 777.600 ;
        RECT 289.950 775.950 292.050 776.400 ;
        RECT 304.950 775.950 307.050 776.400 ;
        RECT 349.950 775.950 352.050 776.400 ;
        RECT 433.950 777.600 436.050 778.050 ;
        RECT 478.950 777.600 481.050 778.050 ;
        RECT 481.950 777.600 484.050 778.050 ;
        RECT 514.950 777.600 517.050 778.050 ;
        RECT 433.950 776.400 517.050 777.600 ;
        RECT 433.950 775.950 436.050 776.400 ;
        RECT 478.950 775.950 481.050 776.400 ;
        RECT 481.950 775.950 484.050 776.400 ;
        RECT 514.950 775.950 517.050 776.400 ;
        RECT 565.950 777.600 568.050 778.050 ;
        RECT 619.950 777.600 622.050 778.050 ;
        RECT 565.950 776.400 622.050 777.600 ;
        RECT 565.950 775.950 568.050 776.400 ;
        RECT 619.950 775.950 622.050 776.400 ;
        RECT 664.950 777.600 667.050 778.050 ;
        RECT 688.950 777.600 691.050 778.050 ;
        RECT 664.950 776.400 691.050 777.600 ;
        RECT 664.950 775.950 667.050 776.400 ;
        RECT 688.950 775.950 691.050 776.400 ;
        RECT 961.950 777.600 964.050 778.050 ;
        RECT 973.950 777.600 976.050 778.050 ;
        RECT 961.950 776.400 976.050 777.600 ;
        RECT 961.950 775.950 964.050 776.400 ;
        RECT 973.950 775.950 976.050 776.400 ;
        RECT 175.950 774.600 178.050 775.050 ;
        RECT 187.950 774.600 190.050 775.050 ;
        RECT 175.950 773.400 190.050 774.600 ;
        RECT 175.950 772.950 178.050 773.400 ;
        RECT 187.950 772.950 190.050 773.400 ;
        RECT 235.950 774.600 238.050 775.050 ;
        RECT 400.950 774.600 403.050 775.050 ;
        RECT 235.950 773.400 403.050 774.600 ;
        RECT 235.950 772.950 238.050 773.400 ;
        RECT 400.950 772.950 403.050 773.400 ;
        RECT 424.950 774.600 427.050 775.050 ;
        RECT 487.950 774.600 490.050 775.050 ;
        RECT 424.950 773.400 490.050 774.600 ;
        RECT 424.950 772.950 427.050 773.400 ;
        RECT 487.950 772.950 490.050 773.400 ;
        RECT 523.950 774.600 526.050 775.050 ;
        RECT 529.950 774.600 532.050 775.050 ;
        RECT 523.950 773.400 532.050 774.600 ;
        RECT 523.950 772.950 526.050 773.400 ;
        RECT 529.950 772.950 532.050 773.400 ;
        RECT 622.950 774.600 625.050 775.050 ;
        RECT 754.950 774.600 757.050 775.050 ;
        RECT 622.950 773.400 757.050 774.600 ;
        RECT 622.950 772.950 625.050 773.400 ;
        RECT 754.950 772.950 757.050 773.400 ;
        RECT 931.950 774.600 934.050 775.050 ;
        RECT 982.950 774.600 985.050 775.050 ;
        RECT 931.950 773.400 985.050 774.600 ;
        RECT 931.950 772.950 934.050 773.400 ;
        RECT 982.950 772.950 985.050 773.400 ;
        RECT 16.950 771.600 19.050 772.050 ;
        RECT 163.950 771.600 166.050 772.050 ;
        RECT 16.950 770.400 166.050 771.600 ;
        RECT 16.950 769.950 19.050 770.400 ;
        RECT 163.950 769.950 166.050 770.400 ;
        RECT 451.950 771.600 454.050 772.050 ;
        RECT 463.950 771.600 466.050 772.050 ;
        RECT 451.950 770.400 466.050 771.600 ;
        RECT 451.950 769.950 454.050 770.400 ;
        RECT 463.950 769.950 466.050 770.400 ;
        RECT 496.950 771.600 499.050 772.050 ;
        RECT 526.950 771.600 529.050 772.050 ;
        RECT 496.950 770.400 529.050 771.600 ;
        RECT 496.950 769.950 499.050 770.400 ;
        RECT 526.950 769.950 529.050 770.400 ;
        RECT 631.950 771.600 634.050 772.050 ;
        RECT 715.950 771.600 718.050 772.050 ;
        RECT 631.950 770.400 718.050 771.600 ;
        RECT 631.950 769.950 634.050 770.400 ;
        RECT 715.950 769.950 718.050 770.400 ;
        RECT 850.950 771.600 853.050 772.050 ;
        RECT 913.950 771.600 916.050 772.050 ;
        RECT 850.950 770.400 916.050 771.600 ;
        RECT 850.950 769.950 853.050 770.400 ;
        RECT 913.950 769.950 916.050 770.400 ;
        RECT 988.950 771.600 991.050 772.050 ;
        RECT 1006.950 771.600 1009.050 772.050 ;
        RECT 988.950 770.400 1009.050 771.600 ;
        RECT 988.950 769.950 991.050 770.400 ;
        RECT 1006.950 769.950 1009.050 770.400 ;
        RECT 241.950 768.600 244.050 769.050 ;
        RECT 253.950 768.600 256.050 769.050 ;
        RECT 241.950 767.400 256.050 768.600 ;
        RECT 241.950 766.950 244.050 767.400 ;
        RECT 253.950 766.950 256.050 767.400 ;
        RECT 325.950 768.600 328.050 769.050 ;
        RECT 337.950 768.600 340.050 769.050 ;
        RECT 325.950 767.400 340.050 768.600 ;
        RECT 325.950 766.950 328.050 767.400 ;
        RECT 337.950 766.950 340.050 767.400 ;
        RECT 487.950 768.600 490.050 769.050 ;
        RECT 535.950 768.600 538.050 769.050 ;
        RECT 550.950 768.600 553.050 769.050 ;
        RECT 586.950 768.600 589.050 769.050 ;
        RECT 622.950 768.600 625.050 769.050 ;
        RECT 487.950 767.400 625.050 768.600 ;
        RECT 487.950 766.950 490.050 767.400 ;
        RECT 535.950 766.950 538.050 767.400 ;
        RECT 550.950 766.950 553.050 767.400 ;
        RECT 586.950 766.950 589.050 767.400 ;
        RECT 622.950 766.950 625.050 767.400 ;
        RECT 649.950 768.600 652.050 769.050 ;
        RECT 670.950 768.600 673.050 769.050 ;
        RECT 649.950 767.400 673.050 768.600 ;
        RECT 649.950 766.950 652.050 767.400 ;
        RECT 670.950 766.950 673.050 767.400 ;
        RECT 712.950 768.600 715.050 769.050 ;
        RECT 736.950 768.600 739.050 769.050 ;
        RECT 712.950 767.400 739.050 768.600 ;
        RECT 712.950 766.950 715.050 767.400 ;
        RECT 736.950 766.950 739.050 767.400 ;
        RECT 748.950 768.600 751.050 769.050 ;
        RECT 787.800 768.600 789.900 769.050 ;
        RECT 748.950 767.400 789.900 768.600 ;
        RECT 748.950 766.950 751.050 767.400 ;
        RECT 787.800 766.950 789.900 767.400 ;
        RECT 790.950 768.600 793.050 769.050 ;
        RECT 814.950 768.600 817.050 769.050 ;
        RECT 790.950 767.400 817.050 768.600 ;
        RECT 790.950 766.950 793.050 767.400 ;
        RECT 814.950 766.950 817.050 767.400 ;
        RECT 937.950 768.600 940.050 769.050 ;
        RECT 967.950 768.600 970.050 769.050 ;
        RECT 937.950 767.400 970.050 768.600 ;
        RECT 937.950 766.950 940.050 767.400 ;
        RECT 967.950 766.950 970.050 767.400 ;
        RECT 991.950 768.600 994.050 769.050 ;
        RECT 997.950 768.600 1000.050 769.050 ;
        RECT 991.950 767.400 1000.050 768.600 ;
        RECT 991.950 766.950 994.050 767.400 ;
        RECT 997.950 766.950 1000.050 767.400 ;
        RECT 190.950 765.600 193.050 766.050 ;
        RECT 205.950 765.600 208.050 766.050 ;
        RECT 271.950 765.600 274.050 766.050 ;
        RECT 190.950 764.400 274.050 765.600 ;
        RECT 190.950 763.950 193.050 764.400 ;
        RECT 205.950 763.950 208.050 764.400 ;
        RECT 271.950 763.950 274.050 764.400 ;
        RECT 415.950 765.600 418.050 766.050 ;
        RECT 421.950 765.600 424.050 766.050 ;
        RECT 415.950 764.400 424.050 765.600 ;
        RECT 415.950 763.950 418.050 764.400 ;
        RECT 421.950 763.950 424.050 764.400 ;
        RECT 472.950 765.600 475.050 766.050 ;
        RECT 493.950 765.600 496.050 766.050 ;
        RECT 472.950 764.400 496.050 765.600 ;
        RECT 472.950 763.950 475.050 764.400 ;
        RECT 493.950 763.950 496.050 764.400 ;
        RECT 682.950 765.600 685.050 766.050 ;
        RECT 697.950 765.600 700.050 766.200 ;
        RECT 682.950 764.400 700.050 765.600 ;
        RECT 682.950 763.950 685.050 764.400 ;
        RECT 697.950 764.100 700.050 764.400 ;
        RECT 781.950 765.600 784.050 766.050 ;
        RECT 838.950 765.600 841.050 766.050 ;
        RECT 853.950 765.600 856.050 766.050 ;
        RECT 781.950 764.400 856.050 765.600 ;
        RECT 781.950 763.950 784.050 764.400 ;
        RECT 838.950 763.950 841.050 764.400 ;
        RECT 853.950 763.950 856.050 764.400 ;
        RECT 859.950 765.600 862.050 766.050 ;
        RECT 868.950 765.600 871.050 766.050 ;
        RECT 859.950 764.400 871.050 765.600 ;
        RECT 859.950 763.950 862.050 764.400 ;
        RECT 868.950 763.950 871.050 764.400 ;
        RECT 10.950 762.600 15.000 763.050 ;
        RECT 22.950 762.750 25.050 763.200 ;
        RECT 28.950 762.750 31.050 763.200 ;
        RECT 10.950 760.950 15.600 762.600 ;
        RECT 22.950 761.550 31.050 762.750 ;
        RECT 22.950 761.100 25.050 761.550 ;
        RECT 28.950 761.100 31.050 761.550 ;
        RECT 52.950 762.750 55.050 763.200 ;
        RECT 58.950 762.750 61.050 763.200 ;
        RECT 52.950 761.550 61.050 762.750 ;
        RECT 52.950 761.100 55.050 761.550 ;
        RECT 58.950 761.100 61.050 761.550 ;
        RECT 64.950 762.600 67.050 763.200 ;
        RECT 94.950 762.600 97.050 763.200 ;
        RECT 64.950 761.400 97.050 762.600 ;
        RECT 64.950 761.100 67.050 761.400 ;
        RECT 94.950 761.100 97.050 761.400 ;
        RECT 100.950 762.600 103.050 763.050 ;
        RECT 121.950 762.600 124.050 763.200 ;
        RECT 139.950 762.600 142.050 763.200 ;
        RECT 100.950 761.400 142.050 762.600 ;
        RECT 100.950 760.950 103.050 761.400 ;
        RECT 121.950 761.100 124.050 761.400 ;
        RECT 139.950 761.100 142.050 761.400 ;
        RECT 145.950 761.100 148.050 763.200 ;
        RECT 184.950 761.100 187.050 763.200 ;
        RECT 241.950 762.600 244.050 763.200 ;
        RECT 250.950 762.600 253.050 763.050 ;
        RECT 241.950 761.400 253.050 762.600 ;
        RECT 241.950 761.100 244.050 761.400 ;
        RECT 14.400 756.900 15.600 760.950 ;
        RECT 13.950 754.800 16.050 756.900 ;
        RECT 19.950 756.600 22.050 756.900 ;
        RECT 31.950 756.600 34.050 757.050 ;
        RECT 19.950 755.400 34.050 756.600 ;
        RECT 19.950 754.800 22.050 755.400 ;
        RECT 31.950 754.950 34.050 755.400 ;
        RECT 46.950 756.600 49.050 757.050 ;
        RECT 52.950 756.600 55.050 757.050 ;
        RECT 79.950 756.600 82.050 756.900 ;
        RECT 46.950 755.400 82.050 756.600 ;
        RECT 46.950 754.950 49.050 755.400 ;
        RECT 52.950 754.950 55.050 755.400 ;
        RECT 79.950 754.800 82.050 755.400 ;
        RECT 115.950 756.600 118.050 756.900 ;
        RECT 146.400 756.600 147.600 761.100 ;
        RECT 185.400 759.600 186.600 761.100 ;
        RECT 250.950 760.950 253.050 761.400 ;
        RECT 277.950 762.750 280.050 763.200 ;
        RECT 286.950 762.750 289.050 763.200 ;
        RECT 277.950 761.550 289.050 762.750 ;
        RECT 277.950 761.100 280.050 761.550 ;
        RECT 286.950 761.100 289.050 761.550 ;
        RECT 292.950 762.750 295.050 763.200 ;
        RECT 298.950 762.750 301.050 763.200 ;
        RECT 292.950 761.550 301.050 762.750 ;
        RECT 292.950 761.100 295.050 761.550 ;
        RECT 298.950 761.100 301.050 761.550 ;
        RECT 337.950 760.950 340.050 763.050 ;
        RECT 343.950 762.750 346.050 763.200 ;
        RECT 352.950 762.750 355.050 763.200 ;
        RECT 343.950 761.550 355.050 762.750 ;
        RECT 343.950 761.100 346.050 761.550 ;
        RECT 352.950 761.100 355.050 761.550 ;
        RECT 382.950 761.100 385.050 763.200 ;
        RECT 388.950 762.600 391.050 763.200 ;
        RECT 403.950 762.600 406.050 763.200 ;
        RECT 388.950 761.400 406.050 762.600 ;
        RECT 388.950 761.100 391.050 761.400 ;
        RECT 403.950 761.100 406.050 761.400 ;
        RECT 430.950 762.750 433.050 763.200 ;
        RECT 436.950 762.750 439.050 763.200 ;
        RECT 430.950 762.600 439.050 762.750 ;
        RECT 460.950 762.600 463.050 763.200 ;
        RECT 430.950 761.550 463.050 762.600 ;
        RECT 430.950 761.100 433.050 761.550 ;
        RECT 436.950 761.400 463.050 761.550 ;
        RECT 436.950 761.100 439.050 761.400 ;
        RECT 460.950 761.100 463.050 761.400 ;
        RECT 490.950 762.600 493.050 763.050 ;
        RECT 502.950 762.600 505.050 763.200 ;
        RECT 490.950 761.400 505.050 762.600 ;
        RECT 226.950 759.600 229.050 760.050 ;
        RECT 185.400 758.400 229.050 759.600 ;
        RECT 226.950 757.950 229.050 758.400 ;
        RECT 115.950 755.400 147.600 756.600 ;
        RECT 166.950 756.600 169.050 756.900 ;
        RECT 175.950 756.600 178.050 757.050 ;
        RECT 166.950 755.400 178.050 756.600 ;
        RECT 115.950 754.800 118.050 755.400 ;
        RECT 166.950 754.800 169.050 755.400 ;
        RECT 175.950 754.950 178.050 755.400 ;
        RECT 238.950 756.450 241.050 756.900 ;
        RECT 247.950 756.450 250.050 757.050 ;
        RECT 253.950 756.450 256.050 756.900 ;
        RECT 238.950 755.250 256.050 756.450 ;
        RECT 238.950 754.800 241.050 755.250 ;
        RECT 247.950 754.950 250.050 755.250 ;
        RECT 253.950 754.800 256.050 755.250 ;
        RECT 283.950 756.450 286.050 756.900 ;
        RECT 304.800 756.450 306.900 756.900 ;
        RECT 313.950 756.600 316.050 756.900 ;
        RECT 283.950 755.250 306.900 756.450 ;
        RECT 308.400 756.000 316.050 756.600 ;
        RECT 283.950 754.800 286.050 755.250 ;
        RECT 304.800 754.800 306.900 755.250 ;
        RECT 307.950 755.400 316.050 756.000 ;
        RECT 16.950 753.600 19.050 754.050 ;
        RECT 34.950 753.600 37.050 754.050 ;
        RECT 16.950 752.400 37.050 753.600 ;
        RECT 16.950 751.950 19.050 752.400 ;
        RECT 34.950 751.950 37.050 752.400 ;
        RECT 43.950 753.600 46.050 754.050 ;
        RECT 49.950 753.600 52.050 754.050 ;
        RECT 43.950 752.400 52.050 753.600 ;
        RECT 43.950 751.950 46.050 752.400 ;
        RECT 49.950 751.950 52.050 752.400 ;
        RECT 307.950 751.950 310.050 755.400 ;
        RECT 313.950 754.800 316.050 755.400 ;
        RECT 331.950 756.600 334.050 757.050 ;
        RECT 338.400 756.600 339.600 760.950 ;
        RECT 331.950 755.400 339.600 756.600 ;
        RECT 349.950 756.600 352.050 757.050 ;
        RECT 361.950 756.600 364.050 756.900 ;
        RECT 349.950 755.400 364.050 756.600 ;
        RECT 331.950 754.950 334.050 755.400 ;
        RECT 349.950 754.950 352.050 755.400 ;
        RECT 361.950 754.800 364.050 755.400 ;
        RECT 373.950 756.450 376.050 756.900 ;
        RECT 379.950 756.450 382.050 756.900 ;
        RECT 373.950 755.250 382.050 756.450 ;
        RECT 373.950 754.800 376.050 755.250 ;
        RECT 379.950 754.800 382.050 755.250 ;
        RECT 383.400 754.050 384.600 761.100 ;
        RECT 490.950 760.950 493.050 761.400 ;
        RECT 502.950 761.100 505.050 761.400 ;
        RECT 538.950 762.750 541.050 763.200 ;
        RECT 544.950 762.750 547.050 763.200 ;
        RECT 538.950 761.550 547.050 762.750 ;
        RECT 538.950 761.100 541.050 761.550 ;
        RECT 544.950 761.100 547.050 761.550 ;
        RECT 556.950 762.750 559.050 763.200 ;
        RECT 565.950 762.750 568.050 763.200 ;
        RECT 556.950 761.550 568.050 762.750 ;
        RECT 556.950 761.100 559.050 761.550 ;
        RECT 565.950 761.100 568.050 761.550 ;
        RECT 571.950 762.600 574.050 763.200 ;
        RECT 595.950 762.600 598.050 763.200 ;
        RECT 571.950 761.400 598.050 762.600 ;
        RECT 571.950 761.100 574.050 761.400 ;
        RECT 595.950 761.100 598.050 761.400 ;
        RECT 613.950 762.600 616.050 763.200 ;
        RECT 643.950 762.600 646.050 763.200 ;
        RECT 613.950 761.400 646.050 762.600 ;
        RECT 613.950 761.100 616.050 761.400 ;
        RECT 643.950 761.100 646.050 761.400 ;
        RECT 649.950 762.600 652.050 763.200 ;
        RECT 676.950 762.600 679.050 763.200 ;
        RECT 697.950 762.600 700.050 763.050 ;
        RECT 649.950 761.400 700.050 762.600 ;
        RECT 649.950 761.100 652.050 761.400 ;
        RECT 676.950 761.100 679.050 761.400 ;
        RECT 697.950 760.950 700.050 761.400 ;
        RECT 703.950 762.750 706.050 763.200 ;
        RECT 712.950 762.750 715.050 763.200 ;
        RECT 703.950 761.550 715.050 762.750 ;
        RECT 703.950 761.100 706.050 761.550 ;
        RECT 712.950 761.100 715.050 761.550 ;
        RECT 718.950 762.600 721.050 763.200 ;
        RECT 733.950 762.600 736.050 763.050 ;
        RECT 718.950 761.400 736.050 762.600 ;
        RECT 718.950 761.100 721.050 761.400 ;
        RECT 733.950 760.950 736.050 761.400 ;
        RECT 763.950 762.600 766.050 763.200 ;
        RECT 796.950 762.750 799.050 763.200 ;
        RECT 802.950 762.750 805.050 763.200 ;
        RECT 796.950 762.600 805.050 762.750 ;
        RECT 820.950 762.600 823.050 763.200 ;
        RECT 763.950 761.400 789.600 762.600 ;
        RECT 763.950 761.100 766.050 761.400 ;
        RECT 394.950 756.450 397.050 756.900 ;
        RECT 406.950 756.450 409.050 756.900 ;
        RECT 394.950 755.250 409.050 756.450 ;
        RECT 394.950 754.800 397.050 755.250 ;
        RECT 406.950 754.800 409.050 755.250 ;
        RECT 424.950 756.450 427.050 756.900 ;
        RECT 442.950 756.450 445.050 756.900 ;
        RECT 424.950 755.250 445.050 756.450 ;
        RECT 424.950 754.800 427.050 755.250 ;
        RECT 442.950 754.800 445.050 755.250 ;
        RECT 547.950 756.600 550.050 756.900 ;
        RECT 556.800 756.600 558.900 757.050 ;
        RECT 547.950 755.400 558.900 756.600 ;
        RECT 547.950 754.800 550.050 755.400 ;
        RECT 556.800 754.950 558.900 755.400 ;
        RECT 559.950 756.600 562.050 757.050 ;
        RECT 568.950 756.600 571.050 756.900 ;
        RECT 559.950 755.400 571.050 756.600 ;
        RECT 559.950 754.950 562.050 755.400 ;
        RECT 568.950 754.800 571.050 755.400 ;
        RECT 607.950 756.600 610.050 757.050 ;
        RECT 646.950 756.600 649.050 756.900 ;
        RECT 673.950 756.600 676.050 756.900 ;
        RECT 607.950 755.400 645.600 756.600 ;
        RECT 607.950 754.950 610.050 755.400 ;
        RECT 382.950 751.950 385.050 754.050 ;
        RECT 535.950 753.600 538.050 754.050 ;
        RECT 544.950 753.600 547.050 754.050 ;
        RECT 535.950 752.400 547.050 753.600 ;
        RECT 535.950 751.950 538.050 752.400 ;
        RECT 544.950 751.950 547.050 752.400 ;
        RECT 628.950 753.600 631.050 754.050 ;
        RECT 640.950 753.600 643.050 754.050 ;
        RECT 628.950 752.400 643.050 753.600 ;
        RECT 644.400 753.600 645.600 755.400 ;
        RECT 646.950 755.400 676.050 756.600 ;
        RECT 646.950 754.800 649.050 755.400 ;
        RECT 673.950 754.800 676.050 755.400 ;
        RECT 721.950 756.600 724.050 756.900 ;
        RECT 733.950 756.600 736.050 757.050 ;
        RECT 721.950 755.400 736.050 756.600 ;
        RECT 721.950 754.800 724.050 755.400 ;
        RECT 733.950 754.950 736.050 755.400 ;
        RECT 772.950 756.600 775.050 756.900 ;
        RECT 781.950 756.600 784.050 757.050 ;
        RECT 788.400 756.900 789.600 761.400 ;
        RECT 796.950 761.550 823.050 762.600 ;
        RECT 796.950 761.100 799.050 761.550 ;
        RECT 802.950 761.400 823.050 761.550 ;
        RECT 802.950 761.100 805.050 761.400 ;
        RECT 820.950 761.100 823.050 761.400 ;
        RECT 844.950 761.100 847.050 763.200 ;
        RECT 845.400 759.600 846.600 761.100 ;
        RECT 883.950 760.950 886.050 763.050 ;
        RECT 895.950 761.100 898.050 763.200 ;
        RECT 824.400 758.400 846.600 759.600 ;
        RECT 824.400 756.900 825.600 758.400 ;
        RECT 772.950 755.400 784.050 756.600 ;
        RECT 772.950 754.800 775.050 755.400 ;
        RECT 781.950 754.950 784.050 755.400 ;
        RECT 787.950 754.800 790.050 756.900 ;
        RECT 793.950 756.600 796.050 756.900 ;
        RECT 793.950 756.000 801.600 756.600 ;
        RECT 808.950 756.450 811.050 756.900 ;
        RECT 817.950 756.450 820.050 756.900 ;
        RECT 793.950 755.400 802.050 756.000 ;
        RECT 793.950 754.800 796.050 755.400 ;
        RECT 694.950 753.600 697.050 754.050 ;
        RECT 644.400 752.400 697.050 753.600 ;
        RECT 628.950 751.950 631.050 752.400 ;
        RECT 640.950 751.950 643.050 752.400 ;
        RECT 694.950 751.950 697.050 752.400 ;
        RECT 730.950 753.600 733.050 754.050 ;
        RECT 739.950 753.600 742.050 754.050 ;
        RECT 730.950 752.400 742.050 753.600 ;
        RECT 730.950 751.950 733.050 752.400 ;
        RECT 739.950 751.950 742.050 752.400 ;
        RECT 799.950 751.950 802.050 755.400 ;
        RECT 808.950 755.250 820.050 756.450 ;
        RECT 808.950 754.800 811.050 755.250 ;
        RECT 817.950 754.800 820.050 755.250 ;
        RECT 823.950 754.800 826.050 756.900 ;
        RECT 853.950 756.450 856.050 756.900 ;
        RECT 862.950 756.450 865.050 756.900 ;
        RECT 853.950 755.250 865.050 756.450 ;
        RECT 884.400 756.600 885.600 760.950 ;
        RECT 896.400 757.050 897.600 761.100 ;
        RECT 919.950 760.950 922.050 763.050 ;
        RECT 946.950 762.750 949.050 763.200 ;
        RECT 955.950 762.750 958.050 763.200 ;
        RECT 946.950 761.550 958.050 762.750 ;
        RECT 946.950 761.100 949.050 761.550 ;
        RECT 955.950 761.100 958.050 761.550 ;
        RECT 991.950 761.100 994.050 763.200 ;
        RECT 907.950 759.600 910.050 760.050 ;
        RECT 920.400 759.600 921.600 760.950 ;
        RECT 907.950 758.400 921.600 759.600 ;
        RECT 907.950 757.950 910.050 758.400 ;
        RECT 886.950 756.600 889.050 756.900 ;
        RECT 884.400 755.400 889.050 756.600 ;
        RECT 896.400 755.400 901.050 757.050 ;
        RECT 853.950 754.800 856.050 755.250 ;
        RECT 862.950 754.800 865.050 755.250 ;
        RECT 886.950 754.800 889.050 755.400 ;
        RECT 897.000 754.950 901.050 755.400 ;
        RECT 904.950 756.600 907.050 757.050 ;
        RECT 916.950 756.600 919.050 756.900 ;
        RECT 904.950 755.400 919.050 756.600 ;
        RECT 904.950 754.950 907.050 755.400 ;
        RECT 916.950 754.800 919.050 755.400 ;
        RECT 928.950 756.450 931.050 756.900 ;
        RECT 943.950 756.450 946.050 756.900 ;
        RECT 928.950 755.250 946.050 756.450 ;
        RECT 992.400 756.600 993.600 761.100 ;
        RECT 1003.950 756.600 1006.050 757.050 ;
        RECT 992.400 755.400 1006.050 756.600 ;
        RECT 928.950 754.800 931.050 755.250 ;
        RECT 943.950 754.800 946.050 755.250 ;
        RECT 1003.950 754.950 1006.050 755.400 ;
        RECT 943.950 753.600 946.050 754.050 ;
        RECT 970.950 753.600 973.050 754.050 ;
        RECT 943.950 752.400 973.050 753.600 ;
        RECT 943.950 751.950 946.050 752.400 ;
        RECT 970.950 751.950 973.050 752.400 ;
        RECT 76.950 750.600 79.050 751.050 ;
        RECT 85.950 750.600 88.050 751.050 ;
        RECT 76.950 749.400 88.050 750.600 ;
        RECT 76.950 748.950 79.050 749.400 ;
        RECT 85.950 748.950 88.050 749.400 ;
        RECT 97.950 750.600 100.050 751.050 ;
        RECT 214.950 750.600 217.050 751.050 ;
        RECT 97.950 749.400 217.050 750.600 ;
        RECT 97.950 748.950 100.050 749.400 ;
        RECT 214.950 748.950 217.050 749.400 ;
        RECT 265.950 750.600 268.050 751.050 ;
        RECT 277.950 750.600 280.050 751.050 ;
        RECT 334.950 750.600 337.050 751.050 ;
        RECT 265.950 749.400 337.050 750.600 ;
        RECT 265.950 748.950 268.050 749.400 ;
        RECT 277.950 748.950 280.050 749.400 ;
        RECT 334.950 748.950 337.050 749.400 ;
        RECT 400.950 750.600 403.050 751.050 ;
        RECT 433.950 750.600 436.050 751.050 ;
        RECT 400.950 749.400 436.050 750.600 ;
        RECT 400.950 748.950 403.050 749.400 ;
        RECT 433.950 748.950 436.050 749.400 ;
        RECT 667.950 750.600 670.050 751.050 ;
        RECT 676.950 750.600 679.050 751.050 ;
        RECT 667.950 749.400 679.050 750.600 ;
        RECT 667.950 748.950 670.050 749.400 ;
        RECT 676.950 748.950 679.050 749.400 ;
        RECT 748.950 750.600 751.050 751.050 ;
        RECT 802.950 750.600 805.050 751.050 ;
        RECT 748.950 749.400 805.050 750.600 ;
        RECT 748.950 748.950 751.050 749.400 ;
        RECT 802.950 748.950 805.050 749.400 ;
        RECT 919.950 750.600 922.050 751.050 ;
        RECT 925.950 750.600 928.050 751.050 ;
        RECT 919.950 749.400 928.050 750.600 ;
        RECT 919.950 748.950 922.050 749.400 ;
        RECT 925.950 748.950 928.050 749.400 ;
        RECT 949.950 750.600 952.050 751.050 ;
        RECT 964.950 750.600 967.050 751.050 ;
        RECT 949.950 749.400 967.050 750.600 ;
        RECT 949.950 748.950 952.050 749.400 ;
        RECT 964.950 748.950 967.050 749.400 ;
        RECT 976.950 750.600 979.050 751.050 ;
        RECT 1000.950 750.600 1003.050 751.050 ;
        RECT 976.950 749.400 1003.050 750.600 ;
        RECT 976.950 748.950 979.050 749.400 ;
        RECT 1000.950 748.950 1003.050 749.400 ;
        RECT 271.950 747.600 274.050 748.050 ;
        RECT 289.950 747.600 292.050 748.050 ;
        RECT 271.950 746.400 292.050 747.600 ;
        RECT 271.950 745.950 274.050 746.400 ;
        RECT 289.950 745.950 292.050 746.400 ;
        RECT 301.950 747.600 304.050 748.050 ;
        RECT 331.950 747.600 334.050 748.050 ;
        RECT 301.950 746.400 334.050 747.600 ;
        RECT 301.950 745.950 304.050 746.400 ;
        RECT 331.950 745.950 334.050 746.400 ;
        RECT 436.950 747.600 439.050 748.050 ;
        RECT 460.950 747.600 463.050 748.050 ;
        RECT 436.950 746.400 463.050 747.600 ;
        RECT 436.950 745.950 439.050 746.400 ;
        RECT 460.950 745.950 463.050 746.400 ;
        RECT 493.950 747.600 496.050 748.050 ;
        RECT 538.950 747.600 541.050 748.050 ;
        RECT 493.950 746.400 541.050 747.600 ;
        RECT 493.950 745.950 496.050 746.400 ;
        RECT 538.950 745.950 541.050 746.400 ;
        RECT 556.950 747.600 559.050 748.050 ;
        RECT 568.950 747.600 571.050 748.050 ;
        RECT 574.950 747.600 577.050 748.050 ;
        RECT 556.950 746.400 577.050 747.600 ;
        RECT 556.950 745.950 559.050 746.400 ;
        RECT 568.950 745.950 571.050 746.400 ;
        RECT 574.950 745.950 577.050 746.400 ;
        RECT 724.950 747.600 727.050 748.050 ;
        RECT 745.950 747.600 748.050 748.050 ;
        RECT 724.950 746.400 748.050 747.600 ;
        RECT 724.950 745.950 727.050 746.400 ;
        RECT 745.950 745.950 748.050 746.400 ;
        RECT 805.950 747.600 808.050 748.050 ;
        RECT 901.950 747.600 904.050 748.050 ;
        RECT 922.950 747.600 925.050 748.050 ;
        RECT 805.950 746.400 925.050 747.600 ;
        RECT 805.950 745.950 808.050 746.400 ;
        RECT 901.950 745.950 904.050 746.400 ;
        RECT 922.950 745.950 925.050 746.400 ;
        RECT 382.950 744.600 385.050 745.050 ;
        RECT 394.950 744.600 397.050 745.050 ;
        RECT 418.950 744.600 421.050 745.050 ;
        RECT 382.950 743.400 421.050 744.600 ;
        RECT 539.400 744.600 540.600 745.950 ;
        RECT 598.950 744.600 601.050 745.050 ;
        RECT 616.950 744.600 619.050 745.050 ;
        RECT 539.400 743.400 619.050 744.600 ;
        RECT 382.950 742.950 385.050 743.400 ;
        RECT 394.950 742.950 397.050 743.400 ;
        RECT 418.950 742.950 421.050 743.400 ;
        RECT 598.950 742.950 601.050 743.400 ;
        RECT 616.950 742.950 619.050 743.400 ;
        RECT 733.950 744.600 736.050 745.050 ;
        RECT 766.950 744.600 769.050 745.050 ;
        RECT 733.950 743.400 769.050 744.600 ;
        RECT 733.950 742.950 736.050 743.400 ;
        RECT 766.950 742.950 769.050 743.400 ;
        RECT 952.950 744.600 955.050 745.050 ;
        RECT 973.950 744.600 976.050 745.050 ;
        RECT 952.950 743.400 976.050 744.600 ;
        RECT 952.950 742.950 955.050 743.400 ;
        RECT 973.950 742.950 976.050 743.400 ;
        RECT 982.950 744.600 985.050 745.050 ;
        RECT 1000.950 744.600 1003.050 745.050 ;
        RECT 982.950 743.400 1003.050 744.600 ;
        RECT 982.950 742.950 985.050 743.400 ;
        RECT 1000.950 742.950 1003.050 743.400 ;
        RECT 106.950 741.600 109.050 742.050 ;
        RECT 127.950 741.600 130.050 742.050 ;
        RECT 148.950 741.600 151.050 742.050 ;
        RECT 187.950 741.600 190.050 742.050 ;
        RECT 106.950 740.400 190.050 741.600 ;
        RECT 106.950 739.950 109.050 740.400 ;
        RECT 127.950 739.950 130.050 740.400 ;
        RECT 148.950 739.950 151.050 740.400 ;
        RECT 187.950 739.950 190.050 740.400 ;
        RECT 226.950 741.600 229.050 742.050 ;
        RECT 280.950 741.600 283.050 742.050 ;
        RECT 226.950 740.400 283.050 741.600 ;
        RECT 226.950 739.950 229.050 740.400 ;
        RECT 280.950 739.950 283.050 740.400 ;
        RECT 298.950 741.600 301.050 742.050 ;
        RECT 346.950 741.600 349.050 742.050 ;
        RECT 298.950 740.400 349.050 741.600 ;
        RECT 298.950 739.950 301.050 740.400 ;
        RECT 346.950 739.950 349.050 740.400 ;
        RECT 514.950 741.600 517.050 742.050 ;
        RECT 547.950 741.600 550.050 742.050 ;
        RECT 514.950 740.400 550.050 741.600 ;
        RECT 514.950 739.950 517.050 740.400 ;
        RECT 547.950 739.950 550.050 740.400 ;
        RECT 574.950 741.600 577.050 742.050 ;
        RECT 607.950 741.600 610.050 742.050 ;
        RECT 574.950 740.400 610.050 741.600 ;
        RECT 574.950 739.950 577.050 740.400 ;
        RECT 607.950 739.950 610.050 740.400 ;
        RECT 655.950 741.600 658.050 742.050 ;
        RECT 682.950 741.600 685.050 742.050 ;
        RECT 655.950 740.400 685.050 741.600 ;
        RECT 655.950 739.950 658.050 740.400 ;
        RECT 682.950 739.950 685.050 740.400 ;
        RECT 709.950 741.600 712.050 742.050 ;
        RECT 724.950 741.600 727.050 742.050 ;
        RECT 709.950 740.400 727.050 741.600 ;
        RECT 709.950 739.950 712.050 740.400 ;
        RECT 724.950 739.950 727.050 740.400 ;
        RECT 925.950 741.600 928.050 742.050 ;
        RECT 949.950 741.600 952.050 742.050 ;
        RECT 925.950 740.400 952.050 741.600 ;
        RECT 925.950 739.950 928.050 740.400 ;
        RECT 949.950 739.950 952.050 740.400 ;
        RECT 61.950 738.600 64.050 739.050 ;
        RECT 109.950 738.600 112.050 739.050 ;
        RECT 61.950 737.400 112.050 738.600 ;
        RECT 61.950 736.950 64.050 737.400 ;
        RECT 109.950 736.950 112.050 737.400 ;
        RECT 148.950 738.600 151.050 738.900 ;
        RECT 220.950 738.600 223.050 739.050 ;
        RECT 148.950 737.400 223.050 738.600 ;
        RECT 148.950 736.800 151.050 737.400 ;
        RECT 220.950 736.950 223.050 737.400 ;
        RECT 259.950 738.600 262.050 739.050 ;
        RECT 283.950 738.600 286.050 739.050 ;
        RECT 259.950 737.400 286.050 738.600 ;
        RECT 259.950 736.950 262.050 737.400 ;
        RECT 283.950 736.950 286.050 737.400 ;
        RECT 367.950 738.600 370.050 739.050 ;
        RECT 391.950 738.600 394.050 739.050 ;
        RECT 367.950 737.400 394.050 738.600 ;
        RECT 367.950 736.950 370.050 737.400 ;
        RECT 391.950 736.950 394.050 737.400 ;
        RECT 415.950 738.600 418.050 739.050 ;
        RECT 424.950 738.600 427.050 739.050 ;
        RECT 415.950 737.400 427.050 738.600 ;
        RECT 415.950 736.950 418.050 737.400 ;
        RECT 424.950 736.950 427.050 737.400 ;
        RECT 730.950 738.600 733.050 739.050 ;
        RECT 757.950 738.600 760.050 739.050 ;
        RECT 730.950 737.400 760.050 738.600 ;
        RECT 730.950 736.950 733.050 737.400 ;
        RECT 757.950 736.950 760.050 737.400 ;
        RECT 772.950 738.600 775.050 739.050 ;
        RECT 850.950 738.600 853.050 739.050 ;
        RECT 772.950 737.400 853.050 738.600 ;
        RECT 772.950 736.950 775.050 737.400 ;
        RECT 850.950 736.950 853.050 737.400 ;
        RECT 856.950 738.600 859.050 739.050 ;
        RECT 901.950 738.600 904.050 739.050 ;
        RECT 856.950 737.400 904.050 738.600 ;
        RECT 856.950 736.950 859.050 737.400 ;
        RECT 901.950 736.950 904.050 737.400 ;
        RECT 937.950 738.600 940.050 739.050 ;
        RECT 955.950 738.600 958.050 739.050 ;
        RECT 937.950 737.400 958.050 738.600 ;
        RECT 937.950 736.950 940.050 737.400 ;
        RECT 955.950 736.950 958.050 737.400 ;
        RECT 961.950 738.600 964.050 739.050 ;
        RECT 976.950 738.600 979.050 739.050 ;
        RECT 961.950 737.400 979.050 738.600 ;
        RECT 961.950 736.950 964.050 737.400 ;
        RECT 976.950 736.950 979.050 737.400 ;
        RECT 85.950 735.600 88.050 736.050 ;
        RECT 100.950 735.600 103.050 736.050 ;
        RECT 85.950 734.400 103.050 735.600 ;
        RECT 85.950 733.950 88.050 734.400 ;
        RECT 100.950 733.950 103.050 734.400 ;
        RECT 184.950 735.600 187.050 736.050 ;
        RECT 196.950 735.600 199.050 736.050 ;
        RECT 184.950 734.400 199.050 735.600 ;
        RECT 184.950 733.950 187.050 734.400 ;
        RECT 196.950 733.950 199.050 734.400 ;
        RECT 259.950 735.600 262.050 735.900 ;
        RECT 271.950 735.600 274.050 736.050 ;
        RECT 259.950 734.400 274.050 735.600 ;
        RECT 259.950 733.800 262.050 734.400 ;
        RECT 271.950 733.950 274.050 734.400 ;
        RECT 295.950 735.600 298.050 736.050 ;
        RECT 343.800 735.600 345.900 736.050 ;
        RECT 295.950 734.400 345.900 735.600 ;
        RECT 295.950 733.950 298.050 734.400 ;
        RECT 343.800 733.950 345.900 734.400 ;
        RECT 346.950 735.600 349.050 736.050 ;
        RECT 430.950 735.600 433.050 736.050 ;
        RECT 346.950 734.400 433.050 735.600 ;
        RECT 346.950 733.950 349.050 734.400 ;
        RECT 430.950 733.950 433.050 734.400 ;
        RECT 592.950 735.600 595.050 736.050 ;
        RECT 604.950 735.600 607.050 736.050 ;
        RECT 592.950 734.400 607.050 735.600 ;
        RECT 592.950 733.950 595.050 734.400 ;
        RECT 604.950 733.950 607.050 734.400 ;
        RECT 610.950 735.600 613.050 736.050 ;
        RECT 616.950 735.600 619.050 736.050 ;
        RECT 610.950 734.400 619.050 735.600 ;
        RECT 610.950 733.950 613.050 734.400 ;
        RECT 616.950 733.950 619.050 734.400 ;
        RECT 790.950 735.600 793.050 736.050 ;
        RECT 814.950 735.600 817.050 736.050 ;
        RECT 790.950 734.400 817.050 735.600 ;
        RECT 790.950 733.950 793.050 734.400 ;
        RECT 814.950 733.950 817.050 734.400 ;
        RECT 931.950 735.600 934.050 736.050 ;
        RECT 949.950 735.600 952.050 736.050 ;
        RECT 931.950 734.400 952.050 735.600 ;
        RECT 931.950 733.950 934.050 734.400 ;
        RECT 949.950 733.950 952.050 734.400 ;
        RECT 958.950 735.600 961.050 736.050 ;
        RECT 979.800 735.600 981.900 736.050 ;
        RECT 958.950 734.400 981.900 735.600 ;
        RECT 958.950 733.950 961.050 734.400 ;
        RECT 979.800 733.950 981.900 734.400 ;
        RECT 982.950 735.600 985.050 736.050 ;
        RECT 994.950 735.600 997.050 736.050 ;
        RECT 982.950 734.400 997.050 735.600 ;
        RECT 982.950 733.950 985.050 734.400 ;
        RECT 994.950 733.950 997.050 734.400 ;
        RECT 142.950 732.600 145.050 733.050 ;
        RECT 157.950 732.600 160.050 733.050 ;
        RECT 142.950 731.400 160.050 732.600 ;
        RECT 142.950 730.950 145.050 731.400 ;
        RECT 157.950 730.950 160.050 731.400 ;
        RECT 244.950 732.600 247.050 733.050 ;
        RECT 298.950 732.600 301.050 733.050 ;
        RECT 244.950 731.400 301.050 732.600 ;
        RECT 244.950 730.950 247.050 731.400 ;
        RECT 298.950 730.950 301.050 731.400 ;
        RECT 451.950 732.600 454.050 733.050 ;
        RECT 463.950 732.600 466.050 733.050 ;
        RECT 520.950 732.600 523.050 733.050 ;
        RECT 529.950 732.600 532.050 733.050 ;
        RECT 451.950 731.400 466.050 732.600 ;
        RECT 451.950 730.950 454.050 731.400 ;
        RECT 463.950 730.950 466.050 731.400 ;
        RECT 488.400 731.400 532.050 732.600 ;
        RECT 55.950 729.600 58.050 730.200 ;
        RECT 67.950 729.600 70.050 730.050 ;
        RECT 55.950 728.400 70.050 729.600 ;
        RECT 55.950 728.100 58.050 728.400 ;
        RECT 67.950 727.950 70.050 728.400 ;
        RECT 76.950 729.600 79.050 730.200 ;
        RECT 91.950 729.600 94.050 730.050 ;
        RECT 105.000 729.600 109.050 730.050 ;
        RECT 76.950 728.400 94.050 729.600 ;
        RECT 76.950 728.100 79.050 728.400 ;
        RECT 91.950 727.950 94.050 728.400 ;
        RECT 104.400 727.950 109.050 729.600 ;
        RECT 121.950 729.600 124.050 730.200 ;
        RECT 139.950 729.600 142.050 730.050 ;
        RECT 121.950 728.400 142.050 729.600 ;
        RECT 121.950 728.100 124.050 728.400 ;
        RECT 139.950 727.950 142.050 728.400 ;
        RECT 154.950 729.750 157.050 730.200 ;
        RECT 160.950 729.750 163.050 730.050 ;
        RECT 169.950 729.750 172.050 730.200 ;
        RECT 154.950 729.600 172.050 729.750 ;
        RECT 190.950 729.600 193.050 730.200 ;
        RECT 154.950 728.550 193.050 729.600 ;
        RECT 154.950 728.100 157.050 728.550 ;
        RECT 160.950 727.950 163.050 728.550 ;
        RECT 169.950 728.400 193.050 728.550 ;
        RECT 169.950 728.100 172.050 728.400 ;
        RECT 190.950 728.100 193.050 728.400 ;
        RECT 208.950 729.600 211.050 730.050 ;
        RECT 241.950 729.600 244.050 730.200 ;
        RECT 208.950 728.400 244.050 729.600 ;
        RECT 208.950 727.950 211.050 728.400 ;
        RECT 241.950 728.100 244.050 728.400 ;
        RECT 104.400 723.900 105.600 727.950 ;
        RECT 245.400 723.900 246.600 730.950 ;
        RECT 259.950 729.750 262.050 729.900 ;
        RECT 277.950 729.750 280.050 730.200 ;
        RECT 259.950 728.550 280.050 729.750 ;
        RECT 259.950 727.800 262.050 728.550 ;
        RECT 277.950 728.100 280.050 728.550 ;
        RECT 301.950 729.750 304.050 730.200 ;
        RECT 313.950 729.750 316.050 730.200 ;
        RECT 301.950 728.550 316.050 729.750 ;
        RECT 301.950 728.100 304.050 728.550 ;
        RECT 313.950 728.100 316.050 728.550 ;
        RECT 415.950 728.100 418.050 730.200 ;
        RECT 436.950 729.750 439.050 730.200 ;
        RECT 445.950 729.750 448.050 730.200 ;
        RECT 436.950 728.550 448.050 729.750 ;
        RECT 488.400 729.600 489.600 731.400 ;
        RECT 520.950 730.950 523.050 731.400 ;
        RECT 529.950 730.950 532.050 731.400 ;
        RECT 634.950 732.600 637.050 733.050 ;
        RECT 670.950 732.600 673.050 733.050 ;
        RECT 634.950 731.400 673.050 732.600 ;
        RECT 634.950 730.950 637.050 731.400 ;
        RECT 670.950 730.950 673.050 731.400 ;
        RECT 700.950 732.600 703.050 733.050 ;
        RECT 709.950 732.600 712.050 733.050 ;
        RECT 700.950 731.400 712.050 732.600 ;
        RECT 700.950 730.950 703.050 731.400 ;
        RECT 709.950 730.950 712.050 731.400 ;
        RECT 826.950 732.600 829.050 733.050 ;
        RECT 841.950 732.600 844.050 733.200 ;
        RECT 862.950 732.600 865.050 733.050 ;
        RECT 826.950 731.400 865.050 732.600 ;
        RECT 826.950 730.950 829.050 731.400 ;
        RECT 841.950 731.100 844.050 731.400 ;
        RECT 862.950 730.950 865.050 731.400 ;
        RECT 964.950 730.950 967.050 733.050 ;
        RECT 436.950 728.100 439.050 728.550 ;
        RECT 445.950 728.100 448.050 728.550 ;
        RECT 449.400 728.400 489.600 729.600 ;
        RECT 400.950 726.600 403.050 727.050 ;
        RECT 416.400 726.600 417.600 728.100 ;
        RECT 449.400 726.600 450.600 728.400 ;
        RECT 511.950 728.100 514.050 730.200 ;
        RECT 535.950 729.600 538.050 730.200 ;
        RECT 565.950 729.600 568.050 730.050 ;
        RECT 535.950 728.400 568.050 729.600 ;
        RECT 535.950 728.100 538.050 728.400 ;
        RECT 347.400 725.400 403.050 726.600 ;
        RECT 67.950 723.450 70.050 723.900 ;
        RECT 73.950 723.450 76.050 723.900 ;
        RECT 67.950 722.250 76.050 723.450 ;
        RECT 67.950 721.800 70.050 722.250 ;
        RECT 73.950 721.800 76.050 722.250 ;
        RECT 79.950 723.450 82.050 723.900 ;
        RECT 85.950 723.450 88.050 723.900 ;
        RECT 79.950 722.250 88.050 723.450 ;
        RECT 79.950 721.800 82.050 722.250 ;
        RECT 85.950 721.800 88.050 722.250 ;
        RECT 103.950 721.800 106.050 723.900 ;
        RECT 145.950 723.450 148.050 723.900 ;
        RECT 160.950 723.450 163.050 723.900 ;
        RECT 145.950 722.250 163.050 723.450 ;
        RECT 145.950 721.800 148.050 722.250 ;
        RECT 160.950 721.800 163.050 722.250 ;
        RECT 166.950 723.600 169.050 723.900 ;
        RECT 193.950 723.600 196.050 723.900 ;
        RECT 166.950 722.400 196.050 723.600 ;
        RECT 166.950 721.800 169.050 722.400 ;
        RECT 193.950 721.800 196.050 722.400 ;
        RECT 199.950 723.450 202.050 723.900 ;
        RECT 208.950 723.450 211.050 723.900 ;
        RECT 199.950 722.250 211.050 723.450 ;
        RECT 199.950 721.800 202.050 722.250 ;
        RECT 208.950 721.800 211.050 722.250 ;
        RECT 223.950 723.600 226.050 723.900 ;
        RECT 238.950 723.600 241.050 723.900 ;
        RECT 223.950 722.400 241.050 723.600 ;
        RECT 223.950 721.800 226.050 722.400 ;
        RECT 238.950 721.800 241.050 722.400 ;
        RECT 244.950 721.800 247.050 723.900 ;
        RECT 253.950 723.450 256.050 723.900 ;
        RECT 262.950 723.450 265.050 723.900 ;
        RECT 253.950 722.250 265.050 723.450 ;
        RECT 253.950 721.800 256.050 722.250 ;
        RECT 262.950 721.800 265.050 722.250 ;
        RECT 283.950 723.600 286.050 724.050 ;
        RECT 298.950 723.600 301.050 723.900 ;
        RECT 283.950 722.400 301.050 723.600 ;
        RECT 283.950 721.950 286.050 722.400 ;
        RECT 298.950 721.800 301.050 722.400 ;
        RECT 328.950 723.600 331.050 724.050 ;
        RECT 347.400 723.900 348.600 725.400 ;
        RECT 400.950 724.950 403.050 725.400 ;
        RECT 407.400 725.400 450.600 726.600 ;
        RECT 458.400 725.400 507.600 726.600 ;
        RECT 346.950 723.600 349.050 723.900 ;
        RECT 328.950 722.400 349.050 723.600 ;
        RECT 328.950 721.950 331.050 722.400 ;
        RECT 346.950 721.800 349.050 722.400 ;
        RECT 370.950 723.600 373.050 723.900 ;
        RECT 391.950 723.600 394.050 723.900 ;
        RECT 370.950 722.400 394.050 723.600 ;
        RECT 370.950 721.800 373.050 722.400 ;
        RECT 391.950 721.800 394.050 722.400 ;
        RECT 400.950 723.600 403.050 723.900 ;
        RECT 407.400 723.600 408.600 725.400 ;
        RECT 458.400 723.900 459.600 725.400 ;
        RECT 400.950 722.400 408.600 723.600 ;
        RECT 424.950 723.450 427.050 723.900 ;
        RECT 433.950 723.450 436.050 723.900 ;
        RECT 400.950 721.800 403.050 722.400 ;
        RECT 424.950 722.250 436.050 723.450 ;
        RECT 424.950 721.800 427.050 722.250 ;
        RECT 433.950 721.800 436.050 722.250 ;
        RECT 439.950 723.600 442.050 723.900 ;
        RECT 457.950 723.600 460.050 723.900 ;
        RECT 439.950 722.400 460.050 723.600 ;
        RECT 439.950 721.800 442.050 722.400 ;
        RECT 457.950 721.800 460.050 722.400 ;
        RECT 496.950 723.450 499.050 723.900 ;
        RECT 502.950 723.450 505.050 723.900 ;
        RECT 496.950 722.250 505.050 723.450 ;
        RECT 506.400 723.600 507.600 725.400 ;
        RECT 508.950 723.600 511.050 723.900 ;
        RECT 506.400 722.400 511.050 723.600 ;
        RECT 512.400 723.600 513.600 728.100 ;
        RECT 565.950 727.950 568.050 728.400 ;
        RECT 577.950 729.600 580.050 730.200 ;
        RECT 604.950 729.600 607.050 730.200 ;
        RECT 577.950 728.400 607.050 729.600 ;
        RECT 577.950 728.100 580.050 728.400 ;
        RECT 604.950 728.100 607.050 728.400 ;
        RECT 610.950 729.600 613.050 730.200 ;
        RECT 619.950 729.750 622.050 730.200 ;
        RECT 625.950 729.750 628.050 730.200 ;
        RECT 619.950 729.600 628.050 729.750 ;
        RECT 655.950 729.600 658.050 730.200 ;
        RECT 610.950 728.550 628.050 729.600 ;
        RECT 610.950 728.400 622.050 728.550 ;
        RECT 610.950 728.100 613.050 728.400 ;
        RECT 619.950 728.100 622.050 728.400 ;
        RECT 625.950 728.100 628.050 728.550 ;
        RECT 635.400 728.400 658.050 729.600 ;
        RECT 517.950 723.600 520.050 724.050 ;
        RECT 635.400 723.900 636.600 728.400 ;
        RECT 655.950 728.100 658.050 728.400 ;
        RECT 688.950 729.600 691.050 730.050 ;
        RECT 706.950 729.600 709.050 730.050 ;
        RECT 712.950 729.600 715.050 730.050 ;
        RECT 754.950 729.600 757.050 730.050 ;
        RECT 688.950 728.400 715.050 729.600 ;
        RECT 688.950 727.950 691.050 728.400 ;
        RECT 706.950 727.950 709.050 728.400 ;
        RECT 712.950 727.950 715.050 728.400 ;
        RECT 746.400 728.400 757.050 729.600 ;
        RECT 701.400 725.400 723.600 726.600 ;
        RECT 512.400 722.400 520.050 723.600 ;
        RECT 496.950 721.800 499.050 722.250 ;
        RECT 502.950 721.800 505.050 722.250 ;
        RECT 508.950 721.800 511.050 722.400 ;
        RECT 517.950 721.950 520.050 722.400 ;
        RECT 526.950 723.450 529.050 723.900 ;
        RECT 553.950 723.450 556.050 723.900 ;
        RECT 526.950 722.250 556.050 723.450 ;
        RECT 526.950 721.800 529.050 722.250 ;
        RECT 553.950 721.800 556.050 722.250 ;
        RECT 568.950 723.450 571.050 723.900 ;
        RECT 574.950 723.450 577.050 723.900 ;
        RECT 568.950 722.250 577.050 723.450 ;
        RECT 568.950 721.800 571.050 722.250 ;
        RECT 574.950 721.800 577.050 722.250 ;
        RECT 595.950 723.450 598.050 723.900 ;
        RECT 601.950 723.450 604.050 723.900 ;
        RECT 595.950 722.250 604.050 723.450 ;
        RECT 595.950 721.800 598.050 722.250 ;
        RECT 601.950 721.800 604.050 722.250 ;
        RECT 634.950 721.800 637.050 723.900 ;
        RECT 643.950 723.450 646.050 723.900 ;
        RECT 658.950 723.600 661.050 723.900 ;
        RECT 673.950 723.600 676.050 723.900 ;
        RECT 701.400 723.600 702.600 725.400 ;
        RECT 658.950 723.450 702.600 723.600 ;
        RECT 643.950 722.400 702.600 723.450 ;
        RECT 706.950 723.600 709.050 724.050 ;
        RECT 715.950 723.600 718.050 724.050 ;
        RECT 722.400 723.900 723.600 725.400 ;
        RECT 746.400 723.900 747.600 728.400 ;
        RECT 754.950 727.950 757.050 728.400 ;
        RECT 763.950 729.600 766.050 730.050 ;
        RECT 781.800 729.600 783.900 730.050 ;
        RECT 763.950 728.400 783.900 729.600 ;
        RECT 763.950 727.950 766.050 728.400 ;
        RECT 781.800 727.950 783.900 728.400 ;
        RECT 784.950 729.750 787.050 730.200 ;
        RECT 790.950 729.750 793.050 730.200 ;
        RECT 784.950 728.550 793.050 729.750 ;
        RECT 784.950 728.100 787.050 728.550 ;
        RECT 790.950 728.100 793.050 728.550 ;
        RECT 796.950 729.750 799.050 730.200 ;
        RECT 802.950 729.750 805.050 730.200 ;
        RECT 796.950 729.600 805.050 729.750 ;
        RECT 820.950 729.600 823.050 730.200 ;
        RECT 796.950 728.550 823.050 729.600 ;
        RECT 796.950 728.100 799.050 728.550 ;
        RECT 802.950 728.400 823.050 728.550 ;
        RECT 802.950 728.100 805.050 728.400 ;
        RECT 820.950 728.100 823.050 728.400 ;
        RECT 835.950 728.100 838.050 730.200 ;
        RECT 841.950 729.600 844.050 730.050 ;
        RECT 880.950 729.750 883.050 730.200 ;
        RECT 889.950 729.750 892.050 730.200 ;
        RECT 841.950 728.400 846.600 729.600 ;
        RECT 706.950 722.400 718.050 723.600 ;
        RECT 643.950 722.250 661.050 722.400 ;
        RECT 643.950 721.800 646.050 722.250 ;
        RECT 658.950 721.800 661.050 722.250 ;
        RECT 673.950 721.800 676.050 722.400 ;
        RECT 706.950 721.950 709.050 722.400 ;
        RECT 715.950 721.950 718.050 722.400 ;
        RECT 721.950 721.800 724.050 723.900 ;
        RECT 745.950 721.800 748.050 723.900 ;
        RECT 775.950 723.600 778.050 723.900 ;
        RECT 802.950 723.600 805.050 724.050 ;
        RECT 775.950 722.400 805.050 723.600 ;
        RECT 775.950 721.800 778.050 722.400 ;
        RECT 802.950 721.950 805.050 722.400 ;
        RECT 817.950 723.600 820.050 723.900 ;
        RECT 836.400 723.600 837.600 728.100 ;
        RECT 841.950 727.950 844.050 728.400 ;
        RECT 817.950 722.400 837.600 723.600 ;
        RECT 817.950 721.800 820.050 722.400 ;
        RECT 845.400 721.050 846.600 728.400 ;
        RECT 880.950 728.550 892.050 729.750 ;
        RECT 880.950 728.100 883.050 728.550 ;
        RECT 889.950 728.100 892.050 728.550 ;
        RECT 895.950 729.600 898.050 730.200 ;
        RECT 904.950 729.600 907.050 730.050 ;
        RECT 895.950 728.400 907.050 729.600 ;
        RECT 895.950 728.100 898.050 728.400 ;
        RECT 904.950 727.950 907.050 728.400 ;
        RECT 913.950 728.100 916.050 730.200 ;
        RECT 914.400 726.600 915.600 728.100 ;
        RECT 934.950 727.950 937.050 730.050 ;
        RECT 943.950 729.600 946.050 730.200 ;
        RECT 941.400 728.400 946.050 729.600 ;
        RECT 890.400 725.400 915.600 726.600 ;
        RECT 850.950 723.450 853.050 723.900 ;
        RECT 871.950 723.600 874.050 723.900 ;
        RECT 886.950 723.600 889.050 723.900 ;
        RECT 871.950 723.450 889.050 723.600 ;
        RECT 850.950 722.400 889.050 723.450 ;
        RECT 850.950 722.250 874.050 722.400 ;
        RECT 850.950 721.800 853.050 722.250 ;
        RECT 871.950 721.800 874.050 722.250 ;
        RECT 886.950 721.800 889.050 722.400 ;
        RECT 890.400 721.050 891.600 725.400 ;
        RECT 935.400 724.050 936.600 727.950 ;
        RECT 892.950 723.450 895.050 723.900 ;
        RECT 901.950 723.450 904.050 723.900 ;
        RECT 892.950 722.250 904.050 723.450 ;
        RECT 892.950 721.800 895.050 722.250 ;
        RECT 901.950 721.800 904.050 722.250 ;
        RECT 934.950 721.950 937.050 724.050 ;
        RECT 941.400 721.050 942.600 728.400 ;
        RECT 943.950 728.100 946.050 728.400 ;
        RECT 965.400 723.900 966.600 730.950 ;
        RECT 967.950 729.600 970.050 730.200 ;
        RECT 991.950 729.600 994.050 730.200 ;
        RECT 997.950 729.600 1000.050 733.050 ;
        RECT 967.950 728.400 978.600 729.600 ;
        RECT 967.950 728.100 970.050 728.400 ;
        RECT 964.950 721.800 967.050 723.900 ;
        RECT 91.950 720.600 94.050 721.050 ;
        RECT 97.950 720.600 100.050 721.050 ;
        RECT 91.950 719.400 100.050 720.600 ;
        RECT 91.950 718.950 94.050 719.400 ;
        RECT 97.950 718.950 100.050 719.400 ;
        RECT 112.950 720.600 115.050 721.050 ;
        RECT 124.950 720.600 127.050 721.050 ;
        RECT 112.950 719.400 127.050 720.600 ;
        RECT 112.950 718.950 115.050 719.400 ;
        RECT 124.950 718.950 127.050 719.400 ;
        RECT 355.950 720.600 358.050 721.050 ;
        RECT 412.950 720.600 415.050 721.050 ;
        RECT 472.950 720.600 475.050 721.050 ;
        RECT 478.950 720.600 481.050 721.050 ;
        RECT 355.950 719.400 481.050 720.600 ;
        RECT 355.950 718.950 358.050 719.400 ;
        RECT 412.950 718.950 415.050 719.400 ;
        RECT 472.950 718.950 475.050 719.400 ;
        RECT 478.950 718.950 481.050 719.400 ;
        RECT 538.950 720.600 541.050 721.050 ;
        RECT 544.950 720.600 547.050 721.050 ;
        RECT 538.950 719.400 547.050 720.600 ;
        RECT 538.950 718.950 541.050 719.400 ;
        RECT 544.950 718.950 547.050 719.400 ;
        RECT 832.950 720.600 835.050 721.050 ;
        RECT 838.950 720.600 841.050 721.050 ;
        RECT 832.950 719.400 841.050 720.600 ;
        RECT 832.950 718.950 835.050 719.400 ;
        RECT 838.950 718.950 841.050 719.400 ;
        RECT 844.950 718.950 847.050 721.050 ;
        RECT 889.950 718.950 892.050 721.050 ;
        RECT 937.950 719.400 942.600 721.050 ;
        RECT 977.400 720.600 978.600 728.400 ;
        RECT 991.950 729.000 1000.050 729.600 ;
        RECT 991.950 728.400 999.600 729.000 ;
        RECT 991.950 728.100 994.050 728.400 ;
        RECT 982.950 723.450 985.050 723.900 ;
        RECT 994.800 723.450 996.900 723.900 ;
        RECT 982.950 722.250 996.900 723.450 ;
        RECT 982.950 721.800 985.050 722.250 ;
        RECT 994.800 721.800 996.900 722.250 ;
        RECT 997.950 723.600 1000.050 724.050 ;
        RECT 1003.950 723.600 1006.050 724.050 ;
        RECT 997.950 722.400 1006.050 723.600 ;
        RECT 997.950 721.950 1000.050 722.400 ;
        RECT 1003.950 721.950 1006.050 722.400 ;
        RECT 988.950 720.600 991.050 721.050 ;
        RECT 977.400 719.400 991.050 720.600 ;
        RECT 937.950 718.950 942.000 719.400 ;
        RECT 988.950 718.950 991.050 719.400 ;
        RECT 139.950 717.600 142.050 718.050 ;
        RECT 151.950 717.600 154.050 718.050 ;
        RECT 166.950 717.600 169.050 718.050 ;
        RECT 139.950 716.400 169.050 717.600 ;
        RECT 139.950 715.950 142.050 716.400 ;
        RECT 151.950 715.950 154.050 716.400 ;
        RECT 166.950 715.950 169.050 716.400 ;
        RECT 175.950 717.600 178.050 718.050 ;
        RECT 202.950 717.600 205.050 718.050 ;
        RECT 214.950 717.600 217.050 718.050 ;
        RECT 175.950 716.400 217.050 717.600 ;
        RECT 175.950 715.950 178.050 716.400 ;
        RECT 202.950 715.950 205.050 716.400 ;
        RECT 214.950 715.950 217.050 716.400 ;
        RECT 238.950 717.600 241.050 718.050 ;
        RECT 259.950 717.600 262.050 718.050 ;
        RECT 238.950 716.400 262.050 717.600 ;
        RECT 238.950 715.950 241.050 716.400 ;
        RECT 259.950 715.950 262.050 716.400 ;
        RECT 316.950 717.600 319.050 718.050 ;
        RECT 331.950 717.600 334.050 718.050 ;
        RECT 316.950 716.400 334.050 717.600 ;
        RECT 316.950 715.950 319.050 716.400 ;
        RECT 331.950 715.950 334.050 716.400 ;
        RECT 487.950 717.600 490.050 718.050 ;
        RECT 493.950 717.600 496.050 718.050 ;
        RECT 487.950 716.400 496.050 717.600 ;
        RECT 487.950 715.950 490.050 716.400 ;
        RECT 493.950 715.950 496.050 716.400 ;
        RECT 625.950 717.600 628.050 718.050 ;
        RECT 763.950 717.600 766.050 718.050 ;
        RECT 625.950 716.400 766.050 717.600 ;
        RECT 625.950 715.950 628.050 716.400 ;
        RECT 763.950 715.950 766.050 716.400 ;
        RECT 769.950 717.600 772.050 718.050 ;
        RECT 784.950 717.600 787.050 718.050 ;
        RECT 769.950 716.400 787.050 717.600 ;
        RECT 769.950 715.950 772.050 716.400 ;
        RECT 784.950 715.950 787.050 716.400 ;
        RECT 877.950 717.600 880.050 718.050 ;
        RECT 886.950 717.600 889.050 718.050 ;
        RECT 877.950 716.400 889.050 717.600 ;
        RECT 877.950 715.950 880.050 716.400 ;
        RECT 886.950 715.950 889.050 716.400 ;
        RECT 952.950 717.600 955.050 718.050 ;
        RECT 967.950 717.600 970.050 718.050 ;
        RECT 952.950 716.400 970.050 717.600 ;
        RECT 952.950 715.950 955.050 716.400 ;
        RECT 967.950 715.950 970.050 716.400 ;
        RECT 28.950 714.600 31.050 715.050 ;
        RECT 37.950 714.600 40.050 715.050 ;
        RECT 28.950 713.400 40.050 714.600 ;
        RECT 28.950 712.950 31.050 713.400 ;
        RECT 37.950 712.950 40.050 713.400 ;
        RECT 52.950 714.600 55.050 715.050 ;
        RECT 112.950 714.600 115.050 715.050 ;
        RECT 52.950 713.400 115.050 714.600 ;
        RECT 52.950 712.950 55.050 713.400 ;
        RECT 112.950 712.950 115.050 713.400 ;
        RECT 586.950 714.600 589.050 715.050 ;
        RECT 628.950 714.600 631.050 715.050 ;
        RECT 586.950 713.400 631.050 714.600 ;
        RECT 586.950 712.950 589.050 713.400 ;
        RECT 628.950 712.950 631.050 713.400 ;
        RECT 670.950 714.600 673.050 715.050 ;
        RECT 709.800 714.600 711.900 715.050 ;
        RECT 670.950 713.400 711.900 714.600 ;
        RECT 670.950 712.950 673.050 713.400 ;
        RECT 709.800 712.950 711.900 713.400 ;
        RECT 712.950 714.600 715.050 715.050 ;
        RECT 721.950 714.600 724.050 715.050 ;
        RECT 751.950 714.600 754.050 715.050 ;
        RECT 712.950 713.400 754.050 714.600 ;
        RECT 712.950 712.950 715.050 713.400 ;
        RECT 721.950 712.950 724.050 713.400 ;
        RECT 751.950 712.950 754.050 713.400 ;
        RECT 793.950 714.600 796.050 715.050 ;
        RECT 862.950 714.600 865.050 715.050 ;
        RECT 793.950 713.400 865.050 714.600 ;
        RECT 793.950 712.950 796.050 713.400 ;
        RECT 862.950 712.950 865.050 713.400 ;
        RECT 940.950 714.600 943.050 715.050 ;
        RECT 994.950 714.600 997.050 715.050 ;
        RECT 940.950 713.400 997.050 714.600 ;
        RECT 940.950 712.950 943.050 713.400 ;
        RECT 994.950 712.950 997.050 713.400 ;
        RECT 475.950 711.600 478.050 712.050 ;
        RECT 526.950 711.600 529.050 712.050 ;
        RECT 643.950 711.600 646.050 712.050 ;
        RECT 475.950 710.400 646.050 711.600 ;
        RECT 475.950 709.950 478.050 710.400 ;
        RECT 526.950 709.950 529.050 710.400 ;
        RECT 643.950 709.950 646.050 710.400 ;
        RECT 682.950 711.600 685.050 712.050 ;
        RECT 688.950 711.600 691.050 712.050 ;
        RECT 682.950 710.400 691.050 711.600 ;
        RECT 682.950 709.950 685.050 710.400 ;
        RECT 688.950 709.950 691.050 710.400 ;
        RECT 727.950 711.600 730.050 712.050 ;
        RECT 739.950 711.600 742.050 712.050 ;
        RECT 727.950 710.400 742.050 711.600 ;
        RECT 727.950 709.950 730.050 710.400 ;
        RECT 739.950 709.950 742.050 710.400 ;
        RECT 865.950 711.600 868.050 712.050 ;
        RECT 907.950 711.600 910.050 712.050 ;
        RECT 865.950 710.400 910.050 711.600 ;
        RECT 865.950 709.950 868.050 710.400 ;
        RECT 907.950 709.950 910.050 710.400 ;
        RECT 946.950 711.600 949.050 712.050 ;
        RECT 988.950 711.600 991.050 712.050 ;
        RECT 946.950 710.400 991.050 711.600 ;
        RECT 946.950 709.950 949.050 710.400 ;
        RECT 988.950 709.950 991.050 710.400 ;
        RECT 226.950 708.600 229.050 709.050 ;
        RECT 352.950 708.600 355.050 709.050 ;
        RECT 226.950 707.400 355.050 708.600 ;
        RECT 226.950 706.950 229.050 707.400 ;
        RECT 352.950 706.950 355.050 707.400 ;
        RECT 445.950 708.600 448.050 709.050 ;
        RECT 463.950 708.600 466.050 709.050 ;
        RECT 514.950 708.600 517.050 709.050 ;
        RECT 445.950 707.400 517.050 708.600 ;
        RECT 445.950 706.950 448.050 707.400 ;
        RECT 463.950 706.950 466.050 707.400 ;
        RECT 514.950 706.950 517.050 707.400 ;
        RECT 532.950 708.600 535.050 709.050 ;
        RECT 586.950 708.600 589.050 709.050 ;
        RECT 532.950 707.400 589.050 708.600 ;
        RECT 532.950 706.950 535.050 707.400 ;
        RECT 586.950 706.950 589.050 707.400 ;
        RECT 604.950 708.600 607.050 709.050 ;
        RECT 637.950 708.600 640.050 709.050 ;
        RECT 604.950 707.400 640.050 708.600 ;
        RECT 604.950 706.950 607.050 707.400 ;
        RECT 637.950 706.950 640.050 707.400 ;
        RECT 772.950 708.600 775.050 709.050 ;
        RECT 805.950 708.600 808.050 709.050 ;
        RECT 772.950 707.400 808.050 708.600 ;
        RECT 772.950 706.950 775.050 707.400 ;
        RECT 805.950 706.950 808.050 707.400 ;
        RECT 868.950 708.600 871.050 709.050 ;
        RECT 916.950 708.600 919.050 709.050 ;
        RECT 868.950 707.400 919.050 708.600 ;
        RECT 868.950 706.950 871.050 707.400 ;
        RECT 916.950 706.950 919.050 707.400 ;
        RECT 964.950 708.600 967.050 709.050 ;
        RECT 979.950 708.600 982.050 709.050 ;
        RECT 964.950 707.400 982.050 708.600 ;
        RECT 964.950 706.950 967.050 707.400 ;
        RECT 979.950 706.950 982.050 707.400 ;
        RECT 7.950 705.600 10.050 706.050 ;
        RECT 19.950 705.600 22.050 706.050 ;
        RECT 67.950 705.600 70.050 706.050 ;
        RECT 7.950 704.400 70.050 705.600 ;
        RECT 7.950 703.950 10.050 704.400 ;
        RECT 19.950 703.950 22.050 704.400 ;
        RECT 67.950 703.950 70.050 704.400 ;
        RECT 220.950 705.600 223.050 706.050 ;
        RECT 355.950 705.600 358.050 706.050 ;
        RECT 220.950 704.400 358.050 705.600 ;
        RECT 220.950 703.950 223.050 704.400 ;
        RECT 355.950 703.950 358.050 704.400 ;
        RECT 517.950 705.600 520.050 706.050 ;
        RECT 562.950 705.600 565.050 706.050 ;
        RECT 667.950 705.600 670.050 706.050 ;
        RECT 940.950 705.600 943.050 706.050 ;
        RECT 517.950 704.400 633.600 705.600 ;
        RECT 517.950 703.950 520.050 704.400 ;
        RECT 562.950 703.950 565.050 704.400 ;
        RECT 124.950 702.600 127.050 703.050 ;
        RECT 217.950 702.600 220.050 703.050 ;
        RECT 124.950 701.400 220.050 702.600 ;
        RECT 632.400 702.600 633.600 704.400 ;
        RECT 667.950 704.400 943.050 705.600 ;
        RECT 667.950 703.950 670.050 704.400 ;
        RECT 940.950 703.950 943.050 704.400 ;
        RECT 955.950 705.600 958.050 706.050 ;
        RECT 1003.950 705.600 1006.050 706.050 ;
        RECT 955.950 704.400 1006.050 705.600 ;
        RECT 955.950 703.950 958.050 704.400 ;
        RECT 1003.950 703.950 1006.050 704.400 ;
        RECT 937.950 702.600 940.050 703.050 ;
        RECT 632.400 701.400 940.050 702.600 ;
        RECT 124.950 700.950 127.050 701.400 ;
        RECT 217.950 700.950 220.050 701.400 ;
        RECT 937.950 700.950 940.050 701.400 ;
        RECT 979.950 702.600 982.050 703.050 ;
        RECT 985.950 702.600 988.050 703.050 ;
        RECT 979.950 701.400 988.050 702.600 ;
        RECT 979.950 700.950 982.050 701.400 ;
        RECT 985.950 700.950 988.050 701.400 ;
        RECT 31.950 699.600 34.050 700.050 ;
        RECT 43.950 699.600 46.050 700.050 ;
        RECT 88.950 699.600 91.050 700.050 ;
        RECT 31.950 698.400 91.050 699.600 ;
        RECT 31.950 697.950 34.050 698.400 ;
        RECT 43.950 697.950 46.050 698.400 ;
        RECT 88.950 697.950 91.050 698.400 ;
        RECT 229.950 699.600 232.050 700.050 ;
        RECT 256.950 699.600 259.050 700.050 ;
        RECT 316.950 699.600 319.050 700.050 ;
        RECT 229.950 698.400 319.050 699.600 ;
        RECT 229.950 697.950 232.050 698.400 ;
        RECT 256.950 697.950 259.050 698.400 ;
        RECT 316.950 697.950 319.050 698.400 ;
        RECT 355.950 699.600 358.050 700.050 ;
        RECT 364.950 699.600 367.050 700.050 ;
        RECT 355.950 698.400 367.050 699.600 ;
        RECT 355.950 697.950 358.050 698.400 ;
        RECT 364.950 697.950 367.050 698.400 ;
        RECT 412.950 699.600 415.050 700.050 ;
        RECT 448.950 699.600 451.050 700.050 ;
        RECT 412.950 698.400 451.050 699.600 ;
        RECT 412.950 697.950 415.050 698.400 ;
        RECT 448.950 697.950 451.050 698.400 ;
        RECT 673.950 699.600 676.050 700.050 ;
        RECT 691.950 699.600 694.050 700.050 ;
        RECT 673.950 698.400 694.050 699.600 ;
        RECT 673.950 697.950 676.050 698.400 ;
        RECT 691.950 697.950 694.050 698.400 ;
        RECT 697.950 699.600 700.050 700.050 ;
        RECT 724.950 699.600 727.050 700.050 ;
        RECT 697.950 698.400 727.050 699.600 ;
        RECT 697.950 697.950 700.050 698.400 ;
        RECT 724.950 697.950 727.050 698.400 ;
        RECT 730.950 699.600 733.050 700.050 ;
        RECT 736.950 699.600 739.050 700.050 ;
        RECT 730.950 698.400 739.050 699.600 ;
        RECT 730.950 697.950 733.050 698.400 ;
        RECT 736.950 697.950 739.050 698.400 ;
        RECT 751.950 699.600 754.050 700.050 ;
        RECT 769.950 699.600 772.050 700.050 ;
        RECT 751.950 698.400 772.050 699.600 ;
        RECT 751.950 697.950 754.050 698.400 ;
        RECT 769.950 697.950 772.050 698.400 ;
        RECT 16.950 696.600 19.050 697.050 ;
        RECT 25.950 696.600 28.050 697.050 ;
        RECT 16.950 695.400 28.050 696.600 ;
        RECT 16.950 694.950 19.050 695.400 ;
        RECT 25.950 694.950 28.050 695.400 ;
        RECT 196.950 696.600 199.050 697.050 ;
        RECT 226.950 696.600 229.050 697.050 ;
        RECT 196.950 695.400 229.050 696.600 ;
        RECT 196.950 694.950 199.050 695.400 ;
        RECT 226.950 694.950 229.050 695.400 ;
        RECT 352.950 696.600 355.050 697.050 ;
        RECT 406.950 696.600 409.050 697.050 ;
        RECT 352.950 695.400 409.050 696.600 ;
        RECT 352.950 694.950 355.050 695.400 ;
        RECT 406.950 694.950 409.050 695.400 ;
        RECT 454.950 696.600 457.050 697.050 ;
        RECT 502.950 696.600 505.050 697.050 ;
        RECT 523.950 696.600 526.050 697.050 ;
        RECT 454.950 695.400 526.050 696.600 ;
        RECT 454.950 694.950 457.050 695.400 ;
        RECT 502.950 694.950 505.050 695.400 ;
        RECT 523.950 694.950 526.050 695.400 ;
        RECT 781.950 696.600 784.050 697.050 ;
        RECT 796.950 696.600 799.050 697.050 ;
        RECT 781.950 695.400 799.050 696.600 ;
        RECT 781.950 694.950 784.050 695.400 ;
        RECT 796.950 694.950 799.050 695.400 ;
        RECT 838.950 696.600 841.050 697.050 ;
        RECT 880.950 696.600 883.050 697.050 ;
        RECT 838.950 695.400 883.050 696.600 ;
        RECT 838.950 694.950 841.050 695.400 ;
        RECT 880.950 694.950 883.050 695.400 ;
        RECT 898.950 696.600 901.050 697.050 ;
        RECT 904.950 696.600 907.050 697.050 ;
        RECT 898.950 695.400 907.050 696.600 ;
        RECT 898.950 694.950 901.050 695.400 ;
        RECT 904.950 694.950 907.050 695.400 ;
        RECT 46.950 693.600 49.050 694.050 ;
        RECT 76.950 693.600 79.050 694.050 ;
        RECT 46.950 692.400 79.050 693.600 ;
        RECT 46.950 691.950 49.050 692.400 ;
        RECT 76.950 691.950 79.050 692.400 ;
        RECT 259.950 693.600 262.050 694.050 ;
        RECT 346.950 693.600 349.050 694.050 ;
        RECT 259.950 692.400 349.050 693.600 ;
        RECT 259.950 691.950 262.050 692.400 ;
        RECT 346.950 691.950 349.050 692.400 ;
        RECT 535.950 693.600 538.050 694.050 ;
        RECT 568.950 693.600 571.050 694.050 ;
        RECT 535.950 692.400 571.050 693.600 ;
        RECT 535.950 691.950 538.050 692.400 ;
        RECT 568.950 691.950 571.050 692.400 ;
        RECT 577.950 693.600 580.050 694.050 ;
        RECT 592.950 693.600 595.050 694.050 ;
        RECT 610.950 693.600 613.050 694.050 ;
        RECT 577.950 692.400 613.050 693.600 ;
        RECT 577.950 691.950 580.050 692.400 ;
        RECT 592.950 691.950 595.050 692.400 ;
        RECT 610.950 691.950 613.050 692.400 ;
        RECT 703.950 693.600 706.050 693.900 ;
        RECT 736.950 693.600 739.050 694.050 ;
        RECT 703.950 692.400 739.050 693.600 ;
        RECT 703.950 691.800 706.050 692.400 ;
        RECT 736.950 691.950 739.050 692.400 ;
        RECT 781.950 693.600 784.050 693.900 ;
        RECT 955.950 693.600 958.050 694.050 ;
        RECT 781.950 692.400 958.050 693.600 ;
        RECT 781.950 691.800 784.050 692.400 ;
        RECT 955.950 691.950 958.050 692.400 ;
        RECT 967.950 693.600 970.050 694.050 ;
        RECT 988.950 693.600 991.050 694.050 ;
        RECT 967.950 692.400 991.050 693.600 ;
        RECT 967.950 691.950 970.050 692.400 ;
        RECT 988.950 691.950 991.050 692.400 ;
        RECT 358.950 690.600 361.050 691.050 ;
        RECT 376.950 690.600 379.050 691.050 ;
        RECT 358.950 689.400 379.050 690.600 ;
        RECT 358.950 688.950 361.050 689.400 ;
        RECT 376.950 688.950 379.050 689.400 ;
        RECT 484.950 690.600 487.050 691.050 ;
        RECT 490.950 690.600 493.050 691.050 ;
        RECT 484.950 689.400 493.050 690.600 ;
        RECT 484.950 688.950 487.050 689.400 ;
        RECT 490.950 688.950 493.050 689.400 ;
        RECT 520.950 690.600 523.050 691.050 ;
        RECT 529.950 690.600 532.050 691.050 ;
        RECT 520.950 689.400 532.050 690.600 ;
        RECT 520.950 688.950 523.050 689.400 ;
        RECT 529.950 688.950 532.050 689.400 ;
        RECT 556.950 690.600 559.050 691.050 ;
        RECT 655.950 690.600 658.050 691.050 ;
        RECT 556.950 689.400 658.050 690.600 ;
        RECT 556.950 688.950 559.050 689.400 ;
        RECT 655.950 688.950 658.050 689.400 ;
        RECT 874.950 690.600 877.050 691.050 ;
        RECT 898.950 690.600 901.050 691.050 ;
        RECT 874.950 689.400 901.050 690.600 ;
        RECT 874.950 688.950 877.050 689.400 ;
        RECT 898.950 688.950 901.050 689.400 ;
        RECT 934.950 690.600 937.050 691.050 ;
        RECT 958.950 690.600 961.050 691.050 ;
        RECT 934.950 689.400 961.050 690.600 ;
        RECT 934.950 688.950 937.050 689.400 ;
        RECT 958.950 688.950 961.050 689.400 ;
        RECT 1012.950 690.600 1017.000 691.050 ;
        RECT 1012.950 688.950 1017.600 690.600 ;
        RECT 52.950 687.600 55.050 688.050 ;
        RECT 295.950 687.600 298.050 688.050 ;
        RECT 313.950 687.600 316.050 688.050 ;
        RECT 52.950 686.400 72.600 687.600 ;
        RECT 52.950 685.950 55.050 686.400 ;
        RECT 71.400 685.200 72.600 686.400 ;
        RECT 295.950 686.400 316.050 687.600 ;
        RECT 295.950 685.950 298.050 686.400 ;
        RECT 313.950 685.950 316.050 686.400 ;
        RECT 352.950 687.600 355.050 688.050 ;
        RECT 370.950 687.600 373.050 688.050 ;
        RECT 352.950 686.400 373.050 687.600 ;
        RECT 352.950 685.950 355.050 686.400 ;
        RECT 370.950 685.950 373.050 686.400 ;
        RECT 463.950 687.600 466.050 688.050 ;
        RECT 475.950 687.600 478.050 688.050 ;
        RECT 463.950 686.400 478.050 687.600 ;
        RECT 463.950 685.950 466.050 686.400 ;
        RECT 475.950 685.950 478.050 686.400 ;
        RECT 550.950 687.600 553.050 688.050 ;
        RECT 616.950 687.600 619.050 688.200 ;
        RECT 703.950 687.600 706.050 688.050 ;
        RECT 550.950 686.400 619.050 687.600 ;
        RECT 550.950 685.950 553.050 686.400 ;
        RECT 616.950 686.100 619.050 686.400 ;
        RECT 689.400 686.400 706.050 687.600 ;
        RECT 22.950 683.100 25.050 685.200 ;
        RECT 58.950 684.750 61.050 685.200 ;
        RECT 64.950 684.750 67.050 685.200 ;
        RECT 58.950 683.550 67.050 684.750 ;
        RECT 58.950 683.100 61.050 683.550 ;
        RECT 64.950 683.100 67.050 683.550 ;
        RECT 70.950 684.750 73.050 685.200 ;
        RECT 82.950 684.750 85.050 685.200 ;
        RECT 70.950 683.550 85.050 684.750 ;
        RECT 70.950 683.100 73.050 683.550 ;
        RECT 82.950 683.100 85.050 683.550 ;
        RECT 100.950 684.750 103.050 685.200 ;
        RECT 157.950 684.750 160.050 685.200 ;
        RECT 100.950 683.550 160.050 684.750 ;
        RECT 100.950 683.100 103.050 683.550 ;
        RECT 157.950 683.100 160.050 683.550 ;
        RECT 163.950 684.600 166.050 685.200 ;
        RECT 178.950 684.600 181.050 685.200 ;
        RECT 163.950 683.400 181.050 684.600 ;
        RECT 163.950 683.100 166.050 683.400 ;
        RECT 178.950 683.100 181.050 683.400 ;
        RECT 235.950 684.600 238.050 685.200 ;
        RECT 244.950 684.750 247.050 685.200 ;
        RECT 250.950 684.750 253.050 685.200 ;
        RECT 244.950 684.600 253.050 684.750 ;
        RECT 235.950 683.550 253.050 684.600 ;
        RECT 235.950 683.400 247.050 683.550 ;
        RECT 235.950 683.100 238.050 683.400 ;
        RECT 244.950 683.100 247.050 683.400 ;
        RECT 250.950 683.100 253.050 683.550 ;
        RECT 289.950 684.600 292.050 685.050 ;
        RECT 301.950 684.600 304.050 685.200 ;
        RECT 319.950 684.600 322.050 685.200 ;
        RECT 289.950 683.400 322.050 684.600 ;
        RECT 23.400 681.600 24.600 683.100 ;
        RECT 289.950 682.950 292.050 683.400 ;
        RECT 301.950 683.100 304.050 683.400 ;
        RECT 319.950 683.100 322.050 683.400 ;
        RECT 340.950 683.100 343.050 685.200 ;
        RECT 355.950 684.750 358.050 685.200 ;
        RECT 376.950 684.750 379.050 685.200 ;
        RECT 355.950 683.550 379.050 684.750 ;
        RECT 355.950 683.100 358.050 683.550 ;
        RECT 376.950 683.100 379.050 683.550 ;
        RECT 385.950 684.600 388.050 685.050 ;
        RECT 391.950 684.600 394.050 685.200 ;
        RECT 385.950 683.400 394.050 684.600 ;
        RECT 148.950 681.600 151.050 682.050 ;
        RECT 23.400 680.400 48.600 681.600 ;
        RECT 4.950 678.450 7.050 678.900 ;
        RECT 43.950 678.450 46.050 678.900 ;
        RECT 4.950 677.250 46.050 678.450 ;
        RECT 47.400 678.600 48.600 680.400 ;
        RECT 148.950 680.400 234.600 681.600 ;
        RECT 148.950 679.950 151.050 680.400 ;
        RECT 55.950 678.600 58.050 678.900 ;
        RECT 47.400 677.400 58.050 678.600 ;
        RECT 4.950 676.800 7.050 677.250 ;
        RECT 43.950 676.800 46.050 677.250 ;
        RECT 55.950 676.800 58.050 677.400 ;
        RECT 64.950 678.600 67.050 679.050 ;
        RECT 233.400 678.900 234.600 680.400 ;
        RECT 341.400 679.050 342.600 683.100 ;
        RECT 385.950 682.950 388.050 683.400 ;
        RECT 391.950 683.100 394.050 683.400 ;
        RECT 418.950 684.750 421.050 685.200 ;
        RECT 430.950 684.750 433.050 685.200 ;
        RECT 418.950 683.550 433.050 684.750 ;
        RECT 418.950 683.100 421.050 683.550 ;
        RECT 430.950 683.100 433.050 683.550 ;
        RECT 490.950 683.100 493.050 685.200 ;
        RECT 511.950 684.600 514.050 685.200 ;
        RECT 523.950 684.600 526.050 685.050 ;
        RECT 511.950 683.400 526.050 684.600 ;
        RECT 511.950 683.100 514.050 683.400 ;
        RECT 491.400 681.600 492.600 683.100 ;
        RECT 523.950 682.950 526.050 683.400 ;
        RECT 529.950 684.600 532.050 685.050 ;
        RECT 556.950 684.600 559.050 685.050 ;
        RECT 568.950 684.750 571.050 685.200 ;
        RECT 574.950 684.750 577.050 685.200 ;
        RECT 529.950 683.400 549.600 684.600 ;
        RECT 529.950 682.950 532.050 683.400 ;
        RECT 499.950 681.600 502.050 682.050 ;
        RECT 491.400 680.400 502.050 681.600 ;
        RECT 548.400 681.600 549.600 683.400 ;
        RECT 556.950 683.400 567.600 684.600 ;
        RECT 556.950 682.950 559.050 683.400 ;
        RECT 548.400 680.400 555.600 681.600 ;
        RECT 499.950 679.950 502.050 680.400 ;
        RECT 554.400 679.050 555.600 680.400 ;
        RECT 79.950 678.600 82.050 678.900 ;
        RECT 64.950 677.400 82.050 678.600 ;
        RECT 64.950 676.950 67.050 677.400 ;
        RECT 79.950 676.800 82.050 677.400 ;
        RECT 232.950 676.800 235.050 678.900 ;
        RECT 253.950 678.600 256.050 678.900 ;
        RECT 268.950 678.600 271.050 679.050 ;
        RECT 253.950 677.400 271.050 678.600 ;
        RECT 253.950 676.800 256.050 677.400 ;
        RECT 268.950 676.950 271.050 677.400 ;
        RECT 277.950 678.600 280.050 678.900 ;
        RECT 298.950 678.600 301.050 678.900 ;
        RECT 277.950 677.400 301.050 678.600 ;
        RECT 277.950 676.800 280.050 677.400 ;
        RECT 298.950 676.800 301.050 677.400 ;
        RECT 337.950 677.400 342.600 679.050 ;
        RECT 358.950 678.450 361.050 678.900 ;
        RECT 367.950 678.450 370.050 678.900 ;
        RECT 337.950 676.950 342.000 677.400 ;
        RECT 358.950 677.250 370.050 678.450 ;
        RECT 358.950 676.800 361.050 677.250 ;
        RECT 367.950 676.800 370.050 677.250 ;
        RECT 439.950 678.600 442.050 678.900 ;
        RECT 454.950 678.600 457.050 678.900 ;
        RECT 439.950 678.450 457.050 678.600 ;
        RECT 460.950 678.450 463.050 678.900 ;
        RECT 439.950 677.400 463.050 678.450 ;
        RECT 439.950 676.800 442.050 677.400 ;
        RECT 454.950 677.250 463.050 677.400 ;
        RECT 454.950 676.800 457.050 677.250 ;
        RECT 460.950 676.800 463.050 677.250 ;
        RECT 502.950 678.450 505.050 678.900 ;
        RECT 508.950 678.450 511.050 678.900 ;
        RECT 502.950 677.250 511.050 678.450 ;
        RECT 502.950 676.800 505.050 677.250 ;
        RECT 508.950 676.800 511.050 677.250 ;
        RECT 520.950 678.600 523.050 679.050 ;
        RECT 529.950 678.600 532.050 679.050 ;
        RECT 520.950 677.400 532.050 678.600 ;
        RECT 554.400 677.400 559.050 679.050 ;
        RECT 566.400 678.900 567.600 683.400 ;
        RECT 568.950 683.550 577.050 684.750 ;
        RECT 568.950 683.100 571.050 683.550 ;
        RECT 574.950 683.100 577.050 683.550 ;
        RECT 586.950 683.100 589.050 685.200 ;
        RECT 592.950 684.750 595.050 685.200 ;
        RECT 601.950 684.750 604.050 685.200 ;
        RECT 592.950 684.600 604.050 684.750 ;
        RECT 607.950 684.600 610.050 685.050 ;
        RECT 592.950 683.550 610.050 684.600 ;
        RECT 592.950 683.100 595.050 683.550 ;
        RECT 601.950 683.400 610.050 683.550 ;
        RECT 601.950 683.100 604.050 683.400 ;
        RECT 520.950 676.950 523.050 677.400 ;
        RECT 529.950 676.950 532.050 677.400 ;
        RECT 555.000 676.950 559.050 677.400 ;
        RECT 565.950 676.800 568.050 678.900 ;
        RECT 580.950 678.600 583.050 679.050 ;
        RECT 587.400 678.600 588.600 683.100 ;
        RECT 607.950 682.950 610.050 683.400 ;
        RECT 616.950 684.600 619.050 685.050 ;
        RECT 637.950 684.600 640.050 685.200 ;
        RECT 616.950 683.400 640.050 684.600 ;
        RECT 616.950 682.950 619.050 683.400 ;
        RECT 637.950 683.100 640.050 683.400 ;
        RECT 643.950 684.600 646.050 685.050 ;
        RECT 689.400 684.600 690.600 686.400 ;
        RECT 703.950 685.950 706.050 686.400 ;
        RECT 787.950 687.600 790.050 688.050 ;
        RECT 820.950 687.600 823.050 688.050 ;
        RECT 826.950 687.600 829.050 688.050 ;
        RECT 787.950 686.400 829.050 687.600 ;
        RECT 787.950 685.950 790.050 686.400 ;
        RECT 820.950 685.950 823.050 686.400 ;
        RECT 826.950 685.950 829.050 686.400 ;
        RECT 922.950 685.950 925.050 688.050 ;
        RECT 643.950 683.400 690.600 684.600 ;
        RECT 691.950 684.750 694.050 685.200 ;
        RECT 697.950 684.750 700.050 685.200 ;
        RECT 691.950 683.550 700.050 684.750 ;
        RECT 643.950 682.950 646.050 683.400 ;
        RECT 691.950 683.100 694.050 683.550 ;
        RECT 697.950 683.100 700.050 683.550 ;
        RECT 718.950 683.100 721.050 685.200 ;
        RECT 742.950 684.600 745.050 685.200 ;
        RECT 760.950 684.600 763.050 685.200 ;
        RECT 742.950 683.400 763.050 684.600 ;
        RECT 742.950 683.100 745.050 683.400 ;
        RECT 760.950 683.100 763.050 683.400 ;
        RECT 719.400 681.600 720.600 683.100 ;
        RECT 781.950 682.950 784.050 685.050 ;
        RECT 775.950 681.600 778.050 682.050 ;
        RECT 782.400 681.600 783.600 682.950 ;
        RECT 793.950 681.600 796.050 685.050 ;
        RECT 799.950 684.750 802.050 685.200 ;
        RECT 805.950 684.750 808.050 685.200 ;
        RECT 799.950 683.550 808.050 684.750 ;
        RECT 799.950 683.100 802.050 683.550 ;
        RECT 805.950 683.100 808.050 683.550 ;
        RECT 853.950 684.750 856.050 685.200 ;
        RECT 865.950 684.750 868.050 685.200 ;
        RECT 853.950 684.600 868.050 684.750 ;
        RECT 880.800 684.600 882.900 685.200 ;
        RECT 853.950 683.550 882.900 684.600 ;
        RECT 853.950 683.100 856.050 683.550 ;
        RECT 865.950 683.400 882.900 683.550 ;
        RECT 865.950 683.100 868.050 683.400 ;
        RECT 880.800 683.100 882.900 683.400 ;
        RECT 719.400 680.400 778.050 681.600 ;
        RECT 779.400 681.000 796.050 681.600 ;
        RECT 800.400 681.600 801.600 683.100 ;
        RECT 883.950 682.950 886.050 685.050 ;
        RECT 913.950 684.600 916.050 685.050 ;
        RECT 919.950 684.600 922.050 685.200 ;
        RECT 913.950 683.400 922.050 684.600 ;
        RECT 913.950 682.950 916.050 683.400 ;
        RECT 919.950 683.100 922.050 683.400 ;
        RECT 775.950 679.950 778.050 680.400 ;
        RECT 778.950 680.400 795.600 681.000 ;
        RECT 800.400 680.400 831.600 681.600 ;
        RECT 580.950 677.400 588.600 678.600 ;
        RECT 589.950 678.600 592.050 678.900 ;
        RECT 604.950 678.600 607.050 679.050 ;
        RECT 589.950 677.400 607.050 678.600 ;
        RECT 580.950 676.950 583.050 677.400 ;
        RECT 589.950 676.800 592.050 677.400 ;
        RECT 604.950 676.950 607.050 677.400 ;
        RECT 667.950 678.450 670.050 678.900 ;
        RECT 676.950 678.450 679.050 678.900 ;
        RECT 667.950 677.250 679.050 678.450 ;
        RECT 667.950 676.800 670.050 677.250 ;
        RECT 676.950 676.800 679.050 677.250 ;
        RECT 715.950 678.600 718.050 678.900 ;
        RECT 748.950 678.600 751.050 679.050 ;
        RECT 763.950 678.600 766.050 678.900 ;
        RECT 715.950 677.400 747.600 678.600 ;
        RECT 715.950 676.800 718.050 677.400 ;
        RECT 22.950 675.600 25.050 676.050 ;
        RECT 37.950 675.600 40.050 676.050 ;
        RECT 22.950 674.400 40.050 675.600 ;
        RECT 22.950 673.950 25.050 674.400 ;
        RECT 37.950 673.950 40.050 674.400 ;
        RECT 217.950 675.600 220.050 676.050 ;
        RECT 229.950 675.600 232.050 676.050 ;
        RECT 217.950 674.400 232.050 675.600 ;
        RECT 217.950 673.950 220.050 674.400 ;
        RECT 229.950 673.950 232.050 674.400 ;
        RECT 493.950 675.600 496.050 676.050 ;
        RECT 514.950 675.600 517.050 676.050 ;
        RECT 493.950 674.400 517.050 675.600 ;
        RECT 493.950 673.950 496.050 674.400 ;
        RECT 514.950 673.950 517.050 674.400 ;
        RECT 523.950 675.600 526.050 676.050 ;
        RECT 538.950 675.600 541.050 676.050 ;
        RECT 523.950 674.400 541.050 675.600 ;
        RECT 523.950 673.950 526.050 674.400 ;
        RECT 538.950 673.950 541.050 674.400 ;
        RECT 613.950 675.600 616.050 676.050 ;
        RECT 625.950 675.600 628.050 676.050 ;
        RECT 613.950 674.400 628.050 675.600 ;
        RECT 746.400 675.600 747.600 677.400 ;
        RECT 748.950 678.450 766.050 678.600 ;
        RECT 769.950 678.450 772.050 678.900 ;
        RECT 748.950 677.400 772.050 678.450 ;
        RECT 748.950 676.950 751.050 677.400 ;
        RECT 763.950 677.250 772.050 677.400 ;
        RECT 763.950 676.800 766.050 677.250 ;
        RECT 769.950 676.800 772.050 677.250 ;
        RECT 778.950 676.950 781.050 680.400 ;
        RECT 830.400 678.900 831.600 680.400 ;
        RECT 829.950 676.800 832.050 678.900 ;
        RECT 835.950 678.450 838.050 678.900 ;
        RECT 862.950 678.450 865.050 679.050 ;
        RECT 871.950 678.450 874.050 678.900 ;
        RECT 835.950 677.250 874.050 678.450 ;
        RECT 835.950 676.800 838.050 677.250 ;
        RECT 862.950 676.950 865.050 677.250 ;
        RECT 871.950 676.800 874.050 677.250 ;
        RECT 784.950 675.600 787.050 676.050 ;
        RECT 799.950 675.600 802.050 676.050 ;
        RECT 746.400 674.400 802.050 675.600 ;
        RECT 613.950 673.950 616.050 674.400 ;
        RECT 625.950 673.950 628.050 674.400 ;
        RECT 784.950 673.950 787.050 674.400 ;
        RECT 799.950 673.950 802.050 674.400 ;
        RECT 808.950 675.600 811.050 676.050 ;
        RECT 820.950 675.600 823.050 676.050 ;
        RECT 808.950 674.400 823.050 675.600 ;
        RECT 808.950 673.950 811.050 674.400 ;
        RECT 820.950 673.950 823.050 674.400 ;
        RECT 874.950 675.600 877.050 676.050 ;
        RECT 884.400 675.600 885.600 682.950 ;
        RECT 923.400 678.900 924.600 685.950 ;
        RECT 928.950 684.750 931.050 685.200 ;
        RECT 940.950 684.750 943.050 685.200 ;
        RECT 928.950 683.550 943.050 684.750 ;
        RECT 928.950 683.100 931.050 683.550 ;
        RECT 940.950 683.100 943.050 683.550 ;
        RECT 979.800 684.000 981.900 685.050 ;
        RECT 979.800 682.950 982.050 684.000 ;
        RECT 982.950 683.100 985.050 685.200 ;
        RECT 979.950 681.600 982.050 682.950 ;
        RECT 956.400 681.000 982.050 681.600 ;
        RECT 983.400 681.600 984.600 683.100 ;
        RECT 956.400 680.400 981.450 681.000 ;
        RECT 983.400 680.400 990.600 681.600 ;
        RECT 922.950 676.800 925.050 678.900 ;
        RECT 934.950 678.600 937.050 678.900 ;
        RECT 956.400 678.600 957.600 680.400 ;
        RECT 934.950 677.400 957.600 678.600 ;
        RECT 958.950 678.450 961.050 678.900 ;
        RECT 985.950 678.450 988.050 678.900 ;
        RECT 934.950 676.800 937.050 677.400 ;
        RECT 958.950 677.250 988.050 678.450 ;
        RECT 958.950 676.800 961.050 677.250 ;
        RECT 985.950 676.800 988.050 677.250 ;
        RECT 989.400 676.050 990.600 680.400 ;
        RECT 987.000 675.750 990.600 676.050 ;
        RECT 874.950 674.400 885.600 675.600 ;
        RECT 985.950 674.400 990.600 675.750 ;
        RECT 991.950 675.600 994.050 676.050 ;
        RECT 1016.400 675.600 1017.600 688.950 ;
        RECT 991.950 674.400 1017.600 675.600 ;
        RECT 874.950 673.950 877.050 674.400 ;
        RECT 985.950 673.950 990.000 674.400 ;
        RECT 991.950 673.950 994.050 674.400 ;
        RECT 985.950 673.650 988.050 673.950 ;
        RECT 40.950 672.600 43.050 673.050 ;
        RECT 49.950 672.600 52.050 673.050 ;
        RECT 40.950 671.400 52.050 672.600 ;
        RECT 40.950 670.950 43.050 671.400 ;
        RECT 49.950 670.950 52.050 671.400 ;
        RECT 58.950 672.600 61.050 673.050 ;
        RECT 67.950 672.600 70.050 673.050 ;
        RECT 58.950 671.400 70.050 672.600 ;
        RECT 58.950 670.950 61.050 671.400 ;
        RECT 67.950 670.950 70.050 671.400 ;
        RECT 118.950 672.600 121.050 673.050 ;
        RECT 136.950 672.600 139.050 673.050 ;
        RECT 118.950 671.400 139.050 672.600 ;
        RECT 118.950 670.950 121.050 671.400 ;
        RECT 136.950 670.950 139.050 671.400 ;
        RECT 349.950 672.600 352.050 673.050 ;
        RECT 355.950 672.600 358.050 673.050 ;
        RECT 409.950 672.600 412.050 673.050 ;
        RECT 349.950 671.400 412.050 672.600 ;
        RECT 349.950 670.950 352.050 671.400 ;
        RECT 355.950 670.950 358.050 671.400 ;
        RECT 409.950 670.950 412.050 671.400 ;
        RECT 448.950 672.600 451.050 673.050 ;
        RECT 466.950 672.600 469.050 673.050 ;
        RECT 487.950 672.600 490.050 673.050 ;
        RECT 448.950 671.400 490.050 672.600 ;
        RECT 448.950 670.950 451.050 671.400 ;
        RECT 466.950 670.950 469.050 671.400 ;
        RECT 487.950 670.950 490.050 671.400 ;
        RECT 568.950 672.600 571.050 673.050 ;
        RECT 634.950 672.600 637.050 673.050 ;
        RECT 568.950 671.400 637.050 672.600 ;
        RECT 568.950 670.950 571.050 671.400 ;
        RECT 634.950 670.950 637.050 671.400 ;
        RECT 724.950 672.600 727.050 673.050 ;
        RECT 745.950 672.600 748.050 673.050 ;
        RECT 724.950 671.400 748.050 672.600 ;
        RECT 724.950 670.950 727.050 671.400 ;
        RECT 745.950 670.950 748.050 671.400 ;
        RECT 835.950 672.600 838.050 673.050 ;
        RECT 916.950 672.600 919.050 673.050 ;
        RECT 922.950 672.600 925.050 673.050 ;
        RECT 835.950 671.400 925.050 672.600 ;
        RECT 835.950 670.950 838.050 671.400 ;
        RECT 916.950 670.950 919.050 671.400 ;
        RECT 922.950 670.950 925.050 671.400 ;
        RECT 994.950 672.600 997.050 673.050 ;
        RECT 1009.950 672.600 1012.050 673.050 ;
        RECT 994.950 671.400 1012.050 672.600 ;
        RECT 994.950 670.950 997.050 671.400 ;
        RECT 1009.950 670.950 1012.050 671.400 ;
        RECT 109.950 669.600 112.050 670.050 ;
        RECT 160.950 669.600 163.050 670.050 ;
        RECT 205.950 669.600 208.050 670.050 ;
        RECT 109.950 668.400 208.050 669.600 ;
        RECT 109.950 667.950 112.050 668.400 ;
        RECT 160.950 667.950 163.050 668.400 ;
        RECT 205.950 667.950 208.050 668.400 ;
        RECT 217.950 669.600 220.050 670.050 ;
        RECT 226.950 669.600 229.050 670.050 ;
        RECT 217.950 668.400 229.050 669.600 ;
        RECT 217.950 667.950 220.050 668.400 ;
        RECT 226.950 667.950 229.050 668.400 ;
        RECT 337.950 669.600 340.050 670.050 ;
        RECT 346.950 669.600 349.050 670.050 ;
        RECT 337.950 668.400 349.050 669.600 ;
        RECT 337.950 667.950 340.050 668.400 ;
        RECT 346.950 667.950 349.050 668.400 ;
        RECT 403.950 669.600 406.050 670.050 ;
        RECT 415.950 669.600 418.050 670.050 ;
        RECT 403.950 668.400 418.050 669.600 ;
        RECT 403.950 667.950 406.050 668.400 ;
        RECT 415.950 667.950 418.050 668.400 ;
        RECT 499.950 669.600 502.050 670.050 ;
        RECT 532.950 669.600 535.050 670.050 ;
        RECT 559.950 669.600 562.050 670.050 ;
        RECT 499.950 668.400 562.050 669.600 ;
        RECT 635.400 669.600 636.600 670.950 ;
        RECT 691.950 669.600 694.050 670.050 ;
        RECT 709.950 669.600 712.050 670.050 ;
        RECT 635.400 668.400 712.050 669.600 ;
        RECT 499.950 667.950 502.050 668.400 ;
        RECT 532.950 667.950 535.050 668.400 ;
        RECT 559.950 667.950 562.050 668.400 ;
        RECT 691.950 667.950 694.050 668.400 ;
        RECT 709.950 667.950 712.050 668.400 ;
        RECT 790.950 669.600 793.050 670.050 ;
        RECT 826.950 669.600 829.050 670.050 ;
        RECT 790.950 668.400 829.050 669.600 ;
        RECT 790.950 667.950 793.050 668.400 ;
        RECT 826.950 667.950 829.050 668.400 ;
        RECT 871.950 669.600 874.050 670.050 ;
        RECT 895.950 669.600 898.050 670.050 ;
        RECT 871.950 668.400 898.050 669.600 ;
        RECT 871.950 667.950 874.050 668.400 ;
        RECT 895.950 667.950 898.050 668.400 ;
        RECT 952.950 669.600 955.050 670.050 ;
        RECT 976.950 669.600 979.050 670.050 ;
        RECT 952.950 668.400 979.050 669.600 ;
        RECT 952.950 667.950 955.050 668.400 ;
        RECT 976.950 667.950 979.050 668.400 ;
        RECT 49.950 666.600 52.050 667.050 ;
        RECT 103.950 666.600 106.050 667.050 ;
        RECT 49.950 665.400 106.050 666.600 ;
        RECT 49.950 664.950 52.050 665.400 ;
        RECT 103.950 664.950 106.050 665.400 ;
        RECT 265.950 666.600 268.050 667.050 ;
        RECT 304.950 666.600 307.050 667.050 ;
        RECT 334.950 666.600 337.050 667.050 ;
        RECT 265.950 665.400 337.050 666.600 ;
        RECT 265.950 664.950 268.050 665.400 ;
        RECT 304.950 664.950 307.050 665.400 ;
        RECT 334.950 664.950 337.050 665.400 ;
        RECT 385.950 666.600 388.050 667.050 ;
        RECT 424.950 666.600 427.050 667.050 ;
        RECT 385.950 665.400 427.050 666.600 ;
        RECT 385.950 664.950 388.050 665.400 ;
        RECT 424.950 664.950 427.050 665.400 ;
        RECT 493.950 666.600 496.050 667.050 ;
        RECT 577.950 666.600 580.050 667.050 ;
        RECT 493.950 665.400 580.050 666.600 ;
        RECT 493.950 664.950 496.050 665.400 ;
        RECT 577.950 664.950 580.050 665.400 ;
        RECT 664.950 666.600 667.050 667.050 ;
        RECT 676.950 666.600 679.050 667.050 ;
        RECT 664.950 665.400 679.050 666.600 ;
        RECT 664.950 664.950 667.050 665.400 ;
        RECT 676.950 664.950 679.050 665.400 ;
        RECT 763.950 666.600 766.050 667.050 ;
        RECT 778.950 666.600 781.050 667.050 ;
        RECT 763.950 665.400 781.050 666.600 ;
        RECT 763.950 664.950 766.050 665.400 ;
        RECT 778.950 664.950 781.050 665.400 ;
        RECT 829.950 666.600 832.050 667.050 ;
        RECT 868.950 666.600 871.050 667.050 ;
        RECT 829.950 665.400 871.050 666.600 ;
        RECT 829.950 664.950 832.050 665.400 ;
        RECT 868.950 664.950 871.050 665.400 ;
        RECT 919.950 666.600 922.050 667.050 ;
        RECT 928.950 666.600 931.050 667.050 ;
        RECT 919.950 665.400 931.050 666.600 ;
        RECT 919.950 664.950 922.050 665.400 ;
        RECT 928.950 664.950 931.050 665.400 ;
        RECT 949.950 666.600 952.050 667.050 ;
        RECT 958.950 666.600 961.050 667.050 ;
        RECT 949.950 665.400 961.050 666.600 ;
        RECT 949.950 664.950 952.050 665.400 ;
        RECT 958.950 664.950 961.050 665.400 ;
        RECT 988.950 666.600 991.050 667.050 ;
        RECT 1009.950 666.600 1012.050 667.050 ;
        RECT 988.950 665.400 1012.050 666.600 ;
        RECT 988.950 664.950 991.050 665.400 ;
        RECT 1009.950 664.950 1012.050 665.400 ;
        RECT 97.950 663.600 100.050 664.050 ;
        RECT 124.950 663.600 127.050 664.050 ;
        RECT 97.950 662.400 127.050 663.600 ;
        RECT 97.950 661.950 100.050 662.400 ;
        RECT 124.950 661.950 127.050 662.400 ;
        RECT 181.950 663.600 184.050 664.050 ;
        RECT 211.950 663.600 214.050 664.050 ;
        RECT 181.950 662.400 214.050 663.600 ;
        RECT 181.950 661.950 184.050 662.400 ;
        RECT 211.950 661.950 214.050 662.400 ;
        RECT 361.950 663.600 364.050 664.050 ;
        RECT 370.950 663.600 373.050 664.050 ;
        RECT 361.950 662.400 373.050 663.600 ;
        RECT 361.950 661.950 364.050 662.400 ;
        RECT 370.950 661.950 373.050 662.400 ;
        RECT 382.950 663.600 385.050 664.050 ;
        RECT 394.950 663.600 397.050 664.050 ;
        RECT 382.950 662.400 397.050 663.600 ;
        RECT 382.950 661.950 385.050 662.400 ;
        RECT 394.950 661.950 397.050 662.400 ;
        RECT 406.950 663.600 409.050 664.050 ;
        RECT 439.950 663.600 442.050 664.050 ;
        RECT 406.950 662.400 442.050 663.600 ;
        RECT 406.950 661.950 409.050 662.400 ;
        RECT 439.950 661.950 442.050 662.400 ;
        RECT 514.950 663.600 517.050 664.050 ;
        RECT 541.950 663.600 544.050 664.050 ;
        RECT 550.800 663.600 552.900 664.050 ;
        RECT 514.950 662.400 552.900 663.600 ;
        RECT 514.950 661.950 517.050 662.400 ;
        RECT 541.950 661.950 544.050 662.400 ;
        RECT 550.800 661.950 552.900 662.400 ;
        RECT 598.950 663.600 601.050 664.050 ;
        RECT 622.950 663.600 625.050 664.050 ;
        RECT 598.950 662.400 625.050 663.600 ;
        RECT 598.950 661.950 601.050 662.400 ;
        RECT 622.950 661.950 625.050 662.400 ;
        RECT 628.950 663.600 631.050 664.050 ;
        RECT 652.950 663.600 655.050 664.050 ;
        RECT 628.950 662.400 655.050 663.600 ;
        RECT 628.950 661.950 631.050 662.400 ;
        RECT 652.950 661.950 655.050 662.400 ;
        RECT 814.950 663.600 817.050 664.050 ;
        RECT 820.950 663.600 823.050 664.050 ;
        RECT 850.950 663.600 853.050 664.050 ;
        RECT 814.950 662.400 853.050 663.600 ;
        RECT 814.950 661.950 817.050 662.400 ;
        RECT 820.950 661.950 823.050 662.400 ;
        RECT 850.950 661.950 853.050 662.400 ;
        RECT 964.950 663.600 967.050 664.050 ;
        RECT 970.950 663.600 973.050 664.050 ;
        RECT 964.950 662.400 973.050 663.600 ;
        RECT 964.950 661.950 967.050 662.400 ;
        RECT 970.950 661.950 973.050 662.400 ;
        RECT 49.950 660.600 52.050 661.050 ;
        RECT 70.950 660.600 73.050 661.050 ;
        RECT 49.950 659.400 73.050 660.600 ;
        RECT 49.950 658.950 52.050 659.400 ;
        RECT 70.950 658.950 73.050 659.400 ;
        RECT 244.950 660.600 247.050 661.050 ;
        RECT 250.950 660.600 253.050 661.050 ;
        RECT 274.950 660.600 277.050 661.050 ;
        RECT 244.950 659.400 277.050 660.600 ;
        RECT 244.950 658.950 247.050 659.400 ;
        RECT 250.950 658.950 253.050 659.400 ;
        RECT 274.950 658.950 277.050 659.400 ;
        RECT 445.950 660.600 448.050 661.050 ;
        RECT 475.950 660.600 478.050 661.050 ;
        RECT 445.950 659.400 478.050 660.600 ;
        RECT 445.950 658.950 448.050 659.400 ;
        RECT 475.950 658.950 478.050 659.400 ;
        RECT 625.950 660.600 628.050 661.050 ;
        RECT 640.950 660.600 643.050 661.050 ;
        RECT 733.950 660.600 736.050 661.050 ;
        RECT 625.950 659.400 643.050 660.600 ;
        RECT 625.950 658.950 628.050 659.400 ;
        RECT 640.950 658.950 643.050 659.400 ;
        RECT 683.400 659.400 736.050 660.600 ;
        RECT 145.950 657.600 148.050 658.050 ;
        RECT 193.950 657.600 196.050 658.050 ;
        RECT 145.950 656.400 196.050 657.600 ;
        RECT 145.950 655.950 148.050 656.400 ;
        RECT 193.950 655.950 196.050 656.400 ;
        RECT 427.950 657.600 430.050 658.050 ;
        RECT 502.950 657.600 505.050 658.050 ;
        RECT 427.950 656.400 505.050 657.600 ;
        RECT 427.950 655.950 430.050 656.400 ;
        RECT 502.950 655.950 505.050 656.400 ;
        RECT 556.950 657.600 559.050 658.050 ;
        RECT 583.950 657.600 586.050 658.050 ;
        RECT 556.950 656.400 586.050 657.600 ;
        RECT 556.950 655.950 559.050 656.400 ;
        RECT 583.950 655.950 586.050 656.400 ;
        RECT 616.950 657.600 619.050 658.050 ;
        RECT 631.950 657.600 634.050 658.050 ;
        RECT 616.950 656.400 634.050 657.600 ;
        RECT 616.950 655.950 619.050 656.400 ;
        RECT 631.950 655.950 634.050 656.400 ;
        RECT 652.950 657.600 655.050 658.050 ;
        RECT 683.400 657.600 684.600 659.400 ;
        RECT 733.950 658.950 736.050 659.400 ;
        RECT 739.950 660.600 742.050 661.050 ;
        RECT 745.950 660.600 748.050 661.050 ;
        RECT 844.950 660.600 847.050 661.050 ;
        RECT 739.950 659.400 847.050 660.600 ;
        RECT 739.950 658.950 742.050 659.400 ;
        RECT 745.950 658.950 748.050 659.400 ;
        RECT 844.950 658.950 847.050 659.400 ;
        RECT 904.950 660.600 907.050 661.050 ;
        RECT 922.950 660.600 925.050 661.050 ;
        RECT 904.950 659.400 925.050 660.600 ;
        RECT 904.950 658.950 907.050 659.400 ;
        RECT 922.950 658.950 925.050 659.400 ;
        RECT 934.950 660.600 937.050 661.050 ;
        RECT 955.950 660.600 958.050 661.050 ;
        RECT 934.950 659.400 958.050 660.600 ;
        RECT 934.950 658.950 937.050 659.400 ;
        RECT 955.950 658.950 958.050 659.400 ;
        RECT 976.950 660.600 979.050 661.050 ;
        RECT 991.950 660.600 994.050 661.050 ;
        RECT 976.950 659.400 994.050 660.600 ;
        RECT 976.950 658.950 979.050 659.400 ;
        RECT 991.950 658.950 994.050 659.400 ;
        RECT 652.950 656.400 684.600 657.600 ;
        RECT 811.950 657.600 814.050 658.050 ;
        RECT 838.950 657.600 841.050 658.050 ;
        RECT 811.950 656.400 841.050 657.600 ;
        RECT 652.950 655.950 655.050 656.400 ;
        RECT 811.950 655.950 814.050 656.400 ;
        RECT 838.950 655.950 841.050 656.400 ;
        RECT 877.950 657.600 880.050 658.050 ;
        RECT 889.950 657.600 892.050 657.900 ;
        RECT 877.950 656.400 892.050 657.600 ;
        RECT 877.950 655.950 880.050 656.400 ;
        RECT 889.950 655.800 892.050 656.400 ;
        RECT 901.950 657.600 904.050 658.050 ;
        RECT 910.950 657.600 913.050 658.050 ;
        RECT 931.950 657.600 934.050 658.050 ;
        RECT 943.950 657.600 946.050 658.050 ;
        RECT 901.950 656.400 946.050 657.600 ;
        RECT 901.950 655.950 904.050 656.400 ;
        RECT 910.950 655.950 913.050 656.400 ;
        RECT 931.950 655.950 934.050 656.400 ;
        RECT 943.950 655.950 946.050 656.400 ;
        RECT 967.950 657.600 970.050 657.900 ;
        RECT 982.950 657.600 985.050 658.050 ;
        RECT 967.950 656.400 985.050 657.600 ;
        RECT 967.950 655.800 970.050 656.400 ;
        RECT 982.950 655.950 985.050 656.400 ;
        RECT 4.950 654.600 7.050 655.050 ;
        RECT 16.950 654.600 19.050 655.050 ;
        RECT 28.950 654.600 31.050 655.050 ;
        RECT 4.950 653.400 31.050 654.600 ;
        RECT 4.950 652.950 7.050 653.400 ;
        RECT 16.950 652.950 19.050 653.400 ;
        RECT 28.950 652.950 31.050 653.400 ;
        RECT 133.950 654.600 136.050 655.050 ;
        RECT 139.950 654.600 142.050 655.050 ;
        RECT 133.950 653.400 142.050 654.600 ;
        RECT 133.950 652.950 136.050 653.400 ;
        RECT 139.950 652.950 142.050 653.400 ;
        RECT 271.950 654.600 274.050 655.050 ;
        RECT 283.950 654.600 286.050 655.050 ;
        RECT 400.950 654.600 403.050 655.050 ;
        RECT 271.950 653.400 403.050 654.600 ;
        RECT 271.950 652.950 274.050 653.400 ;
        RECT 283.950 652.950 286.050 653.400 ;
        RECT 400.950 652.950 403.050 653.400 ;
        RECT 430.950 654.600 433.050 655.050 ;
        RECT 463.950 654.600 466.050 655.050 ;
        RECT 643.950 654.600 646.050 655.050 ;
        RECT 430.950 653.400 466.050 654.600 ;
        RECT 430.950 652.950 433.050 653.400 ;
        RECT 463.950 652.950 466.050 653.400 ;
        RECT 620.400 653.400 646.050 654.600 ;
        RECT 37.950 651.600 40.050 652.200 ;
        RECT 46.950 651.600 49.050 652.050 ;
        RECT 37.950 650.400 49.050 651.600 ;
        RECT 37.950 650.100 40.050 650.400 ;
        RECT 46.950 649.950 49.050 650.400 ;
        RECT 58.950 650.100 61.050 652.200 ;
        RECT 64.950 651.600 67.050 652.200 ;
        RECT 85.950 651.600 88.050 652.050 ;
        RECT 64.950 650.400 88.050 651.600 ;
        RECT 64.950 650.100 67.050 650.400 ;
        RECT 59.400 648.600 60.600 650.100 ;
        RECT 85.950 649.950 88.050 650.400 ;
        RECT 106.950 651.750 109.050 652.200 ;
        RECT 118.950 651.750 121.050 652.200 ;
        RECT 106.950 650.550 121.050 651.750 ;
        RECT 106.950 650.100 109.050 650.550 ;
        RECT 118.950 650.100 121.050 650.550 ;
        RECT 124.950 651.750 127.050 652.200 ;
        RECT 130.950 651.750 133.050 652.200 ;
        RECT 124.950 650.550 133.050 651.750 ;
        RECT 124.950 650.100 127.050 650.550 ;
        RECT 130.950 650.100 133.050 650.550 ;
        RECT 154.950 651.600 157.050 652.050 ;
        RECT 169.950 651.600 172.050 652.200 ;
        RECT 205.950 651.600 208.050 652.200 ;
        RECT 217.950 651.600 220.050 652.050 ;
        RECT 223.950 651.600 226.050 652.200 ;
        RECT 154.950 650.400 172.050 651.600 ;
        RECT 107.400 648.600 108.600 650.100 ;
        RECT 154.950 649.950 157.050 650.400 ;
        RECT 169.950 650.100 172.050 650.400 ;
        RECT 173.400 650.400 226.050 651.600 ;
        RECT 59.400 647.400 108.600 648.600 ;
        RECT 28.950 645.450 31.050 645.900 ;
        RECT 34.950 645.450 37.050 645.900 ;
        RECT 28.950 644.250 37.050 645.450 ;
        RECT 28.950 643.800 31.050 644.250 ;
        RECT 34.950 643.800 37.050 644.250 ;
        RECT 40.950 645.600 43.050 645.900 ;
        RECT 49.950 645.600 52.050 646.050 ;
        RECT 173.400 645.900 174.600 650.400 ;
        RECT 205.950 650.100 208.050 650.400 ;
        RECT 217.950 649.950 220.050 650.400 ;
        RECT 223.950 650.100 226.050 650.400 ;
        RECT 241.950 651.600 244.050 652.050 ;
        RECT 259.950 651.600 262.050 652.200 ;
        RECT 241.950 650.400 262.050 651.600 ;
        RECT 241.950 649.950 244.050 650.400 ;
        RECT 259.950 650.100 262.050 650.400 ;
        RECT 295.950 651.750 298.050 652.200 ;
        RECT 331.950 651.750 334.050 652.200 ;
        RECT 295.950 650.550 334.050 651.750 ;
        RECT 402.000 651.600 406.050 652.050 ;
        RECT 295.950 650.100 298.050 650.550 ;
        RECT 331.950 650.100 334.050 650.550 ;
        RECT 401.400 649.950 406.050 651.600 ;
        RECT 418.950 650.100 421.050 652.200 ;
        RECT 328.950 648.600 331.050 649.050 ;
        RECT 314.400 647.400 331.050 648.600 ;
        RECT 40.950 644.400 52.050 645.600 ;
        RECT 40.950 643.800 43.050 644.400 ;
        RECT 49.950 643.950 52.050 644.400 ;
        RECT 79.950 645.450 82.050 645.900 ;
        RECT 85.950 645.450 88.050 645.900 ;
        RECT 121.950 645.600 124.050 645.900 ;
        RECT 79.950 644.250 88.050 645.450 ;
        RECT 79.950 643.800 82.050 644.250 ;
        RECT 85.950 643.800 88.050 644.250 ;
        RECT 89.400 644.400 124.050 645.600 ;
        RECT 13.950 642.600 16.050 643.050 ;
        RECT 22.950 642.600 25.050 643.050 ;
        RECT 13.950 641.400 25.050 642.600 ;
        RECT 13.950 640.950 16.050 641.400 ;
        RECT 22.950 640.950 25.050 641.400 ;
        RECT 61.950 642.600 64.050 643.050 ;
        RECT 89.400 642.600 90.600 644.400 ;
        RECT 121.950 643.800 124.050 644.400 ;
        RECT 148.950 645.450 151.050 645.900 ;
        RECT 154.950 645.450 157.050 645.900 ;
        RECT 148.950 644.250 157.050 645.450 ;
        RECT 148.950 643.800 151.050 644.250 ;
        RECT 154.950 643.800 157.050 644.250 ;
        RECT 172.950 643.800 175.050 645.900 ;
        RECT 187.950 645.450 190.050 645.900 ;
        RECT 193.950 645.450 196.050 645.900 ;
        RECT 187.950 644.250 196.050 645.450 ;
        RECT 187.950 643.800 190.050 644.250 ;
        RECT 193.950 643.800 196.050 644.250 ;
        RECT 250.950 645.450 253.050 645.900 ;
        RECT 256.950 645.450 259.050 645.900 ;
        RECT 250.950 644.250 259.050 645.450 ;
        RECT 250.950 643.800 253.050 644.250 ;
        RECT 256.950 643.800 259.050 644.250 ;
        RECT 274.950 645.600 277.050 646.050 ;
        RECT 314.400 645.900 315.600 647.400 ;
        RECT 328.950 646.950 331.050 647.400 ;
        RECT 401.400 645.900 402.600 649.950 ;
        RECT 419.400 648.600 420.600 650.100 ;
        RECT 430.950 648.600 433.050 649.050 ;
        RECT 419.400 647.400 433.050 648.600 ;
        RECT 433.950 648.600 436.050 652.050 ;
        RECT 517.950 651.600 520.050 652.200 ;
        RECT 529.950 651.600 532.050 652.050 ;
        RECT 517.950 650.400 532.050 651.600 ;
        RECT 517.950 650.100 520.050 650.400 ;
        RECT 529.950 649.950 532.050 650.400 ;
        RECT 589.950 651.750 592.050 652.200 ;
        RECT 598.950 651.750 601.050 652.200 ;
        RECT 589.950 650.550 601.050 651.750 ;
        RECT 589.950 650.100 592.050 650.550 ;
        RECT 598.950 650.100 601.050 650.550 ;
        RECT 604.950 651.600 607.050 652.050 ;
        RECT 620.400 651.600 621.600 653.400 ;
        RECT 643.950 652.950 646.050 653.400 ;
        RECT 670.950 654.600 673.050 655.050 ;
        RECT 685.950 654.600 688.050 655.050 ;
        RECT 670.950 653.400 688.050 654.600 ;
        RECT 670.950 652.950 673.050 653.400 ;
        RECT 685.950 652.950 688.050 653.400 ;
        RECT 730.950 654.600 733.050 655.050 ;
        RECT 742.950 654.600 745.050 655.050 ;
        RECT 730.950 653.400 745.050 654.600 ;
        RECT 730.950 652.950 733.050 653.400 ;
        RECT 742.950 652.950 745.050 653.400 ;
        RECT 757.950 654.600 760.050 655.050 ;
        RECT 784.950 654.600 787.050 655.050 ;
        RECT 757.950 653.400 787.050 654.600 ;
        RECT 757.950 652.950 760.050 653.400 ;
        RECT 784.950 652.950 787.050 653.400 ;
        RECT 907.950 652.950 910.050 655.050 ;
        RECT 928.950 652.950 931.050 655.050 ;
        RECT 964.950 654.600 967.050 655.050 ;
        RECT 959.400 653.400 967.050 654.600 ;
        RECT 604.950 650.400 621.600 651.600 ;
        RECT 622.950 651.750 625.050 652.200 ;
        RECT 628.950 651.750 631.050 652.200 ;
        RECT 622.950 650.550 631.050 651.750 ;
        RECT 604.950 649.950 607.050 650.400 ;
        RECT 622.950 650.100 625.050 650.550 ;
        RECT 628.950 650.100 631.050 650.550 ;
        RECT 646.950 650.100 649.050 652.200 ;
        RECT 658.950 651.600 661.050 652.050 ;
        RECT 682.950 651.600 685.050 652.050 ;
        RECT 658.950 650.400 685.050 651.600 ;
        RECT 433.950 648.000 444.600 648.600 ;
        RECT 434.400 647.400 444.600 648.000 ;
        RECT 430.950 646.950 433.050 647.400 ;
        RECT 443.400 645.900 444.600 647.400 ;
        RECT 286.950 645.600 289.050 645.900 ;
        RECT 274.950 644.400 289.050 645.600 ;
        RECT 274.950 643.950 277.050 644.400 ;
        RECT 286.950 643.800 289.050 644.400 ;
        RECT 313.950 643.800 316.050 645.900 ;
        RECT 331.950 645.450 334.050 645.900 ;
        RECT 343.950 645.450 346.050 645.900 ;
        RECT 331.950 644.250 346.050 645.450 ;
        RECT 331.950 643.800 334.050 644.250 ;
        RECT 343.950 643.800 346.050 644.250 ;
        RECT 364.950 645.450 367.050 645.900 ;
        RECT 370.950 645.450 373.050 645.900 ;
        RECT 364.950 644.250 373.050 645.450 ;
        RECT 364.950 643.800 367.050 644.250 ;
        RECT 370.950 643.800 373.050 644.250 ;
        RECT 400.950 643.800 403.050 645.900 ;
        RECT 442.950 643.800 445.050 645.900 ;
        RECT 490.950 645.450 493.050 645.900 ;
        RECT 505.950 645.450 508.050 645.900 ;
        RECT 490.950 644.250 508.050 645.450 ;
        RECT 490.950 643.800 493.050 644.250 ;
        RECT 505.950 643.800 508.050 644.250 ;
        RECT 514.950 645.450 517.050 645.900 ;
        RECT 532.950 645.450 535.050 645.900 ;
        RECT 514.950 644.250 535.050 645.450 ;
        RECT 514.950 643.800 517.050 644.250 ;
        RECT 532.950 643.800 535.050 644.250 ;
        RECT 592.950 645.450 595.050 645.900 ;
        RECT 607.950 645.450 610.050 645.900 ;
        RECT 592.950 644.250 610.050 645.450 ;
        RECT 592.950 643.800 595.050 644.250 ;
        RECT 607.950 643.800 610.050 644.250 ;
        RECT 61.950 641.400 90.600 642.600 ;
        RECT 142.950 642.600 145.050 643.050 ;
        RECT 166.950 642.600 169.050 643.050 ;
        RECT 142.950 641.400 169.050 642.600 ;
        RECT 61.950 640.950 64.050 641.400 ;
        RECT 142.950 640.950 145.050 641.400 ;
        RECT 166.950 640.950 169.050 641.400 ;
        RECT 640.950 642.600 643.050 643.050 ;
        RECT 647.400 642.600 648.600 650.100 ;
        RECT 658.950 649.950 661.050 650.400 ;
        RECT 682.950 649.950 685.050 650.400 ;
        RECT 712.950 651.600 715.050 652.200 ;
        RECT 724.950 651.600 727.050 652.050 ;
        RECT 712.950 650.400 727.050 651.600 ;
        RECT 712.950 650.100 715.050 650.400 ;
        RECT 724.950 649.950 727.050 650.400 ;
        RECT 751.950 649.950 754.050 652.050 ;
        RECT 766.950 651.600 769.050 652.050 ;
        RECT 778.950 651.600 781.050 652.200 ;
        RECT 766.950 650.400 781.050 651.600 ;
        RECT 766.950 649.950 769.050 650.400 ;
        RECT 778.950 650.100 781.050 650.400 ;
        RECT 784.950 651.750 787.050 652.200 ;
        RECT 793.950 651.750 796.050 652.200 ;
        RECT 784.950 651.600 796.050 651.750 ;
        RECT 805.950 651.600 808.050 652.200 ;
        RECT 784.950 650.550 808.050 651.600 ;
        RECT 784.950 650.100 787.050 650.550 ;
        RECT 793.950 650.400 808.050 650.550 ;
        RECT 793.950 650.100 796.050 650.400 ;
        RECT 805.950 650.100 808.050 650.400 ;
        RECT 752.400 645.600 753.600 649.950 ;
        RECT 823.950 648.600 826.050 652.050 ;
        RECT 841.950 651.750 844.050 652.200 ;
        RECT 856.950 651.750 859.050 652.200 ;
        RECT 841.950 650.550 859.050 651.750 ;
        RECT 841.950 650.100 844.050 650.550 ;
        RECT 856.950 650.100 859.050 650.550 ;
        RECT 862.950 651.600 865.050 652.200 ;
        RECT 871.950 651.600 874.050 652.050 ;
        RECT 880.950 651.600 883.050 652.200 ;
        RECT 862.950 650.400 883.050 651.600 ;
        RECT 862.950 650.100 865.050 650.400 ;
        RECT 871.950 649.950 874.050 650.400 ;
        RECT 880.950 650.100 883.050 650.400 ;
        RECT 886.950 651.600 889.050 652.200 ;
        RECT 898.950 651.600 901.050 652.050 ;
        RECT 886.950 650.400 901.050 651.600 ;
        RECT 886.950 650.100 889.050 650.400 ;
        RECT 898.950 649.950 901.050 650.400 ;
        RECT 815.400 648.000 826.050 648.600 ;
        RECT 814.950 647.400 825.600 648.000 ;
        RECT 760.950 645.600 763.050 645.900 ;
        RECT 752.400 644.400 763.050 645.600 ;
        RECT 760.950 643.800 763.050 644.400 ;
        RECT 787.950 645.600 790.050 645.900 ;
        RECT 802.950 645.600 805.050 645.900 ;
        RECT 787.950 644.400 805.050 645.600 ;
        RECT 787.950 643.800 790.050 644.400 ;
        RECT 802.950 643.800 805.050 644.400 ;
        RECT 814.950 643.950 817.050 647.400 ;
        RECT 820.950 645.450 823.050 645.900 ;
        RECT 826.950 645.450 829.050 645.900 ;
        RECT 820.950 644.250 829.050 645.450 ;
        RECT 820.950 643.800 823.050 644.250 ;
        RECT 826.950 643.800 829.050 644.250 ;
        RECT 832.950 645.450 835.050 645.900 ;
        RECT 841.950 645.450 844.050 645.900 ;
        RECT 832.950 644.250 844.050 645.450 ;
        RECT 832.950 643.800 835.050 644.250 ;
        RECT 841.950 643.800 844.050 644.250 ;
        RECT 847.950 645.450 850.050 645.900 ;
        RECT 853.950 645.450 856.050 645.900 ;
        RECT 847.950 644.250 856.050 645.450 ;
        RECT 847.950 643.800 850.050 644.250 ;
        RECT 853.950 643.800 856.050 644.250 ;
        RECT 859.950 645.450 862.050 645.900 ;
        RECT 871.950 645.600 874.050 645.900 ;
        RECT 908.400 645.600 909.600 652.950 ;
        RECT 915.000 651.600 919.050 652.050 ;
        RECT 914.400 649.950 919.050 651.600 ;
        RECT 914.400 645.900 915.600 649.950 ;
        RECT 929.400 648.600 930.600 652.950 ;
        RECT 937.950 651.600 940.050 652.200 ;
        RECT 959.400 651.600 960.600 653.400 ;
        RECT 964.950 652.950 967.050 653.400 ;
        RECT 985.950 652.950 988.050 655.050 ;
        RECT 967.950 651.600 970.050 652.050 ;
        RECT 937.950 650.400 960.600 651.600 ;
        RECT 962.400 650.400 970.050 651.600 ;
        RECT 937.950 650.100 940.050 650.400 ;
        RECT 962.400 648.600 963.600 650.400 ;
        RECT 967.950 649.950 970.050 650.400 ;
        RECT 976.950 649.950 979.050 652.050 ;
        RECT 929.400 647.400 933.600 648.600 ;
        RECT 953.400 648.000 963.600 648.600 ;
        RECT 871.950 645.450 909.600 645.600 ;
        RECT 859.950 644.400 909.600 645.450 ;
        RECT 913.950 645.600 916.050 645.900 ;
        RECT 928.950 645.600 931.050 645.900 ;
        RECT 913.950 644.400 931.050 645.600 ;
        RECT 859.950 644.250 874.050 644.400 ;
        RECT 859.950 643.800 862.050 644.250 ;
        RECT 871.950 643.800 874.050 644.250 ;
        RECT 913.950 643.800 916.050 644.400 ;
        RECT 928.950 643.800 931.050 644.400 ;
        RECT 640.950 641.400 648.600 642.600 ;
        RECT 730.950 642.600 733.050 643.050 ;
        RECT 745.950 642.600 748.050 643.050 ;
        RECT 730.950 641.400 748.050 642.600 ;
        RECT 640.950 640.950 643.050 641.400 ;
        RECT 730.950 640.950 733.050 641.400 ;
        RECT 745.950 640.950 748.050 641.400 ;
        RECT 862.950 642.600 865.050 643.050 ;
        RECT 868.950 642.600 871.050 643.050 ;
        RECT 862.950 641.400 871.050 642.600 ;
        RECT 862.950 640.950 865.050 641.400 ;
        RECT 868.950 640.950 871.050 641.400 ;
        RECT 883.950 642.600 886.050 643.050 ;
        RECT 892.950 642.600 895.050 643.050 ;
        RECT 883.950 641.400 895.050 642.600 ;
        RECT 932.400 642.600 933.600 647.400 ;
        RECT 952.950 647.400 963.600 648.000 ;
        RECT 940.950 645.600 943.050 646.050 ;
        RECT 946.950 645.600 949.050 646.050 ;
        RECT 940.950 644.400 949.050 645.600 ;
        RECT 940.950 643.950 943.050 644.400 ;
        RECT 946.950 643.950 949.050 644.400 ;
        RECT 952.950 643.950 955.050 647.400 ;
        RECT 977.400 645.600 978.600 649.950 ;
        RECT 965.400 644.400 978.600 645.600 ;
        RECT 937.950 642.600 940.050 643.050 ;
        RECT 932.400 641.400 940.050 642.600 ;
        RECT 883.950 640.950 886.050 641.400 ;
        RECT 892.950 640.950 895.050 641.400 ;
        RECT 937.950 640.950 940.050 641.400 ;
        RECT 958.950 642.600 961.050 643.050 ;
        RECT 965.400 642.600 966.600 644.400 ;
        RECT 979.950 643.800 982.050 645.900 ;
        RECT 986.400 645.600 987.600 652.950 ;
        RECT 988.950 651.600 991.050 652.200 ;
        RECT 1003.950 651.600 1006.050 652.200 ;
        RECT 988.950 650.400 1006.050 651.600 ;
        RECT 1006.950 651.600 1009.050 655.050 ;
        RECT 1006.950 651.000 1011.600 651.600 ;
        RECT 1007.400 650.400 1011.600 651.000 ;
        RECT 988.950 650.100 991.050 650.400 ;
        RECT 1003.950 650.100 1006.050 650.400 ;
        RECT 1006.950 645.600 1009.050 645.900 ;
        RECT 986.400 644.400 1009.050 645.600 ;
        RECT 1006.950 643.800 1009.050 644.400 ;
        RECT 958.950 641.400 966.600 642.600 ;
        RECT 980.400 643.050 981.600 643.800 ;
        RECT 1010.400 643.050 1011.600 650.400 ;
        RECT 1015.950 649.950 1018.050 652.050 ;
        RECT 1016.400 646.050 1017.600 649.950 ;
        RECT 1015.950 643.950 1018.050 646.050 ;
        RECT 980.400 641.400 985.050 643.050 ;
        RECT 958.950 640.950 961.050 641.400 ;
        RECT 981.000 640.950 985.050 641.400 ;
        RECT 1009.950 640.950 1012.050 643.050 ;
        RECT 190.950 639.600 193.050 640.050 ;
        RECT 304.950 639.600 307.050 640.050 ;
        RECT 322.950 639.600 325.050 640.050 ;
        RECT 355.950 639.600 358.050 640.050 ;
        RECT 373.950 639.600 376.050 640.050 ;
        RECT 391.950 639.600 394.050 640.050 ;
        RECT 190.950 638.400 394.050 639.600 ;
        RECT 190.950 637.950 193.050 638.400 ;
        RECT 304.950 637.950 307.050 638.400 ;
        RECT 322.950 637.950 325.050 638.400 ;
        RECT 355.950 637.950 358.050 638.400 ;
        RECT 373.950 637.950 376.050 638.400 ;
        RECT 391.950 637.950 394.050 638.400 ;
        RECT 430.950 639.600 433.050 640.050 ;
        RECT 460.950 639.600 463.050 640.050 ;
        RECT 430.950 638.400 463.050 639.600 ;
        RECT 430.950 637.950 433.050 638.400 ;
        RECT 460.950 637.950 463.050 638.400 ;
        RECT 679.950 639.600 682.050 640.050 ;
        RECT 715.950 639.600 718.050 640.050 ;
        RECT 742.950 639.600 745.050 640.050 ;
        RECT 679.950 638.400 745.050 639.600 ;
        RECT 679.950 637.950 682.050 638.400 ;
        RECT 715.950 637.950 718.050 638.400 ;
        RECT 742.950 637.950 745.050 638.400 ;
        RECT 907.950 639.600 910.050 639.900 ;
        RECT 925.950 639.600 928.050 640.050 ;
        RECT 907.950 638.400 928.050 639.600 ;
        RECT 907.950 637.800 910.050 638.400 ;
        RECT 925.950 637.950 928.050 638.400 ;
        RECT 949.950 639.600 952.050 640.050 ;
        RECT 967.950 639.600 970.050 640.050 ;
        RECT 949.950 638.400 970.050 639.600 ;
        RECT 949.950 637.950 952.050 638.400 ;
        RECT 967.950 637.950 970.050 638.400 ;
        RECT 994.950 639.600 997.050 640.050 ;
        RECT 1012.950 639.600 1015.050 640.050 ;
        RECT 994.950 638.400 1015.050 639.600 ;
        RECT 994.950 637.950 997.050 638.400 ;
        RECT 1012.950 637.950 1015.050 638.400 ;
        RECT 16.950 636.600 19.050 637.050 ;
        RECT 124.950 636.600 127.050 637.050 ;
        RECT 16.950 635.400 127.050 636.600 ;
        RECT 16.950 634.950 19.050 635.400 ;
        RECT 124.950 634.950 127.050 635.400 ;
        RECT 130.950 636.600 133.050 637.050 ;
        RECT 427.950 636.600 430.050 637.050 ;
        RECT 130.950 635.400 430.050 636.600 ;
        RECT 130.950 634.950 133.050 635.400 ;
        RECT 427.950 634.950 430.050 635.400 ;
        RECT 505.950 636.600 508.050 637.050 ;
        RECT 565.950 636.600 568.050 637.050 ;
        RECT 505.950 635.400 568.050 636.600 ;
        RECT 505.950 634.950 508.050 635.400 ;
        RECT 565.950 634.950 568.050 635.400 ;
        RECT 604.950 636.600 607.050 637.050 ;
        RECT 625.950 636.600 628.050 637.050 ;
        RECT 604.950 635.400 628.050 636.600 ;
        RECT 604.950 634.950 607.050 635.400 ;
        RECT 625.950 634.950 628.050 635.400 ;
        RECT 793.950 636.600 796.050 636.900 ;
        RECT 817.950 636.600 820.050 637.050 ;
        RECT 793.950 635.400 820.050 636.600 ;
        RECT 793.950 634.800 796.050 635.400 ;
        RECT 817.950 634.950 820.050 635.400 ;
        RECT 844.950 636.600 847.050 637.050 ;
        RECT 943.950 636.600 946.050 637.050 ;
        RECT 844.950 635.400 946.050 636.600 ;
        RECT 844.950 634.950 847.050 635.400 ;
        RECT 943.950 634.950 946.050 635.400 ;
        RECT 1000.950 636.600 1003.050 637.050 ;
        RECT 1006.950 636.600 1009.050 637.050 ;
        RECT 1000.950 635.400 1009.050 636.600 ;
        RECT 1000.950 634.950 1003.050 635.400 ;
        RECT 1006.950 634.950 1009.050 635.400 ;
        RECT 43.950 633.600 46.050 634.050 ;
        RECT 55.950 633.600 58.050 634.050 ;
        RECT 43.950 632.400 58.050 633.600 ;
        RECT 43.950 631.950 46.050 632.400 ;
        RECT 55.950 631.950 58.050 632.400 ;
        RECT 70.950 633.600 73.050 634.050 ;
        RECT 88.950 633.600 91.050 634.050 ;
        RECT 178.950 633.600 181.050 634.050 ;
        RECT 70.950 632.400 181.050 633.600 ;
        RECT 70.950 631.950 73.050 632.400 ;
        RECT 88.950 631.950 91.050 632.400 ;
        RECT 178.950 631.950 181.050 632.400 ;
        RECT 211.950 633.600 214.050 634.050 ;
        RECT 274.950 633.600 277.050 634.050 ;
        RECT 211.950 632.400 277.050 633.600 ;
        RECT 211.950 631.950 214.050 632.400 ;
        RECT 274.950 631.950 277.050 632.400 ;
        RECT 451.950 633.600 454.050 634.050 ;
        RECT 466.950 633.600 469.050 634.050 ;
        RECT 451.950 632.400 469.050 633.600 ;
        RECT 451.950 631.950 454.050 632.400 ;
        RECT 466.950 631.950 469.050 632.400 ;
        RECT 535.950 633.600 538.050 634.050 ;
        RECT 547.950 633.600 550.050 634.050 ;
        RECT 586.950 633.600 589.050 634.050 ;
        RECT 610.950 633.600 613.050 634.050 ;
        RECT 535.950 632.400 613.050 633.600 ;
        RECT 535.950 631.950 538.050 632.400 ;
        RECT 547.950 631.950 550.050 632.400 ;
        RECT 586.950 631.950 589.050 632.400 ;
        RECT 610.950 631.950 613.050 632.400 ;
        RECT 661.950 633.600 664.050 634.050 ;
        RECT 679.950 633.600 682.050 634.050 ;
        RECT 661.950 632.400 682.050 633.600 ;
        RECT 661.950 631.950 664.050 632.400 ;
        RECT 679.950 631.950 682.050 632.400 ;
        RECT 688.950 633.600 691.050 634.050 ;
        RECT 733.950 633.600 736.050 634.050 ;
        RECT 688.950 632.400 736.050 633.600 ;
        RECT 688.950 631.950 691.050 632.400 ;
        RECT 733.950 631.950 736.050 632.400 ;
        RECT 877.950 633.600 880.050 634.050 ;
        RECT 889.950 633.600 892.050 634.050 ;
        RECT 877.950 632.400 892.050 633.600 ;
        RECT 877.950 631.950 880.050 632.400 ;
        RECT 889.950 631.950 892.050 632.400 ;
        RECT 910.950 633.600 913.050 634.050 ;
        RECT 949.950 633.600 952.050 634.050 ;
        RECT 910.950 632.400 952.050 633.600 ;
        RECT 910.950 631.950 913.050 632.400 ;
        RECT 949.950 631.950 952.050 632.400 ;
        RECT 961.950 633.600 964.050 634.050 ;
        RECT 970.950 633.600 973.050 634.050 ;
        RECT 961.950 632.400 973.050 633.600 ;
        RECT 961.950 631.950 964.050 632.400 ;
        RECT 970.950 631.950 973.050 632.400 ;
        RECT 349.950 630.600 352.050 631.050 ;
        RECT 409.950 630.600 412.050 631.050 ;
        RECT 454.950 630.600 457.050 631.050 ;
        RECT 349.950 629.400 457.050 630.600 ;
        RECT 349.950 628.950 352.050 629.400 ;
        RECT 409.950 628.950 412.050 629.400 ;
        RECT 454.950 628.950 457.050 629.400 ;
        RECT 469.950 630.600 472.050 631.050 ;
        RECT 526.950 630.600 529.050 631.050 ;
        RECT 469.950 629.400 529.050 630.600 ;
        RECT 469.950 628.950 472.050 629.400 ;
        RECT 526.950 628.950 529.050 629.400 ;
        RECT 553.950 630.600 556.050 631.050 ;
        RECT 559.950 630.600 562.050 631.050 ;
        RECT 553.950 629.400 562.050 630.600 ;
        RECT 553.950 628.950 556.050 629.400 ;
        RECT 559.950 628.950 562.050 629.400 ;
        RECT 580.950 630.600 583.050 631.050 ;
        RECT 625.950 630.600 628.050 631.050 ;
        RECT 580.950 629.400 628.050 630.600 ;
        RECT 580.950 628.950 583.050 629.400 ;
        RECT 625.950 628.950 628.050 629.400 ;
        RECT 898.950 630.600 901.050 631.050 ;
        RECT 958.950 630.600 961.050 631.050 ;
        RECT 964.950 630.600 967.050 631.050 ;
        RECT 898.950 629.400 967.050 630.600 ;
        RECT 898.950 628.950 901.050 629.400 ;
        RECT 958.950 628.950 961.050 629.400 ;
        RECT 964.950 628.950 967.050 629.400 ;
        RECT 973.950 630.600 976.050 631.050 ;
        RECT 985.950 630.600 988.050 631.050 ;
        RECT 1009.950 630.600 1012.050 631.050 ;
        RECT 973.950 629.400 1012.050 630.600 ;
        RECT 973.950 628.950 976.050 629.400 ;
        RECT 985.950 628.950 988.050 629.400 ;
        RECT 1009.950 628.950 1012.050 629.400 ;
        RECT 262.950 627.600 265.050 628.050 ;
        RECT 358.950 627.600 361.050 628.050 ;
        RECT 262.950 626.400 361.050 627.600 ;
        RECT 262.950 625.950 265.050 626.400 ;
        RECT 358.950 625.950 361.050 626.400 ;
        RECT 460.950 627.600 463.050 628.050 ;
        RECT 472.950 627.600 475.050 628.050 ;
        RECT 460.950 626.400 475.050 627.600 ;
        RECT 460.950 625.950 463.050 626.400 ;
        RECT 472.950 625.950 475.050 626.400 ;
        RECT 478.950 627.600 481.050 628.050 ;
        RECT 484.950 627.600 487.050 628.050 ;
        RECT 554.400 627.600 555.600 628.950 ;
        RECT 478.950 626.400 555.600 627.600 ;
        RECT 733.950 627.600 736.050 628.050 ;
        RECT 760.950 627.600 763.050 628.050 ;
        RECT 733.950 626.400 763.050 627.600 ;
        RECT 478.950 625.950 481.050 626.400 ;
        RECT 484.950 625.950 487.050 626.400 ;
        RECT 733.950 625.950 736.050 626.400 ;
        RECT 760.950 625.950 763.050 626.400 ;
        RECT 931.950 627.600 934.050 628.050 ;
        RECT 940.950 627.600 943.050 628.050 ;
        RECT 931.950 626.400 943.050 627.600 ;
        RECT 931.950 625.950 934.050 626.400 ;
        RECT 940.950 625.950 943.050 626.400 ;
        RECT 985.950 627.600 988.050 627.900 ;
        RECT 991.950 627.600 994.050 628.050 ;
        RECT 985.950 626.400 994.050 627.600 ;
        RECT 985.950 625.800 988.050 626.400 ;
        RECT 991.950 625.950 994.050 626.400 ;
        RECT 859.950 624.600 862.050 625.050 ;
        RECT 895.950 624.600 898.050 625.050 ;
        RECT 859.950 623.400 898.050 624.600 ;
        RECT 859.950 622.950 862.050 623.400 ;
        RECT 895.950 622.950 898.050 623.400 ;
        RECT 967.950 624.600 970.050 625.050 ;
        RECT 997.950 624.600 1000.050 625.050 ;
        RECT 967.950 623.400 1000.050 624.600 ;
        RECT 967.950 622.950 970.050 623.400 ;
        RECT 997.950 622.950 1000.050 623.400 ;
        RECT 64.950 621.600 67.050 622.050 ;
        RECT 196.950 621.600 199.050 622.050 ;
        RECT 64.950 620.400 199.050 621.600 ;
        RECT 64.950 619.950 67.050 620.400 ;
        RECT 196.950 619.950 199.050 620.400 ;
        RECT 436.950 621.600 439.050 622.050 ;
        RECT 478.950 621.600 481.050 622.050 ;
        RECT 436.950 620.400 481.050 621.600 ;
        RECT 436.950 619.950 439.050 620.400 ;
        RECT 478.950 619.950 481.050 620.400 ;
        RECT 505.950 621.600 508.050 622.050 ;
        RECT 556.950 621.600 559.050 622.050 ;
        RECT 505.950 620.400 559.050 621.600 ;
        RECT 505.950 619.950 508.050 620.400 ;
        RECT 556.950 619.950 559.050 620.400 ;
        RECT 562.950 621.600 565.050 622.050 ;
        RECT 826.950 621.600 829.050 622.050 ;
        RECT 844.950 621.600 847.050 622.050 ;
        RECT 562.950 620.400 847.050 621.600 ;
        RECT 562.950 619.950 565.050 620.400 ;
        RECT 826.950 619.950 829.050 620.400 ;
        RECT 844.950 619.950 847.050 620.400 ;
        RECT 970.950 621.600 973.050 622.050 ;
        RECT 979.950 621.600 982.050 622.050 ;
        RECT 970.950 620.400 982.050 621.600 ;
        RECT 970.950 619.950 973.050 620.400 ;
        RECT 979.950 619.950 982.050 620.400 ;
        RECT 40.950 618.600 43.050 619.050 ;
        RECT 52.950 618.600 55.050 619.050 ;
        RECT 40.950 617.400 55.050 618.600 ;
        RECT 40.950 616.950 43.050 617.400 ;
        RECT 52.950 616.950 55.050 617.400 ;
        RECT 202.950 618.600 205.050 619.050 ;
        RECT 259.950 618.600 262.050 619.050 ;
        RECT 202.950 617.400 262.050 618.600 ;
        RECT 479.400 618.600 480.600 619.950 ;
        RECT 520.950 618.600 523.050 619.050 ;
        RECT 479.400 617.400 523.050 618.600 ;
        RECT 202.950 616.950 205.050 617.400 ;
        RECT 259.950 616.950 262.050 617.400 ;
        RECT 520.950 616.950 523.050 617.400 ;
        RECT 583.950 618.600 586.050 619.050 ;
        RECT 619.950 618.600 622.050 619.050 ;
        RECT 703.950 618.600 706.050 619.050 ;
        RECT 712.950 618.600 715.050 619.050 ;
        RECT 583.950 617.400 622.050 618.600 ;
        RECT 583.950 616.950 586.050 617.400 ;
        RECT 619.950 616.950 622.050 617.400 ;
        RECT 659.400 617.400 715.050 618.600 ;
        RECT 82.950 615.600 85.050 616.050 ;
        RECT 130.950 615.600 133.050 616.050 ;
        RECT 82.950 614.400 133.050 615.600 ;
        RECT 82.950 613.950 85.050 614.400 ;
        RECT 130.950 613.950 133.050 614.400 ;
        RECT 415.950 615.600 418.050 616.050 ;
        RECT 436.950 615.600 439.050 616.050 ;
        RECT 415.950 614.400 439.050 615.600 ;
        RECT 415.950 613.950 418.050 614.400 ;
        RECT 436.950 613.950 439.050 614.400 ;
        RECT 559.950 615.600 562.050 616.050 ;
        RECT 598.950 615.600 601.050 616.050 ;
        RECT 559.950 614.400 601.050 615.600 ;
        RECT 559.950 613.950 562.050 614.400 ;
        RECT 598.950 613.950 601.050 614.400 ;
        RECT 610.950 615.600 613.050 616.050 ;
        RECT 659.400 615.600 660.600 617.400 ;
        RECT 703.950 616.950 706.050 617.400 ;
        RECT 712.950 616.950 715.050 617.400 ;
        RECT 871.950 618.600 874.050 619.050 ;
        RECT 913.950 618.600 916.050 619.050 ;
        RECT 871.950 617.400 916.050 618.600 ;
        RECT 871.950 616.950 874.050 617.400 ;
        RECT 913.950 616.950 916.050 617.400 ;
        RECT 610.950 614.400 660.600 615.600 ;
        RECT 673.950 615.600 676.050 616.050 ;
        RECT 754.950 615.600 757.050 616.050 ;
        RECT 760.950 615.600 763.050 616.050 ;
        RECT 787.950 615.600 790.050 616.050 ;
        RECT 820.950 615.600 823.050 616.050 ;
        RECT 841.950 615.600 844.050 616.050 ;
        RECT 673.950 614.400 844.050 615.600 ;
        RECT 610.950 613.950 613.050 614.400 ;
        RECT 673.950 613.950 676.050 614.400 ;
        RECT 754.950 613.950 757.050 614.400 ;
        RECT 760.950 613.950 763.050 614.400 ;
        RECT 787.950 613.950 790.050 614.400 ;
        RECT 820.950 613.950 823.050 614.400 ;
        RECT 841.950 613.950 844.050 614.400 ;
        RECT 922.950 615.600 925.050 616.050 ;
        RECT 928.950 615.600 931.050 616.050 ;
        RECT 922.950 614.400 931.050 615.600 ;
        RECT 922.950 613.950 925.050 614.400 ;
        RECT 928.950 613.950 931.050 614.400 ;
        RECT 937.950 615.600 940.050 616.050 ;
        RECT 979.950 615.600 982.050 616.050 ;
        RECT 937.950 614.400 982.050 615.600 ;
        RECT 937.950 613.950 940.050 614.400 ;
        RECT 979.950 613.950 982.050 614.400 ;
        RECT 46.950 612.600 49.050 613.050 ;
        RECT 58.950 612.600 61.050 613.050 ;
        RECT 46.950 611.400 61.050 612.600 ;
        RECT 46.950 610.950 49.050 611.400 ;
        RECT 58.950 610.950 61.050 611.400 ;
        RECT 217.950 612.600 220.050 613.050 ;
        RECT 289.950 612.600 292.050 613.050 ;
        RECT 217.950 611.400 292.050 612.600 ;
        RECT 217.950 610.950 220.050 611.400 ;
        RECT 289.950 610.950 292.050 611.400 ;
        RECT 526.950 612.600 529.050 613.050 ;
        RECT 547.950 612.600 550.050 613.050 ;
        RECT 526.950 611.400 550.050 612.600 ;
        RECT 526.950 610.950 529.050 611.400 ;
        RECT 547.950 610.950 550.050 611.400 ;
        RECT 556.950 612.600 559.050 613.050 ;
        RECT 574.950 612.600 577.050 612.900 ;
        RECT 556.950 611.400 577.050 612.600 ;
        RECT 556.950 610.950 559.050 611.400 ;
        RECT 574.950 610.800 577.050 611.400 ;
        RECT 586.950 612.600 589.050 613.050 ;
        RECT 592.950 612.600 595.050 613.050 ;
        RECT 586.950 611.400 595.050 612.600 ;
        RECT 586.950 610.950 589.050 611.400 ;
        RECT 592.950 610.950 595.050 611.400 ;
        RECT 661.950 612.600 664.050 613.050 ;
        RECT 685.950 612.600 688.050 613.050 ;
        RECT 661.950 611.400 688.050 612.600 ;
        RECT 661.950 610.950 664.050 611.400 ;
        RECT 685.950 610.950 688.050 611.400 ;
        RECT 868.950 612.600 871.050 613.050 ;
        RECT 880.950 612.600 883.050 613.050 ;
        RECT 925.950 612.600 928.050 613.050 ;
        RECT 868.950 611.400 928.050 612.600 ;
        RECT 868.950 610.950 871.050 611.400 ;
        RECT 880.950 610.950 883.050 611.400 ;
        RECT 925.950 610.950 928.050 611.400 ;
        RECT 991.950 612.600 994.050 613.050 ;
        RECT 1003.950 612.600 1006.050 613.050 ;
        RECT 991.950 611.400 1006.050 612.600 ;
        RECT 991.950 610.950 994.050 611.400 ;
        RECT 1003.950 610.950 1006.050 611.400 ;
        RECT 4.950 607.950 7.050 610.050 ;
        RECT 70.950 609.600 73.050 610.050 ;
        RECT 88.950 609.600 91.050 610.050 ;
        RECT 343.950 609.600 346.050 610.050 ;
        RECT 400.950 609.600 403.050 610.050 ;
        RECT 38.400 608.400 91.050 609.600 ;
        RECT 5.400 600.900 6.600 607.950 ;
        RECT 38.400 607.200 39.600 608.400 ;
        RECT 70.950 607.950 73.050 608.400 ;
        RECT 88.950 607.950 91.050 608.400 ;
        RECT 92.400 608.400 141.600 609.600 ;
        RECT 16.950 606.750 19.050 607.200 ;
        RECT 22.950 606.750 25.050 607.200 ;
        RECT 16.950 605.550 25.050 606.750 ;
        RECT 16.950 605.100 19.050 605.550 ;
        RECT 22.950 605.100 25.050 605.550 ;
        RECT 31.950 606.750 34.050 607.200 ;
        RECT 37.950 606.750 40.050 607.200 ;
        RECT 31.950 605.550 40.050 606.750 ;
        RECT 31.950 605.100 34.050 605.550 ;
        RECT 37.950 605.100 40.050 605.550 ;
        RECT 52.950 606.600 55.050 607.200 ;
        RECT 76.950 606.600 79.050 607.200 ;
        RECT 92.400 606.600 93.600 608.400 ;
        RECT 52.950 605.400 93.600 606.600 ;
        RECT 52.950 605.100 55.050 605.400 ;
        RECT 76.950 605.100 79.050 605.400 ;
        RECT 97.950 605.100 100.050 607.200 ;
        RECT 124.950 606.600 127.050 607.050 ;
        RECT 136.950 606.600 139.050 607.200 ;
        RECT 124.950 605.400 139.050 606.600 ;
        RECT 140.400 606.600 141.600 608.400 ;
        RECT 343.950 608.400 403.050 609.600 ;
        RECT 343.950 607.950 346.050 608.400 ;
        RECT 400.950 607.950 403.050 608.400 ;
        RECT 430.950 609.600 433.050 610.050 ;
        RECT 436.950 609.600 439.050 610.050 ;
        RECT 430.950 608.400 439.050 609.600 ;
        RECT 430.950 607.950 433.050 608.400 ;
        RECT 436.950 607.950 439.050 608.400 ;
        RECT 454.950 609.600 457.050 610.050 ;
        RECT 496.950 609.600 499.050 610.050 ;
        RECT 454.950 608.400 499.050 609.600 ;
        RECT 454.950 607.950 457.050 608.400 ;
        RECT 496.950 607.950 499.050 608.400 ;
        RECT 508.950 609.600 511.050 610.050 ;
        RECT 523.950 609.600 526.050 610.050 ;
        RECT 508.950 608.400 526.050 609.600 ;
        RECT 508.950 607.950 511.050 608.400 ;
        RECT 523.950 607.950 526.050 608.400 ;
        RECT 580.950 609.600 583.050 610.050 ;
        RECT 589.950 609.600 592.050 610.050 ;
        RECT 580.950 608.400 592.050 609.600 ;
        RECT 580.950 607.950 583.050 608.400 ;
        RECT 589.950 607.950 592.050 608.400 ;
        RECT 613.950 609.600 616.050 610.050 ;
        RECT 631.950 609.600 634.050 610.050 ;
        RECT 613.950 608.400 634.050 609.600 ;
        RECT 613.950 607.950 616.050 608.400 ;
        RECT 631.950 607.950 634.050 608.400 ;
        RECT 889.950 609.600 892.050 610.200 ;
        RECT 895.950 609.600 898.050 610.050 ;
        RECT 889.950 608.400 898.050 609.600 ;
        RECT 889.950 608.100 892.050 608.400 ;
        RECT 895.950 607.950 898.050 608.400 ;
        RECT 142.950 606.750 145.050 607.200 ;
        RECT 148.950 606.750 151.050 607.200 ;
        RECT 142.950 606.600 151.050 606.750 ;
        RECT 140.400 605.550 151.050 606.600 ;
        RECT 140.400 605.400 145.050 605.550 ;
        RECT 4.950 598.800 7.050 600.900 ;
        RECT 13.950 600.600 16.050 601.050 ;
        RECT 19.950 600.600 22.050 601.050 ;
        RECT 13.950 599.400 22.050 600.600 ;
        RECT 13.950 598.950 16.050 599.400 ;
        RECT 19.950 598.950 22.050 599.400 ;
        RECT 43.950 600.600 46.050 601.050 ;
        RECT 49.950 600.600 52.050 600.900 ;
        RECT 43.950 599.400 52.050 600.600 ;
        RECT 43.950 598.950 46.050 599.400 ;
        RECT 49.950 598.800 52.050 599.400 ;
        RECT 79.950 600.600 82.050 600.900 ;
        RECT 98.400 600.600 99.600 605.100 ;
        RECT 124.950 604.950 127.050 605.400 ;
        RECT 136.950 605.100 139.050 605.400 ;
        RECT 142.950 605.100 145.050 605.400 ;
        RECT 148.950 605.100 151.050 605.550 ;
        RECT 154.950 606.600 157.050 607.050 ;
        RECT 163.950 606.600 166.050 607.200 ;
        RECT 190.950 606.600 193.050 607.200 ;
        RECT 154.950 605.400 193.050 606.600 ;
        RECT 154.950 604.950 157.050 605.400 ;
        RECT 163.950 605.100 166.050 605.400 ;
        RECT 190.950 605.100 193.050 605.400 ;
        RECT 238.950 606.600 241.050 607.200 ;
        RECT 244.800 606.600 246.900 607.050 ;
        RECT 238.950 605.400 246.900 606.600 ;
        RECT 238.950 605.100 241.050 605.400 ;
        RECT 244.800 604.950 246.900 605.400 ;
        RECT 247.950 606.750 250.050 607.200 ;
        RECT 253.950 606.750 256.050 607.200 ;
        RECT 247.950 605.550 256.050 606.750 ;
        RECT 247.950 605.100 250.050 605.550 ;
        RECT 253.950 605.100 256.050 605.550 ;
        RECT 265.950 606.600 268.050 607.200 ;
        RECT 280.950 606.600 283.050 607.200 ;
        RECT 265.950 605.400 283.050 606.600 ;
        RECT 265.950 605.100 268.050 605.400 ;
        RECT 280.950 605.100 283.050 605.400 ;
        RECT 307.950 606.600 310.050 607.050 ;
        RECT 313.950 606.600 316.050 607.200 ;
        RECT 307.950 605.400 316.050 606.600 ;
        RECT 307.950 604.950 310.050 605.400 ;
        RECT 313.950 605.100 316.050 605.400 ;
        RECT 367.950 606.750 370.050 607.200 ;
        RECT 382.950 606.750 385.050 607.200 ;
        RECT 367.950 605.550 385.050 606.750 ;
        RECT 367.950 605.100 370.050 605.550 ;
        RECT 382.950 605.100 385.050 605.550 ;
        RECT 412.950 606.600 415.050 607.050 ;
        RECT 448.950 606.600 451.050 607.200 ;
        RECT 412.950 605.400 451.050 606.600 ;
        RECT 412.950 604.950 415.050 605.400 ;
        RECT 448.950 605.100 451.050 605.400 ;
        RECT 553.950 604.950 556.050 607.050 ;
        RECT 568.950 606.600 571.050 607.200 ;
        RECT 595.950 606.600 598.050 607.200 ;
        RECT 640.950 606.600 643.050 607.200 ;
        RECT 568.950 605.400 643.050 606.600 ;
        RECT 568.950 605.100 571.050 605.400 ;
        RECT 595.950 605.100 598.050 605.400 ;
        RECT 554.400 601.050 555.600 604.950 ;
        RECT 79.950 599.400 99.600 600.600 ;
        RECT 115.950 600.450 118.050 600.900 ;
        RECT 124.950 600.450 127.050 600.900 ;
        RECT 79.950 598.800 82.050 599.400 ;
        RECT 115.950 599.250 127.050 600.450 ;
        RECT 115.950 598.800 118.050 599.250 ;
        RECT 124.950 598.800 127.050 599.250 ;
        RECT 130.950 600.600 133.050 601.050 ;
        RECT 139.950 600.600 142.050 600.900 ;
        RECT 130.950 599.400 142.050 600.600 ;
        RECT 130.950 598.950 133.050 599.400 ;
        RECT 139.950 598.800 142.050 599.400 ;
        RECT 217.950 600.600 220.050 600.900 ;
        RECT 235.950 600.600 238.050 600.900 ;
        RECT 217.950 599.400 238.050 600.600 ;
        RECT 217.950 598.800 220.050 599.400 ;
        RECT 235.950 598.800 238.050 599.400 ;
        RECT 244.950 600.450 247.050 600.900 ;
        RECT 256.950 600.450 259.050 600.900 ;
        RECT 244.950 599.250 259.050 600.450 ;
        RECT 244.950 598.800 247.050 599.250 ;
        RECT 256.950 598.800 259.050 599.250 ;
        RECT 262.950 600.450 265.050 600.900 ;
        RECT 274.950 600.450 277.050 600.900 ;
        RECT 262.950 599.250 277.050 600.450 ;
        RECT 262.950 598.800 265.050 599.250 ;
        RECT 274.950 598.800 277.050 599.250 ;
        RECT 340.950 600.600 343.050 600.900 ;
        RECT 349.950 600.600 352.050 600.900 ;
        RECT 340.950 599.400 352.050 600.600 ;
        RECT 340.950 598.800 343.050 599.400 ;
        RECT 349.950 598.800 352.050 599.400 ;
        RECT 382.950 600.600 385.050 601.050 ;
        RECT 403.950 600.600 406.050 600.900 ;
        RECT 382.950 599.400 406.050 600.600 ;
        RECT 382.950 598.950 385.050 599.400 ;
        RECT 403.950 598.800 406.050 599.400 ;
        RECT 436.950 600.600 439.050 601.050 ;
        RECT 451.950 600.600 454.050 600.900 ;
        RECT 436.950 599.400 454.050 600.600 ;
        RECT 436.950 598.950 439.050 599.400 ;
        RECT 451.950 598.800 454.050 599.400 ;
        RECT 502.950 600.600 505.050 600.900 ;
        RECT 520.950 600.600 523.050 600.900 ;
        RECT 502.950 599.400 523.050 600.600 ;
        RECT 502.950 598.800 505.050 599.400 ;
        RECT 520.950 598.800 523.050 599.400 ;
        RECT 529.950 600.450 532.050 600.900 ;
        RECT 541.950 600.450 544.050 600.900 ;
        RECT 529.950 599.250 544.050 600.450 ;
        RECT 529.950 598.800 532.050 599.250 ;
        RECT 541.950 598.800 544.050 599.250 ;
        RECT 553.950 598.950 556.050 601.050 ;
        RECT 583.950 600.600 586.050 601.050 ;
        RECT 611.400 600.900 612.600 605.400 ;
        RECT 640.950 605.100 643.050 605.400 ;
        RECT 649.950 606.750 652.050 607.200 ;
        RECT 655.950 606.750 658.050 607.200 ;
        RECT 649.950 606.600 658.050 606.750 ;
        RECT 679.950 606.600 682.050 607.200 ;
        RECT 649.950 605.550 682.050 606.600 ;
        RECT 649.950 605.100 652.050 605.550 ;
        RECT 655.950 605.400 682.050 605.550 ;
        RECT 655.950 605.100 658.050 605.400 ;
        RECT 679.950 605.100 682.050 605.400 ;
        RECT 685.950 606.750 688.050 607.200 ;
        RECT 694.950 606.750 697.050 607.200 ;
        RECT 685.950 605.550 697.050 606.750 ;
        RECT 685.950 605.100 688.050 605.550 ;
        RECT 694.950 605.100 697.050 605.550 ;
        RECT 721.950 606.750 724.050 607.200 ;
        RECT 733.950 606.750 736.050 607.200 ;
        RECT 721.950 605.550 736.050 606.750 ;
        RECT 721.950 605.100 724.050 605.550 ;
        RECT 733.950 605.100 736.050 605.550 ;
        RECT 742.950 606.750 745.050 607.200 ;
        RECT 775.950 606.750 778.050 607.200 ;
        RECT 742.950 605.550 778.050 606.750 ;
        RECT 742.950 605.100 745.050 605.550 ;
        RECT 775.950 605.100 778.050 605.550 ;
        RECT 802.950 606.600 805.050 607.200 ;
        RECT 811.950 606.600 814.050 607.050 ;
        RECT 850.950 606.600 853.050 607.200 ;
        RECT 802.950 605.400 853.050 606.600 ;
        RECT 802.950 605.100 805.050 605.400 ;
        RECT 811.950 604.950 814.050 605.400 ;
        RECT 850.950 605.100 853.050 605.400 ;
        RECT 865.950 604.950 868.050 607.050 ;
        RECT 874.950 606.600 877.050 607.050 ;
        RECT 883.950 606.600 886.050 607.050 ;
        RECT 889.950 606.600 892.050 607.050 ;
        RECT 874.950 605.400 879.600 606.600 ;
        RECT 874.950 604.950 877.050 605.400 ;
        RECT 662.400 602.400 684.600 603.600 ;
        RECT 592.950 600.600 595.050 600.900 ;
        RECT 583.950 599.400 595.050 600.600 ;
        RECT 583.950 598.950 586.050 599.400 ;
        RECT 592.950 598.800 595.050 599.400 ;
        RECT 610.950 598.800 613.050 600.900 ;
        RECT 637.950 600.600 640.050 600.900 ;
        RECT 632.400 600.000 640.050 600.600 ;
        RECT 631.950 599.400 640.050 600.000 ;
        RECT 88.950 597.600 91.050 598.050 ;
        RECT 106.950 597.600 109.050 598.050 ;
        RECT 88.950 596.400 109.050 597.600 ;
        RECT 88.950 595.950 91.050 596.400 ;
        RECT 106.950 595.950 109.050 596.400 ;
        RECT 556.950 597.600 559.050 598.050 ;
        RECT 571.950 597.600 574.050 598.050 ;
        RECT 556.950 596.400 574.050 597.600 ;
        RECT 556.950 595.950 559.050 596.400 ;
        RECT 571.950 595.950 574.050 596.400 ;
        RECT 631.950 595.950 634.050 599.400 ;
        RECT 637.950 598.800 640.050 599.400 ;
        RECT 658.950 600.600 661.050 600.900 ;
        RECT 662.400 600.600 663.600 602.400 ;
        RECT 658.950 599.400 663.600 600.600 ;
        RECT 664.950 600.600 667.050 600.900 ;
        RECT 673.950 600.600 676.050 601.050 ;
        RECT 683.400 600.900 684.600 602.400 ;
        RECT 664.950 599.400 676.050 600.600 ;
        RECT 658.950 598.800 661.050 599.400 ;
        RECT 664.950 598.800 667.050 599.400 ;
        RECT 673.950 598.950 676.050 599.400 ;
        RECT 682.950 598.800 685.050 600.900 ;
        RECT 757.950 600.600 760.050 600.900 ;
        RECT 769.950 600.600 772.050 601.050 ;
        RECT 757.950 599.400 772.050 600.600 ;
        RECT 757.950 598.800 760.050 599.400 ;
        RECT 769.950 598.950 772.050 599.400 ;
        RECT 811.950 600.450 814.050 600.900 ;
        RECT 823.950 600.450 826.050 600.900 ;
        RECT 811.950 599.250 826.050 600.450 ;
        RECT 811.950 598.800 814.050 599.250 ;
        RECT 823.950 598.800 826.050 599.250 ;
        RECT 838.950 600.450 841.050 600.900 ;
        RECT 847.950 600.450 850.050 600.900 ;
        RECT 838.950 599.250 850.050 600.450 ;
        RECT 838.950 598.800 841.050 599.250 ;
        RECT 847.950 598.800 850.050 599.250 ;
        RECT 685.950 597.600 688.050 598.050 ;
        RECT 694.950 597.600 697.050 598.050 ;
        RECT 685.950 596.400 697.050 597.600 ;
        RECT 685.950 595.950 688.050 596.400 ;
        RECT 694.950 595.950 697.050 596.400 ;
        RECT 730.950 597.600 733.050 598.050 ;
        RECT 739.950 597.600 742.050 598.050 ;
        RECT 730.950 596.400 742.050 597.600 ;
        RECT 730.950 595.950 733.050 596.400 ;
        RECT 739.950 595.950 742.050 596.400 ;
        RECT 808.950 597.600 811.050 598.050 ;
        RECT 829.950 597.600 832.050 598.050 ;
        RECT 808.950 596.400 832.050 597.600 ;
        RECT 808.950 595.950 811.050 596.400 ;
        RECT 829.950 595.950 832.050 596.400 ;
        RECT 850.950 597.600 853.050 598.050 ;
        RECT 866.400 597.600 867.600 604.950 ;
        RECT 878.400 603.600 879.600 605.400 ;
        RECT 883.950 605.400 892.050 606.600 ;
        RECT 883.950 604.950 886.050 605.400 ;
        RECT 889.950 604.950 892.050 605.400 ;
        RECT 940.950 605.100 943.050 607.200 ;
        RECT 904.950 603.600 907.050 604.050 ;
        RECT 878.400 602.400 907.050 603.600 ;
        RECT 904.950 601.950 907.050 602.400 ;
        RECT 941.400 601.050 942.600 605.100 ;
        RECT 946.950 604.950 949.050 607.050 ;
        RECT 976.950 605.100 979.050 607.200 ;
        RECT 991.950 605.100 994.050 607.200 ;
        RECT 871.950 600.600 874.050 600.900 ;
        RECT 883.950 600.600 886.050 601.050 ;
        RECT 871.950 599.400 886.050 600.600 ;
        RECT 871.950 598.800 874.050 599.400 ;
        RECT 883.950 598.950 886.050 599.400 ;
        RECT 937.950 599.400 942.600 601.050 ;
        RECT 947.400 603.600 948.600 604.950 ;
        RECT 977.400 603.600 978.600 605.100 ;
        RECT 947.400 602.400 978.600 603.600 ;
        RECT 947.400 600.600 948.600 602.400 ;
        RECT 952.950 600.600 955.050 601.050 ;
        RECT 947.400 599.400 955.050 600.600 ;
        RECT 937.950 598.950 942.000 599.400 ;
        RECT 952.950 598.950 955.050 599.400 ;
        RECT 958.950 600.450 961.050 600.900 ;
        RECT 967.950 600.450 970.050 600.900 ;
        RECT 958.950 599.250 970.050 600.450 ;
        RECT 958.950 598.800 961.050 599.250 ;
        RECT 967.950 598.800 970.050 599.250 ;
        RECT 850.950 596.400 867.600 597.600 ;
        RECT 886.950 597.600 889.050 598.050 ;
        RECT 892.950 597.600 895.050 598.050 ;
        RECT 886.950 596.400 895.050 597.600 ;
        RECT 850.950 595.950 853.050 596.400 ;
        RECT 886.950 595.950 889.050 596.400 ;
        RECT 892.950 595.950 895.050 596.400 ;
        RECT 898.950 597.600 901.050 598.050 ;
        RECT 904.950 597.600 907.050 598.050 ;
        RECT 919.950 597.600 922.050 598.050 ;
        RECT 898.950 596.400 922.050 597.600 ;
        RECT 898.950 595.950 901.050 596.400 ;
        RECT 904.950 595.950 907.050 596.400 ;
        RECT 919.950 595.950 922.050 596.400 ;
        RECT 970.950 597.600 973.050 598.050 ;
        RECT 982.950 597.600 985.050 598.050 ;
        RECT 970.950 596.400 985.050 597.600 ;
        RECT 992.400 597.600 993.600 605.100 ;
        RECT 1003.950 604.950 1006.050 607.050 ;
        RECT 1004.400 601.050 1005.600 604.950 ;
        RECT 1003.950 598.950 1006.050 601.050 ;
        RECT 997.950 597.600 1000.050 598.050 ;
        RECT 992.400 596.400 1000.050 597.600 ;
        RECT 970.950 595.950 973.050 596.400 ;
        RECT 982.950 595.950 985.050 596.400 ;
        RECT 997.950 595.950 1000.050 596.400 ;
        RECT 16.950 594.600 19.050 595.050 ;
        RECT 55.950 594.600 58.050 595.050 ;
        RECT 16.950 593.400 58.050 594.600 ;
        RECT 16.950 592.950 19.050 593.400 ;
        RECT 55.950 592.950 58.050 593.400 ;
        RECT 142.950 594.600 145.050 595.050 ;
        RECT 148.950 594.600 151.050 595.050 ;
        RECT 142.950 593.400 151.050 594.600 ;
        RECT 142.950 592.950 145.050 593.400 ;
        RECT 148.950 592.950 151.050 593.400 ;
        RECT 205.950 594.600 208.050 595.050 ;
        RECT 247.950 594.600 250.050 595.050 ;
        RECT 421.950 594.600 424.050 595.050 ;
        RECT 205.950 593.400 424.050 594.600 ;
        RECT 205.950 592.950 208.050 593.400 ;
        RECT 247.950 592.950 250.050 593.400 ;
        RECT 421.950 592.950 424.050 593.400 ;
        RECT 580.950 594.600 583.050 595.050 ;
        RECT 601.950 594.600 604.050 595.050 ;
        RECT 580.950 593.400 604.050 594.600 ;
        RECT 580.950 592.950 583.050 593.400 ;
        RECT 601.950 592.950 604.050 593.400 ;
        RECT 637.950 594.600 640.050 595.050 ;
        RECT 658.950 594.600 661.050 595.050 ;
        RECT 637.950 593.400 661.050 594.600 ;
        RECT 637.950 592.950 640.050 593.400 ;
        RECT 658.950 592.950 661.050 593.400 ;
        RECT 748.950 594.600 751.050 595.050 ;
        RECT 799.950 594.600 802.050 595.050 ;
        RECT 748.950 593.400 802.050 594.600 ;
        RECT 748.950 592.950 751.050 593.400 ;
        RECT 799.950 592.950 802.050 593.400 ;
        RECT 859.950 594.600 862.050 595.050 ;
        RECT 871.950 594.600 874.050 595.050 ;
        RECT 859.950 593.400 874.050 594.600 ;
        RECT 859.950 592.950 862.050 593.400 ;
        RECT 871.950 592.950 874.050 593.400 ;
        RECT 928.950 594.600 931.050 595.050 ;
        RECT 940.800 594.600 942.900 595.050 ;
        RECT 928.950 593.400 942.900 594.600 ;
        RECT 928.950 592.950 931.050 593.400 ;
        RECT 940.800 592.950 942.900 593.400 ;
        RECT 943.950 594.600 946.050 595.050 ;
        RECT 964.950 594.600 967.050 595.050 ;
        RECT 943.950 593.400 967.050 594.600 ;
        RECT 943.950 592.950 946.050 593.400 ;
        RECT 964.950 592.950 967.050 593.400 ;
        RECT 58.950 591.600 61.050 592.050 ;
        RECT 73.950 591.600 76.050 592.050 ;
        RECT 58.950 590.400 76.050 591.600 ;
        RECT 58.950 589.950 61.050 590.400 ;
        RECT 73.950 589.950 76.050 590.400 ;
        RECT 247.950 591.600 250.050 591.900 ;
        RECT 307.950 591.600 310.050 592.050 ;
        RECT 247.950 590.400 310.050 591.600 ;
        RECT 247.950 589.800 250.050 590.400 ;
        RECT 307.950 589.950 310.050 590.400 ;
        RECT 559.950 591.600 562.050 592.050 ;
        RECT 574.950 591.600 577.050 592.050 ;
        RECT 559.950 590.400 577.050 591.600 ;
        RECT 559.950 589.950 562.050 590.400 ;
        RECT 574.950 589.950 577.050 590.400 ;
        RECT 661.950 591.600 664.050 592.050 ;
        RECT 736.950 591.600 739.050 592.050 ;
        RECT 661.950 590.400 739.050 591.600 ;
        RECT 661.950 589.950 664.050 590.400 ;
        RECT 736.950 589.950 739.050 590.400 ;
        RECT 910.950 591.600 913.050 592.050 ;
        RECT 919.950 591.600 922.050 592.050 ;
        RECT 910.950 590.400 922.050 591.600 ;
        RECT 910.950 589.950 913.050 590.400 ;
        RECT 919.950 589.950 922.050 590.400 ;
        RECT 967.950 591.600 970.050 592.050 ;
        RECT 985.950 591.600 988.050 592.050 ;
        RECT 967.950 590.400 988.050 591.600 ;
        RECT 967.950 589.950 970.050 590.400 ;
        RECT 985.950 589.950 988.050 590.400 ;
        RECT 106.950 588.600 109.050 589.050 ;
        RECT 163.950 588.600 166.050 589.050 ;
        RECT 106.950 587.400 166.050 588.600 ;
        RECT 106.950 586.950 109.050 587.400 ;
        RECT 163.950 586.950 166.050 587.400 ;
        RECT 211.950 588.600 214.050 589.050 ;
        RECT 244.950 588.600 247.050 589.050 ;
        RECT 295.950 588.600 298.050 589.050 ;
        RECT 211.950 587.400 247.050 588.600 ;
        RECT 211.950 586.950 214.050 587.400 ;
        RECT 244.950 586.950 247.050 587.400 ;
        RECT 248.400 587.400 298.050 588.600 ;
        RECT 139.950 585.600 142.050 586.050 ;
        RECT 154.950 585.600 157.050 586.050 ;
        RECT 139.950 584.400 157.050 585.600 ;
        RECT 139.950 583.950 142.050 584.400 ;
        RECT 154.950 583.950 157.050 584.400 ;
        RECT 220.950 585.600 223.050 586.050 ;
        RECT 248.400 585.600 249.600 587.400 ;
        RECT 295.950 586.950 298.050 587.400 ;
        RECT 319.950 588.600 322.050 589.050 ;
        RECT 331.950 588.600 334.050 589.050 ;
        RECT 319.950 587.400 334.050 588.600 ;
        RECT 319.950 586.950 322.050 587.400 ;
        RECT 331.950 586.950 334.050 587.400 ;
        RECT 376.950 588.600 379.050 589.050 ;
        RECT 475.950 588.600 478.050 589.050 ;
        RECT 376.950 587.400 478.050 588.600 ;
        RECT 376.950 586.950 379.050 587.400 ;
        RECT 475.950 586.950 478.050 587.400 ;
        RECT 487.950 588.600 490.050 589.050 ;
        RECT 547.950 588.600 550.050 589.050 ;
        RECT 487.950 587.400 550.050 588.600 ;
        RECT 487.950 586.950 490.050 587.400 ;
        RECT 547.950 586.950 550.050 587.400 ;
        RECT 589.950 588.600 592.050 589.050 ;
        RECT 640.950 588.600 643.050 589.050 ;
        RECT 589.950 587.400 643.050 588.600 ;
        RECT 589.950 586.950 592.050 587.400 ;
        RECT 640.950 586.950 643.050 587.400 ;
        RECT 670.950 588.600 673.050 589.050 ;
        RECT 682.950 588.600 685.050 589.050 ;
        RECT 670.950 587.400 685.050 588.600 ;
        RECT 670.950 586.950 673.050 587.400 ;
        RECT 682.950 586.950 685.050 587.400 ;
        RECT 688.950 588.600 691.050 589.050 ;
        RECT 745.950 588.600 748.050 589.050 ;
        RECT 688.950 587.400 748.050 588.600 ;
        RECT 688.950 586.950 691.050 587.400 ;
        RECT 745.950 586.950 748.050 587.400 ;
        RECT 901.950 588.600 904.050 589.050 ;
        RECT 922.950 588.600 925.050 589.050 ;
        RECT 937.950 588.600 940.050 589.050 ;
        RECT 901.950 587.400 940.050 588.600 ;
        RECT 901.950 586.950 904.050 587.400 ;
        RECT 922.950 586.950 925.050 587.400 ;
        RECT 937.950 586.950 940.050 587.400 ;
        RECT 988.950 588.600 991.050 589.050 ;
        RECT 1003.950 588.600 1006.050 589.050 ;
        RECT 988.950 587.400 1006.050 588.600 ;
        RECT 988.950 586.950 991.050 587.400 ;
        RECT 1003.950 586.950 1006.050 587.400 ;
        RECT 220.950 584.400 249.600 585.600 ;
        RECT 298.950 585.600 301.050 586.050 ;
        RECT 304.950 585.600 307.050 586.050 ;
        RECT 298.950 584.400 307.050 585.600 ;
        RECT 220.950 583.950 223.050 584.400 ;
        RECT 298.950 583.950 301.050 584.400 ;
        RECT 304.950 583.950 307.050 584.400 ;
        RECT 394.950 585.600 397.050 586.050 ;
        RECT 427.950 585.600 430.050 586.050 ;
        RECT 394.950 584.400 430.050 585.600 ;
        RECT 394.950 583.950 397.050 584.400 ;
        RECT 427.950 583.950 430.050 584.400 ;
        RECT 451.950 585.600 454.050 586.050 ;
        RECT 541.950 585.600 544.050 586.050 ;
        RECT 451.950 584.400 544.050 585.600 ;
        RECT 451.950 583.950 454.050 584.400 ;
        RECT 541.950 583.950 544.050 584.400 ;
        RECT 604.950 585.600 607.050 586.050 ;
        RECT 610.950 585.600 613.050 586.050 ;
        RECT 604.950 584.400 613.050 585.600 ;
        RECT 604.950 583.950 607.050 584.400 ;
        RECT 610.950 583.950 613.050 584.400 ;
        RECT 718.950 585.600 721.050 586.050 ;
        RECT 724.950 585.600 727.050 586.050 ;
        RECT 718.950 584.400 727.050 585.600 ;
        RECT 718.950 583.950 721.050 584.400 ;
        RECT 724.950 583.950 727.050 584.400 ;
        RECT 730.950 585.600 733.050 586.050 ;
        RECT 742.950 585.600 745.050 586.050 ;
        RECT 730.950 584.400 745.050 585.600 ;
        RECT 730.950 583.950 733.050 584.400 ;
        RECT 742.950 583.950 745.050 584.400 ;
        RECT 862.950 585.600 865.050 586.050 ;
        RECT 877.950 585.600 880.050 586.050 ;
        RECT 862.950 584.400 880.050 585.600 ;
        RECT 862.950 583.950 865.050 584.400 ;
        RECT 877.950 583.950 880.050 584.400 ;
        RECT 949.950 585.600 952.050 586.050 ;
        RECT 961.950 585.600 964.050 586.050 ;
        RECT 994.950 585.600 997.050 586.050 ;
        RECT 949.950 584.400 997.050 585.600 ;
        RECT 949.950 583.950 952.050 584.400 ;
        RECT 961.950 583.950 964.050 584.400 ;
        RECT 994.950 583.950 997.050 584.400 ;
        RECT 145.950 582.600 148.050 583.050 ;
        RECT 199.950 582.600 202.050 583.050 ;
        RECT 145.950 581.400 202.050 582.600 ;
        RECT 145.950 580.950 148.050 581.400 ;
        RECT 199.950 580.950 202.050 581.400 ;
        RECT 364.950 582.600 367.050 583.050 ;
        RECT 415.950 582.600 418.050 583.050 ;
        RECT 364.950 581.400 418.050 582.600 ;
        RECT 364.950 580.950 367.050 581.400 ;
        RECT 415.950 580.950 418.050 581.400 ;
        RECT 547.950 582.600 550.050 583.050 ;
        RECT 616.950 582.600 619.050 583.050 ;
        RECT 547.950 581.400 619.050 582.600 ;
        RECT 547.950 580.950 550.050 581.400 ;
        RECT 616.950 580.950 619.050 581.400 ;
        RECT 670.950 582.600 673.050 583.050 ;
        RECT 694.950 582.600 697.050 583.050 ;
        RECT 670.950 581.400 697.050 582.600 ;
        RECT 670.950 580.950 673.050 581.400 ;
        RECT 694.950 580.950 697.050 581.400 ;
        RECT 718.950 582.600 721.050 582.900 ;
        RECT 751.950 582.600 754.050 583.050 ;
        RECT 790.950 582.600 793.050 583.050 ;
        RECT 718.950 581.400 793.050 582.600 ;
        RECT 718.950 580.800 721.050 581.400 ;
        RECT 751.950 580.950 754.050 581.400 ;
        RECT 790.950 580.950 793.050 581.400 ;
        RECT 901.950 582.600 904.050 583.050 ;
        RECT 907.950 582.600 910.050 583.050 ;
        RECT 901.950 581.400 910.050 582.600 ;
        RECT 901.950 580.950 904.050 581.400 ;
        RECT 907.950 580.950 910.050 581.400 ;
        RECT 976.950 582.600 979.050 583.050 ;
        RECT 1003.950 582.600 1006.050 583.050 ;
        RECT 976.950 581.400 1006.050 582.600 ;
        RECT 976.950 580.950 979.050 581.400 ;
        RECT 1003.950 580.950 1006.050 581.400 ;
        RECT 229.950 579.600 232.050 580.050 ;
        RECT 271.950 579.600 274.050 580.050 ;
        RECT 229.950 578.400 274.050 579.600 ;
        RECT 229.950 577.950 232.050 578.400 ;
        RECT 271.950 577.950 274.050 578.400 ;
        RECT 277.950 579.600 280.050 580.050 ;
        RECT 340.950 579.600 343.050 580.050 ;
        RECT 277.950 578.400 343.050 579.600 ;
        RECT 277.950 577.950 280.050 578.400 ;
        RECT 340.950 577.950 343.050 578.400 ;
        RECT 349.950 579.600 352.050 580.050 ;
        RECT 370.950 579.600 373.050 580.050 ;
        RECT 349.950 578.400 373.050 579.600 ;
        RECT 349.950 577.950 352.050 578.400 ;
        RECT 370.950 577.950 373.050 578.400 ;
        RECT 505.950 579.600 508.050 580.050 ;
        RECT 511.950 579.600 514.050 580.050 ;
        RECT 505.950 578.400 514.050 579.600 ;
        RECT 505.950 577.950 508.050 578.400 ;
        RECT 511.950 577.950 514.050 578.400 ;
        RECT 541.950 579.600 544.050 580.050 ;
        RECT 613.950 579.600 616.050 580.050 ;
        RECT 649.950 579.600 652.050 580.050 ;
        RECT 541.950 578.400 616.050 579.600 ;
        RECT 541.950 577.950 544.050 578.400 ;
        RECT 613.950 577.950 616.050 578.400 ;
        RECT 638.400 578.400 652.050 579.600 ;
        RECT 52.950 576.600 55.050 577.050 ;
        RECT 64.950 576.600 67.050 577.050 ;
        RECT 52.950 575.400 67.050 576.600 ;
        RECT 52.950 574.950 55.050 575.400 ;
        RECT 64.950 574.950 67.050 575.400 ;
        RECT 187.950 576.600 190.050 577.050 ;
        RECT 205.950 576.600 208.050 577.050 ;
        RECT 187.950 575.400 208.050 576.600 ;
        RECT 187.950 574.950 190.050 575.400 ;
        RECT 205.950 574.950 208.050 575.400 ;
        RECT 214.950 576.600 217.050 577.050 ;
        RECT 223.950 576.600 226.050 577.050 ;
        RECT 214.950 575.400 226.050 576.600 ;
        RECT 214.950 574.950 217.050 575.400 ;
        RECT 223.950 574.950 226.050 575.400 ;
        RECT 466.950 576.600 469.050 577.050 ;
        RECT 493.950 576.600 496.050 577.050 ;
        RECT 502.950 576.600 505.050 577.050 ;
        RECT 466.950 575.400 492.600 576.600 ;
        RECT 466.950 574.950 469.050 575.400 ;
        RECT 97.950 572.100 100.050 574.200 ;
        RECT 103.950 573.600 106.050 574.050 ;
        RECT 115.950 573.600 118.050 574.050 ;
        RECT 103.950 572.400 118.050 573.600 ;
        RECT 22.950 567.450 25.050 567.900 ;
        RECT 28.950 567.450 31.050 567.900 ;
        RECT 22.950 566.250 31.050 567.450 ;
        RECT 98.400 567.600 99.600 572.100 ;
        RECT 103.950 571.950 106.050 572.400 ;
        RECT 115.950 571.950 118.050 572.400 ;
        RECT 151.950 572.100 154.050 574.200 ;
        RECT 157.950 573.600 160.050 574.200 ;
        RECT 169.950 573.600 172.050 574.050 ;
        RECT 157.950 572.400 172.050 573.600 ;
        RECT 157.950 572.100 160.050 572.400 ;
        RECT 103.950 567.600 106.050 568.050 ;
        RECT 98.400 566.400 106.050 567.600 ;
        RECT 22.950 565.800 25.050 566.250 ;
        RECT 28.950 565.800 31.050 566.250 ;
        RECT 103.950 565.950 106.050 566.400 ;
        RECT 124.950 567.450 127.050 567.900 ;
        RECT 145.950 567.450 148.050 567.900 ;
        RECT 124.950 566.250 148.050 567.450 ;
        RECT 124.950 565.800 127.050 566.250 ;
        RECT 145.950 565.800 148.050 566.250 ;
        RECT 152.400 565.050 153.600 572.100 ;
        RECT 169.950 571.950 172.050 572.400 ;
        RECT 178.950 573.600 181.050 574.200 ;
        RECT 190.950 573.600 193.050 574.050 ;
        RECT 178.950 572.400 193.050 573.600 ;
        RECT 178.950 572.100 181.050 572.400 ;
        RECT 190.950 571.950 193.050 572.400 ;
        RECT 238.950 573.750 241.050 574.200 ;
        RECT 253.800 573.750 255.900 574.200 ;
        RECT 238.950 572.550 255.900 573.750 ;
        RECT 238.950 572.100 241.050 572.550 ;
        RECT 253.800 572.100 255.900 572.550 ;
        RECT 256.950 573.600 259.050 574.050 ;
        RECT 268.950 573.600 271.050 574.200 ;
        RECT 256.950 572.400 271.050 573.600 ;
        RECT 256.950 571.950 259.050 572.400 ;
        RECT 268.950 572.100 271.050 572.400 ;
        RECT 280.950 573.600 283.050 574.050 ;
        RECT 292.950 573.600 295.050 574.200 ;
        RECT 280.950 572.400 295.050 573.600 ;
        RECT 280.950 571.950 283.050 572.400 ;
        RECT 292.950 572.100 295.050 572.400 ;
        RECT 298.950 573.600 303.000 574.050 ;
        RECT 328.950 573.600 331.050 574.200 ;
        RECT 340.950 573.600 343.050 574.050 ;
        RECT 346.950 573.600 349.050 574.200 ;
        RECT 375.000 573.600 379.050 574.050 ;
        RECT 391.950 573.600 394.050 574.050 ;
        RECT 298.950 571.950 303.600 573.600 ;
        RECT 328.950 572.400 349.050 573.600 ;
        RECT 328.950 572.100 331.050 572.400 ;
        RECT 340.950 571.950 343.050 572.400 ;
        RECT 346.950 572.100 349.050 572.400 ;
        RECT 374.400 571.950 379.050 573.600 ;
        RECT 380.400 572.400 394.050 573.600 ;
        RECT 302.400 567.900 303.600 571.950 ;
        RECT 374.400 567.900 375.600 571.950 ;
        RECT 380.400 567.900 381.600 572.400 ;
        RECT 391.950 571.950 394.050 572.400 ;
        RECT 406.950 573.750 409.050 574.200 ;
        RECT 412.950 573.750 415.050 574.200 ;
        RECT 406.950 573.600 415.050 573.750 ;
        RECT 418.950 573.600 421.050 574.050 ;
        RECT 406.950 572.550 421.050 573.600 ;
        RECT 406.950 572.100 409.050 572.550 ;
        RECT 412.950 572.400 421.050 572.550 ;
        RECT 412.950 572.100 415.050 572.400 ;
        RECT 418.950 571.950 421.050 572.400 ;
        RECT 430.950 573.600 433.050 574.200 ;
        RECT 439.950 573.750 442.050 574.200 ;
        RECT 448.950 573.750 451.050 574.200 ;
        RECT 430.950 572.400 438.600 573.600 ;
        RECT 430.950 572.100 433.050 572.400 ;
        RECT 437.400 568.050 438.600 572.400 ;
        RECT 439.950 572.550 451.050 573.750 ;
        RECT 486.000 573.600 490.050 574.050 ;
        RECT 439.950 572.100 442.050 572.550 ;
        RECT 448.950 572.100 451.050 572.550 ;
        RECT 485.400 571.950 490.050 573.600 ;
        RECT 190.950 567.450 193.050 567.900 ;
        RECT 196.950 567.450 199.050 567.900 ;
        RECT 190.950 566.250 199.050 567.450 ;
        RECT 190.950 565.800 193.050 566.250 ;
        RECT 196.950 565.800 199.050 566.250 ;
        RECT 202.950 567.450 205.050 567.900 ;
        RECT 211.950 567.450 214.050 567.900 ;
        RECT 202.950 566.250 214.050 567.450 ;
        RECT 202.950 565.800 205.050 566.250 ;
        RECT 211.950 565.800 214.050 566.250 ;
        RECT 223.950 567.600 226.050 567.900 ;
        RECT 241.950 567.600 244.050 567.900 ;
        RECT 223.950 566.400 244.050 567.600 ;
        RECT 223.950 565.800 226.050 566.400 ;
        RECT 241.950 565.800 244.050 566.400 ;
        RECT 247.950 567.450 250.050 567.900 ;
        RECT 256.950 567.450 259.050 567.900 ;
        RECT 247.950 566.250 259.050 567.450 ;
        RECT 247.950 565.800 250.050 566.250 ;
        RECT 256.950 565.800 259.050 566.250 ;
        RECT 271.950 567.450 274.050 567.900 ;
        RECT 277.950 567.450 280.050 567.900 ;
        RECT 271.950 566.250 280.050 567.450 ;
        RECT 271.950 565.800 274.050 566.250 ;
        RECT 277.950 565.800 280.050 566.250 ;
        RECT 301.950 565.800 304.050 567.900 ;
        RECT 310.950 567.450 313.050 567.900 ;
        RECT 337.950 567.450 340.050 567.900 ;
        RECT 310.950 566.250 340.050 567.450 ;
        RECT 310.950 565.800 313.050 566.250 ;
        RECT 337.950 565.800 340.050 566.250 ;
        RECT 349.950 567.600 352.050 567.900 ;
        RECT 367.950 567.600 370.050 567.900 ;
        RECT 349.950 566.400 370.050 567.600 ;
        RECT 349.950 565.800 352.050 566.400 ;
        RECT 367.950 565.800 370.050 566.400 ;
        RECT 373.950 565.800 376.050 567.900 ;
        RECT 379.950 565.800 382.050 567.900 ;
        RECT 388.950 567.450 391.050 567.900 ;
        RECT 394.950 567.450 397.050 567.900 ;
        RECT 388.950 566.250 397.050 567.450 ;
        RECT 388.950 565.800 391.050 566.250 ;
        RECT 394.950 565.800 397.050 566.250 ;
        RECT 436.950 565.950 439.050 568.050 ;
        RECT 485.400 567.900 486.600 571.950 ;
        RECT 451.950 567.450 454.050 567.900 ;
        RECT 457.950 567.450 460.050 567.900 ;
        RECT 451.950 566.250 460.050 567.450 ;
        RECT 451.950 565.800 454.050 566.250 ;
        RECT 457.950 565.800 460.050 566.250 ;
        RECT 466.950 567.600 469.050 567.900 ;
        RECT 475.950 567.600 478.050 567.900 ;
        RECT 466.950 566.400 478.050 567.600 ;
        RECT 466.950 565.800 469.050 566.400 ;
        RECT 475.950 565.800 478.050 566.400 ;
        RECT 484.950 565.800 487.050 567.900 ;
        RECT 37.950 564.600 40.050 565.050 ;
        RECT 43.950 564.600 46.050 565.050 ;
        RECT 70.950 564.600 73.050 565.050 ;
        RECT 37.950 563.400 73.050 564.600 ;
        RECT 37.950 562.950 40.050 563.400 ;
        RECT 43.950 562.950 46.050 563.400 ;
        RECT 70.950 562.950 73.050 563.400 ;
        RECT 151.950 562.950 154.050 565.050 ;
        RECT 253.950 564.600 256.050 565.050 ;
        RECT 265.950 564.600 268.050 565.050 ;
        RECT 283.950 564.600 286.050 565.050 ;
        RECT 289.950 564.600 292.050 565.050 ;
        RECT 253.950 563.400 292.050 564.600 ;
        RECT 253.950 562.950 256.050 563.400 ;
        RECT 265.950 562.950 268.050 563.400 ;
        RECT 283.950 562.950 286.050 563.400 ;
        RECT 289.950 562.950 292.050 563.400 ;
        RECT 397.950 564.600 400.050 565.050 ;
        RECT 412.950 564.600 415.050 565.050 ;
        RECT 397.950 563.400 415.050 564.600 ;
        RECT 491.400 564.600 492.600 575.400 ;
        RECT 493.950 575.400 505.050 576.600 ;
        RECT 493.950 574.950 496.050 575.400 ;
        RECT 502.950 574.950 505.050 575.400 ;
        RECT 613.950 576.600 616.050 576.900 ;
        RECT 638.400 576.600 639.600 578.400 ;
        RECT 649.950 577.950 652.050 578.400 ;
        RECT 709.950 579.600 712.050 580.050 ;
        RECT 748.950 579.600 751.050 580.050 ;
        RECT 709.950 578.400 751.050 579.600 ;
        RECT 709.950 577.950 712.050 578.400 ;
        RECT 748.950 577.950 751.050 578.400 ;
        RECT 889.950 579.600 892.050 580.050 ;
        RECT 931.800 579.600 933.900 580.050 ;
        RECT 889.950 578.400 933.900 579.600 ;
        RECT 889.950 577.950 892.050 578.400 ;
        RECT 931.800 577.950 933.900 578.400 ;
        RECT 934.950 579.600 937.050 580.050 ;
        RECT 940.950 579.600 943.050 580.050 ;
        RECT 934.950 578.400 943.050 579.600 ;
        RECT 934.950 577.950 937.050 578.400 ;
        RECT 940.950 577.950 943.050 578.400 ;
        RECT 1009.950 577.950 1012.050 580.050 ;
        RECT 613.950 575.400 639.600 576.600 ;
        RECT 835.950 576.600 838.050 577.050 ;
        RECT 853.950 576.600 856.050 577.050 ;
        RECT 859.950 576.600 862.050 577.050 ;
        RECT 835.950 575.400 862.050 576.600 ;
        RECT 613.950 574.800 616.050 575.400 ;
        RECT 835.950 574.950 838.050 575.400 ;
        RECT 853.950 574.950 856.050 575.400 ;
        RECT 859.950 574.950 862.050 575.400 ;
        RECT 958.950 576.600 961.050 577.050 ;
        RECT 973.950 576.600 976.050 577.050 ;
        RECT 982.950 576.600 985.050 577.050 ;
        RECT 958.950 575.400 985.050 576.600 ;
        RECT 958.950 574.950 961.050 575.400 ;
        RECT 973.950 574.950 976.050 575.400 ;
        RECT 982.950 574.950 985.050 575.400 ;
        RECT 514.950 573.600 517.050 574.050 ;
        RECT 520.950 573.600 523.050 574.200 ;
        RECT 514.950 572.400 523.050 573.600 ;
        RECT 514.950 571.950 517.050 572.400 ;
        RECT 520.950 572.100 523.050 572.400 ;
        RECT 541.950 573.750 544.050 574.200 ;
        RECT 553.950 573.750 556.050 574.200 ;
        RECT 541.950 572.550 556.050 573.750 ;
        RECT 589.950 573.600 592.050 574.200 ;
        RECT 609.000 573.600 613.050 574.050 ;
        RECT 541.950 572.100 544.050 572.550 ;
        RECT 553.950 572.100 556.050 572.550 ;
        RECT 569.400 572.400 592.050 573.600 ;
        RECT 529.950 565.950 532.050 568.050 ;
        RECT 544.950 567.600 547.050 567.900 ;
        RECT 550.950 567.600 553.050 568.050 ;
        RECT 569.400 567.900 570.600 572.400 ;
        RECT 589.950 572.100 592.050 572.400 ;
        RECT 608.400 571.950 613.050 573.600 ;
        RECT 640.950 571.950 643.050 574.050 ;
        RECT 646.950 573.600 649.050 574.200 ;
        RECT 670.950 573.600 673.050 574.200 ;
        RECT 646.950 572.400 673.050 573.600 ;
        RECT 646.950 572.100 649.050 572.400 ;
        RECT 670.950 572.100 673.050 572.400 ;
        RECT 676.950 573.600 679.050 574.200 ;
        RECT 700.950 573.600 703.050 574.200 ;
        RECT 676.950 572.400 690.600 573.600 ;
        RECT 676.950 572.100 679.050 572.400 ;
        RECT 608.400 567.900 609.600 571.950 ;
        RECT 544.950 566.400 553.050 567.600 ;
        RECT 502.950 564.600 505.050 565.050 ;
        RECT 491.400 563.400 505.050 564.600 ;
        RECT 397.950 562.950 400.050 563.400 ;
        RECT 412.950 562.950 415.050 563.400 ;
        RECT 502.950 562.950 505.050 563.400 ;
        RECT 295.950 561.600 298.050 562.050 ;
        RECT 319.950 561.600 322.050 562.050 ;
        RECT 295.950 560.400 322.050 561.600 ;
        RECT 295.950 559.950 298.050 560.400 ;
        RECT 319.950 559.950 322.050 560.400 ;
        RECT 523.950 561.600 526.050 562.050 ;
        RECT 530.400 561.600 531.600 565.950 ;
        RECT 544.950 565.800 547.050 566.400 ;
        RECT 550.950 565.950 553.050 566.400 ;
        RECT 568.950 565.800 571.050 567.900 ;
        RECT 607.950 565.800 610.050 567.900 ;
        RECT 641.400 567.600 642.600 571.950 ;
        RECT 643.950 567.600 646.050 567.900 ;
        RECT 641.400 566.400 646.050 567.600 ;
        RECT 643.950 565.800 646.050 566.400 ;
        RECT 538.950 564.600 541.050 565.050 ;
        RECT 577.950 564.600 580.050 565.050 ;
        RECT 538.950 563.400 580.050 564.600 ;
        RECT 538.950 562.950 541.050 563.400 ;
        RECT 577.950 562.950 580.050 563.400 ;
        RECT 523.950 560.400 531.600 561.600 ;
        RECT 580.950 561.600 583.050 562.050 ;
        RECT 589.950 561.600 592.050 562.050 ;
        RECT 580.950 560.400 592.050 561.600 ;
        RECT 523.950 559.950 526.050 560.400 ;
        RECT 580.950 559.950 583.050 560.400 ;
        RECT 589.950 559.950 592.050 560.400 ;
        RECT 616.950 561.600 619.050 562.050 ;
        RECT 667.950 561.600 670.050 562.050 ;
        RECT 679.950 561.600 682.050 562.050 ;
        RECT 616.950 560.400 682.050 561.600 ;
        RECT 689.400 561.600 690.600 572.400 ;
        RECT 700.950 572.400 714.600 573.600 ;
        RECT 700.950 572.100 703.050 572.400 ;
        RECT 713.400 570.600 714.600 572.400 ;
        RECT 724.950 571.950 727.050 574.050 ;
        RECT 736.950 573.600 739.050 574.200 ;
        RECT 748.950 573.600 751.050 574.050 ;
        RECT 736.950 572.400 751.050 573.600 ;
        RECT 736.950 572.100 739.050 572.400 ;
        RECT 748.950 571.950 751.050 572.400 ;
        RECT 754.950 573.750 757.050 574.200 ;
        RECT 763.950 573.750 766.050 574.200 ;
        RECT 754.950 572.550 766.050 573.750 ;
        RECT 754.950 572.100 757.050 572.550 ;
        RECT 763.950 572.100 766.050 572.550 ;
        RECT 769.950 573.600 772.050 574.200 ;
        RECT 781.950 573.600 784.050 574.050 ;
        RECT 769.950 572.400 784.050 573.600 ;
        RECT 769.950 572.100 772.050 572.400 ;
        RECT 781.950 571.950 784.050 572.400 ;
        RECT 811.950 573.750 814.050 574.200 ;
        RECT 826.950 573.750 829.050 574.200 ;
        RECT 811.950 572.550 829.050 573.750 ;
        RECT 811.950 572.100 814.050 572.550 ;
        RECT 826.950 572.100 829.050 572.550 ;
        RECT 841.950 573.600 844.050 574.200 ;
        RECT 865.950 573.600 868.050 574.200 ;
        RECT 874.950 573.600 877.050 574.050 ;
        RECT 841.950 573.000 855.600 573.600 ;
        RECT 841.950 572.400 856.050 573.000 ;
        RECT 841.950 572.100 844.050 572.400 ;
        RECT 713.400 569.400 723.600 570.600 ;
        RECT 691.950 564.600 694.050 565.050 ;
        RECT 709.950 564.600 712.050 565.050 ;
        RECT 691.950 563.400 712.050 564.600 ;
        RECT 722.400 564.600 723.600 569.400 ;
        RECT 725.400 568.050 726.600 571.950 ;
        RECT 853.950 568.950 856.050 572.400 ;
        RECT 865.950 572.400 877.050 573.600 ;
        RECT 865.950 572.100 868.050 572.400 ;
        RECT 874.950 571.950 877.050 572.400 ;
        RECT 910.950 572.100 913.050 574.200 ;
        RECT 922.950 573.600 927.000 574.050 ;
        RECT 934.950 573.600 937.050 574.200 ;
        RECT 946.950 573.600 949.050 574.050 ;
        RECT 911.400 568.050 912.600 572.100 ;
        RECT 922.950 571.950 927.600 573.600 ;
        RECT 934.950 572.400 949.050 573.600 ;
        RECT 934.950 572.100 937.050 572.400 ;
        RECT 946.950 571.950 949.050 572.400 ;
        RECT 952.950 573.600 955.050 574.200 ;
        RECT 1010.400 573.600 1011.600 577.950 ;
        RECT 952.950 572.400 1011.600 573.600 ;
        RECT 952.950 572.100 955.050 572.400 ;
        RECT 1012.950 571.950 1015.050 574.050 ;
        RECT 724.950 565.950 727.050 568.050 ;
        RECT 745.950 567.450 748.050 567.900 ;
        RECT 751.950 567.600 754.050 567.900 ;
        RECT 766.950 567.600 769.050 567.900 ;
        RECT 751.950 567.450 769.050 567.600 ;
        RECT 745.950 566.400 769.050 567.450 ;
        RECT 745.950 566.250 754.050 566.400 ;
        RECT 745.950 565.800 748.050 566.250 ;
        RECT 751.950 565.800 754.050 566.250 ;
        RECT 766.950 565.800 769.050 566.400 ;
        RECT 778.950 567.450 781.050 567.900 ;
        RECT 814.950 567.450 817.050 567.900 ;
        RECT 778.950 566.250 817.050 567.450 ;
        RECT 778.950 565.800 781.050 566.250 ;
        RECT 814.950 565.800 817.050 566.250 ;
        RECT 823.950 567.450 826.050 567.900 ;
        RECT 838.950 567.600 841.050 567.900 ;
        RECT 862.950 567.600 865.050 567.900 ;
        RECT 838.950 567.450 865.050 567.600 ;
        RECT 823.950 566.400 865.050 567.450 ;
        RECT 823.950 566.250 841.050 566.400 ;
        RECT 823.950 565.800 826.050 566.250 ;
        RECT 838.950 565.800 841.050 566.250 ;
        RECT 862.950 565.800 865.050 566.400 ;
        RECT 886.950 567.600 889.050 567.900 ;
        RECT 898.950 567.600 901.050 568.050 ;
        RECT 886.950 566.400 901.050 567.600 ;
        RECT 911.400 566.400 916.050 568.050 ;
        RECT 926.400 567.900 927.600 571.950 ;
        RECT 1013.400 568.050 1014.600 571.950 ;
        RECT 886.950 565.800 889.050 566.400 ;
        RECT 898.950 565.950 901.050 566.400 ;
        RECT 912.000 565.950 916.050 566.400 ;
        RECT 925.950 565.800 928.050 567.900 ;
        RECT 961.950 567.600 964.050 567.900 ;
        RECT 979.950 567.600 982.050 567.900 ;
        RECT 961.950 566.400 982.050 567.600 ;
        RECT 961.950 565.800 964.050 566.400 ;
        RECT 979.950 565.800 982.050 566.400 ;
        RECT 997.950 567.450 1000.050 567.900 ;
        RECT 1006.950 567.450 1009.050 567.900 ;
        RECT 997.950 566.250 1009.050 567.450 ;
        RECT 997.950 565.800 1000.050 566.250 ;
        RECT 1006.950 565.800 1009.050 566.250 ;
        RECT 1012.950 565.950 1015.050 568.050 ;
        RECT 763.950 564.600 766.050 565.050 ;
        RECT 722.400 563.400 766.050 564.600 ;
        RECT 691.950 562.950 694.050 563.400 ;
        RECT 709.950 562.950 712.050 563.400 ;
        RECT 763.950 562.950 766.050 563.400 ;
        RECT 946.950 564.600 949.050 565.050 ;
        RECT 961.950 564.600 964.050 565.050 ;
        RECT 946.950 563.400 964.050 564.600 ;
        RECT 946.950 562.950 949.050 563.400 ;
        RECT 961.950 562.950 964.050 563.400 ;
        RECT 823.950 561.600 826.050 562.050 ;
        RECT 689.400 560.400 826.050 561.600 ;
        RECT 616.950 559.950 619.050 560.400 ;
        RECT 667.950 559.950 670.050 560.400 ;
        RECT 679.950 559.950 682.050 560.400 ;
        RECT 823.950 559.950 826.050 560.400 ;
        RECT 844.950 561.600 847.050 562.050 ;
        RECT 913.950 561.600 916.050 562.050 ;
        RECT 844.950 560.400 916.050 561.600 ;
        RECT 844.950 559.950 847.050 560.400 ;
        RECT 913.950 559.950 916.050 560.400 ;
        RECT 967.950 561.600 970.050 562.050 ;
        RECT 973.950 561.600 976.050 562.050 ;
        RECT 967.950 560.400 976.050 561.600 ;
        RECT 967.950 559.950 970.050 560.400 ;
        RECT 973.950 559.950 976.050 560.400 ;
        RECT 28.950 558.600 31.050 559.050 ;
        RECT 88.950 558.600 91.050 559.050 ;
        RECT 154.950 558.600 157.050 559.050 ;
        RECT 28.950 557.400 157.050 558.600 ;
        RECT 28.950 556.950 31.050 557.400 ;
        RECT 88.950 556.950 91.050 557.400 ;
        RECT 154.950 556.950 157.050 557.400 ;
        RECT 433.950 558.600 436.050 559.050 ;
        RECT 448.950 558.600 451.050 559.050 ;
        RECT 538.950 558.600 541.050 559.050 ;
        RECT 433.950 557.400 541.050 558.600 ;
        RECT 433.950 556.950 436.050 557.400 ;
        RECT 448.950 556.950 451.050 557.400 ;
        RECT 538.950 556.950 541.050 557.400 ;
        RECT 559.950 558.600 562.050 559.050 ;
        RECT 592.950 558.600 595.050 559.050 ;
        RECT 613.950 558.600 616.050 559.050 ;
        RECT 559.950 557.400 616.050 558.600 ;
        RECT 559.950 556.950 562.050 557.400 ;
        RECT 592.950 556.950 595.050 557.400 ;
        RECT 613.950 556.950 616.050 557.400 ;
        RECT 727.950 558.600 730.050 559.050 ;
        RECT 760.950 558.600 763.050 559.050 ;
        RECT 727.950 557.400 763.050 558.600 ;
        RECT 727.950 556.950 730.050 557.400 ;
        RECT 760.950 556.950 763.050 557.400 ;
        RECT 829.950 558.600 832.050 559.050 ;
        RECT 925.950 558.600 928.050 559.050 ;
        RECT 829.950 557.400 928.050 558.600 ;
        RECT 829.950 556.950 832.050 557.400 ;
        RECT 925.950 556.950 928.050 557.400 ;
        RECT 931.950 558.600 934.050 559.050 ;
        RECT 967.950 558.600 970.050 558.900 ;
        RECT 931.950 557.400 970.050 558.600 ;
        RECT 931.950 556.950 934.050 557.400 ;
        RECT 967.950 556.800 970.050 557.400 ;
        RECT 334.950 555.600 337.050 556.050 ;
        RECT 376.950 555.600 379.050 556.050 ;
        RECT 532.950 555.600 535.050 556.050 ;
        RECT 334.950 554.400 535.050 555.600 ;
        RECT 334.950 553.950 337.050 554.400 ;
        RECT 376.950 553.950 379.050 554.400 ;
        RECT 532.950 553.950 535.050 554.400 ;
        RECT 553.950 555.600 556.050 556.050 ;
        RECT 586.950 555.600 589.050 556.050 ;
        RECT 592.950 555.600 595.050 555.900 ;
        RECT 553.950 554.400 595.050 555.600 ;
        RECT 553.950 553.950 556.050 554.400 ;
        RECT 586.950 553.950 589.050 554.400 ;
        RECT 592.950 553.800 595.050 554.400 ;
        RECT 673.950 555.600 676.050 556.050 ;
        RECT 691.950 555.600 694.050 556.050 ;
        RECT 673.950 554.400 694.050 555.600 ;
        RECT 673.950 553.950 676.050 554.400 ;
        RECT 691.950 553.950 694.050 554.400 ;
        RECT 784.950 555.600 787.050 556.050 ;
        RECT 814.950 555.600 817.050 556.050 ;
        RECT 820.950 555.600 823.050 556.050 ;
        RECT 838.950 555.600 841.050 556.050 ;
        RECT 784.950 554.400 841.050 555.600 ;
        RECT 784.950 553.950 787.050 554.400 ;
        RECT 814.950 553.950 817.050 554.400 ;
        RECT 820.950 553.950 823.050 554.400 ;
        RECT 838.950 553.950 841.050 554.400 ;
        RECT 868.950 555.600 871.050 556.050 ;
        RECT 907.950 555.600 910.050 556.050 ;
        RECT 868.950 554.400 910.050 555.600 ;
        RECT 868.950 553.950 871.050 554.400 ;
        RECT 907.950 553.950 910.050 554.400 ;
        RECT 991.950 555.600 994.050 556.050 ;
        RECT 1009.950 555.600 1012.050 556.050 ;
        RECT 991.950 554.400 1012.050 555.600 ;
        RECT 991.950 553.950 994.050 554.400 ;
        RECT 1009.950 553.950 1012.050 554.400 ;
        RECT 163.950 552.600 166.050 553.050 ;
        RECT 175.950 552.600 178.050 553.050 ;
        RECT 232.950 552.600 235.050 553.050 ;
        RECT 163.950 551.400 235.050 552.600 ;
        RECT 163.950 550.950 166.050 551.400 ;
        RECT 175.950 550.950 178.050 551.400 ;
        RECT 232.950 550.950 235.050 551.400 ;
        RECT 337.950 552.600 340.050 553.050 ;
        RECT 463.950 552.600 466.050 553.050 ;
        RECT 466.950 552.600 469.050 553.050 ;
        RECT 337.950 551.400 469.050 552.600 ;
        RECT 337.950 550.950 340.050 551.400 ;
        RECT 463.950 550.950 466.050 551.400 ;
        RECT 466.950 550.950 469.050 551.400 ;
        RECT 562.950 552.600 565.050 553.050 ;
        RECT 646.950 552.600 649.050 553.050 ;
        RECT 562.950 551.400 649.050 552.600 ;
        RECT 562.950 550.950 565.050 551.400 ;
        RECT 646.950 550.950 649.050 551.400 ;
        RECT 916.950 552.600 919.050 553.050 ;
        RECT 946.950 552.600 949.050 553.050 ;
        RECT 916.950 551.400 949.050 552.600 ;
        RECT 916.950 550.950 919.050 551.400 ;
        RECT 946.950 550.950 949.050 551.400 ;
        RECT 952.950 552.600 955.050 553.050 ;
        RECT 988.950 552.600 991.050 553.050 ;
        RECT 952.950 551.400 991.050 552.600 ;
        RECT 952.950 550.950 955.050 551.400 ;
        RECT 988.950 550.950 991.050 551.400 ;
        RECT 139.950 549.600 142.050 550.050 ;
        RECT 334.950 549.600 337.050 550.050 ;
        RECT 139.950 548.400 337.050 549.600 ;
        RECT 139.950 547.950 142.050 548.400 ;
        RECT 334.950 547.950 337.050 548.400 ;
        RECT 421.950 549.600 424.050 550.050 ;
        RECT 472.950 549.600 475.050 550.050 ;
        RECT 421.950 548.400 475.050 549.600 ;
        RECT 421.950 547.950 424.050 548.400 ;
        RECT 472.950 547.950 475.050 548.400 ;
        RECT 532.950 549.600 535.050 550.050 ;
        RECT 574.950 549.600 577.050 550.050 ;
        RECT 532.950 548.400 577.050 549.600 ;
        RECT 647.400 549.600 648.600 550.950 ;
        RECT 685.950 549.600 688.050 550.050 ;
        RECT 647.400 548.400 688.050 549.600 ;
        RECT 532.950 547.950 535.050 548.400 ;
        RECT 574.950 547.950 577.050 548.400 ;
        RECT 685.950 547.950 688.050 548.400 ;
        RECT 955.950 549.600 958.050 550.050 ;
        RECT 982.950 549.600 985.050 550.050 ;
        RECT 955.950 548.400 985.050 549.600 ;
        RECT 955.950 547.950 958.050 548.400 ;
        RECT 982.950 547.950 985.050 548.400 ;
        RECT 103.950 546.600 106.050 547.050 ;
        RECT 124.950 546.600 127.050 547.050 ;
        RECT 259.950 546.600 262.050 547.050 ;
        RECT 103.950 545.400 262.050 546.600 ;
        RECT 103.950 544.950 106.050 545.400 ;
        RECT 124.950 544.950 127.050 545.400 ;
        RECT 259.950 544.950 262.050 545.400 ;
        RECT 289.950 546.600 292.050 547.050 ;
        RECT 412.950 546.600 415.050 547.050 ;
        RECT 289.950 545.400 415.050 546.600 ;
        RECT 289.950 544.950 292.050 545.400 ;
        RECT 412.950 544.950 415.050 545.400 ;
        RECT 739.950 546.600 742.050 547.050 ;
        RECT 748.950 546.600 751.050 547.050 ;
        RECT 754.950 546.600 757.050 547.050 ;
        RECT 739.950 545.400 757.050 546.600 ;
        RECT 739.950 544.950 742.050 545.400 ;
        RECT 748.950 544.950 751.050 545.400 ;
        RECT 754.950 544.950 757.050 545.400 ;
        RECT 829.950 546.600 832.050 547.050 ;
        RECT 844.950 546.600 847.050 547.050 ;
        RECT 829.950 545.400 847.050 546.600 ;
        RECT 829.950 544.950 832.050 545.400 ;
        RECT 844.950 544.950 847.050 545.400 ;
        RECT 985.950 546.600 988.050 547.050 ;
        RECT 1015.950 546.600 1018.050 547.050 ;
        RECT 985.950 545.400 1018.050 546.600 ;
        RECT 985.950 544.950 988.050 545.400 ;
        RECT 1015.950 544.950 1018.050 545.400 ;
        RECT 358.950 543.600 361.050 544.050 ;
        RECT 373.950 543.600 376.050 544.050 ;
        RECT 358.950 542.400 376.050 543.600 ;
        RECT 358.950 541.950 361.050 542.400 ;
        RECT 373.950 541.950 376.050 542.400 ;
        RECT 502.950 543.600 505.050 544.050 ;
        RECT 514.950 543.600 517.050 544.050 ;
        RECT 502.950 542.400 517.050 543.600 ;
        RECT 502.950 541.950 505.050 542.400 ;
        RECT 514.950 541.950 517.050 542.400 ;
        RECT 535.950 543.600 538.050 544.050 ;
        RECT 559.950 543.600 562.050 544.050 ;
        RECT 535.950 542.400 562.050 543.600 ;
        RECT 535.950 541.950 538.050 542.400 ;
        RECT 559.950 541.950 562.050 542.400 ;
        RECT 730.950 543.600 733.050 544.050 ;
        RECT 736.950 543.600 739.050 544.050 ;
        RECT 730.950 542.400 739.050 543.600 ;
        RECT 730.950 541.950 733.050 542.400 ;
        RECT 736.950 541.950 739.050 542.400 ;
        RECT 784.950 543.600 787.050 544.050 ;
        RECT 928.950 543.600 931.050 544.050 ;
        RECT 940.950 543.600 943.050 544.050 ;
        RECT 784.950 542.400 888.600 543.600 ;
        RECT 784.950 541.950 787.050 542.400 ;
        RECT 887.400 541.050 888.600 542.400 ;
        RECT 928.950 542.400 943.050 543.600 ;
        RECT 928.950 541.950 931.050 542.400 ;
        RECT 940.950 541.950 943.050 542.400 ;
        RECT 187.950 540.600 190.050 541.050 ;
        RECT 223.950 540.600 226.050 541.050 ;
        RECT 187.950 539.400 226.050 540.600 ;
        RECT 187.950 538.950 190.050 539.400 ;
        RECT 223.950 538.950 226.050 539.400 ;
        RECT 364.950 540.600 367.050 541.050 ;
        RECT 433.950 540.600 436.050 541.050 ;
        RECT 517.950 540.600 520.050 541.050 ;
        RECT 562.950 540.600 565.050 541.050 ;
        RECT 364.950 539.400 436.050 540.600 ;
        RECT 364.950 538.950 367.050 539.400 ;
        RECT 433.950 538.950 436.050 539.400 ;
        RECT 455.400 539.400 565.050 540.600 ;
        RECT 169.950 537.600 172.050 538.050 ;
        RECT 196.950 537.600 199.050 538.050 ;
        RECT 169.950 536.400 199.050 537.600 ;
        RECT 169.950 535.950 172.050 536.400 ;
        RECT 196.950 535.950 199.050 536.400 ;
        RECT 259.950 537.600 262.050 538.050 ;
        RECT 455.400 537.600 456.600 539.400 ;
        RECT 517.950 538.950 520.050 539.400 ;
        RECT 562.950 538.950 565.050 539.400 ;
        RECT 604.950 540.600 607.050 541.050 ;
        RECT 631.950 540.600 634.050 541.050 ;
        RECT 604.950 539.400 634.050 540.600 ;
        RECT 604.950 538.950 607.050 539.400 ;
        RECT 631.950 538.950 634.050 539.400 ;
        RECT 685.950 540.600 688.050 541.050 ;
        RECT 712.950 540.600 715.050 541.050 ;
        RECT 685.950 539.400 715.050 540.600 ;
        RECT 685.950 538.950 688.050 539.400 ;
        RECT 712.950 538.950 715.050 539.400 ;
        RECT 724.950 540.600 727.050 541.050 ;
        RECT 754.950 540.600 757.050 541.050 ;
        RECT 724.950 539.400 757.050 540.600 ;
        RECT 724.950 538.950 727.050 539.400 ;
        RECT 754.950 538.950 757.050 539.400 ;
        RECT 799.950 540.600 802.050 541.050 ;
        RECT 832.950 540.600 835.050 541.050 ;
        RECT 799.950 539.400 835.050 540.600 ;
        RECT 887.400 539.400 892.050 541.050 ;
        RECT 799.950 538.950 802.050 539.400 ;
        RECT 832.950 538.950 835.050 539.400 ;
        RECT 888.000 538.950 892.050 539.400 ;
        RECT 907.950 540.600 910.050 541.050 ;
        RECT 913.950 540.600 916.050 541.050 ;
        RECT 907.950 539.400 916.050 540.600 ;
        RECT 907.950 538.950 910.050 539.400 ;
        RECT 913.950 538.950 916.050 539.400 ;
        RECT 259.950 536.400 456.600 537.600 ;
        RECT 508.950 537.600 511.050 538.050 ;
        RECT 520.950 537.600 523.050 538.050 ;
        RECT 508.950 536.400 523.050 537.600 ;
        RECT 259.950 535.950 262.050 536.400 ;
        RECT 508.950 535.950 511.050 536.400 ;
        RECT 520.950 535.950 523.050 536.400 ;
        RECT 682.950 537.600 685.050 538.050 ;
        RECT 703.950 537.600 706.050 538.050 ;
        RECT 682.950 536.400 706.050 537.600 ;
        RECT 682.950 535.950 685.050 536.400 ;
        RECT 703.950 535.950 706.050 536.400 ;
        RECT 757.950 537.600 760.050 538.050 ;
        RECT 787.950 537.600 790.050 538.050 ;
        RECT 943.950 537.600 946.050 538.050 ;
        RECT 757.950 536.400 790.050 537.600 ;
        RECT 757.950 535.950 760.050 536.400 ;
        RECT 787.950 535.950 790.050 536.400 ;
        RECT 917.400 536.400 946.050 537.600 ;
        RECT 37.950 534.600 40.050 535.050 ;
        RECT 58.950 534.600 61.050 535.050 ;
        RECT 67.950 534.600 70.050 535.050 ;
        RECT 37.950 533.400 70.050 534.600 ;
        RECT 37.950 532.950 40.050 533.400 ;
        RECT 58.950 532.950 61.050 533.400 ;
        RECT 67.950 532.950 70.050 533.400 ;
        RECT 85.950 534.600 88.050 535.050 ;
        RECT 415.950 534.600 418.050 535.050 ;
        RECT 427.950 534.600 430.050 535.050 ;
        RECT 85.950 533.400 219.600 534.600 ;
        RECT 85.950 532.950 88.050 533.400 ;
        RECT 218.400 532.050 219.600 533.400 ;
        RECT 415.950 533.400 430.050 534.600 ;
        RECT 415.950 532.950 418.050 533.400 ;
        RECT 427.950 532.950 430.050 533.400 ;
        RECT 433.950 534.600 436.050 535.050 ;
        RECT 484.950 534.600 487.050 535.050 ;
        RECT 526.950 534.600 529.050 535.050 ;
        RECT 433.950 533.400 529.050 534.600 ;
        RECT 433.950 532.950 436.050 533.400 ;
        RECT 484.950 532.950 487.050 533.400 ;
        RECT 526.950 532.950 529.050 533.400 ;
        RECT 568.950 534.600 571.050 535.050 ;
        RECT 598.950 534.600 601.050 535.050 ;
        RECT 568.950 533.400 601.050 534.600 ;
        RECT 568.950 532.950 571.050 533.400 ;
        RECT 598.950 532.950 601.050 533.400 ;
        RECT 613.950 534.600 616.050 535.050 ;
        RECT 763.950 534.600 766.050 535.050 ;
        RECT 799.950 534.600 802.050 535.050 ;
        RECT 613.950 533.400 696.600 534.600 ;
        RECT 613.950 532.950 616.050 533.400 ;
        RECT 695.400 532.050 696.600 533.400 ;
        RECT 763.950 533.400 802.050 534.600 ;
        RECT 763.950 532.950 766.050 533.400 ;
        RECT 799.950 532.950 802.050 533.400 ;
        RECT 805.950 534.600 808.050 535.050 ;
        RECT 868.950 534.600 871.050 535.050 ;
        RECT 805.950 533.400 871.050 534.600 ;
        RECT 805.950 532.950 808.050 533.400 ;
        RECT 868.950 532.950 871.050 533.400 ;
        RECT 874.950 534.600 877.050 535.050 ;
        RECT 917.400 534.600 918.600 536.400 ;
        RECT 943.950 535.950 946.050 536.400 ;
        RECT 874.950 533.400 918.600 534.600 ;
        RECT 940.950 534.600 943.050 535.050 ;
        RECT 958.950 534.600 961.050 535.050 ;
        RECT 940.950 533.400 961.050 534.600 ;
        RECT 874.950 532.950 877.050 533.400 ;
        RECT 940.950 532.950 943.050 533.400 ;
        RECT 958.950 532.950 961.050 533.400 ;
        RECT 964.950 534.600 967.050 535.050 ;
        RECT 991.950 534.600 994.050 535.050 ;
        RECT 964.950 533.400 994.050 534.600 ;
        RECT 964.950 532.950 967.050 533.400 ;
        RECT 991.950 532.950 994.050 533.400 ;
        RECT 1003.950 534.600 1006.050 535.050 ;
        RECT 1015.950 534.600 1018.050 535.050 ;
        RECT 1003.950 533.400 1018.050 534.600 ;
        RECT 1003.950 532.950 1006.050 533.400 ;
        RECT 1015.950 532.950 1018.050 533.400 ;
        RECT 217.950 531.600 220.050 532.050 ;
        RECT 229.950 531.600 232.050 532.050 ;
        RECT 217.950 530.400 232.050 531.600 ;
        RECT 217.950 529.950 220.050 530.400 ;
        RECT 229.950 529.950 232.050 530.400 ;
        RECT 430.950 531.600 433.050 532.050 ;
        RECT 436.950 531.600 439.050 532.050 ;
        RECT 430.950 530.400 439.050 531.600 ;
        RECT 430.950 529.950 433.050 530.400 ;
        RECT 436.950 529.950 439.050 530.400 ;
        RECT 598.950 531.600 601.050 531.900 ;
        RECT 610.950 531.600 613.050 532.050 ;
        RECT 598.950 530.400 613.050 531.600 ;
        RECT 695.400 531.600 700.050 532.050 ;
        RECT 727.950 531.600 730.050 532.050 ;
        RECT 739.950 531.600 742.050 532.050 ;
        RECT 695.400 530.400 742.050 531.600 ;
        RECT 598.950 529.800 601.050 530.400 ;
        RECT 610.950 529.950 613.050 530.400 ;
        RECT 696.000 529.950 700.050 530.400 ;
        RECT 727.950 529.950 730.050 530.400 ;
        RECT 739.950 529.950 742.050 530.400 ;
        RECT 769.950 531.600 772.050 532.050 ;
        RECT 778.950 531.600 781.050 532.050 ;
        RECT 769.950 530.400 781.050 531.600 ;
        RECT 769.950 529.950 772.050 530.400 ;
        RECT 778.950 529.950 781.050 530.400 ;
        RECT 886.950 531.600 891.000 532.050 ;
        RECT 886.950 529.950 891.600 531.600 ;
        RECT 892.950 529.950 895.050 532.050 ;
        RECT 976.950 531.600 979.050 532.050 ;
        RECT 985.950 531.600 988.050 532.050 ;
        RECT 976.950 530.400 988.050 531.600 ;
        RECT 976.950 529.950 979.050 530.400 ;
        RECT 985.950 529.950 988.050 530.400 ;
        RECT 52.950 528.600 55.050 529.200 ;
        RECT 50.400 527.400 55.050 528.600 ;
        RECT 50.400 523.050 51.600 527.400 ;
        RECT 52.950 527.100 55.050 527.400 ;
        RECT 58.950 527.100 61.050 529.200 ;
        RECT 64.950 528.750 67.050 529.200 ;
        RECT 73.950 528.750 76.050 529.200 ;
        RECT 64.950 527.550 76.050 528.750 ;
        RECT 64.950 527.100 67.050 527.550 ;
        RECT 73.950 527.100 76.050 527.550 ;
        RECT 79.950 528.750 82.050 529.200 ;
        RECT 85.950 528.750 88.050 529.200 ;
        RECT 79.950 527.550 88.050 528.750 ;
        RECT 79.950 527.100 82.050 527.550 ;
        RECT 85.950 527.100 88.050 527.550 ;
        RECT 91.950 528.750 94.050 529.200 ;
        RECT 100.950 528.750 103.050 529.200 ;
        RECT 91.950 527.550 103.050 528.750 ;
        RECT 91.950 527.100 94.050 527.550 ;
        RECT 100.950 527.100 103.050 527.550 ;
        RECT 106.950 528.750 109.050 529.200 ;
        RECT 115.950 528.750 118.050 529.200 ;
        RECT 106.950 527.550 118.050 528.750 ;
        RECT 106.950 527.100 109.050 527.550 ;
        RECT 115.950 527.100 118.050 527.550 ;
        RECT 130.950 527.100 133.050 529.200 ;
        RECT 151.950 528.600 154.050 529.200 ;
        RECT 157.950 528.600 160.050 529.050 ;
        RECT 151.950 527.400 160.050 528.600 ;
        RECT 151.950 527.100 154.050 527.400 ;
        RECT 59.400 525.600 60.600 527.100 ;
        RECT 131.400 525.600 132.600 527.100 ;
        RECT 157.950 526.950 160.050 527.400 ;
        RECT 163.950 528.600 166.050 529.050 ;
        RECT 169.950 528.600 172.050 529.200 ;
        RECT 163.950 527.400 172.050 528.600 ;
        RECT 163.950 526.950 166.050 527.400 ;
        RECT 169.950 527.100 172.050 527.400 ;
        RECT 175.950 527.100 178.050 529.200 ;
        RECT 181.950 527.100 184.050 529.200 ;
        RECT 190.950 528.600 193.050 529.200 ;
        RECT 241.950 528.750 244.050 529.200 ;
        RECT 253.950 528.750 256.050 529.200 ;
        RECT 190.950 527.400 195.600 528.600 ;
        RECT 190.950 527.100 193.050 527.400 ;
        RECT 160.950 525.600 163.050 525.900 ;
        RECT 59.400 524.400 81.600 525.600 ;
        RECT 131.400 524.400 163.050 525.600 ;
        RECT 19.950 522.600 22.050 522.900 ;
        RECT 43.950 522.600 46.050 523.050 ;
        RECT 19.950 521.400 46.050 522.600 ;
        RECT 19.950 520.800 22.050 521.400 ;
        RECT 43.950 520.950 46.050 521.400 ;
        RECT 49.950 520.950 52.050 523.050 ;
        RECT 55.950 522.600 58.050 522.900 ;
        RECT 55.950 522.000 63.600 522.600 ;
        RECT 64.950 522.450 67.050 522.900 ;
        RECT 76.950 522.450 79.050 522.900 ;
        RECT 55.950 521.400 64.050 522.000 ;
        RECT 55.950 520.800 58.050 521.400 ;
        RECT 61.950 517.950 64.050 521.400 ;
        RECT 64.950 521.250 79.050 522.450 ;
        RECT 80.400 522.600 81.600 524.400 ;
        RECT 160.950 523.800 163.050 524.400 ;
        RECT 82.950 522.600 85.050 522.900 ;
        RECT 80.400 521.400 85.050 522.600 ;
        RECT 64.950 520.800 67.050 521.250 ;
        RECT 76.950 520.800 79.050 521.250 ;
        RECT 82.950 520.800 85.050 521.400 ;
        RECT 88.950 522.600 91.050 523.050 ;
        RECT 103.950 522.600 106.050 522.900 ;
        RECT 88.950 521.400 106.050 522.600 ;
        RECT 88.950 520.950 91.050 521.400 ;
        RECT 103.950 520.800 106.050 521.400 ;
        RECT 115.950 522.600 118.050 523.050 ;
        RECT 127.950 522.600 130.050 522.900 ;
        RECT 115.950 521.400 130.050 522.600 ;
        RECT 115.950 520.950 118.050 521.400 ;
        RECT 127.950 520.800 130.050 521.400 ;
        RECT 142.950 522.600 145.050 523.050 ;
        RECT 166.950 522.600 169.050 522.900 ;
        RECT 142.950 521.400 169.050 522.600 ;
        RECT 142.950 520.950 145.050 521.400 ;
        RECT 166.950 520.800 169.050 521.400 ;
        RECT 176.400 519.600 177.600 527.100 ;
        RECT 182.400 523.050 183.600 527.100 ;
        RECT 194.400 523.050 195.600 527.400 ;
        RECT 241.950 527.550 256.050 528.750 ;
        RECT 241.950 527.100 244.050 527.550 ;
        RECT 253.950 527.100 256.050 527.550 ;
        RECT 277.950 528.600 280.050 529.200 ;
        RECT 298.950 528.600 301.050 529.200 ;
        RECT 277.950 527.400 301.050 528.600 ;
        RECT 277.950 527.100 280.050 527.400 ;
        RECT 298.950 527.100 301.050 527.400 ;
        RECT 325.950 528.750 328.050 529.200 ;
        RECT 358.950 528.750 361.050 529.200 ;
        RECT 325.950 528.600 361.050 528.750 ;
        RECT 382.950 528.600 385.050 529.200 ;
        RECT 325.950 527.550 385.050 528.600 ;
        RECT 325.950 527.100 328.050 527.550 ;
        RECT 358.950 527.400 385.050 527.550 ;
        RECT 358.950 527.100 361.050 527.400 ;
        RECT 382.950 527.100 385.050 527.400 ;
        RECT 388.950 528.600 391.050 529.200 ;
        RECT 397.950 528.600 400.050 529.050 ;
        RECT 403.950 528.600 406.050 529.200 ;
        RECT 388.950 527.400 406.050 528.600 ;
        RECT 388.950 527.100 391.050 527.400 ;
        RECT 383.400 525.600 384.600 527.100 ;
        RECT 397.950 526.950 400.050 527.400 ;
        RECT 403.950 527.100 406.050 527.400 ;
        RECT 424.950 527.100 427.050 529.200 ;
        RECT 454.950 528.600 457.050 529.200 ;
        RECT 440.400 527.400 457.050 528.600 ;
        RECT 394.950 525.600 397.050 526.050 ;
        RECT 383.400 524.400 397.050 525.600 ;
        RECT 394.950 523.950 397.050 524.400 ;
        RECT 178.950 521.400 183.600 523.050 ;
        RECT 178.950 520.950 183.000 521.400 ;
        RECT 193.950 520.950 196.050 523.050 ;
        RECT 244.950 522.600 247.050 523.050 ;
        RECT 256.950 522.600 259.050 522.900 ;
        RECT 244.950 521.400 259.050 522.600 ;
        RECT 244.950 520.950 247.050 521.400 ;
        RECT 256.950 520.800 259.050 521.400 ;
        RECT 274.950 522.450 277.050 522.900 ;
        RECT 289.950 522.450 292.050 522.900 ;
        RECT 274.950 521.250 292.050 522.450 ;
        RECT 274.950 520.800 277.050 521.250 ;
        RECT 289.950 520.800 292.050 521.250 ;
        RECT 415.950 522.600 418.050 523.050 ;
        RECT 421.950 522.600 424.050 522.900 ;
        RECT 415.950 521.400 424.050 522.600 ;
        RECT 415.950 520.950 418.050 521.400 ;
        RECT 421.950 520.800 424.050 521.400 ;
        RECT 425.400 520.050 426.600 527.100 ;
        RECT 440.400 525.600 441.600 527.400 ;
        RECT 454.950 527.100 457.050 527.400 ;
        RECT 463.950 528.600 466.050 529.200 ;
        RECT 469.950 528.600 472.050 529.050 ;
        RECT 463.950 527.400 472.050 528.600 ;
        RECT 463.950 527.100 466.050 527.400 ;
        RECT 469.950 526.950 472.050 527.400 ;
        RECT 490.950 528.750 493.050 529.200 ;
        RECT 496.950 528.750 499.050 529.200 ;
        RECT 490.950 527.550 499.050 528.750 ;
        RECT 490.950 527.100 493.050 527.550 ;
        RECT 496.950 527.100 499.050 527.550 ;
        RECT 505.950 527.100 508.050 529.200 ;
        RECT 428.400 524.400 441.600 525.600 ;
        RECT 428.400 522.900 429.600 524.400 ;
        RECT 427.950 520.800 430.050 522.900 ;
        RECT 481.950 522.600 484.050 522.900 ;
        RECT 506.400 522.600 507.600 527.100 ;
        RECT 523.950 526.950 526.050 529.050 ;
        RECT 547.950 528.600 550.050 529.050 ;
        RECT 553.950 528.600 556.050 529.200 ;
        RECT 547.950 527.400 556.050 528.600 ;
        RECT 547.950 526.950 550.050 527.400 ;
        RECT 553.950 527.100 556.050 527.400 ;
        RECT 625.950 528.750 628.050 529.200 ;
        RECT 631.950 528.750 634.050 529.200 ;
        RECT 625.950 527.550 634.050 528.750 ;
        RECT 625.950 527.100 628.050 527.550 ;
        RECT 631.950 527.100 634.050 527.550 ;
        RECT 643.950 527.100 646.050 529.200 ;
        RECT 649.950 527.100 652.050 529.200 ;
        RECT 673.950 528.750 676.050 529.200 ;
        RECT 685.950 528.750 688.050 529.200 ;
        RECT 673.950 527.550 688.050 528.750 ;
        RECT 673.950 527.100 676.050 527.550 ;
        RECT 685.950 527.100 688.050 527.550 ;
        RECT 481.950 521.400 507.600 522.600 ;
        RECT 514.950 522.600 517.050 523.050 ;
        RECT 524.400 522.600 525.600 526.950 ;
        RECT 514.950 521.400 525.600 522.600 ;
        RECT 583.950 522.600 586.050 522.900 ;
        RECT 589.950 522.600 592.050 523.050 ;
        RECT 583.950 521.400 592.050 522.600 ;
        RECT 481.950 520.800 484.050 521.400 ;
        RECT 514.950 520.950 517.050 521.400 ;
        RECT 583.950 520.800 586.050 521.400 ;
        RECT 589.950 520.950 592.050 521.400 ;
        RECT 613.950 522.600 616.050 523.050 ;
        RECT 622.950 522.600 625.050 522.900 ;
        RECT 613.950 521.400 625.050 522.600 ;
        RECT 613.950 520.950 616.050 521.400 ;
        RECT 622.950 520.800 625.050 521.400 ;
        RECT 631.950 522.600 634.050 523.050 ;
        RECT 640.950 522.600 643.050 523.050 ;
        RECT 631.950 521.400 643.050 522.600 ;
        RECT 631.950 520.950 634.050 521.400 ;
        RECT 640.950 520.950 643.050 521.400 ;
        RECT 644.400 520.050 645.600 527.100 ;
        RECT 650.400 522.600 651.600 527.100 ;
        RECT 718.950 526.950 721.050 529.050 ;
        RECT 760.950 528.750 763.050 529.200 ;
        RECT 769.950 528.750 772.050 529.200 ;
        RECT 760.950 527.550 772.050 528.750 ;
        RECT 760.950 527.100 763.050 527.550 ;
        RECT 769.950 527.100 772.050 527.550 ;
        RECT 787.950 528.600 792.000 529.050 ;
        RECT 787.950 526.950 792.600 528.600 ;
        RECT 799.950 527.100 802.050 529.200 ;
        RECT 808.950 528.750 811.050 529.200 ;
        RECT 820.950 528.750 823.050 529.200 ;
        RECT 808.950 527.550 823.050 528.750 ;
        RECT 808.950 527.100 811.050 527.550 ;
        RECT 820.950 527.100 823.050 527.550 ;
        RECT 844.950 527.100 847.050 529.200 ;
        RECT 719.400 523.050 720.600 526.950 ;
        RECT 655.950 522.600 658.050 523.050 ;
        RECT 650.400 521.400 658.050 522.600 ;
        RECT 655.950 520.950 658.050 521.400 ;
        RECT 661.950 522.600 664.050 523.050 ;
        RECT 667.950 522.600 670.050 523.050 ;
        RECT 661.950 521.400 670.050 522.600 ;
        RECT 661.950 520.950 664.050 521.400 ;
        RECT 667.950 520.950 670.050 521.400 ;
        RECT 676.950 522.600 679.050 522.900 ;
        RECT 700.950 522.600 703.050 522.900 ;
        RECT 676.950 521.400 703.050 522.600 ;
        RECT 676.950 520.800 679.050 521.400 ;
        RECT 700.950 520.800 703.050 521.400 ;
        RECT 718.950 520.950 721.050 523.050 ;
        RECT 739.950 522.450 742.050 522.900 ;
        RECT 745.950 522.450 748.050 522.900 ;
        RECT 739.950 521.250 748.050 522.450 ;
        RECT 739.950 520.800 742.050 521.250 ;
        RECT 745.950 520.800 748.050 521.250 ;
        RECT 772.950 522.600 775.050 522.900 ;
        RECT 784.950 522.600 787.050 523.050 ;
        RECT 791.400 522.900 792.600 526.950 ;
        RECT 772.950 521.400 787.050 522.600 ;
        RECT 772.950 520.800 775.050 521.400 ;
        RECT 784.950 520.950 787.050 521.400 ;
        RECT 790.950 520.800 793.050 522.900 ;
        RECT 199.950 519.600 202.050 520.050 ;
        RECT 176.400 518.400 202.050 519.600 ;
        RECT 199.950 517.950 202.050 518.400 ;
        RECT 406.950 519.600 409.050 520.050 ;
        RECT 412.950 519.600 415.050 520.050 ;
        RECT 406.950 518.400 415.050 519.600 ;
        RECT 406.950 517.950 409.050 518.400 ;
        RECT 412.950 517.950 415.050 518.400 ;
        RECT 424.950 517.950 427.050 520.050 ;
        RECT 643.950 517.950 646.050 520.050 ;
        RECT 700.950 519.600 703.050 520.050 ;
        RECT 712.950 519.600 715.050 520.050 ;
        RECT 700.950 518.400 715.050 519.600 ;
        RECT 700.950 517.950 703.050 518.400 ;
        RECT 712.950 517.950 715.050 518.400 ;
        RECT 730.950 519.600 733.050 520.050 ;
        RECT 760.950 519.600 763.050 520.050 ;
        RECT 730.950 518.400 763.050 519.600 ;
        RECT 730.950 517.950 733.050 518.400 ;
        RECT 760.950 517.950 763.050 518.400 ;
        RECT 793.950 519.600 796.050 520.050 ;
        RECT 800.400 519.600 801.600 527.100 ;
        RECT 817.950 522.600 820.050 522.900 ;
        RECT 841.950 522.600 844.050 522.900 ;
        RECT 817.950 521.400 844.050 522.600 ;
        RECT 817.950 520.800 820.050 521.400 ;
        RECT 841.950 520.800 844.050 521.400 ;
        RECT 845.400 519.600 846.600 527.100 ;
        RECT 850.950 526.950 853.050 529.050 ;
        RECT 856.950 528.750 859.050 529.200 ;
        RECT 862.950 528.750 865.050 529.200 ;
        RECT 856.950 527.550 865.050 528.750 ;
        RECT 856.950 527.100 859.050 527.550 ;
        RECT 862.950 527.100 865.050 527.550 ;
        RECT 851.400 523.050 852.600 526.950 ;
        RECT 890.400 525.600 891.600 529.950 ;
        RECT 887.400 524.400 891.600 525.600 ;
        RECT 850.950 520.950 853.050 523.050 ;
        RECT 874.950 522.600 877.050 523.050 ;
        RECT 880.950 522.600 883.050 523.050 ;
        RECT 887.400 522.900 888.600 524.400 ;
        RECT 893.400 522.900 894.600 529.950 ;
        RECT 895.950 528.750 898.050 529.200 ;
        RECT 901.950 528.750 904.050 529.200 ;
        RECT 895.950 527.550 904.050 528.750 ;
        RECT 895.950 527.100 898.050 527.550 ;
        RECT 901.950 527.100 904.050 527.550 ;
        RECT 919.950 528.750 922.050 529.200 ;
        RECT 931.950 528.750 934.050 529.200 ;
        RECT 919.950 527.550 934.050 528.750 ;
        RECT 942.000 528.600 946.050 529.050 ;
        RECT 919.950 527.100 922.050 527.550 ;
        RECT 931.950 527.100 934.050 527.550 ;
        RECT 941.400 526.950 946.050 528.600 ;
        RECT 952.950 526.950 955.050 529.050 ;
        RECT 941.400 523.050 942.600 526.950 ;
        RECT 874.950 521.400 883.050 522.600 ;
        RECT 874.950 520.950 877.050 521.400 ;
        RECT 880.950 520.950 883.050 521.400 ;
        RECT 886.950 520.800 889.050 522.900 ;
        RECT 892.950 520.800 895.050 522.900 ;
        RECT 916.950 522.450 919.050 522.900 ;
        RECT 925.950 522.450 928.050 522.900 ;
        RECT 916.950 521.250 928.050 522.450 ;
        RECT 941.400 521.400 946.050 523.050 ;
        RECT 916.950 520.800 919.050 521.250 ;
        RECT 925.950 520.800 928.050 521.250 ;
        RECT 942.000 520.950 946.050 521.400 ;
        RECT 953.400 520.050 954.600 526.950 ;
        RECT 967.950 525.600 970.050 529.050 ;
        RECT 997.950 528.600 1002.000 529.050 ;
        RECT 997.950 526.950 1002.600 528.600 ;
        RECT 1009.800 527.100 1011.900 529.200 ;
        RECT 1012.950 528.600 1017.000 529.050 ;
        RECT 1001.400 525.600 1002.600 526.950 ;
        RECT 967.950 525.000 999.600 525.600 ;
        RECT 968.400 524.400 999.600 525.000 ;
        RECT 1001.400 524.400 1008.600 525.600 ;
        RECT 985.950 522.600 988.050 522.900 ;
        RECT 994.950 522.600 997.050 523.050 ;
        RECT 985.950 521.400 997.050 522.600 ;
        RECT 998.400 522.600 999.600 524.400 ;
        RECT 1007.400 522.900 1008.600 524.400 ;
        RECT 998.400 521.400 1002.600 522.600 ;
        RECT 985.950 520.800 988.050 521.400 ;
        RECT 994.950 520.950 997.050 521.400 ;
        RECT 1001.400 520.050 1002.600 521.400 ;
        RECT 1006.950 520.800 1009.050 522.900 ;
        RECT 1010.250 520.050 1011.450 527.100 ;
        RECT 1012.950 526.950 1017.600 528.600 ;
        RECT 1016.400 520.050 1017.600 526.950 ;
        RECT 892.950 519.600 895.050 520.050 ;
        RECT 793.950 518.400 846.600 519.600 ;
        RECT 878.400 518.400 895.050 519.600 ;
        RECT 953.400 518.400 958.050 520.050 ;
        RECT 793.950 517.950 796.050 518.400 ;
        RECT 43.950 516.600 46.050 517.050 ;
        RECT 64.800 516.600 66.900 517.050 ;
        RECT 43.950 515.400 66.900 516.600 ;
        RECT 43.950 514.950 46.050 515.400 ;
        RECT 64.800 514.950 66.900 515.400 ;
        RECT 67.950 516.600 70.050 517.050 ;
        RECT 97.950 516.600 100.050 517.050 ;
        RECT 67.950 515.400 100.050 516.600 ;
        RECT 67.950 514.950 70.050 515.400 ;
        RECT 97.950 514.950 100.050 515.400 ;
        RECT 148.950 516.600 151.050 517.050 ;
        RECT 229.950 516.600 232.050 517.050 ;
        RECT 259.950 516.600 262.050 517.050 ;
        RECT 265.950 516.600 268.050 517.050 ;
        RECT 325.950 516.600 328.050 517.050 ;
        RECT 148.950 515.400 328.050 516.600 ;
        RECT 148.950 514.950 151.050 515.400 ;
        RECT 229.950 514.950 232.050 515.400 ;
        RECT 259.950 514.950 262.050 515.400 ;
        RECT 265.950 514.950 268.050 515.400 ;
        RECT 325.950 514.950 328.050 515.400 ;
        RECT 394.950 516.600 397.050 517.050 ;
        RECT 430.950 516.600 433.050 517.050 ;
        RECT 448.950 516.600 451.050 517.050 ;
        RECT 394.950 515.400 451.050 516.600 ;
        RECT 394.950 514.950 397.050 515.400 ;
        RECT 430.950 514.950 433.050 515.400 ;
        RECT 448.950 514.950 451.050 515.400 ;
        RECT 481.950 516.600 484.050 517.050 ;
        RECT 499.950 516.600 502.050 517.050 ;
        RECT 481.950 515.400 502.050 516.600 ;
        RECT 481.950 514.950 484.050 515.400 ;
        RECT 499.950 514.950 502.050 515.400 ;
        RECT 508.950 516.600 511.050 517.050 ;
        RECT 520.950 516.600 523.050 517.050 ;
        RECT 571.950 516.600 574.050 517.050 ;
        RECT 508.950 515.400 523.050 516.600 ;
        RECT 508.950 514.950 511.050 515.400 ;
        RECT 520.950 514.950 523.050 515.400 ;
        RECT 551.400 515.400 574.050 516.600 ;
        RECT 49.950 513.600 52.050 514.050 ;
        RECT 58.950 513.600 61.050 514.050 ;
        RECT 49.950 512.400 61.050 513.600 ;
        RECT 49.950 511.950 52.050 512.400 ;
        RECT 58.950 511.950 61.050 512.400 ;
        RECT 79.950 513.600 82.050 514.050 ;
        RECT 91.950 513.600 94.050 514.050 ;
        RECT 79.950 512.400 94.050 513.600 ;
        RECT 79.950 511.950 82.050 512.400 ;
        RECT 91.950 511.950 94.050 512.400 ;
        RECT 337.950 513.600 340.050 514.050 ;
        RECT 361.950 513.600 364.050 514.050 ;
        RECT 337.950 512.400 364.050 513.600 ;
        RECT 337.950 511.950 340.050 512.400 ;
        RECT 361.950 511.950 364.050 512.400 ;
        RECT 397.950 513.600 400.050 514.050 ;
        RECT 424.950 513.600 427.050 514.050 ;
        RECT 397.950 512.400 427.050 513.600 ;
        RECT 397.950 511.950 400.050 512.400 ;
        RECT 424.950 511.950 427.050 512.400 ;
        RECT 535.950 513.600 538.050 514.050 ;
        RECT 551.400 513.600 552.600 515.400 ;
        RECT 571.950 514.950 574.050 515.400 ;
        RECT 742.950 516.600 745.050 517.050 ;
        RECT 754.950 516.600 757.050 517.050 ;
        RECT 742.950 515.400 757.050 516.600 ;
        RECT 742.950 514.950 745.050 515.400 ;
        RECT 754.950 514.950 757.050 515.400 ;
        RECT 796.950 516.600 799.050 517.050 ;
        RECT 805.950 516.600 808.050 517.050 ;
        RECT 796.950 515.400 808.050 516.600 ;
        RECT 796.950 514.950 799.050 515.400 ;
        RECT 805.950 514.950 808.050 515.400 ;
        RECT 868.950 516.600 871.050 517.050 ;
        RECT 878.400 516.600 879.600 518.400 ;
        RECT 892.950 517.950 895.050 518.400 ;
        RECT 954.000 517.950 958.050 518.400 ;
        RECT 970.950 519.600 973.050 520.050 ;
        RECT 997.950 519.600 1000.050 520.050 ;
        RECT 970.950 518.400 1000.050 519.600 ;
        RECT 1001.400 518.400 1006.050 520.050 ;
        RECT 970.950 517.950 973.050 518.400 ;
        RECT 997.950 517.950 1000.050 518.400 ;
        RECT 1002.000 517.950 1006.050 518.400 ;
        RECT 1009.800 517.950 1011.900 520.050 ;
        RECT 1015.950 517.950 1018.050 520.050 ;
        RECT 868.950 515.400 879.600 516.600 ;
        RECT 868.950 514.950 871.050 515.400 ;
        RECT 535.950 512.400 552.600 513.600 ;
        RECT 592.950 513.600 595.050 514.050 ;
        RECT 622.950 513.600 625.050 514.050 ;
        RECT 637.950 513.600 640.050 514.050 ;
        RECT 592.950 512.400 640.050 513.600 ;
        RECT 535.950 511.950 538.050 512.400 ;
        RECT 592.950 511.950 595.050 512.400 ;
        RECT 622.950 511.950 625.050 512.400 ;
        RECT 637.950 511.950 640.050 512.400 ;
        RECT 706.950 513.600 709.050 514.050 ;
        RECT 817.950 513.600 820.050 514.050 ;
        RECT 706.950 512.400 820.050 513.600 ;
        RECT 706.950 511.950 709.050 512.400 ;
        RECT 817.950 511.950 820.050 512.400 ;
        RECT 823.950 513.600 826.050 514.050 ;
        RECT 865.950 513.600 868.050 514.050 ;
        RECT 823.950 512.400 868.050 513.600 ;
        RECT 823.950 511.950 826.050 512.400 ;
        RECT 865.950 511.950 868.050 512.400 ;
        RECT 880.950 513.600 883.050 514.050 ;
        RECT 901.950 513.600 904.050 514.050 ;
        RECT 880.950 512.400 904.050 513.600 ;
        RECT 880.950 511.950 883.050 512.400 ;
        RECT 901.950 511.950 904.050 512.400 ;
        RECT 907.950 513.600 910.050 514.050 ;
        RECT 949.950 513.600 952.050 514.050 ;
        RECT 907.950 512.400 952.050 513.600 ;
        RECT 907.950 511.950 910.050 512.400 ;
        RECT 949.950 511.950 952.050 512.400 ;
        RECT 82.950 510.600 85.050 511.050 ;
        RECT 133.950 510.600 136.050 511.050 ;
        RECT 82.950 509.400 136.050 510.600 ;
        RECT 82.950 508.950 85.050 509.400 ;
        RECT 133.950 508.950 136.050 509.400 ;
        RECT 301.950 510.600 304.050 511.050 ;
        RECT 307.950 510.600 310.050 511.050 ;
        RECT 319.950 510.600 322.050 511.050 ;
        RECT 301.950 509.400 322.050 510.600 ;
        RECT 301.950 508.950 304.050 509.400 ;
        RECT 307.950 508.950 310.050 509.400 ;
        RECT 319.950 508.950 322.050 509.400 ;
        RECT 487.950 510.600 490.050 511.050 ;
        RECT 547.950 510.600 550.050 511.050 ;
        RECT 487.950 509.400 550.050 510.600 ;
        RECT 487.950 508.950 490.050 509.400 ;
        RECT 547.950 508.950 550.050 509.400 ;
        RECT 559.950 510.600 562.050 511.050 ;
        RECT 565.950 510.600 568.050 511.050 ;
        RECT 559.950 509.400 568.050 510.600 ;
        RECT 559.950 508.950 562.050 509.400 ;
        RECT 565.950 508.950 568.050 509.400 ;
        RECT 652.950 510.600 655.050 511.050 ;
        RECT 703.950 510.600 706.050 511.050 ;
        RECT 652.950 509.400 706.050 510.600 ;
        RECT 652.950 508.950 655.050 509.400 ;
        RECT 703.950 508.950 706.050 509.400 ;
        RECT 709.950 510.600 712.050 511.050 ;
        RECT 781.950 510.600 784.050 511.050 ;
        RECT 808.950 510.600 811.050 511.050 ;
        RECT 709.950 509.400 811.050 510.600 ;
        RECT 709.950 508.950 712.050 509.400 ;
        RECT 781.950 508.950 784.050 509.400 ;
        RECT 808.950 508.950 811.050 509.400 ;
        RECT 832.950 510.600 835.050 511.050 ;
        RECT 871.950 510.600 874.050 511.050 ;
        RECT 832.950 509.400 874.050 510.600 ;
        RECT 832.950 508.950 835.050 509.400 ;
        RECT 871.950 508.950 874.050 509.400 ;
        RECT 889.950 510.600 892.050 511.050 ;
        RECT 925.950 510.600 928.050 511.050 ;
        RECT 889.950 509.400 928.050 510.600 ;
        RECT 889.950 508.950 892.050 509.400 ;
        RECT 925.950 508.950 928.050 509.400 ;
        RECT 19.950 507.600 22.050 508.050 ;
        RECT 235.950 507.600 238.050 508.050 ;
        RECT 19.950 506.400 238.050 507.600 ;
        RECT 19.950 505.950 22.050 506.400 ;
        RECT 235.950 505.950 238.050 506.400 ;
        RECT 271.950 507.600 274.050 508.050 ;
        RECT 352.950 507.600 355.050 508.050 ;
        RECT 271.950 506.400 355.050 507.600 ;
        RECT 271.950 505.950 274.050 506.400 ;
        RECT 352.950 505.950 355.050 506.400 ;
        RECT 421.950 507.600 424.050 508.050 ;
        RECT 568.950 507.600 571.050 508.050 ;
        RECT 610.950 507.600 613.050 508.050 ;
        RECT 616.950 507.600 619.050 508.050 ;
        RECT 421.950 506.400 474.600 507.600 ;
        RECT 421.950 505.950 424.050 506.400 ;
        RECT 190.950 504.600 193.050 505.050 ;
        RECT 196.950 504.600 199.050 505.050 ;
        RECT 220.950 504.600 223.050 505.050 ;
        RECT 229.950 504.600 232.050 505.050 ;
        RECT 190.950 503.400 232.050 504.600 ;
        RECT 190.950 502.950 193.050 503.400 ;
        RECT 196.950 502.950 199.050 503.400 ;
        RECT 220.950 502.950 223.050 503.400 ;
        RECT 229.950 502.950 232.050 503.400 ;
        RECT 379.950 504.600 382.050 505.050 ;
        RECT 388.950 504.600 391.050 505.050 ;
        RECT 379.950 503.400 391.050 504.600 ;
        RECT 379.950 502.950 382.050 503.400 ;
        RECT 388.950 502.950 391.050 503.400 ;
        RECT 409.950 504.600 412.050 505.050 ;
        RECT 436.950 504.600 439.050 505.050 ;
        RECT 409.950 503.400 439.050 504.600 ;
        RECT 473.400 504.600 474.600 506.400 ;
        RECT 568.950 506.400 619.050 507.600 ;
        RECT 568.950 505.950 571.050 506.400 ;
        RECT 610.950 505.950 613.050 506.400 ;
        RECT 616.950 505.950 619.050 506.400 ;
        RECT 643.950 507.600 646.050 508.050 ;
        RECT 778.950 507.600 781.050 508.050 ;
        RECT 643.950 506.400 781.050 507.600 ;
        RECT 643.950 505.950 646.050 506.400 ;
        RECT 778.950 505.950 781.050 506.400 ;
        RECT 847.950 507.600 850.050 508.050 ;
        RECT 868.950 507.600 871.050 508.050 ;
        RECT 847.950 506.400 871.050 507.600 ;
        RECT 847.950 505.950 850.050 506.400 ;
        RECT 868.950 505.950 871.050 506.400 ;
        RECT 883.950 507.600 886.050 508.050 ;
        RECT 916.950 507.600 919.050 508.050 ;
        RECT 883.950 506.400 919.050 507.600 ;
        RECT 883.950 505.950 886.050 506.400 ;
        RECT 916.950 505.950 919.050 506.400 ;
        RECT 949.950 507.600 952.050 508.050 ;
        RECT 1000.950 507.600 1003.050 508.050 ;
        RECT 949.950 506.400 1003.050 507.600 ;
        RECT 949.950 505.950 952.050 506.400 ;
        RECT 1000.950 505.950 1003.050 506.400 ;
        RECT 511.950 504.600 514.050 505.050 ;
        RECT 473.400 503.400 514.050 504.600 ;
        RECT 409.950 502.950 412.050 503.400 ;
        RECT 436.950 502.950 439.050 503.400 ;
        RECT 511.950 502.950 514.050 503.400 ;
        RECT 691.950 504.600 694.050 505.050 ;
        RECT 724.950 504.600 727.050 505.050 ;
        RECT 739.950 504.600 742.050 505.050 ;
        RECT 691.950 503.400 742.050 504.600 ;
        RECT 691.950 502.950 694.050 503.400 ;
        RECT 724.950 502.950 727.050 503.400 ;
        RECT 739.950 502.950 742.050 503.400 ;
        RECT 925.950 504.600 928.050 505.050 ;
        RECT 937.950 504.600 940.050 505.050 ;
        RECT 925.950 503.400 940.050 504.600 ;
        RECT 925.950 502.950 928.050 503.400 ;
        RECT 937.950 502.950 940.050 503.400 ;
        RECT 1003.950 504.600 1006.050 505.050 ;
        RECT 1009.950 504.600 1012.050 508.050 ;
        RECT 1003.950 504.000 1012.050 504.600 ;
        RECT 1003.950 503.400 1011.600 504.000 ;
        RECT 1003.950 502.950 1006.050 503.400 ;
        RECT 127.950 501.600 130.050 502.050 ;
        RECT 148.950 501.600 151.050 502.050 ;
        RECT 127.950 500.400 151.050 501.600 ;
        RECT 127.950 499.950 130.050 500.400 ;
        RECT 148.950 499.950 151.050 500.400 ;
        RECT 154.950 501.600 157.050 502.050 ;
        RECT 181.950 501.600 184.050 502.050 ;
        RECT 154.950 500.400 184.050 501.600 ;
        RECT 154.950 499.950 157.050 500.400 ;
        RECT 181.950 499.950 184.050 500.400 ;
        RECT 199.950 501.600 202.050 502.050 ;
        RECT 271.950 501.600 274.050 502.050 ;
        RECT 199.950 500.400 274.050 501.600 ;
        RECT 199.950 499.950 202.050 500.400 ;
        RECT 271.950 499.950 274.050 500.400 ;
        RECT 340.950 501.600 343.050 502.050 ;
        RECT 358.950 501.600 361.050 502.050 ;
        RECT 340.950 500.400 361.050 501.600 ;
        RECT 340.950 499.950 343.050 500.400 ;
        RECT 358.950 499.950 361.050 500.400 ;
        RECT 367.950 501.600 370.050 502.050 ;
        RECT 415.950 501.600 418.050 502.050 ;
        RECT 463.950 501.600 466.050 502.050 ;
        RECT 367.950 500.400 466.050 501.600 ;
        RECT 367.950 499.950 370.050 500.400 ;
        RECT 415.950 499.950 418.050 500.400 ;
        RECT 463.950 499.950 466.050 500.400 ;
        RECT 469.950 501.600 472.050 502.050 ;
        RECT 544.950 501.600 547.050 502.050 ;
        RECT 559.950 501.600 562.050 502.050 ;
        RECT 469.950 500.400 562.050 501.600 ;
        RECT 469.950 499.950 472.050 500.400 ;
        RECT 544.950 499.950 547.050 500.400 ;
        RECT 559.950 499.950 562.050 500.400 ;
        RECT 601.950 501.600 604.050 502.050 ;
        RECT 631.950 501.600 634.050 502.050 ;
        RECT 601.950 500.400 634.050 501.600 ;
        RECT 601.950 499.950 604.050 500.400 ;
        RECT 631.950 499.950 634.050 500.400 ;
        RECT 643.950 501.600 646.050 502.050 ;
        RECT 655.950 501.600 658.050 502.050 ;
        RECT 643.950 500.400 658.050 501.600 ;
        RECT 643.950 499.950 646.050 500.400 ;
        RECT 655.950 499.950 658.050 500.400 ;
        RECT 664.950 501.600 667.050 502.050 ;
        RECT 679.950 501.600 682.050 502.050 ;
        RECT 664.950 500.400 682.050 501.600 ;
        RECT 664.950 499.950 667.050 500.400 ;
        RECT 679.950 499.950 682.050 500.400 ;
        RECT 778.950 501.600 781.050 502.050 ;
        RECT 805.950 501.600 808.050 502.050 ;
        RECT 778.950 500.400 808.050 501.600 ;
        RECT 778.950 499.950 781.050 500.400 ;
        RECT 805.950 499.950 808.050 500.400 ;
        RECT 820.950 501.600 823.050 502.050 ;
        RECT 859.950 501.600 862.050 502.050 ;
        RECT 820.950 500.400 862.050 501.600 ;
        RECT 820.950 499.950 823.050 500.400 ;
        RECT 859.950 499.950 862.050 500.400 ;
        RECT 871.950 501.600 874.050 502.050 ;
        RECT 877.950 501.600 880.050 502.050 ;
        RECT 871.950 500.400 880.050 501.600 ;
        RECT 871.950 499.950 874.050 500.400 ;
        RECT 877.950 499.950 880.050 500.400 ;
        RECT 904.950 501.600 907.050 502.050 ;
        RECT 910.950 501.600 913.050 502.050 ;
        RECT 904.950 500.400 913.050 501.600 ;
        RECT 904.950 499.950 907.050 500.400 ;
        RECT 910.950 499.950 913.050 500.400 ;
        RECT 943.950 501.600 946.050 502.050 ;
        RECT 961.950 501.600 964.050 502.050 ;
        RECT 964.950 501.600 967.050 502.050 ;
        RECT 943.950 500.400 967.050 501.600 ;
        RECT 943.950 499.950 946.050 500.400 ;
        RECT 961.950 499.950 964.050 500.400 ;
        RECT 964.950 499.950 967.050 500.400 ;
        RECT 991.950 501.600 994.050 502.050 ;
        RECT 1000.950 501.600 1003.050 502.050 ;
        RECT 991.950 500.400 1003.050 501.600 ;
        RECT 991.950 499.950 994.050 500.400 ;
        RECT 1000.950 499.950 1003.050 500.400 ;
        RECT 193.950 498.600 196.050 499.050 ;
        RECT 208.950 498.600 211.050 499.050 ;
        RECT 193.950 497.400 211.050 498.600 ;
        RECT 193.950 496.950 196.050 497.400 ;
        RECT 208.950 496.950 211.050 497.400 ;
        RECT 232.950 496.950 235.050 499.050 ;
        RECT 280.950 498.600 283.050 499.050 ;
        RECT 280.950 497.400 291.600 498.600 ;
        RECT 280.950 496.950 283.050 497.400 ;
        RECT 91.950 495.600 94.050 496.200 ;
        RECT 133.950 495.750 136.050 496.200 ;
        RECT 148.950 495.750 151.050 496.200 ;
        RECT 91.950 494.400 99.600 495.600 ;
        RECT 91.950 494.100 94.050 494.400 ;
        RECT 73.950 489.450 76.050 489.900 ;
        RECT 82.950 489.450 85.050 489.900 ;
        RECT 73.950 488.250 85.050 489.450 ;
        RECT 98.400 489.600 99.600 494.400 ;
        RECT 133.950 494.550 151.050 495.750 ;
        RECT 133.950 494.100 136.050 494.550 ;
        RECT 148.950 494.100 151.050 494.550 ;
        RECT 154.950 494.100 157.050 496.200 ;
        RECT 163.950 495.750 166.050 496.200 ;
        RECT 169.950 495.750 172.050 496.200 ;
        RECT 163.950 494.550 172.050 495.750 ;
        RECT 163.950 494.100 166.050 494.550 ;
        RECT 169.950 494.100 172.050 494.550 ;
        RECT 109.950 489.600 112.050 489.900 ;
        RECT 98.400 488.400 112.050 489.600 ;
        RECT 155.400 489.600 156.600 494.100 ;
        RECT 233.400 489.900 234.600 496.950 ;
        RECT 290.400 489.900 291.600 497.400 ;
        RECT 385.950 496.950 388.050 499.050 ;
        RECT 445.950 498.600 448.050 499.050 ;
        RECT 457.950 498.600 460.050 499.050 ;
        RECT 670.950 498.600 673.050 499.050 ;
        RECT 445.950 497.400 460.050 498.600 ;
        RECT 445.950 496.950 448.050 497.400 ;
        RECT 457.950 496.950 460.050 497.400 ;
        RECT 653.400 497.400 673.050 498.600 ;
        RECT 316.950 495.600 319.050 496.050 ;
        RECT 331.950 495.600 334.050 496.200 ;
        RECT 336.000 495.600 340.050 496.050 ;
        RECT 351.000 495.600 355.050 496.050 ;
        RECT 316.950 494.400 334.050 495.600 ;
        RECT 316.950 493.950 319.050 494.400 ;
        RECT 331.950 494.100 334.050 494.400 ;
        RECT 335.400 493.950 340.050 495.600 ;
        RECT 350.400 493.950 355.050 495.600 ;
        RECT 335.400 489.900 336.600 493.950 ;
        RECT 350.400 489.900 351.600 493.950 ;
        RECT 386.400 489.900 387.600 496.950 ;
        RECT 418.950 495.600 421.050 496.050 ;
        RECT 436.950 495.600 439.050 496.200 ;
        RECT 418.950 494.400 439.050 495.600 ;
        RECT 418.950 493.950 421.050 494.400 ;
        RECT 436.950 494.100 439.050 494.400 ;
        RECT 463.950 495.750 466.050 496.200 ;
        RECT 499.950 495.750 502.050 496.200 ;
        RECT 463.950 494.550 502.050 495.750 ;
        RECT 463.950 494.100 466.050 494.550 ;
        RECT 499.950 494.100 502.050 494.550 ;
        RECT 511.950 495.750 514.050 496.200 ;
        RECT 529.950 495.750 532.050 496.200 ;
        RECT 511.950 494.550 532.050 495.750 ;
        RECT 511.950 494.100 514.050 494.550 ;
        RECT 529.950 494.100 532.050 494.550 ;
        RECT 553.950 495.600 556.050 496.200 ;
        RECT 559.950 495.600 562.050 496.200 ;
        RECT 610.950 495.600 613.050 496.200 ;
        RECT 553.950 494.400 562.050 495.600 ;
        RECT 553.950 494.100 556.050 494.400 ;
        RECT 559.950 494.100 562.050 494.400 ;
        RECT 599.400 494.400 613.050 495.600 ;
        RECT 599.400 492.600 600.600 494.400 ;
        RECT 610.950 494.100 613.050 494.400 ;
        RECT 649.950 495.600 652.050 496.200 ;
        RECT 653.400 495.600 654.600 497.400 ;
        RECT 670.950 496.950 673.050 497.400 ;
        RECT 676.950 498.600 679.050 499.050 ;
        RECT 691.950 498.600 694.050 499.050 ;
        RECT 676.950 497.400 694.050 498.600 ;
        RECT 676.950 496.950 679.050 497.400 ;
        RECT 691.950 496.950 694.050 497.400 ;
        RECT 925.950 498.600 928.050 499.050 ;
        RECT 940.950 498.600 943.050 499.050 ;
        RECT 925.950 497.400 943.050 498.600 ;
        RECT 925.950 496.950 928.050 497.400 ;
        RECT 940.950 496.950 943.050 497.400 ;
        RECT 952.950 498.600 955.050 499.050 ;
        RECT 958.950 498.600 961.050 499.050 ;
        RECT 952.950 497.400 961.050 498.600 ;
        RECT 965.400 498.600 966.600 499.950 ;
        RECT 988.950 498.600 991.050 499.050 ;
        RECT 965.400 497.400 991.050 498.600 ;
        RECT 952.950 496.950 955.050 497.400 ;
        RECT 958.950 496.950 961.050 497.400 ;
        RECT 988.950 496.950 991.050 497.400 ;
        RECT 649.950 494.400 654.600 495.600 ;
        RECT 655.950 495.750 658.050 496.200 ;
        RECT 664.800 495.750 666.900 496.200 ;
        RECT 655.950 494.550 666.900 495.750 ;
        RECT 649.950 494.100 652.050 494.400 ;
        RECT 655.950 494.100 658.050 494.550 ;
        RECT 664.800 494.100 666.900 494.550 ;
        RECT 650.400 492.600 651.600 494.100 ;
        RECT 667.950 493.950 670.050 496.050 ;
        RECT 679.950 495.750 682.050 496.200 ;
        RECT 700.950 495.750 703.050 496.200 ;
        RECT 679.950 494.550 703.050 495.750 ;
        RECT 679.950 494.100 682.050 494.550 ;
        RECT 700.950 494.100 703.050 494.550 ;
        RECT 751.950 495.600 754.050 496.200 ;
        RECT 763.950 495.750 766.050 496.200 ;
        RECT 769.950 495.750 772.050 496.200 ;
        RECT 763.950 495.600 772.050 495.750 ;
        RECT 787.950 495.600 790.050 496.200 ;
        RECT 751.950 494.400 759.600 495.600 ;
        RECT 751.950 494.100 754.050 494.400 ;
        RECT 587.400 491.400 600.600 492.600 ;
        RECT 638.400 492.000 651.600 492.600 ;
        RECT 637.950 491.400 651.600 492.000 ;
        RECT 172.950 489.600 175.050 489.900 ;
        RECT 155.400 488.400 175.050 489.600 ;
        RECT 73.950 487.800 76.050 488.250 ;
        RECT 82.950 487.800 85.050 488.250 ;
        RECT 109.950 487.800 112.050 488.400 ;
        RECT 172.950 487.800 175.050 488.400 ;
        RECT 181.950 489.450 184.050 489.900 ;
        RECT 187.950 489.450 190.050 489.900 ;
        RECT 181.950 488.250 190.050 489.450 ;
        RECT 181.950 487.800 184.050 488.250 ;
        RECT 187.950 487.800 190.050 488.250 ;
        RECT 232.950 487.800 235.050 489.900 ;
        RECT 238.950 489.450 241.050 489.900 ;
        RECT 262.950 489.450 265.050 489.900 ;
        RECT 238.950 488.250 265.050 489.450 ;
        RECT 238.950 487.800 241.050 488.250 ;
        RECT 262.950 487.800 265.050 488.250 ;
        RECT 289.950 487.800 292.050 489.900 ;
        RECT 319.950 489.450 322.050 489.900 ;
        RECT 328.950 489.450 331.050 489.900 ;
        RECT 319.950 488.250 331.050 489.450 ;
        RECT 319.950 487.800 322.050 488.250 ;
        RECT 328.950 487.800 331.050 488.250 ;
        RECT 334.950 487.800 337.050 489.900 ;
        RECT 349.950 487.800 352.050 489.900 ;
        RECT 385.950 487.800 388.050 489.900 ;
        RECT 421.950 489.450 424.050 489.900 ;
        RECT 433.950 489.450 436.050 489.900 ;
        RECT 421.950 488.250 436.050 489.450 ;
        RECT 421.950 487.800 424.050 488.250 ;
        RECT 433.950 487.800 436.050 488.250 ;
        RECT 439.950 489.450 442.050 489.900 ;
        RECT 445.950 489.450 448.050 489.900 ;
        RECT 439.950 488.250 448.050 489.450 ;
        RECT 439.950 487.800 442.050 488.250 ;
        RECT 445.950 487.800 448.050 488.250 ;
        RECT 505.950 489.600 508.050 489.900 ;
        RECT 511.950 489.600 514.050 490.050 ;
        RECT 505.950 488.400 514.050 489.600 ;
        RECT 505.950 487.800 508.050 488.400 ;
        RECT 511.950 487.950 514.050 488.400 ;
        RECT 577.950 489.600 580.050 489.900 ;
        RECT 587.400 489.600 588.600 491.400 ;
        RECT 577.950 488.400 588.600 489.600 ;
        RECT 598.950 489.450 601.050 489.900 ;
        RECT 607.950 489.450 610.050 489.900 ;
        RECT 577.950 487.800 580.050 488.400 ;
        RECT 598.950 488.250 610.050 489.450 ;
        RECT 598.950 487.800 601.050 488.250 ;
        RECT 607.950 487.800 610.050 488.250 ;
        RECT 637.950 487.950 640.050 491.400 ;
        RECT 668.400 490.050 669.600 493.950 ;
        RECT 758.400 493.050 759.600 494.400 ;
        RECT 763.950 494.550 790.050 495.600 ;
        RECT 763.950 494.100 766.050 494.550 ;
        RECT 769.950 494.400 790.050 494.550 ;
        RECT 769.950 494.100 772.050 494.400 ;
        RECT 787.950 494.100 790.050 494.400 ;
        RECT 802.950 495.750 805.050 496.200 ;
        RECT 814.950 495.750 817.050 496.200 ;
        RECT 802.950 494.550 817.050 495.750 ;
        RECT 802.950 494.100 805.050 494.550 ;
        RECT 814.950 494.100 817.050 494.550 ;
        RECT 841.950 494.100 844.050 496.200 ;
        RECT 895.950 495.600 898.050 496.200 ;
        RECT 895.950 494.400 906.600 495.600 ;
        RECT 895.950 494.100 898.050 494.400 ;
        RECT 712.950 492.600 715.050 493.050 ;
        RECT 712.950 491.400 750.600 492.600 ;
        RECT 758.400 491.400 763.050 493.050 ;
        RECT 712.950 490.950 715.050 491.400 ;
        RECT 643.950 489.600 646.050 490.050 ;
        RECT 652.950 489.600 655.050 489.900 ;
        RECT 643.950 488.400 655.050 489.600 ;
        RECT 643.950 487.950 646.050 488.400 ;
        RECT 652.950 487.800 655.050 488.400 ;
        RECT 667.950 487.950 670.050 490.050 ;
        RECT 749.400 489.900 750.600 491.400 ;
        RECT 759.000 490.950 763.050 491.400 ;
        RECT 748.950 487.800 751.050 489.900 ;
        RECT 805.950 489.450 808.050 489.900 ;
        RECT 811.950 489.450 814.050 489.900 ;
        RECT 805.950 488.250 814.050 489.450 ;
        RECT 842.400 489.600 843.600 494.100 ;
        RECT 901.950 490.950 904.050 493.050 ;
        RECT 847.950 489.600 850.050 490.050 ;
        RECT 859.950 489.600 862.050 490.050 ;
        RECT 842.400 489.000 846.600 489.600 ;
        RECT 842.400 488.400 847.050 489.000 ;
        RECT 805.950 487.800 808.050 488.250 ;
        RECT 811.950 487.800 814.050 488.250 ;
        RECT 55.950 486.600 58.050 487.050 ;
        RECT 64.950 486.600 67.050 487.050 ;
        RECT 55.950 485.400 67.050 486.600 ;
        RECT 55.950 484.950 58.050 485.400 ;
        RECT 64.950 484.950 67.050 485.400 ;
        RECT 151.950 486.600 154.050 487.050 ;
        RECT 160.950 486.600 163.050 487.050 ;
        RECT 151.950 485.400 163.050 486.600 ;
        RECT 151.950 484.950 154.050 485.400 ;
        RECT 160.950 484.950 163.050 485.400 ;
        RECT 358.950 486.600 361.050 487.050 ;
        RECT 391.950 486.600 394.050 487.050 ;
        RECT 358.950 485.400 394.050 486.600 ;
        RECT 358.950 484.950 361.050 485.400 ;
        RECT 391.950 484.950 394.050 485.400 ;
        RECT 694.950 486.600 697.050 487.050 ;
        RECT 730.950 486.600 733.050 487.050 ;
        RECT 694.950 485.400 733.050 486.600 ;
        RECT 694.950 484.950 697.050 485.400 ;
        RECT 730.950 484.950 733.050 485.400 ;
        RECT 760.950 486.600 763.050 487.050 ;
        RECT 796.950 486.600 799.050 487.050 ;
        RECT 760.950 485.400 799.050 486.600 ;
        RECT 760.950 484.950 763.050 485.400 ;
        RECT 796.950 484.950 799.050 485.400 ;
        RECT 844.950 484.950 847.050 488.400 ;
        RECT 847.950 488.400 862.050 489.600 ;
        RECT 847.950 487.950 850.050 488.400 ;
        RECT 859.950 487.950 862.050 488.400 ;
        RECT 877.950 489.450 880.050 490.050 ;
        RECT 886.950 489.450 889.050 489.900 ;
        RECT 877.950 488.250 889.050 489.450 ;
        RECT 877.950 487.950 880.050 488.250 ;
        RECT 886.950 487.800 889.050 488.250 ;
        RECT 856.950 486.600 859.050 487.050 ;
        RECT 865.950 486.600 868.050 487.050 ;
        RECT 856.950 485.400 868.050 486.600 ;
        RECT 856.950 484.950 859.050 485.400 ;
        RECT 865.950 484.950 868.050 485.400 ;
        RECT 883.950 486.600 886.050 487.050 ;
        RECT 902.400 486.600 903.600 490.950 ;
        RECT 883.950 485.400 903.600 486.600 ;
        RECT 905.400 486.600 906.600 494.400 ;
        RECT 910.950 494.100 913.050 496.200 ;
        RECT 931.950 495.600 936.000 496.050 ;
        RECT 994.950 495.600 997.050 496.200 ;
        RECT 911.400 490.050 912.600 494.100 ;
        RECT 931.950 493.950 936.600 495.600 ;
        RECT 907.950 488.400 912.600 490.050 ;
        RECT 919.950 489.450 922.050 489.900 ;
        RECT 925.950 489.450 928.050 490.050 ;
        RECT 907.950 487.950 912.000 488.400 ;
        RECT 919.950 488.250 928.050 489.450 ;
        RECT 935.400 489.600 936.600 493.950 ;
        RECT 992.400 494.400 997.050 495.600 ;
        RECT 979.950 492.600 982.050 493.050 ;
        RECT 992.400 492.600 993.600 494.400 ;
        RECT 994.950 494.100 997.050 494.400 ;
        RECT 979.950 491.400 993.600 492.600 ;
        RECT 979.950 490.950 982.050 491.400 ;
        RECT 940.950 489.600 943.050 489.900 ;
        RECT 935.400 488.400 943.050 489.600 ;
        RECT 919.950 487.800 922.050 488.250 ;
        RECT 925.950 487.950 928.050 488.250 ;
        RECT 940.950 487.800 943.050 488.400 ;
        RECT 949.950 489.600 952.050 490.050 ;
        RECT 955.950 489.600 958.050 490.050 ;
        RECT 949.950 488.400 958.050 489.600 ;
        RECT 949.950 487.950 952.050 488.400 ;
        RECT 955.950 487.950 958.050 488.400 ;
        RECT 967.950 489.600 970.050 489.900 ;
        RECT 985.950 489.600 988.050 489.900 ;
        RECT 967.950 488.400 988.050 489.600 ;
        RECT 967.950 487.800 970.050 488.400 ;
        RECT 985.950 487.800 988.050 488.400 ;
        RECT 913.950 486.600 916.050 487.050 ;
        RECT 905.400 485.400 916.050 486.600 ;
        RECT 883.950 484.950 886.050 485.400 ;
        RECT 913.950 484.950 916.050 485.400 ;
        RECT 112.950 483.600 115.050 484.050 ;
        RECT 172.950 483.600 175.050 484.050 ;
        RECT 112.950 482.400 175.050 483.600 ;
        RECT 112.950 481.950 115.050 482.400 ;
        RECT 172.950 481.950 175.050 482.400 ;
        RECT 496.950 483.600 499.050 484.050 ;
        RECT 505.950 483.600 508.050 484.050 ;
        RECT 523.950 483.600 526.050 484.050 ;
        RECT 496.950 482.400 526.050 483.600 ;
        RECT 496.950 481.950 499.050 482.400 ;
        RECT 505.950 481.950 508.050 482.400 ;
        RECT 523.950 481.950 526.050 482.400 ;
        RECT 742.950 483.600 745.050 484.050 ;
        RECT 754.950 483.600 757.050 484.050 ;
        RECT 742.950 482.400 757.050 483.600 ;
        RECT 742.950 481.950 745.050 482.400 ;
        RECT 754.950 481.950 757.050 482.400 ;
        RECT 64.950 480.600 67.050 481.050 ;
        RECT 100.950 480.600 103.050 481.050 ;
        RECT 64.950 479.400 103.050 480.600 ;
        RECT 64.950 478.950 67.050 479.400 ;
        RECT 100.950 478.950 103.050 479.400 ;
        RECT 220.950 480.600 223.050 481.050 ;
        RECT 298.950 480.600 301.050 481.050 ;
        RECT 382.950 480.600 385.050 481.050 ;
        RECT 220.950 479.400 385.050 480.600 ;
        RECT 220.950 478.950 223.050 479.400 ;
        RECT 298.950 478.950 301.050 479.400 ;
        RECT 382.950 478.950 385.050 479.400 ;
        RECT 511.950 480.600 514.050 481.050 ;
        RECT 604.950 480.600 607.050 481.050 ;
        RECT 511.950 479.400 607.050 480.600 ;
        RECT 511.950 478.950 514.050 479.400 ;
        RECT 604.950 478.950 607.050 479.400 ;
        RECT 703.950 480.600 706.050 481.050 ;
        RECT 730.950 480.600 733.050 481.050 ;
        RECT 703.950 479.400 733.050 480.600 ;
        RECT 703.950 478.950 706.050 479.400 ;
        RECT 730.950 478.950 733.050 479.400 ;
        RECT 757.950 480.600 760.050 481.050 ;
        RECT 790.950 480.600 793.050 481.050 ;
        RECT 757.950 479.400 793.050 480.600 ;
        RECT 757.950 478.950 760.050 479.400 ;
        RECT 790.950 478.950 793.050 479.400 ;
        RECT 838.950 480.600 841.050 481.050 ;
        RECT 874.950 480.600 877.050 481.050 ;
        RECT 838.950 479.400 877.050 480.600 ;
        RECT 838.950 478.950 841.050 479.400 ;
        RECT 874.950 478.950 877.050 479.400 ;
        RECT 886.950 480.600 889.050 481.050 ;
        RECT 940.950 480.600 943.050 481.050 ;
        RECT 886.950 479.400 943.050 480.600 ;
        RECT 886.950 478.950 889.050 479.400 ;
        RECT 940.950 478.950 943.050 479.400 ;
        RECT 217.950 477.600 220.050 478.050 ;
        RECT 244.950 477.600 247.050 478.050 ;
        RECT 280.950 477.600 283.050 478.050 ;
        RECT 340.950 477.600 343.050 478.050 ;
        RECT 217.950 476.400 343.050 477.600 ;
        RECT 217.950 475.950 220.050 476.400 ;
        RECT 244.950 475.950 247.050 476.400 ;
        RECT 280.950 475.950 283.050 476.400 ;
        RECT 340.950 475.950 343.050 476.400 ;
        RECT 616.950 477.600 619.050 478.050 ;
        RECT 631.950 477.600 634.050 478.050 ;
        RECT 649.950 477.600 652.050 478.050 ;
        RECT 682.950 477.600 685.050 478.050 ;
        RECT 616.950 476.400 685.050 477.600 ;
        RECT 616.950 475.950 619.050 476.400 ;
        RECT 631.950 475.950 634.050 476.400 ;
        RECT 649.950 475.950 652.050 476.400 ;
        RECT 682.950 475.950 685.050 476.400 ;
        RECT 892.950 477.600 895.050 478.050 ;
        RECT 934.950 477.600 937.050 478.050 ;
        RECT 892.950 476.400 937.050 477.600 ;
        RECT 892.950 475.950 895.050 476.400 ;
        RECT 934.950 475.950 937.050 476.400 ;
        RECT 460.950 474.600 463.050 475.050 ;
        RECT 550.950 474.600 553.050 475.050 ;
        RECT 613.950 474.600 616.050 475.050 ;
        RECT 460.950 473.400 616.050 474.600 ;
        RECT 460.950 472.950 463.050 473.400 ;
        RECT 550.950 472.950 553.050 473.400 ;
        RECT 613.950 472.950 616.050 473.400 ;
        RECT 796.950 474.600 799.050 475.050 ;
        RECT 826.950 474.600 829.050 475.050 ;
        RECT 841.950 474.600 844.050 475.050 ;
        RECT 796.950 473.400 844.050 474.600 ;
        RECT 796.950 472.950 799.050 473.400 ;
        RECT 826.950 472.950 829.050 473.400 ;
        RECT 841.950 472.950 844.050 473.400 ;
        RECT 871.950 474.600 874.050 475.050 ;
        RECT 961.950 474.600 964.050 475.050 ;
        RECT 991.950 474.600 994.050 475.050 ;
        RECT 1000.950 474.600 1003.050 475.050 ;
        RECT 871.950 473.400 1003.050 474.600 ;
        RECT 871.950 472.950 874.050 473.400 ;
        RECT 961.950 472.950 964.050 473.400 ;
        RECT 991.950 472.950 994.050 473.400 ;
        RECT 1000.950 472.950 1003.050 473.400 ;
        RECT 79.950 471.600 82.050 472.050 ;
        RECT 124.950 471.600 127.050 472.050 ;
        RECT 79.950 470.400 127.050 471.600 ;
        RECT 79.950 469.950 82.050 470.400 ;
        RECT 124.950 469.950 127.050 470.400 ;
        RECT 223.950 471.600 226.050 472.050 ;
        RECT 256.950 471.600 259.050 472.050 ;
        RECT 292.950 471.600 295.050 472.050 ;
        RECT 223.950 470.400 295.050 471.600 ;
        RECT 223.950 469.950 226.050 470.400 ;
        RECT 256.950 469.950 259.050 470.400 ;
        RECT 292.950 469.950 295.050 470.400 ;
        RECT 508.950 471.600 511.050 472.050 ;
        RECT 631.950 471.600 634.050 472.050 ;
        RECT 508.950 470.400 634.050 471.600 ;
        RECT 508.950 469.950 511.050 470.400 ;
        RECT 631.950 469.950 634.050 470.400 ;
        RECT 646.950 471.600 649.050 472.050 ;
        RECT 670.950 471.600 673.050 472.050 ;
        RECT 646.950 470.400 673.050 471.600 ;
        RECT 646.950 469.950 649.050 470.400 ;
        RECT 670.950 469.950 673.050 470.400 ;
        RECT 844.950 471.600 847.050 472.050 ;
        RECT 895.950 471.600 898.050 472.050 ;
        RECT 907.950 471.600 910.050 472.050 ;
        RECT 844.950 470.400 910.050 471.600 ;
        RECT 844.950 469.950 847.050 470.400 ;
        RECT 895.950 469.950 898.050 470.400 ;
        RECT 907.950 469.950 910.050 470.400 ;
        RECT 919.950 471.600 922.050 472.050 ;
        RECT 967.950 471.600 970.050 472.050 ;
        RECT 919.950 470.400 970.050 471.600 ;
        RECT 919.950 469.950 922.050 470.400 ;
        RECT 967.950 469.950 970.050 470.400 ;
        RECT 181.950 468.600 184.050 469.050 ;
        RECT 217.950 468.600 220.050 469.050 ;
        RECT 181.950 467.400 220.050 468.600 ;
        RECT 181.950 466.950 184.050 467.400 ;
        RECT 217.950 466.950 220.050 467.400 ;
        RECT 262.950 468.600 265.050 469.050 ;
        RECT 340.950 468.600 343.050 469.050 ;
        RECT 262.950 467.400 343.050 468.600 ;
        RECT 262.950 466.950 265.050 467.400 ;
        RECT 340.950 466.950 343.050 467.400 ;
        RECT 517.950 468.600 520.050 469.050 ;
        RECT 595.950 468.600 598.050 469.050 ;
        RECT 517.950 467.400 598.050 468.600 ;
        RECT 517.950 466.950 520.050 467.400 ;
        RECT 595.950 466.950 598.050 467.400 ;
        RECT 604.950 468.600 607.050 469.050 ;
        RECT 616.950 468.600 619.050 469.050 ;
        RECT 604.950 467.400 619.050 468.600 ;
        RECT 604.950 466.950 607.050 467.400 ;
        RECT 616.950 466.950 619.050 467.400 ;
        RECT 640.950 468.600 643.050 469.050 ;
        RECT 691.950 468.600 694.050 469.050 ;
        RECT 640.950 467.400 694.050 468.600 ;
        RECT 640.950 466.950 643.050 467.400 ;
        RECT 691.950 466.950 694.050 467.400 ;
        RECT 700.950 468.600 703.050 469.050 ;
        RECT 760.950 468.600 763.050 469.050 ;
        RECT 700.950 467.400 763.050 468.600 ;
        RECT 700.950 466.950 703.050 467.400 ;
        RECT 760.950 466.950 763.050 467.400 ;
        RECT 862.950 468.600 865.050 469.050 ;
        RECT 892.950 468.600 895.050 469.050 ;
        RECT 862.950 467.400 895.050 468.600 ;
        RECT 862.950 466.950 865.050 467.400 ;
        RECT 892.950 466.950 895.050 467.400 ;
        RECT 970.950 468.600 973.050 469.050 ;
        RECT 1015.950 468.600 1018.050 469.050 ;
        RECT 970.950 467.400 1018.050 468.600 ;
        RECT 970.950 466.950 973.050 467.400 ;
        RECT 1015.950 466.950 1018.050 467.400 ;
        RECT 97.950 465.600 100.050 466.050 ;
        RECT 157.950 465.600 160.050 466.050 ;
        RECT 97.950 464.400 160.050 465.600 ;
        RECT 97.950 463.950 100.050 464.400 ;
        RECT 157.950 463.950 160.050 464.400 ;
        RECT 169.950 465.600 172.050 466.050 ;
        RECT 253.950 465.600 256.050 466.050 ;
        RECT 169.950 464.400 256.050 465.600 ;
        RECT 169.950 463.950 172.050 464.400 ;
        RECT 253.950 463.950 256.050 464.400 ;
        RECT 355.950 465.600 358.050 466.050 ;
        RECT 469.950 465.600 472.050 466.050 ;
        RECT 355.950 464.400 472.050 465.600 ;
        RECT 355.950 463.950 358.050 464.400 ;
        RECT 469.950 463.950 472.050 464.400 ;
        RECT 625.950 465.600 628.050 466.050 ;
        RECT 697.950 465.600 700.050 466.050 ;
        RECT 838.950 465.600 841.050 466.050 ;
        RECT 863.400 465.600 864.600 466.950 ;
        RECT 625.950 464.400 700.050 465.600 ;
        RECT 625.950 463.950 628.050 464.400 ;
        RECT 697.950 463.950 700.050 464.400 ;
        RECT 725.400 464.400 841.050 465.600 ;
        RECT 725.400 463.050 726.600 464.400 ;
        RECT 838.950 463.950 841.050 464.400 ;
        RECT 845.400 464.400 864.600 465.600 ;
        RECT 82.950 462.600 85.050 463.050 ;
        RECT 121.950 462.600 124.050 463.050 ;
        RECT 82.950 461.400 124.050 462.600 ;
        RECT 82.950 460.950 85.050 461.400 ;
        RECT 121.950 460.950 124.050 461.400 ;
        RECT 373.950 462.600 376.050 463.050 ;
        RECT 511.950 462.600 514.050 463.050 ;
        RECT 373.950 461.400 514.050 462.600 ;
        RECT 373.950 460.950 376.050 461.400 ;
        RECT 511.950 460.950 514.050 461.400 ;
        RECT 544.950 462.600 547.050 463.050 ;
        RECT 550.950 462.600 553.050 463.050 ;
        RECT 586.950 462.600 589.050 463.050 ;
        RECT 598.950 462.600 601.050 463.050 ;
        RECT 544.950 461.400 601.050 462.600 ;
        RECT 544.950 460.950 547.050 461.400 ;
        RECT 550.950 460.950 553.050 461.400 ;
        RECT 586.950 460.950 589.050 461.400 ;
        RECT 598.950 460.950 601.050 461.400 ;
        RECT 631.950 462.600 634.050 463.050 ;
        RECT 661.950 462.600 664.050 463.050 ;
        RECT 631.950 461.400 664.050 462.600 ;
        RECT 631.950 460.950 634.050 461.400 ;
        RECT 661.950 460.950 664.050 461.400 ;
        RECT 721.950 461.400 726.600 463.050 ;
        RECT 727.950 462.600 730.050 463.050 ;
        RECT 799.950 462.600 802.050 463.050 ;
        RECT 727.950 461.400 802.050 462.600 ;
        RECT 721.950 460.950 726.000 461.400 ;
        RECT 727.950 460.950 730.050 461.400 ;
        RECT 799.950 460.950 802.050 461.400 ;
        RECT 829.950 462.600 832.050 463.050 ;
        RECT 845.400 462.600 846.600 464.400 ;
        RECT 829.950 461.400 846.600 462.600 ;
        RECT 886.950 462.600 889.050 463.050 ;
        RECT 901.950 462.600 904.050 463.050 ;
        RECT 886.950 461.400 904.050 462.600 ;
        RECT 829.950 460.950 832.050 461.400 ;
        RECT 886.950 460.950 889.050 461.400 ;
        RECT 901.950 460.950 904.050 461.400 ;
        RECT 907.950 462.600 910.050 463.050 ;
        RECT 952.950 462.600 955.050 463.050 ;
        RECT 907.950 461.400 955.050 462.600 ;
        RECT 907.950 460.950 910.050 461.400 ;
        RECT 952.950 460.950 955.050 461.400 ;
        RECT 976.950 462.600 979.050 463.050 ;
        RECT 1015.950 462.600 1018.050 463.050 ;
        RECT 976.950 461.400 1018.050 462.600 ;
        RECT 976.950 460.950 979.050 461.400 ;
        RECT 1015.950 460.950 1018.050 461.400 ;
        RECT 109.950 459.600 112.050 460.050 ;
        RECT 139.950 459.600 142.050 460.050 ;
        RECT 109.950 458.400 142.050 459.600 ;
        RECT 109.950 457.950 112.050 458.400 ;
        RECT 139.950 457.950 142.050 458.400 ;
        RECT 172.950 459.600 175.050 460.050 ;
        RECT 250.950 459.600 253.050 460.050 ;
        RECT 172.950 458.400 253.050 459.600 ;
        RECT 172.950 457.950 175.050 458.400 ;
        RECT 250.950 457.950 253.050 458.400 ;
        RECT 514.950 459.600 517.050 460.050 ;
        RECT 520.950 459.600 523.050 460.050 ;
        RECT 514.950 458.400 523.050 459.600 ;
        RECT 514.950 457.950 517.050 458.400 ;
        RECT 520.950 457.950 523.050 458.400 ;
        RECT 958.950 459.600 961.050 460.050 ;
        RECT 964.950 459.600 967.050 460.050 ;
        RECT 979.950 459.600 982.050 460.050 ;
        RECT 958.950 458.400 982.050 459.600 ;
        RECT 958.950 457.950 961.050 458.400 ;
        RECT 964.950 457.950 967.050 458.400 ;
        RECT 979.950 457.950 982.050 458.400 ;
        RECT 61.950 456.600 64.050 457.050 ;
        RECT 82.950 456.600 85.050 457.050 ;
        RECT 61.950 455.400 85.050 456.600 ;
        RECT 61.950 454.950 64.050 455.400 ;
        RECT 82.950 454.950 85.050 455.400 ;
        RECT 319.950 456.600 322.050 457.050 ;
        RECT 367.950 456.600 370.050 457.050 ;
        RECT 319.950 455.400 370.050 456.600 ;
        RECT 319.950 454.950 322.050 455.400 ;
        RECT 367.950 454.950 370.050 455.400 ;
        RECT 433.950 456.600 436.050 457.050 ;
        RECT 451.950 456.600 454.050 457.050 ;
        RECT 433.950 455.400 454.050 456.600 ;
        RECT 433.950 454.950 436.050 455.400 ;
        RECT 451.950 454.950 454.050 455.400 ;
        RECT 595.950 456.600 598.050 457.050 ;
        RECT 646.950 456.600 649.050 457.050 ;
        RECT 595.950 455.400 649.050 456.600 ;
        RECT 595.950 454.950 598.050 455.400 ;
        RECT 646.950 454.950 649.050 455.400 ;
        RECT 691.950 456.600 694.050 457.050 ;
        RECT 769.950 456.600 772.050 457.050 ;
        RECT 781.950 456.600 784.050 457.050 ;
        RECT 823.950 456.600 826.050 457.050 ;
        RECT 832.950 456.600 835.050 457.050 ;
        RECT 691.950 455.400 784.050 456.600 ;
        RECT 691.950 454.950 694.050 455.400 ;
        RECT 769.950 454.950 772.050 455.400 ;
        RECT 781.950 454.950 784.050 455.400 ;
        RECT 815.400 455.400 835.050 456.600 ;
        RECT 76.950 453.600 79.050 454.050 ;
        RECT 103.950 453.600 106.050 454.050 ;
        RECT 76.950 452.400 106.050 453.600 ;
        RECT 76.950 451.950 79.050 452.400 ;
        RECT 103.950 451.950 106.050 452.400 ;
        RECT 124.950 453.600 127.050 454.050 ;
        RECT 151.950 453.600 154.050 454.050 ;
        RECT 172.950 453.600 175.050 454.050 ;
        RECT 124.950 452.400 175.050 453.600 ;
        RECT 124.950 451.950 127.050 452.400 ;
        RECT 151.950 451.950 154.050 452.400 ;
        RECT 172.950 451.950 175.050 452.400 ;
        RECT 88.950 450.750 91.050 451.200 ;
        RECT 94.950 450.750 97.050 451.200 ;
        RECT 88.950 449.550 97.050 450.750 ;
        RECT 88.950 449.100 91.050 449.550 ;
        RECT 94.950 449.100 97.050 449.550 ;
        RECT 115.950 450.600 118.050 451.050 ;
        RECT 139.950 450.600 142.050 451.050 ;
        RECT 115.950 449.400 142.050 450.600 ;
        RECT 115.950 448.950 118.050 449.400 ;
        RECT 139.950 448.950 142.050 449.400 ;
        RECT 157.950 450.600 160.050 451.200 ;
        RECT 190.950 450.750 193.050 451.200 ;
        RECT 196.950 450.750 199.050 451.200 ;
        RECT 157.950 449.400 168.600 450.600 ;
        RECT 157.950 449.100 160.050 449.400 ;
        RECT 167.400 447.600 168.600 449.400 ;
        RECT 190.950 449.550 199.050 450.750 ;
        RECT 208.950 450.600 211.050 454.050 ;
        RECT 226.950 453.600 229.050 454.050 ;
        RECT 235.950 453.600 238.050 454.050 ;
        RECT 226.950 452.400 238.050 453.600 ;
        RECT 226.950 451.950 229.050 452.400 ;
        RECT 235.950 451.950 238.050 452.400 ;
        RECT 334.950 453.600 337.050 454.050 ;
        RECT 373.950 453.600 376.050 454.050 ;
        RECT 334.950 452.400 376.050 453.600 ;
        RECT 334.950 451.950 337.050 452.400 ;
        RECT 373.950 451.950 376.050 452.400 ;
        RECT 379.950 453.600 382.050 454.050 ;
        RECT 391.950 453.600 394.050 454.050 ;
        RECT 541.950 453.600 544.050 454.050 ;
        RECT 379.950 452.400 394.050 453.600 ;
        RECT 379.950 451.950 382.050 452.400 ;
        RECT 391.950 451.950 394.050 452.400 ;
        RECT 494.400 452.400 544.050 453.600 ;
        RECT 190.950 449.100 193.050 449.550 ;
        RECT 196.950 449.100 199.050 449.550 ;
        RECT 206.400 450.000 211.050 450.600 ;
        RECT 206.400 449.400 210.600 450.000 ;
        RECT 41.400 446.400 108.600 447.600 ;
        RECT 167.400 446.400 171.600 447.600 ;
        RECT 22.950 444.600 25.050 444.900 ;
        RECT 41.400 444.600 42.600 446.400 ;
        RECT 22.950 443.400 42.600 444.600 ;
        RECT 43.950 444.600 46.050 444.900 ;
        RECT 97.950 444.600 100.050 445.050 ;
        RECT 107.400 444.900 108.600 446.400 ;
        RECT 43.950 443.400 100.050 444.600 ;
        RECT 22.950 442.800 25.050 443.400 ;
        RECT 43.950 442.800 46.050 443.400 ;
        RECT 97.950 442.950 100.050 443.400 ;
        RECT 106.950 442.800 109.050 444.900 ;
        RECT 118.950 444.450 121.050 444.900 ;
        RECT 148.950 444.450 151.050 444.900 ;
        RECT 118.950 443.250 151.050 444.450 ;
        RECT 170.400 444.600 171.600 446.400 ;
        RECT 206.400 445.050 207.600 449.400 ;
        RECT 211.950 448.950 214.050 451.050 ;
        RECT 265.950 450.600 268.050 451.200 ;
        RECT 260.400 449.400 268.050 450.600 ;
        RECT 178.950 444.600 181.050 445.050 ;
        RECT 170.400 443.400 181.050 444.600 ;
        RECT 118.950 442.800 121.050 443.250 ;
        RECT 148.950 442.800 151.050 443.250 ;
        RECT 178.950 442.950 181.050 443.400 ;
        RECT 205.950 442.950 208.050 445.050 ;
        RECT 76.950 441.600 79.050 442.050 ;
        RECT 85.950 441.600 88.050 442.050 ;
        RECT 76.950 440.400 88.050 441.600 ;
        RECT 76.950 439.950 79.050 440.400 ;
        RECT 85.950 439.950 88.050 440.400 ;
        RECT 193.950 441.600 196.050 442.050 ;
        RECT 212.400 441.600 213.600 448.950 ;
        RECT 232.950 447.600 235.050 448.050 ;
        RECT 260.400 447.600 261.600 449.400 ;
        RECT 265.950 449.100 268.050 449.400 ;
        RECT 271.950 449.100 274.050 451.200 ;
        RECT 277.950 450.600 280.050 451.050 ;
        RECT 286.950 450.600 289.050 451.200 ;
        RECT 277.950 449.400 289.050 450.600 ;
        RECT 232.950 446.400 261.600 447.600 ;
        RECT 232.950 445.950 235.050 446.400 ;
        RECT 256.950 444.450 259.050 444.900 ;
        RECT 262.950 444.450 265.050 444.900 ;
        RECT 256.950 443.250 265.050 444.450 ;
        RECT 272.400 444.600 273.600 449.100 ;
        RECT 277.950 448.950 280.050 449.400 ;
        RECT 286.950 449.100 289.050 449.400 ;
        RECT 325.950 450.750 328.050 451.200 ;
        RECT 334.950 450.750 337.050 451.200 ;
        RECT 325.950 449.550 337.050 450.750 ;
        RECT 325.950 449.100 328.050 449.550 ;
        RECT 334.950 449.100 337.050 449.550 ;
        RECT 346.950 450.600 349.050 451.200 ;
        RECT 361.950 450.600 364.050 451.200 ;
        RECT 346.950 449.400 364.050 450.600 ;
        RECT 346.950 449.100 349.050 449.400 ;
        RECT 361.950 449.100 364.050 449.400 ;
        RECT 397.950 450.750 400.050 451.200 ;
        RECT 403.950 450.750 406.050 451.200 ;
        RECT 397.950 449.550 406.050 450.750 ;
        RECT 397.950 449.100 400.050 449.550 ;
        RECT 403.950 449.100 406.050 449.550 ;
        RECT 430.950 450.750 433.050 451.200 ;
        RECT 439.950 450.750 442.050 451.200 ;
        RECT 430.950 449.550 442.050 450.750 ;
        RECT 430.950 449.100 433.050 449.550 ;
        RECT 439.950 449.100 442.050 449.550 ;
        RECT 475.950 450.750 478.050 451.200 ;
        RECT 484.950 450.750 487.050 451.200 ;
        RECT 475.950 449.550 487.050 450.750 ;
        RECT 475.950 449.100 478.050 449.550 ;
        RECT 484.950 449.100 487.050 449.550 ;
        RECT 328.950 447.600 331.050 448.050 ;
        RECT 347.400 447.600 348.600 449.100 ;
        RECT 328.950 446.400 348.600 447.600 ;
        RECT 328.950 445.950 331.050 446.400 ;
        RECT 289.950 444.600 292.050 444.900 ;
        RECT 272.400 443.400 292.050 444.600 ;
        RECT 256.950 442.800 259.050 443.250 ;
        RECT 262.950 442.800 265.050 443.250 ;
        RECT 289.950 442.800 292.050 443.400 ;
        RECT 298.950 444.450 301.050 444.900 ;
        RECT 310.950 444.450 313.050 444.900 ;
        RECT 298.950 443.250 313.050 444.450 ;
        RECT 298.950 442.800 301.050 443.250 ;
        RECT 310.950 442.800 313.050 443.250 ;
        RECT 382.950 444.450 385.050 444.900 ;
        RECT 388.950 444.600 391.050 444.900 ;
        RECT 412.950 444.600 415.050 444.900 ;
        RECT 388.950 444.450 415.050 444.600 ;
        RECT 382.950 443.400 415.050 444.450 ;
        RECT 382.950 443.250 391.050 443.400 ;
        RECT 382.950 442.800 385.050 443.250 ;
        RECT 388.950 442.800 391.050 443.250 ;
        RECT 412.950 442.800 415.050 443.400 ;
        RECT 418.950 444.450 421.050 444.900 ;
        RECT 424.950 444.450 427.050 444.900 ;
        RECT 418.950 443.250 427.050 444.450 ;
        RECT 418.950 442.800 421.050 443.250 ;
        RECT 424.950 442.800 427.050 443.250 ;
        RECT 472.950 444.600 475.050 444.900 ;
        RECT 481.950 444.600 484.050 445.050 ;
        RECT 494.400 444.900 495.600 452.400 ;
        RECT 541.950 451.950 544.050 452.400 ;
        RECT 697.950 453.600 700.050 454.050 ;
        RECT 727.950 453.600 730.050 454.050 ;
        RECT 697.950 452.400 730.050 453.600 ;
        RECT 697.950 451.950 700.050 452.400 ;
        RECT 727.950 451.950 730.050 452.400 ;
        RECT 787.950 453.600 790.050 454.050 ;
        RECT 815.400 453.600 816.600 455.400 ;
        RECT 823.950 454.950 826.050 455.400 ;
        RECT 832.950 454.950 835.050 455.400 ;
        RECT 853.950 456.600 856.050 457.050 ;
        RECT 889.950 456.600 892.050 457.050 ;
        RECT 919.950 456.600 922.050 457.050 ;
        RECT 853.950 455.400 922.050 456.600 ;
        RECT 853.950 454.950 856.050 455.400 ;
        RECT 889.950 454.950 892.050 455.400 ;
        RECT 919.950 454.950 922.050 455.400 ;
        RECT 937.950 456.600 940.050 457.050 ;
        RECT 946.950 456.600 949.050 457.050 ;
        RECT 976.950 456.600 979.050 457.050 ;
        RECT 997.950 456.600 1000.050 457.050 ;
        RECT 937.950 455.400 979.050 456.600 ;
        RECT 937.950 454.950 940.050 455.400 ;
        RECT 946.950 454.950 949.050 455.400 ;
        RECT 976.950 454.950 979.050 455.400 ;
        RECT 989.400 455.400 1000.050 456.600 ;
        RECT 787.950 452.400 816.600 453.600 ;
        RECT 979.950 453.600 982.050 454.050 ;
        RECT 989.400 453.600 990.600 455.400 ;
        RECT 997.950 454.950 1000.050 455.400 ;
        RECT 979.950 452.400 990.600 453.600 ;
        RECT 787.950 451.950 790.050 452.400 ;
        RECT 979.950 451.950 982.050 452.400 ;
        RECT 520.950 447.600 523.050 451.050 ;
        RECT 571.950 450.600 574.050 451.050 ;
        RECT 577.950 450.600 580.050 451.200 ;
        RECT 571.950 449.400 580.050 450.600 ;
        RECT 571.950 448.950 574.050 449.400 ;
        RECT 577.950 449.100 580.050 449.400 ;
        RECT 664.950 450.600 667.050 451.050 ;
        RECT 676.950 450.600 679.050 451.200 ;
        RECT 664.950 449.400 679.050 450.600 ;
        RECT 664.950 448.950 667.050 449.400 ;
        RECT 671.400 447.600 672.600 449.400 ;
        RECT 676.950 449.100 679.050 449.400 ;
        RECT 682.950 449.100 685.050 451.200 ;
        RECT 691.950 450.750 694.050 451.200 ;
        RECT 706.950 450.750 709.050 451.200 ;
        RECT 691.950 449.550 709.050 450.750 ;
        RECT 691.950 449.100 694.050 449.550 ;
        RECT 706.950 449.100 709.050 449.550 ;
        RECT 512.400 447.000 523.050 447.600 ;
        RECT 511.950 446.400 522.600 447.000 ;
        RECT 665.400 446.400 672.600 447.600 ;
        RECT 683.400 447.600 684.600 449.100 ;
        RECT 712.950 447.600 715.050 451.050 ;
        RECT 721.950 448.950 724.050 451.050 ;
        RECT 730.950 450.750 733.050 451.200 ;
        RECT 742.950 450.750 745.050 451.200 ;
        RECT 730.950 449.550 745.050 450.750 ;
        RECT 730.950 449.100 733.050 449.550 ;
        RECT 742.950 449.100 745.050 449.550 ;
        RECT 817.950 449.100 820.050 451.200 ;
        RECT 847.950 450.750 850.050 451.200 ;
        RECT 853.950 450.750 856.050 451.200 ;
        RECT 847.950 450.600 856.050 450.750 ;
        RECT 874.950 450.600 877.050 451.200 ;
        RECT 847.950 449.550 877.050 450.600 ;
        RECT 847.950 449.100 850.050 449.550 ;
        RECT 853.950 449.400 877.050 449.550 ;
        RECT 853.950 449.100 856.050 449.400 ;
        RECT 874.950 449.100 877.050 449.400 ;
        RECT 683.400 447.000 715.050 447.600 ;
        RECT 683.400 446.400 714.600 447.000 ;
        RECT 472.950 443.400 484.050 444.600 ;
        RECT 472.950 442.800 475.050 443.400 ;
        RECT 481.950 442.950 484.050 443.400 ;
        RECT 493.950 442.800 496.050 444.900 ;
        RECT 511.950 442.950 514.050 446.400 ;
        RECT 517.950 444.600 520.050 444.900 ;
        RECT 523.950 444.600 526.050 444.900 ;
        RECT 517.950 443.400 526.050 444.600 ;
        RECT 517.950 442.800 520.050 443.400 ;
        RECT 523.950 442.800 526.050 443.400 ;
        RECT 553.950 444.600 556.050 445.050 ;
        RECT 568.950 444.600 571.050 445.050 ;
        RECT 553.950 443.400 571.050 444.600 ;
        RECT 553.950 442.950 556.050 443.400 ;
        RECT 568.950 442.950 571.050 443.400 ;
        RECT 610.950 444.600 613.050 444.900 ;
        RECT 658.950 444.600 661.050 444.900 ;
        RECT 665.400 444.600 666.600 446.400 ;
        RECT 610.950 444.000 618.600 444.600 ;
        RECT 610.950 443.400 619.050 444.000 ;
        RECT 610.950 442.800 613.050 443.400 ;
        RECT 193.950 440.400 213.600 441.600 ;
        RECT 244.950 441.600 247.050 442.050 ;
        RECT 277.950 441.600 280.050 442.050 ;
        RECT 355.950 441.600 358.050 442.050 ;
        RECT 244.950 440.400 358.050 441.600 ;
        RECT 193.950 439.950 196.050 440.400 ;
        RECT 244.950 439.950 247.050 440.400 ;
        RECT 277.950 439.950 280.050 440.400 ;
        RECT 355.950 439.950 358.050 440.400 ;
        RECT 394.950 441.600 397.050 442.050 ;
        RECT 400.950 441.600 403.050 442.050 ;
        RECT 394.950 440.400 403.050 441.600 ;
        RECT 394.950 439.950 397.050 440.400 ;
        RECT 400.950 439.950 403.050 440.400 ;
        RECT 616.950 439.950 619.050 443.400 ;
        RECT 658.950 443.400 666.600 444.600 ;
        RECT 667.950 444.600 670.050 445.050 ;
        RECT 673.950 444.600 676.050 445.050 ;
        RECT 667.950 443.400 676.050 444.600 ;
        RECT 658.950 442.800 661.050 443.400 ;
        RECT 667.950 442.950 670.050 443.400 ;
        RECT 673.950 442.950 676.050 443.400 ;
        RECT 679.950 444.600 682.050 444.900 ;
        RECT 691.950 444.600 694.050 445.050 ;
        RECT 679.950 443.400 694.050 444.600 ;
        RECT 679.950 442.800 682.050 443.400 ;
        RECT 691.950 442.950 694.050 443.400 ;
        RECT 695.400 441.600 696.600 446.400 ;
        RECT 709.950 444.600 712.050 444.900 ;
        RECT 722.400 444.600 723.600 448.950 ;
        RECT 808.950 447.600 811.050 448.050 ;
        RECT 818.400 447.600 819.600 449.100 ;
        RECT 886.950 448.950 889.050 451.050 ;
        RECT 895.950 450.600 898.050 451.200 ;
        RECT 913.950 450.600 916.050 451.200 ;
        RECT 895.950 449.400 916.050 450.600 ;
        RECT 895.950 449.100 898.050 449.400 ;
        RECT 913.950 449.100 916.050 449.400 ;
        RECT 937.950 448.950 940.050 451.050 ;
        RECT 946.950 450.600 949.050 451.200 ;
        RECT 970.950 450.600 973.050 451.050 ;
        RECT 946.950 449.400 973.050 450.600 ;
        RECT 946.950 449.100 949.050 449.400 ;
        RECT 970.950 448.950 973.050 449.400 ;
        RECT 976.950 450.750 979.050 451.200 ;
        RECT 991.950 450.750 994.050 451.200 ;
        RECT 976.950 449.550 994.050 450.750 ;
        RECT 976.950 449.100 979.050 449.550 ;
        RECT 808.950 446.400 819.600 447.600 ;
        RECT 808.950 445.950 811.050 446.400 ;
        RECT 887.400 445.050 888.600 448.950 ;
        RECT 709.950 443.400 723.600 444.600 ;
        RECT 727.950 444.600 730.050 444.900 ;
        RECT 739.950 444.600 742.050 445.050 ;
        RECT 727.950 443.400 742.050 444.600 ;
        RECT 709.950 442.800 712.050 443.400 ;
        RECT 727.950 442.800 730.050 443.400 ;
        RECT 739.950 442.950 742.050 443.400 ;
        RECT 751.950 444.600 754.050 444.900 ;
        RECT 760.950 444.600 763.050 445.050 ;
        RECT 751.950 443.400 763.050 444.600 ;
        RECT 751.950 442.800 754.050 443.400 ;
        RECT 760.950 442.950 763.050 443.400 ;
        RECT 772.950 444.600 775.050 444.900 ;
        RECT 787.950 444.600 790.050 445.050 ;
        RECT 772.950 443.400 790.050 444.600 ;
        RECT 772.950 442.800 775.050 443.400 ;
        RECT 787.950 442.950 790.050 443.400 ;
        RECT 832.950 444.450 835.050 444.900 ;
        RECT 838.950 444.450 841.050 444.900 ;
        RECT 832.950 443.250 841.050 444.450 ;
        RECT 832.950 442.800 835.050 443.250 ;
        RECT 838.950 442.800 841.050 443.250 ;
        RECT 844.950 444.600 847.050 444.900 ;
        RECT 880.950 444.600 883.050 445.050 ;
        RECT 844.950 443.400 883.050 444.600 ;
        RECT 844.950 442.800 847.050 443.400 ;
        RECT 880.950 442.950 883.050 443.400 ;
        RECT 886.950 442.950 889.050 445.050 ;
        RECT 904.950 444.450 907.050 444.900 ;
        RECT 916.950 444.450 919.050 444.900 ;
        RECT 904.950 443.250 919.050 444.450 ;
        RECT 904.950 442.800 907.050 443.250 ;
        RECT 916.950 442.800 919.050 443.250 ;
        RECT 922.950 444.600 925.050 444.900 ;
        RECT 931.950 444.600 934.050 445.050 ;
        RECT 922.950 443.400 934.050 444.600 ;
        RECT 938.400 444.600 939.600 448.950 ;
        RECT 989.400 445.050 990.600 449.550 ;
        RECT 991.950 449.100 994.050 449.550 ;
        RECT 1003.950 448.950 1006.050 451.050 ;
        RECT 949.950 444.600 952.050 444.900 ;
        RECT 938.400 443.400 952.050 444.600 ;
        RECT 922.950 442.800 925.050 443.400 ;
        RECT 931.950 442.950 934.050 443.400 ;
        RECT 949.950 442.800 952.050 443.400 ;
        RECT 955.950 444.600 960.000 445.050 ;
        RECT 955.950 442.950 960.600 444.600 ;
        RECT 988.950 442.950 991.050 445.050 ;
        RECT 706.950 441.600 709.050 442.050 ;
        RECT 695.400 440.400 709.050 441.600 ;
        RECT 706.950 439.950 709.050 440.400 ;
        RECT 775.950 441.600 778.050 442.050 ;
        RECT 781.950 441.600 784.050 442.050 ;
        RECT 775.950 440.400 784.050 441.600 ;
        RECT 775.950 439.950 778.050 440.400 ;
        RECT 781.950 439.950 784.050 440.400 ;
        RECT 892.950 441.600 895.050 442.050 ;
        RECT 905.400 441.600 906.600 442.800 ;
        RECT 892.950 440.400 906.600 441.600 ;
        RECT 934.950 441.600 937.050 442.050 ;
        RECT 940.950 441.600 943.050 442.050 ;
        RECT 934.950 440.400 943.050 441.600 ;
        RECT 959.400 441.600 960.600 442.950 ;
        RECT 1004.400 442.050 1005.600 448.950 ;
        RECT 964.950 441.600 967.050 442.050 ;
        RECT 959.400 440.400 967.050 441.600 ;
        RECT 892.950 439.950 895.050 440.400 ;
        RECT 934.950 439.950 937.050 440.400 ;
        RECT 940.950 439.950 943.050 440.400 ;
        RECT 964.950 439.950 967.050 440.400 ;
        RECT 982.950 441.600 985.050 442.050 ;
        RECT 997.950 441.600 1000.050 442.050 ;
        RECT 982.950 440.400 1000.050 441.600 ;
        RECT 1004.400 440.400 1009.050 442.050 ;
        RECT 982.950 439.950 985.050 440.400 ;
        RECT 997.950 439.950 1000.050 440.400 ;
        RECT 1005.000 439.950 1009.050 440.400 ;
        RECT 127.950 438.600 130.050 439.050 ;
        RECT 148.950 438.600 151.050 439.050 ;
        RECT 68.400 437.400 151.050 438.600 ;
        RECT 68.400 436.050 69.600 437.400 ;
        RECT 127.950 436.950 130.050 437.400 ;
        RECT 148.950 436.950 151.050 437.400 ;
        RECT 280.950 438.600 283.050 439.050 ;
        RECT 289.950 438.600 292.050 439.050 ;
        RECT 280.950 437.400 292.050 438.600 ;
        RECT 280.950 436.950 283.050 437.400 ;
        RECT 289.950 436.950 292.050 437.400 ;
        RECT 364.950 438.600 367.050 439.050 ;
        RECT 421.950 438.600 424.050 439.050 ;
        RECT 364.950 437.400 424.050 438.600 ;
        RECT 364.950 436.950 367.050 437.400 ;
        RECT 421.950 436.950 424.050 437.400 ;
        RECT 484.950 438.600 487.050 439.050 ;
        RECT 493.950 438.600 496.050 439.050 ;
        RECT 484.950 437.400 496.050 438.600 ;
        RECT 484.950 436.950 487.050 437.400 ;
        RECT 493.950 436.950 496.050 437.400 ;
        RECT 535.950 438.600 538.050 439.050 ;
        RECT 550.950 438.600 553.050 439.050 ;
        RECT 535.950 437.400 553.050 438.600 ;
        RECT 535.950 436.950 538.050 437.400 ;
        RECT 550.950 436.950 553.050 437.400 ;
        RECT 559.950 438.600 562.050 439.050 ;
        RECT 586.950 438.600 589.050 439.050 ;
        RECT 559.950 437.400 589.050 438.600 ;
        RECT 559.950 436.950 562.050 437.400 ;
        RECT 586.950 436.950 589.050 437.400 ;
        RECT 610.950 438.600 613.050 439.050 ;
        RECT 622.950 438.600 625.050 439.050 ;
        RECT 610.950 437.400 625.050 438.600 ;
        RECT 610.950 436.950 613.050 437.400 ;
        RECT 622.950 436.950 625.050 437.400 ;
        RECT 745.950 438.600 748.050 439.050 ;
        RECT 808.950 438.600 811.050 439.050 ;
        RECT 745.950 437.400 811.050 438.600 ;
        RECT 745.950 436.950 748.050 437.400 ;
        RECT 808.950 436.950 811.050 437.400 ;
        RECT 922.950 438.600 925.050 439.050 ;
        RECT 928.800 438.600 930.900 439.050 ;
        RECT 922.950 437.400 930.900 438.600 ;
        RECT 922.950 436.950 925.050 437.400 ;
        RECT 928.800 436.950 930.900 437.400 ;
        RECT 931.950 438.600 934.050 439.050 ;
        RECT 973.950 438.600 976.050 439.050 ;
        RECT 979.950 438.600 982.050 439.050 ;
        RECT 931.950 437.400 963.600 438.600 ;
        RECT 931.950 436.950 934.050 437.400 ;
        RECT 31.950 435.600 34.050 436.050 ;
        RECT 67.950 435.600 70.050 436.050 ;
        RECT 31.950 434.400 70.050 435.600 ;
        RECT 31.950 433.950 34.050 434.400 ;
        RECT 67.950 433.950 70.050 434.400 ;
        RECT 175.950 435.600 178.050 436.050 ;
        RECT 193.950 435.600 196.050 436.050 ;
        RECT 175.950 434.400 196.050 435.600 ;
        RECT 175.950 433.950 178.050 434.400 ;
        RECT 193.950 433.950 196.050 434.400 ;
        RECT 235.950 435.600 238.050 436.050 ;
        RECT 268.950 435.600 271.050 436.050 ;
        RECT 235.950 434.400 271.050 435.600 ;
        RECT 235.950 433.950 238.050 434.400 ;
        RECT 268.950 433.950 271.050 434.400 ;
        RECT 337.950 435.600 340.050 436.050 ;
        RECT 385.950 435.600 388.050 436.050 ;
        RECT 337.950 434.400 388.050 435.600 ;
        RECT 337.950 433.950 340.050 434.400 ;
        RECT 385.950 433.950 388.050 434.400 ;
        RECT 442.950 435.600 445.050 436.050 ;
        RECT 517.950 435.600 520.050 436.050 ;
        RECT 595.950 435.600 598.050 436.050 ;
        RECT 442.950 434.400 520.050 435.600 ;
        RECT 442.950 433.950 445.050 434.400 ;
        RECT 517.950 433.950 520.050 434.400 ;
        RECT 590.400 434.400 598.050 435.600 ;
        RECT 154.950 432.600 157.050 433.050 ;
        RECT 196.950 432.600 199.050 433.050 ;
        RECT 154.950 431.400 199.050 432.600 ;
        RECT 154.950 430.950 157.050 431.400 ;
        RECT 196.950 430.950 199.050 431.400 ;
        RECT 202.950 432.600 205.050 433.050 ;
        RECT 208.950 432.600 211.050 433.050 ;
        RECT 202.950 431.400 211.050 432.600 ;
        RECT 202.950 430.950 205.050 431.400 ;
        RECT 208.950 430.950 211.050 431.400 ;
        RECT 238.950 432.600 241.050 433.050 ;
        RECT 250.800 432.600 252.900 433.050 ;
        RECT 238.950 431.400 252.900 432.600 ;
        RECT 238.950 430.950 241.050 431.400 ;
        RECT 250.800 430.950 252.900 431.400 ;
        RECT 253.950 432.600 256.050 433.050 ;
        RECT 316.950 432.600 319.050 433.050 ;
        RECT 253.950 431.400 319.050 432.600 ;
        RECT 253.950 430.950 256.050 431.400 ;
        RECT 316.950 430.950 319.050 431.400 ;
        RECT 445.950 432.600 448.050 433.050 ;
        RECT 559.950 432.600 562.050 433.050 ;
        RECT 445.950 431.400 562.050 432.600 ;
        RECT 445.950 430.950 448.050 431.400 ;
        RECT 559.950 430.950 562.050 431.400 ;
        RECT 580.950 432.600 583.050 433.050 ;
        RECT 590.400 432.600 591.600 434.400 ;
        RECT 595.950 433.950 598.050 434.400 ;
        RECT 640.950 435.600 643.050 436.050 ;
        RECT 673.950 435.600 676.050 436.050 ;
        RECT 811.950 435.600 814.050 436.050 ;
        RECT 814.950 435.600 817.050 436.050 ;
        RECT 640.950 434.400 672.600 435.600 ;
        RECT 640.950 433.950 643.050 434.400 ;
        RECT 580.950 431.400 591.600 432.600 ;
        RECT 671.400 432.600 672.600 434.400 ;
        RECT 673.950 434.400 817.050 435.600 ;
        RECT 673.950 433.950 676.050 434.400 ;
        RECT 811.950 433.950 814.050 434.400 ;
        RECT 814.950 433.950 817.050 434.400 ;
        RECT 910.950 435.600 913.050 436.050 ;
        RECT 919.950 435.600 922.050 436.050 ;
        RECT 910.950 434.400 922.050 435.600 ;
        RECT 910.950 433.950 913.050 434.400 ;
        RECT 919.950 433.950 922.050 434.400 ;
        RECT 943.950 435.600 946.050 436.050 ;
        RECT 952.950 435.600 955.050 436.050 ;
        RECT 958.950 435.600 961.050 436.050 ;
        RECT 943.950 434.400 961.050 435.600 ;
        RECT 962.400 435.600 963.600 437.400 ;
        RECT 973.950 437.400 982.050 438.600 ;
        RECT 973.950 436.950 976.050 437.400 ;
        RECT 979.950 436.950 982.050 437.400 ;
        RECT 967.950 435.600 970.050 436.050 ;
        RECT 962.400 434.400 970.050 435.600 ;
        RECT 943.950 433.950 946.050 434.400 ;
        RECT 952.950 433.950 955.050 434.400 ;
        RECT 958.950 433.950 961.050 434.400 ;
        RECT 967.950 433.950 970.050 434.400 ;
        RECT 979.950 435.600 982.050 435.900 ;
        RECT 1000.950 435.600 1003.050 436.050 ;
        RECT 979.950 434.400 1003.050 435.600 ;
        RECT 979.950 433.800 982.050 434.400 ;
        RECT 1000.950 433.950 1003.050 434.400 ;
        RECT 703.950 432.600 706.050 433.050 ;
        RECT 671.400 431.400 706.050 432.600 ;
        RECT 580.950 430.950 583.050 431.400 ;
        RECT 703.950 430.950 706.050 431.400 ;
        RECT 838.950 432.600 841.050 433.050 ;
        RECT 847.950 432.600 850.050 433.050 ;
        RECT 853.950 432.600 856.050 433.050 ;
        RECT 838.950 431.400 856.050 432.600 ;
        RECT 838.950 430.950 841.050 431.400 ;
        RECT 847.950 430.950 850.050 431.400 ;
        RECT 853.950 430.950 856.050 431.400 ;
        RECT 859.950 432.600 862.050 433.050 ;
        RECT 892.950 432.600 895.050 433.050 ;
        RECT 859.950 431.400 895.050 432.600 ;
        RECT 859.950 430.950 862.050 431.400 ;
        RECT 892.950 430.950 895.050 431.400 ;
        RECT 19.950 429.600 22.050 430.050 ;
        RECT 46.950 429.600 49.050 430.050 ;
        RECT 85.950 429.600 88.050 430.050 ;
        RECT 19.950 428.400 88.050 429.600 ;
        RECT 19.950 427.950 22.050 428.400 ;
        RECT 46.950 427.950 49.050 428.400 ;
        RECT 85.950 427.950 88.050 428.400 ;
        RECT 115.950 429.600 118.050 430.050 ;
        RECT 124.950 429.600 127.050 430.050 ;
        RECT 115.950 428.400 127.050 429.600 ;
        RECT 115.950 427.950 118.050 428.400 ;
        RECT 124.950 427.950 127.050 428.400 ;
        RECT 166.950 429.600 169.050 430.050 ;
        RECT 214.950 429.600 217.050 430.050 ;
        RECT 265.950 429.600 268.050 430.050 ;
        RECT 298.950 429.600 301.050 430.050 ;
        RECT 166.950 428.400 301.050 429.600 ;
        RECT 166.950 427.950 169.050 428.400 ;
        RECT 214.950 427.950 217.050 428.400 ;
        RECT 265.950 427.950 268.050 428.400 ;
        RECT 298.950 427.950 301.050 428.400 ;
        RECT 379.950 429.600 382.050 430.050 ;
        RECT 487.950 429.600 490.050 430.050 ;
        RECT 379.950 428.400 490.050 429.600 ;
        RECT 379.950 427.950 382.050 428.400 ;
        RECT 487.950 427.950 490.050 428.400 ;
        RECT 583.950 429.600 586.050 430.050 ;
        RECT 592.950 429.600 595.050 430.050 ;
        RECT 583.950 428.400 595.050 429.600 ;
        RECT 583.950 427.950 586.050 428.400 ;
        RECT 592.950 427.950 595.050 428.400 ;
        RECT 613.950 429.600 616.050 430.050 ;
        RECT 640.950 429.600 643.050 430.050 ;
        RECT 613.950 428.400 643.050 429.600 ;
        RECT 613.950 427.950 616.050 428.400 ;
        RECT 640.950 427.950 643.050 428.400 ;
        RECT 694.950 429.600 697.050 430.050 ;
        RECT 703.950 429.600 706.050 429.900 ;
        RECT 694.950 428.400 706.050 429.600 ;
        RECT 694.950 427.950 697.050 428.400 ;
        RECT 703.950 427.800 706.050 428.400 ;
        RECT 736.950 429.600 739.050 430.050 ;
        RECT 769.950 429.600 772.050 430.050 ;
        RECT 736.950 428.400 772.050 429.600 ;
        RECT 736.950 427.950 739.050 428.400 ;
        RECT 769.950 427.950 772.050 428.400 ;
        RECT 820.950 429.600 823.050 430.050 ;
        RECT 865.950 429.600 868.050 430.050 ;
        RECT 874.950 429.600 877.050 430.050 ;
        RECT 820.950 428.400 877.050 429.600 ;
        RECT 820.950 427.950 823.050 428.400 ;
        RECT 865.950 427.950 868.050 428.400 ;
        RECT 874.950 427.950 877.050 428.400 ;
        RECT 883.950 429.600 886.050 430.050 ;
        RECT 919.950 429.600 922.050 430.050 ;
        RECT 883.950 428.400 922.050 429.600 ;
        RECT 883.950 427.950 886.050 428.400 ;
        RECT 919.950 427.950 922.050 428.400 ;
        RECT 970.950 429.600 973.050 430.050 ;
        RECT 985.950 429.600 988.050 430.050 ;
        RECT 994.950 429.600 997.050 430.050 ;
        RECT 970.950 428.400 997.050 429.600 ;
        RECT 970.950 427.950 973.050 428.400 ;
        RECT 985.950 427.950 988.050 428.400 ;
        RECT 994.950 427.950 997.050 428.400 ;
        RECT 148.950 426.600 151.050 427.050 ;
        RECT 175.800 426.600 177.900 427.050 ;
        RECT 148.950 425.400 177.900 426.600 ;
        RECT 148.950 424.950 151.050 425.400 ;
        RECT 175.800 424.950 177.900 425.400 ;
        RECT 178.950 426.600 181.050 427.050 ;
        RECT 223.950 426.600 226.050 427.050 ;
        RECT 178.950 425.400 226.050 426.600 ;
        RECT 178.950 424.950 181.050 425.400 ;
        RECT 223.950 424.950 226.050 425.400 ;
        RECT 373.950 426.600 376.050 427.050 ;
        RECT 445.950 426.600 448.050 427.050 ;
        RECT 373.950 425.400 448.050 426.600 ;
        RECT 373.950 424.950 376.050 425.400 ;
        RECT 445.950 424.950 448.050 425.400 ;
        RECT 526.950 426.600 529.050 427.050 ;
        RECT 604.950 426.600 607.050 427.050 ;
        RECT 526.950 425.400 607.050 426.600 ;
        RECT 526.950 424.950 529.050 425.400 ;
        RECT 604.950 424.950 607.050 425.400 ;
        RECT 784.950 426.600 787.050 427.050 ;
        RECT 835.950 426.600 838.050 427.050 ;
        RECT 868.950 426.600 871.050 427.050 ;
        RECT 784.950 425.400 871.050 426.600 ;
        RECT 784.950 424.950 787.050 425.400 ;
        RECT 835.950 424.950 838.050 425.400 ;
        RECT 868.950 424.950 871.050 425.400 ;
        RECT 937.950 426.600 940.050 427.050 ;
        RECT 991.950 426.600 994.050 427.050 ;
        RECT 937.950 425.400 994.050 426.600 ;
        RECT 937.950 424.950 940.050 425.400 ;
        RECT 991.950 424.950 994.050 425.400 ;
        RECT 76.950 423.600 79.050 424.050 ;
        RECT 94.950 423.600 97.050 424.050 ;
        RECT 76.950 422.400 97.050 423.600 ;
        RECT 76.950 421.950 79.050 422.400 ;
        RECT 94.950 421.950 97.050 422.400 ;
        RECT 136.950 423.600 139.050 424.050 ;
        RECT 229.950 423.600 232.050 424.050 ;
        RECT 271.950 423.600 274.050 424.050 ;
        RECT 304.950 423.600 307.050 424.050 ;
        RECT 328.950 423.600 331.050 424.050 ;
        RECT 418.950 423.600 421.050 424.050 ;
        RECT 430.950 423.600 433.050 424.050 ;
        RECT 136.950 422.400 433.050 423.600 ;
        RECT 136.950 421.950 139.050 422.400 ;
        RECT 229.950 421.950 232.050 422.400 ;
        RECT 271.950 421.950 274.050 422.400 ;
        RECT 304.950 421.950 307.050 422.400 ;
        RECT 328.950 421.950 331.050 422.400 ;
        RECT 418.950 421.950 421.050 422.400 ;
        RECT 430.950 421.950 433.050 422.400 ;
        RECT 463.950 423.600 466.050 424.050 ;
        RECT 469.950 423.600 472.050 424.050 ;
        RECT 496.950 423.600 499.050 424.050 ;
        RECT 463.950 422.400 499.050 423.600 ;
        RECT 463.950 421.950 466.050 422.400 ;
        RECT 469.950 421.950 472.050 422.400 ;
        RECT 496.950 421.950 499.050 422.400 ;
        RECT 571.950 423.600 574.050 424.050 ;
        RECT 613.950 423.600 616.050 424.050 ;
        RECT 571.950 422.400 616.050 423.600 ;
        RECT 571.950 421.950 574.050 422.400 ;
        RECT 613.950 421.950 616.050 422.400 ;
        RECT 907.950 423.600 910.050 424.050 ;
        RECT 913.950 423.600 916.050 424.050 ;
        RECT 907.950 422.400 916.050 423.600 ;
        RECT 907.950 421.950 910.050 422.400 ;
        RECT 913.950 421.950 916.050 422.400 ;
        RECT 973.950 423.600 976.050 424.050 ;
        RECT 988.950 423.600 991.050 424.050 ;
        RECT 973.950 422.400 991.050 423.600 ;
        RECT 973.950 421.950 976.050 422.400 ;
        RECT 988.950 421.950 991.050 422.400 ;
        RECT 343.950 420.600 346.050 421.050 ;
        RECT 373.950 420.600 376.050 421.050 ;
        RECT 394.950 420.600 397.050 421.050 ;
        RECT 343.950 419.400 397.050 420.600 ;
        RECT 343.950 418.950 346.050 419.400 ;
        RECT 373.950 418.950 376.050 419.400 ;
        RECT 394.950 418.950 397.050 419.400 ;
        RECT 541.950 420.600 544.050 421.050 ;
        RECT 556.950 420.600 559.050 421.050 ;
        RECT 541.950 419.400 559.050 420.600 ;
        RECT 541.950 418.950 544.050 419.400 ;
        RECT 556.950 418.950 559.050 419.400 ;
        RECT 598.950 420.600 601.050 421.050 ;
        RECT 604.950 420.600 607.050 421.050 ;
        RECT 598.950 419.400 607.050 420.600 ;
        RECT 598.950 418.950 601.050 419.400 ;
        RECT 604.950 418.950 607.050 419.400 ;
        RECT 898.950 420.600 901.050 421.050 ;
        RECT 922.950 420.600 925.050 421.050 ;
        RECT 898.950 419.400 925.050 420.600 ;
        RECT 898.950 418.950 901.050 419.400 ;
        RECT 922.950 418.950 925.050 419.400 ;
        RECT 928.950 420.600 931.050 421.050 ;
        RECT 970.950 420.600 973.050 421.050 ;
        RECT 928.950 419.400 973.050 420.600 ;
        RECT 928.950 418.950 931.050 419.400 ;
        RECT 970.950 418.950 973.050 419.400 ;
        RECT 31.950 417.600 34.050 418.200 ;
        RECT 58.950 417.750 61.050 418.200 ;
        RECT 67.950 417.750 70.050 418.200 ;
        RECT 31.950 416.400 54.600 417.600 ;
        RECT 31.950 416.100 34.050 416.400 ;
        RECT 53.400 412.050 54.600 416.400 ;
        RECT 58.950 416.550 70.050 417.750 ;
        RECT 58.950 416.100 61.050 416.550 ;
        RECT 67.950 416.100 70.050 416.550 ;
        RECT 73.950 417.600 76.050 418.050 ;
        RECT 91.950 417.600 94.050 418.200 ;
        RECT 73.950 416.400 94.050 417.600 ;
        RECT 73.950 415.950 76.050 416.400 ;
        RECT 91.950 416.100 94.050 416.400 ;
        RECT 127.950 417.750 130.050 418.200 ;
        RECT 133.950 417.750 136.050 418.200 ;
        RECT 127.950 416.550 136.050 417.750 ;
        RECT 127.950 416.100 130.050 416.550 ;
        RECT 133.950 416.100 136.050 416.550 ;
        RECT 139.950 417.600 142.050 418.050 ;
        RECT 151.950 417.600 154.050 418.200 ;
        RECT 139.950 416.400 154.050 417.600 ;
        RECT 139.950 415.950 142.050 416.400 ;
        RECT 151.950 416.100 154.050 416.400 ;
        RECT 157.950 416.100 160.050 418.200 ;
        RECT 241.950 417.750 244.050 418.200 ;
        RECT 247.950 417.750 250.050 418.200 ;
        RECT 241.950 416.550 250.050 417.750 ;
        RECT 241.950 416.100 244.050 416.550 ;
        RECT 247.950 416.100 250.050 416.550 ;
        RECT 253.950 417.600 256.050 418.200 ;
        RECT 262.950 417.600 265.050 418.050 ;
        RECT 253.950 416.400 265.050 417.600 ;
        RECT 253.950 416.100 256.050 416.400 ;
        RECT 52.950 409.950 55.050 412.050 ;
        RECT 88.950 411.450 91.050 411.900 ;
        RECT 115.950 411.450 118.050 411.900 ;
        RECT 88.950 410.250 118.050 411.450 ;
        RECT 88.950 409.800 91.050 410.250 ;
        RECT 115.950 409.800 118.050 410.250 ;
        RECT 133.950 411.450 136.050 411.900 ;
        RECT 148.950 411.450 151.050 411.900 ;
        RECT 133.950 410.250 151.050 411.450 ;
        RECT 158.400 411.600 159.600 416.100 ;
        RECT 262.950 415.950 265.050 416.400 ;
        RECT 277.950 417.600 280.050 418.200 ;
        RECT 286.950 417.600 289.050 418.050 ;
        RECT 277.950 416.400 289.050 417.600 ;
        RECT 277.950 416.100 280.050 416.400 ;
        RECT 286.950 415.950 289.050 416.400 ;
        RECT 292.950 417.600 295.050 418.050 ;
        RECT 328.950 417.750 331.050 418.200 ;
        RECT 337.950 417.750 340.050 418.200 ;
        RECT 328.950 417.600 340.050 417.750 ;
        RECT 292.950 416.550 340.050 417.600 ;
        RECT 292.950 416.400 331.050 416.550 ;
        RECT 292.950 415.950 295.050 416.400 ;
        RECT 328.950 416.100 331.050 416.400 ;
        RECT 337.950 416.100 340.050 416.550 ;
        RECT 403.950 417.600 406.050 418.050 ;
        RECT 457.950 417.750 460.050 418.200 ;
        RECT 472.950 417.750 475.050 418.200 ;
        RECT 403.950 416.400 423.600 417.600 ;
        RECT 403.950 415.950 406.050 416.400 ;
        RECT 422.400 414.600 423.600 416.400 ;
        RECT 446.400 416.400 453.600 417.600 ;
        RECT 446.400 414.600 447.600 416.400 ;
        RECT 422.400 413.400 447.600 414.600 ;
        RECT 160.950 411.600 163.050 412.050 ;
        RECT 181.950 411.600 184.050 411.900 ;
        RECT 158.400 410.400 184.050 411.600 ;
        RECT 133.950 409.800 136.050 410.250 ;
        RECT 148.950 409.800 151.050 410.250 ;
        RECT 160.950 409.950 163.050 410.400 ;
        RECT 181.950 409.800 184.050 410.400 ;
        RECT 193.950 411.450 196.050 411.900 ;
        RECT 205.950 411.450 208.050 411.900 ;
        RECT 193.950 410.250 208.050 411.450 ;
        RECT 193.950 409.800 196.050 410.250 ;
        RECT 205.950 409.800 208.050 410.250 ;
        RECT 214.950 411.450 217.050 411.900 ;
        RECT 226.950 411.450 229.050 411.900 ;
        RECT 214.950 410.250 229.050 411.450 ;
        RECT 214.950 409.800 217.050 410.250 ;
        RECT 226.950 409.800 229.050 410.250 ;
        RECT 238.950 411.450 241.050 411.900 ;
        RECT 250.950 411.450 253.050 411.900 ;
        RECT 238.950 410.250 253.050 411.450 ;
        RECT 238.950 409.800 241.050 410.250 ;
        RECT 250.950 409.800 253.050 410.250 ;
        RECT 265.950 411.450 268.050 411.900 ;
        RECT 274.950 411.450 277.050 411.900 ;
        RECT 265.950 410.250 277.050 411.450 ;
        RECT 265.950 409.800 268.050 410.250 ;
        RECT 274.950 409.800 277.050 410.250 ;
        RECT 280.950 411.450 283.050 411.900 ;
        RECT 292.950 411.450 295.050 411.900 ;
        RECT 280.950 410.250 295.050 411.450 ;
        RECT 280.950 409.800 283.050 410.250 ;
        RECT 292.950 409.800 295.050 410.250 ;
        RECT 418.950 411.450 421.050 411.900 ;
        RECT 448.950 411.450 451.050 411.900 ;
        RECT 418.950 410.250 451.050 411.450 ;
        RECT 452.400 411.600 453.600 416.400 ;
        RECT 457.950 416.550 475.050 417.750 ;
        RECT 457.950 416.100 460.050 416.550 ;
        RECT 472.950 416.100 475.050 416.550 ;
        RECT 481.950 417.600 484.050 418.200 ;
        RECT 505.950 417.750 508.050 418.200 ;
        RECT 517.950 417.750 520.050 418.200 ;
        RECT 505.950 417.600 520.050 417.750 ;
        RECT 481.950 416.550 520.050 417.600 ;
        RECT 481.950 416.400 508.050 416.550 ;
        RECT 481.950 416.100 484.050 416.400 ;
        RECT 505.950 416.100 508.050 416.400 ;
        RECT 517.950 416.100 520.050 416.550 ;
        RECT 547.950 417.750 550.050 418.200 ;
        RECT 553.950 417.750 556.050 418.200 ;
        RECT 547.950 416.550 556.050 417.750 ;
        RECT 565.950 417.600 568.050 418.200 ;
        RECT 571.950 417.600 574.050 418.200 ;
        RECT 547.950 416.100 550.050 416.550 ;
        RECT 553.950 416.100 556.050 416.550 ;
        RECT 560.400 416.400 574.050 417.600 ;
        RECT 560.400 415.050 561.600 416.400 ;
        RECT 565.950 416.100 568.050 416.400 ;
        RECT 571.950 416.100 574.050 416.400 ;
        RECT 558.000 414.900 561.600 415.050 ;
        RECT 556.950 413.400 561.600 414.900 ;
        RECT 586.950 414.600 589.050 418.050 ;
        RECT 619.950 417.600 622.050 418.200 ;
        RECT 631.950 417.600 634.050 418.050 ;
        RECT 619.950 416.400 634.050 417.600 ;
        RECT 619.950 416.100 622.050 416.400 ;
        RECT 631.950 415.950 634.050 416.400 ;
        RECT 646.950 417.750 649.050 418.200 ;
        RECT 652.950 417.750 655.050 417.900 ;
        RECT 646.950 416.550 655.050 417.750 ;
        RECT 646.950 416.100 649.050 416.550 ;
        RECT 652.950 415.800 655.050 416.550 ;
        RECT 664.950 417.600 667.050 418.200 ;
        RECT 805.950 417.600 808.050 418.200 ;
        RECT 814.950 417.600 817.050 418.050 ;
        RECT 664.950 416.400 672.600 417.600 ;
        RECT 664.950 416.100 667.050 416.400 ;
        RECT 586.950 414.000 597.600 414.600 ;
        RECT 587.400 413.400 597.600 414.000 ;
        RECT 556.950 412.950 561.000 413.400 ;
        RECT 556.950 412.800 559.050 412.950 ;
        RECT 454.950 411.600 457.050 411.900 ;
        RECT 475.950 411.600 478.050 411.900 ;
        RECT 452.400 410.400 457.050 411.600 ;
        RECT 418.950 409.800 421.050 410.250 ;
        RECT 448.950 409.800 451.050 410.250 ;
        RECT 454.950 409.800 457.050 410.400 ;
        RECT 458.400 410.400 478.050 411.600 ;
        RECT 31.950 408.600 34.050 409.050 ;
        RECT 49.950 408.600 52.050 409.050 ;
        RECT 31.950 407.400 52.050 408.600 ;
        RECT 31.950 406.950 34.050 407.400 ;
        RECT 49.950 406.950 52.050 407.400 ;
        RECT 73.950 405.600 76.050 406.050 ;
        RECT 109.950 405.600 112.050 409.050 ;
        RECT 298.950 408.600 301.050 409.050 ;
        RECT 310.950 408.600 313.050 409.050 ;
        RECT 346.950 408.600 349.050 409.050 ;
        RECT 298.950 407.400 349.050 408.600 ;
        RECT 298.950 406.950 301.050 407.400 ;
        RECT 310.950 406.950 313.050 407.400 ;
        RECT 346.950 406.950 349.050 407.400 ;
        RECT 379.950 408.600 382.050 409.050 ;
        RECT 458.400 408.600 459.600 410.400 ;
        RECT 475.950 409.800 478.050 410.400 ;
        RECT 493.950 411.600 496.050 412.050 ;
        RECT 502.950 411.600 505.050 411.900 ;
        RECT 553.950 411.600 556.050 412.050 ;
        RECT 589.950 411.600 592.050 411.900 ;
        RECT 493.950 410.400 556.050 411.600 ;
        RECT 560.400 411.000 592.050 411.600 ;
        RECT 493.950 409.950 496.050 410.400 ;
        RECT 502.950 409.800 505.050 410.400 ;
        RECT 553.950 409.950 556.050 410.400 ;
        RECT 559.950 410.400 592.050 411.000 ;
        RECT 379.950 407.400 459.600 408.600 ;
        RECT 508.950 408.600 511.050 409.050 ;
        RECT 517.950 408.600 520.050 409.050 ;
        RECT 508.950 407.400 520.050 408.600 ;
        RECT 379.950 406.950 382.050 407.400 ;
        RECT 508.950 406.950 511.050 407.400 ;
        RECT 517.950 406.950 520.050 407.400 ;
        RECT 535.950 408.600 538.050 409.050 ;
        RECT 550.950 408.600 553.050 409.050 ;
        RECT 535.950 407.400 553.050 408.600 ;
        RECT 535.950 406.950 538.050 407.400 ;
        RECT 550.950 406.950 553.050 407.400 ;
        RECT 559.950 406.950 562.050 410.400 ;
        RECT 589.950 409.800 592.050 410.400 ;
        RECT 596.400 408.600 597.600 413.400 ;
        RECT 671.400 412.050 672.600 416.400 ;
        RECT 805.950 416.400 817.050 417.600 ;
        RECT 805.950 416.100 808.050 416.400 ;
        RECT 814.950 415.950 817.050 416.400 ;
        RECT 820.950 417.750 823.050 418.200 ;
        RECT 826.950 417.750 829.050 418.200 ;
        RECT 820.950 416.550 829.050 417.750 ;
        RECT 820.950 416.100 823.050 416.550 ;
        RECT 826.950 416.100 829.050 416.550 ;
        RECT 841.950 417.750 844.050 418.200 ;
        RECT 853.950 417.750 856.050 418.200 ;
        RECT 841.950 416.550 856.050 417.750 ;
        RECT 841.950 416.100 844.050 416.550 ;
        RECT 853.950 416.100 856.050 416.550 ;
        RECT 880.950 417.600 883.050 418.200 ;
        RECT 904.950 417.600 907.050 418.200 ;
        RECT 916.950 417.600 919.050 418.050 ;
        RECT 880.950 416.400 897.600 417.600 ;
        RECT 880.950 416.100 883.050 416.400 ;
        RECT 896.400 412.050 897.600 416.400 ;
        RECT 904.950 416.400 919.050 417.600 ;
        RECT 904.950 416.100 907.050 416.400 ;
        RECT 916.950 415.950 919.050 416.400 ;
        RECT 973.950 417.600 976.050 418.200 ;
        RECT 973.950 416.400 996.600 417.600 ;
        RECT 973.950 416.100 976.050 416.400 ;
        RECT 937.950 414.600 940.050 415.050 ;
        RECT 937.950 413.400 951.600 414.600 ;
        RECT 937.950 412.950 940.050 413.400 ;
        RECT 598.950 411.450 601.050 411.900 ;
        RECT 604.950 411.450 607.050 411.900 ;
        RECT 598.950 410.250 607.050 411.450 ;
        RECT 598.950 409.800 601.050 410.250 ;
        RECT 604.950 409.800 607.050 410.250 ;
        RECT 631.950 411.450 634.050 411.900 ;
        RECT 637.950 411.450 640.050 411.900 ;
        RECT 631.950 410.250 640.050 411.450 ;
        RECT 631.950 409.800 634.050 410.250 ;
        RECT 637.950 409.800 640.050 410.250 ;
        RECT 670.950 409.950 673.050 412.050 ;
        RECT 703.950 411.600 706.050 412.050 ;
        RECT 742.950 411.600 745.050 411.900 ;
        RECT 703.950 410.400 745.050 411.600 ;
        RECT 703.950 409.950 706.050 410.400 ;
        RECT 742.950 409.800 745.050 410.400 ;
        RECT 766.950 411.600 769.050 411.900 ;
        RECT 781.950 411.600 784.050 411.900 ;
        RECT 802.950 411.600 805.050 411.900 ;
        RECT 766.950 410.400 805.050 411.600 ;
        RECT 766.950 409.800 769.050 410.400 ;
        RECT 781.950 409.800 784.050 410.400 ;
        RECT 802.950 409.800 805.050 410.400 ;
        RECT 835.950 411.450 838.050 411.900 ;
        RECT 850.950 411.450 853.050 411.900 ;
        RECT 835.950 410.250 853.050 411.450 ;
        RECT 835.950 409.800 838.050 410.250 ;
        RECT 850.950 409.800 853.050 410.250 ;
        RECT 856.950 411.450 859.050 411.900 ;
        RECT 865.950 411.450 868.050 411.900 ;
        RECT 856.950 410.250 868.050 411.450 ;
        RECT 856.950 409.800 859.050 410.250 ;
        RECT 865.950 409.800 868.050 410.250 ;
        RECT 895.950 409.950 898.050 412.050 ;
        RECT 950.400 411.900 951.600 413.400 ;
        RECT 913.950 411.450 916.050 411.900 ;
        RECT 925.950 411.450 928.050 411.900 ;
        RECT 913.950 410.250 928.050 411.450 ;
        RECT 913.950 409.800 916.050 410.250 ;
        RECT 925.950 409.800 928.050 410.250 ;
        RECT 949.950 409.800 952.050 411.900 ;
        RECT 958.950 411.600 961.050 412.050 ;
        RECT 964.950 411.600 967.050 412.050 ;
        RECT 958.950 410.400 967.050 411.600 ;
        RECT 958.950 409.950 961.050 410.400 ;
        RECT 964.950 409.950 967.050 410.400 ;
        RECT 970.950 411.600 973.050 411.900 ;
        RECT 991.950 411.600 994.050 411.900 ;
        RECT 970.950 410.400 994.050 411.600 ;
        RECT 995.400 411.600 996.600 416.400 ;
        RECT 1000.950 411.600 1003.050 412.050 ;
        RECT 995.400 410.400 1003.050 411.600 ;
        RECT 970.950 409.800 973.050 410.400 ;
        RECT 991.950 409.800 994.050 410.400 ;
        RECT 1000.950 409.950 1003.050 410.400 ;
        RECT 616.950 408.600 619.050 409.050 ;
        RECT 596.400 407.400 619.050 408.600 ;
        RECT 616.950 406.950 619.050 407.400 ;
        RECT 667.950 408.600 670.050 409.050 ;
        RECT 706.950 408.600 709.050 409.050 ;
        RECT 712.950 408.600 715.050 409.050 ;
        RECT 667.950 407.400 684.600 408.600 ;
        RECT 667.950 406.950 670.050 407.400 ;
        RECT 683.400 406.050 684.600 407.400 ;
        RECT 706.950 407.400 715.050 408.600 ;
        RECT 706.950 406.950 709.050 407.400 ;
        RECT 712.950 406.950 715.050 407.400 ;
        RECT 730.950 408.600 733.050 409.050 ;
        RECT 739.950 408.600 742.050 409.050 ;
        RECT 730.950 407.400 742.050 408.600 ;
        RECT 730.950 406.950 733.050 407.400 ;
        RECT 739.950 406.950 742.050 407.400 ;
        RECT 886.950 408.600 889.050 409.050 ;
        RECT 892.950 408.600 895.050 409.050 ;
        RECT 886.950 407.400 895.050 408.600 ;
        RECT 886.950 406.950 889.050 407.400 ;
        RECT 892.950 406.950 895.050 407.400 ;
        RECT 907.950 408.600 910.050 409.050 ;
        RECT 934.950 408.600 937.050 409.050 ;
        RECT 940.950 408.600 943.050 409.050 ;
        RECT 907.950 407.400 943.050 408.600 ;
        RECT 907.950 406.950 910.050 407.400 ;
        RECT 934.950 406.950 937.050 407.400 ;
        RECT 940.950 406.950 943.050 407.400 ;
        RECT 73.950 405.000 112.050 405.600 ;
        RECT 136.950 405.600 139.050 406.050 ;
        RECT 241.950 405.600 244.050 406.050 ;
        RECT 73.950 404.400 111.600 405.000 ;
        RECT 136.950 404.400 244.050 405.600 ;
        RECT 73.950 403.950 76.050 404.400 ;
        RECT 136.950 403.950 139.050 404.400 ;
        RECT 241.950 403.950 244.050 404.400 ;
        RECT 256.950 405.600 259.050 406.050 ;
        RECT 286.950 405.600 289.050 406.050 ;
        RECT 256.950 404.400 289.050 405.600 ;
        RECT 256.950 403.950 259.050 404.400 ;
        RECT 286.950 403.950 289.050 404.400 ;
        RECT 295.950 405.600 298.050 405.900 ;
        RECT 322.950 405.600 325.050 406.050 ;
        RECT 295.950 404.400 325.050 405.600 ;
        RECT 295.950 403.800 298.050 404.400 ;
        RECT 322.950 403.950 325.050 404.400 ;
        RECT 472.950 405.600 475.050 406.050 ;
        RECT 556.950 405.600 559.050 406.050 ;
        RECT 472.950 404.400 559.050 405.600 ;
        RECT 472.950 403.950 475.050 404.400 ;
        RECT 556.950 403.950 559.050 404.400 ;
        RECT 622.950 405.600 625.050 406.050 ;
        RECT 652.950 405.600 655.050 406.050 ;
        RECT 622.950 404.400 655.050 405.600 ;
        RECT 622.950 403.950 625.050 404.400 ;
        RECT 652.950 403.950 655.050 404.400 ;
        RECT 667.950 405.600 670.050 405.900 ;
        RECT 673.950 405.600 676.050 406.050 ;
        RECT 667.950 404.400 676.050 405.600 ;
        RECT 667.950 403.800 670.050 404.400 ;
        RECT 673.950 403.950 676.050 404.400 ;
        RECT 682.950 405.600 685.050 406.050 ;
        RECT 694.950 405.600 697.050 406.050 ;
        RECT 682.950 404.400 697.050 405.600 ;
        RECT 682.950 403.950 685.050 404.400 ;
        RECT 694.950 403.950 697.050 404.400 ;
        RECT 829.950 405.600 832.050 406.050 ;
        RECT 841.950 405.600 844.050 406.050 ;
        RECT 877.950 405.600 880.050 406.050 ;
        RECT 829.950 404.400 880.050 405.600 ;
        RECT 829.950 403.950 832.050 404.400 ;
        RECT 841.950 403.950 844.050 404.400 ;
        RECT 877.950 403.950 880.050 404.400 ;
        RECT 919.950 405.600 922.050 406.050 ;
        RECT 952.950 405.600 955.050 406.050 ;
        RECT 919.950 404.400 955.050 405.600 ;
        RECT 919.950 403.950 922.050 404.400 ;
        RECT 952.950 403.950 955.050 404.400 ;
        RECT 997.950 405.600 1000.050 406.050 ;
        RECT 1006.950 405.600 1009.050 406.050 ;
        RECT 997.950 404.400 1009.050 405.600 ;
        RECT 997.950 403.950 1000.050 404.400 ;
        RECT 1006.950 403.950 1009.050 404.400 ;
        RECT 4.950 402.600 7.050 403.050 ;
        RECT 40.950 402.600 43.050 403.050 ;
        RECT 55.950 402.600 58.050 403.050 ;
        RECT 4.950 401.400 58.050 402.600 ;
        RECT 4.950 400.950 7.050 401.400 ;
        RECT 40.950 400.950 43.050 401.400 ;
        RECT 55.950 400.950 58.050 401.400 ;
        RECT 340.950 402.600 343.050 403.050 ;
        RECT 481.950 402.600 484.050 403.050 ;
        RECT 340.950 401.400 484.050 402.600 ;
        RECT 340.950 400.950 343.050 401.400 ;
        RECT 481.950 400.950 484.050 401.400 ;
        RECT 544.950 402.600 547.050 403.050 ;
        RECT 562.950 402.600 565.050 403.050 ;
        RECT 544.950 401.400 565.050 402.600 ;
        RECT 544.950 400.950 547.050 401.400 ;
        RECT 562.950 400.950 565.050 401.400 ;
        RECT 715.950 402.600 718.050 403.050 ;
        RECT 745.950 402.600 748.050 403.050 ;
        RECT 808.950 402.600 811.050 403.050 ;
        RECT 715.950 401.400 811.050 402.600 ;
        RECT 715.950 400.950 718.050 401.400 ;
        RECT 745.950 400.950 748.050 401.400 ;
        RECT 808.950 400.950 811.050 401.400 ;
        RECT 901.950 402.600 904.050 403.050 ;
        RECT 913.950 402.600 916.050 403.050 ;
        RECT 901.950 401.400 916.050 402.600 ;
        RECT 901.950 400.950 904.050 401.400 ;
        RECT 913.950 400.950 916.050 401.400 ;
        RECT 964.950 402.600 967.050 403.050 ;
        RECT 994.950 402.600 997.050 403.050 ;
        RECT 964.950 401.400 997.050 402.600 ;
        RECT 964.950 400.950 967.050 401.400 ;
        RECT 994.950 400.950 997.050 401.400 ;
        RECT 76.950 399.600 79.050 400.050 ;
        RECT 109.950 399.600 112.050 400.050 ;
        RECT 76.950 398.400 112.050 399.600 ;
        RECT 76.950 397.950 79.050 398.400 ;
        RECT 109.950 397.950 112.050 398.400 ;
        RECT 205.950 399.600 208.050 400.050 ;
        RECT 268.950 399.600 271.050 400.050 ;
        RECT 301.950 399.600 304.050 400.050 ;
        RECT 325.950 399.600 328.050 400.050 ;
        RECT 433.950 399.600 436.050 400.050 ;
        RECT 445.950 399.600 448.050 400.050 ;
        RECT 460.950 399.600 463.050 400.050 ;
        RECT 205.950 398.400 463.050 399.600 ;
        RECT 205.950 397.950 208.050 398.400 ;
        RECT 268.950 397.950 271.050 398.400 ;
        RECT 301.950 397.950 304.050 398.400 ;
        RECT 325.950 397.950 328.050 398.400 ;
        RECT 433.950 397.950 436.050 398.400 ;
        RECT 445.950 397.950 448.050 398.400 ;
        RECT 460.950 397.950 463.050 398.400 ;
        RECT 487.950 399.600 490.050 400.050 ;
        RECT 541.950 399.600 544.050 400.050 ;
        RECT 487.950 398.400 544.050 399.600 ;
        RECT 487.950 397.950 490.050 398.400 ;
        RECT 541.950 397.950 544.050 398.400 ;
        RECT 616.950 399.600 619.050 400.050 ;
        RECT 643.950 399.600 646.050 400.050 ;
        RECT 616.950 398.400 646.050 399.600 ;
        RECT 616.950 397.950 619.050 398.400 ;
        RECT 643.950 397.950 646.050 398.400 ;
        RECT 733.950 399.600 736.050 400.050 ;
        RECT 787.950 399.600 790.050 400.050 ;
        RECT 793.950 399.600 796.050 400.050 ;
        RECT 733.950 398.400 796.050 399.600 ;
        RECT 733.950 397.950 736.050 398.400 ;
        RECT 787.950 397.950 790.050 398.400 ;
        RECT 793.950 397.950 796.050 398.400 ;
        RECT 961.950 399.600 964.050 400.050 ;
        RECT 1006.950 399.600 1009.050 400.050 ;
        RECT 961.950 398.400 1009.050 399.600 ;
        RECT 961.950 397.950 964.050 398.400 ;
        RECT 1006.950 397.950 1009.050 398.400 ;
        RECT 1.950 396.600 4.050 397.050 ;
        RECT 58.950 396.600 61.050 397.050 ;
        RECT 1.950 395.400 61.050 396.600 ;
        RECT 1.950 394.950 4.050 395.400 ;
        RECT 58.950 394.950 61.050 395.400 ;
        RECT 94.950 396.600 97.050 397.050 ;
        RECT 139.950 396.600 142.050 397.050 ;
        RECT 94.950 395.400 142.050 396.600 ;
        RECT 94.950 394.950 97.050 395.400 ;
        RECT 139.950 394.950 142.050 395.400 ;
        RECT 211.950 396.600 214.050 397.050 ;
        RECT 220.950 396.600 223.050 397.050 ;
        RECT 340.950 396.600 343.050 397.050 ;
        RECT 211.950 395.400 343.050 396.600 ;
        RECT 211.950 394.950 214.050 395.400 ;
        RECT 220.950 394.950 223.050 395.400 ;
        RECT 340.950 394.950 343.050 395.400 ;
        RECT 466.950 396.600 469.050 397.050 ;
        RECT 475.950 396.600 478.050 397.050 ;
        RECT 466.950 395.400 478.050 396.600 ;
        RECT 466.950 394.950 469.050 395.400 ;
        RECT 475.950 394.950 478.050 395.400 ;
        RECT 889.950 396.600 892.050 397.050 ;
        RECT 904.950 396.600 907.050 397.050 ;
        RECT 889.950 395.400 907.050 396.600 ;
        RECT 889.950 394.950 892.050 395.400 ;
        RECT 904.950 394.950 907.050 395.400 ;
        RECT 64.950 393.600 67.050 394.050 ;
        RECT 88.950 393.600 91.050 394.050 ;
        RECT 64.950 392.400 91.050 393.600 ;
        RECT 64.950 391.950 67.050 392.400 ;
        RECT 88.950 391.950 91.050 392.400 ;
        RECT 511.950 393.600 514.050 394.050 ;
        RECT 538.950 393.600 541.050 394.050 ;
        RECT 625.950 393.600 628.050 394.050 ;
        RECT 511.950 392.400 628.050 393.600 ;
        RECT 511.950 391.950 514.050 392.400 ;
        RECT 538.950 391.950 541.050 392.400 ;
        RECT 625.950 391.950 628.050 392.400 ;
        RECT 691.950 393.600 694.050 394.050 ;
        RECT 757.950 393.600 760.050 394.050 ;
        RECT 775.950 393.600 778.050 394.050 ;
        RECT 787.950 393.600 790.050 394.050 ;
        RECT 691.950 392.400 790.050 393.600 ;
        RECT 691.950 391.950 694.050 392.400 ;
        RECT 757.950 391.950 760.050 392.400 ;
        RECT 775.950 391.950 778.050 392.400 ;
        RECT 787.950 391.950 790.050 392.400 ;
        RECT 430.950 390.600 433.050 391.050 ;
        RECT 490.950 390.600 493.050 391.050 ;
        RECT 430.950 389.400 493.050 390.600 ;
        RECT 430.950 388.950 433.050 389.400 ;
        RECT 490.950 388.950 493.050 389.400 ;
        RECT 526.950 390.600 529.050 391.050 ;
        RECT 556.950 390.600 559.050 391.050 ;
        RECT 526.950 389.400 559.050 390.600 ;
        RECT 526.950 388.950 529.050 389.400 ;
        RECT 556.950 388.950 559.050 389.400 ;
        RECT 655.950 390.600 658.050 391.050 ;
        RECT 727.950 390.600 730.050 391.050 ;
        RECT 655.950 389.400 730.050 390.600 ;
        RECT 655.950 388.950 658.050 389.400 ;
        RECT 727.950 388.950 730.050 389.400 ;
        RECT 838.950 390.600 841.050 391.050 ;
        RECT 868.950 390.600 871.050 391.050 ;
        RECT 838.950 389.400 871.050 390.600 ;
        RECT 838.950 388.950 841.050 389.400 ;
        RECT 868.950 388.950 871.050 389.400 ;
        RECT 916.950 390.600 919.050 391.050 ;
        RECT 961.950 390.600 964.050 391.050 ;
        RECT 916.950 389.400 964.050 390.600 ;
        RECT 916.950 388.950 919.050 389.400 ;
        RECT 961.950 388.950 964.050 389.400 ;
        RECT 367.950 387.600 370.050 388.050 ;
        RECT 391.950 387.600 394.050 388.050 ;
        RECT 367.950 386.400 394.050 387.600 ;
        RECT 367.950 385.950 370.050 386.400 ;
        RECT 391.950 385.950 394.050 386.400 ;
        RECT 448.950 387.600 451.050 388.050 ;
        RECT 469.950 387.600 472.050 388.050 ;
        RECT 448.950 386.400 472.050 387.600 ;
        RECT 448.950 385.950 451.050 386.400 ;
        RECT 469.950 385.950 472.050 386.400 ;
        RECT 481.950 387.600 484.050 388.050 ;
        RECT 511.950 387.600 514.050 388.050 ;
        RECT 481.950 386.400 514.050 387.600 ;
        RECT 481.950 385.950 484.050 386.400 ;
        RECT 511.950 385.950 514.050 386.400 ;
        RECT 607.950 387.600 610.050 387.900 ;
        RECT 631.950 387.600 634.050 388.050 ;
        RECT 607.950 386.400 634.050 387.600 ;
        RECT 607.950 385.800 610.050 386.400 ;
        RECT 631.950 385.950 634.050 386.400 ;
        RECT 670.950 387.600 673.050 388.050 ;
        RECT 796.950 387.600 799.050 388.050 ;
        RECT 820.950 387.600 823.050 388.050 ;
        RECT 826.950 387.600 829.050 388.050 ;
        RECT 670.950 386.400 829.050 387.600 ;
        RECT 670.950 385.950 673.050 386.400 ;
        RECT 796.950 385.950 799.050 386.400 ;
        RECT 820.950 385.950 823.050 386.400 ;
        RECT 826.950 385.950 829.050 386.400 ;
        RECT 910.950 387.600 913.050 388.050 ;
        RECT 949.950 387.600 952.050 388.050 ;
        RECT 910.950 386.400 952.050 387.600 ;
        RECT 910.950 385.950 913.050 386.400 ;
        RECT 949.950 385.950 952.050 386.400 ;
        RECT 85.950 384.600 88.050 385.050 ;
        RECT 118.950 384.600 121.050 385.050 ;
        RECT 85.950 383.400 121.050 384.600 ;
        RECT 85.950 382.950 88.050 383.400 ;
        RECT 118.950 382.950 121.050 383.400 ;
        RECT 514.950 384.600 517.050 385.050 ;
        RECT 595.950 384.600 598.050 385.050 ;
        RECT 514.950 383.400 598.050 384.600 ;
        RECT 514.950 382.950 517.050 383.400 ;
        RECT 595.950 382.950 598.050 383.400 ;
        RECT 688.950 384.600 691.050 385.050 ;
        RECT 811.950 384.600 814.050 385.050 ;
        RECT 688.950 383.400 814.050 384.600 ;
        RECT 688.950 382.950 691.050 383.400 ;
        RECT 811.950 382.950 814.050 383.400 ;
        RECT 835.950 384.600 838.050 385.050 ;
        RECT 874.950 384.600 877.050 385.050 ;
        RECT 907.950 384.600 910.050 385.050 ;
        RECT 835.950 383.400 910.050 384.600 ;
        RECT 835.950 382.950 838.050 383.400 ;
        RECT 874.950 382.950 877.050 383.400 ;
        RECT 907.950 382.950 910.050 383.400 ;
        RECT 997.950 384.600 1002.000 385.050 ;
        RECT 997.950 382.950 1002.600 384.600 ;
        RECT 37.950 381.600 40.050 382.050 ;
        RECT 49.950 381.600 52.050 382.050 ;
        RECT 37.950 380.400 52.050 381.600 ;
        RECT 37.950 379.950 40.050 380.400 ;
        RECT 49.950 379.950 52.050 380.400 ;
        RECT 472.950 381.600 475.050 382.050 ;
        RECT 511.950 381.600 514.050 382.050 ;
        RECT 472.950 380.400 514.050 381.600 ;
        RECT 472.950 379.950 475.050 380.400 ;
        RECT 511.950 379.950 514.050 380.400 ;
        RECT 625.950 381.600 628.050 382.050 ;
        RECT 652.950 381.600 655.050 382.050 ;
        RECT 676.950 381.600 679.050 382.050 ;
        RECT 625.950 380.400 679.050 381.600 ;
        RECT 625.950 379.950 628.050 380.400 ;
        RECT 652.950 379.950 655.050 380.400 ;
        RECT 676.950 379.950 679.050 380.400 ;
        RECT 865.950 381.600 868.050 382.050 ;
        RECT 931.950 381.600 934.050 382.050 ;
        RECT 997.950 381.600 1000.050 381.900 ;
        RECT 865.950 380.400 1000.050 381.600 ;
        RECT 865.950 379.950 868.050 380.400 ;
        RECT 931.950 379.950 934.050 380.400 ;
        RECT 997.950 379.800 1000.050 380.400 ;
        RECT 55.950 378.600 58.050 379.050 ;
        RECT 70.950 378.600 73.050 379.050 ;
        RECT 100.950 378.600 103.050 379.050 ;
        RECT 55.950 377.400 103.050 378.600 ;
        RECT 55.950 376.950 58.050 377.400 ;
        RECT 70.950 376.950 73.050 377.400 ;
        RECT 100.950 376.950 103.050 377.400 ;
        RECT 190.950 378.600 193.050 379.050 ;
        RECT 310.950 378.600 313.050 379.050 ;
        RECT 190.950 377.400 313.050 378.600 ;
        RECT 190.950 376.950 193.050 377.400 ;
        RECT 310.950 376.950 313.050 377.400 ;
        RECT 550.950 378.600 553.050 379.050 ;
        RECT 610.950 378.600 613.050 379.050 ;
        RECT 619.950 378.600 622.050 379.050 ;
        RECT 550.950 377.400 622.050 378.600 ;
        RECT 550.950 376.950 553.050 377.400 ;
        RECT 610.950 376.950 613.050 377.400 ;
        RECT 619.950 376.950 622.050 377.400 ;
        RECT 685.950 378.600 688.050 379.050 ;
        RECT 691.950 378.600 694.050 379.050 ;
        RECT 685.950 377.400 694.050 378.600 ;
        RECT 685.950 376.950 688.050 377.400 ;
        RECT 691.950 376.950 694.050 377.400 ;
        RECT 703.950 378.600 706.050 379.050 ;
        RECT 742.950 378.600 745.050 379.050 ;
        RECT 775.950 378.600 778.050 379.050 ;
        RECT 703.950 377.400 778.050 378.600 ;
        RECT 703.950 376.950 706.050 377.400 ;
        RECT 742.950 376.950 745.050 377.400 ;
        RECT 775.950 376.950 778.050 377.400 ;
        RECT 790.950 378.600 793.050 379.050 ;
        RECT 820.950 378.600 823.050 379.050 ;
        RECT 790.950 377.400 823.050 378.600 ;
        RECT 790.950 376.950 793.050 377.400 ;
        RECT 820.950 376.950 823.050 377.400 ;
        RECT 907.950 378.600 910.050 379.050 ;
        RECT 925.950 378.600 928.050 379.050 ;
        RECT 907.950 377.400 928.050 378.600 ;
        RECT 907.950 376.950 910.050 377.400 ;
        RECT 925.950 376.950 928.050 377.400 ;
        RECT 943.950 378.600 946.050 379.050 ;
        RECT 970.950 378.600 973.050 379.050 ;
        RECT 943.950 377.400 973.050 378.600 ;
        RECT 943.950 376.950 946.050 377.400 ;
        RECT 970.950 376.950 973.050 377.400 ;
        RECT 481.950 375.600 486.000 376.050 ;
        RECT 526.950 375.600 529.050 376.050 ;
        RECT 553.950 375.600 556.050 376.050 ;
        RECT 481.950 373.950 486.600 375.600 ;
        RECT 526.950 374.400 556.050 375.600 ;
        RECT 526.950 373.950 529.050 374.400 ;
        RECT 553.950 373.950 556.050 374.400 ;
        RECT 601.950 375.600 604.050 376.050 ;
        RECT 622.950 375.600 625.050 376.050 ;
        RECT 682.950 375.600 685.050 376.050 ;
        RECT 865.950 375.600 868.050 376.050 ;
        RECT 601.950 374.400 625.050 375.600 ;
        RECT 601.950 373.950 604.050 374.400 ;
        RECT 622.950 373.950 625.050 374.400 ;
        RECT 662.400 374.400 685.050 375.600 ;
        RECT 43.950 371.100 46.050 373.200 ;
        RECT 79.950 372.750 82.050 373.200 ;
        RECT 103.950 372.750 106.050 373.200 ;
        RECT 79.950 371.550 106.050 372.750 ;
        RECT 79.950 371.100 82.050 371.550 ;
        RECT 103.950 371.100 106.050 371.550 ;
        RECT 124.950 372.750 127.050 373.200 ;
        RECT 151.950 372.750 154.050 373.050 ;
        RECT 160.950 372.750 163.050 373.200 ;
        RECT 124.950 372.600 163.050 372.750 ;
        RECT 175.950 372.600 178.050 373.050 ;
        RECT 124.950 371.550 178.050 372.600 ;
        RECT 124.950 371.100 127.050 371.550 ;
        RECT 28.950 366.600 31.050 367.050 ;
        RECT 40.950 366.600 43.050 366.900 ;
        RECT 28.950 365.400 43.050 366.600 ;
        RECT 44.400 366.600 45.600 371.100 ;
        RECT 151.950 370.950 154.050 371.550 ;
        RECT 160.950 371.400 178.050 371.550 ;
        RECT 160.950 371.100 163.050 371.400 ;
        RECT 175.950 370.950 178.050 371.400 ;
        RECT 181.950 372.600 184.050 373.200 ;
        RECT 190.950 372.600 193.050 373.200 ;
        RECT 181.950 371.400 193.050 372.600 ;
        RECT 181.950 371.100 184.050 371.400 ;
        RECT 190.950 371.100 193.050 371.400 ;
        RECT 199.950 372.750 202.050 373.200 ;
        RECT 208.950 372.750 211.050 373.200 ;
        RECT 199.950 371.550 211.050 372.750 ;
        RECT 199.950 371.100 202.050 371.550 ;
        RECT 208.950 371.100 211.050 371.550 ;
        RECT 226.950 372.750 229.050 373.200 ;
        RECT 238.950 372.750 241.050 373.200 ;
        RECT 226.950 371.550 241.050 372.750 ;
        RECT 226.950 371.100 229.050 371.550 ;
        RECT 238.950 371.100 241.050 371.550 ;
        RECT 244.950 372.750 247.050 373.200 ;
        RECT 256.950 372.750 259.050 373.200 ;
        RECT 244.950 371.550 259.050 372.750 ;
        RECT 244.950 371.100 247.050 371.550 ;
        RECT 256.950 371.100 259.050 371.550 ;
        RECT 283.950 372.600 286.050 373.200 ;
        RECT 292.950 372.600 295.050 373.200 ;
        RECT 283.950 371.400 295.050 372.600 ;
        RECT 283.950 371.100 286.050 371.400 ;
        RECT 292.950 371.100 295.050 371.400 ;
        RECT 301.950 372.600 304.050 373.200 ;
        RECT 334.950 372.600 337.050 373.050 ;
        RECT 301.950 371.400 337.050 372.600 ;
        RECT 301.950 371.100 304.050 371.400 ;
        RECT 334.950 370.950 337.050 371.400 ;
        RECT 340.950 371.100 343.050 373.200 ;
        RECT 346.950 372.750 349.050 373.200 ;
        RECT 352.800 372.750 354.900 373.200 ;
        RECT 346.950 371.550 354.900 372.750 ;
        RECT 346.950 371.100 349.050 371.550 ;
        RECT 352.800 371.100 354.900 371.550 ;
        RECT 355.950 372.750 358.050 373.200 ;
        RECT 385.950 372.750 388.050 373.200 ;
        RECT 355.950 371.550 388.050 372.750 ;
        RECT 355.950 371.100 358.050 371.550 ;
        RECT 385.950 371.100 388.050 371.550 ;
        RECT 391.950 371.100 394.050 373.200 ;
        RECT 397.950 372.750 400.050 373.200 ;
        RECT 406.950 372.750 409.050 373.200 ;
        RECT 397.950 371.550 409.050 372.750 ;
        RECT 397.950 371.100 400.050 371.550 ;
        RECT 406.950 371.100 409.050 371.550 ;
        RECT 412.950 371.100 415.050 373.200 ;
        RECT 430.950 371.100 433.050 373.200 ;
        RECT 442.950 372.600 447.000 373.050 ;
        RECT 341.400 369.600 342.600 371.100 ;
        RECT 341.400 368.400 360.600 369.600 ;
        RECT 61.950 366.600 64.050 366.900 ;
        RECT 44.400 365.400 64.050 366.600 ;
        RECT 28.950 364.950 31.050 365.400 ;
        RECT 40.950 364.800 43.050 365.400 ;
        RECT 61.950 364.800 64.050 365.400 ;
        RECT 88.950 366.600 91.050 367.050 ;
        RECT 139.950 366.600 142.050 366.900 ;
        RECT 88.950 366.450 142.050 366.600 ;
        RECT 151.950 366.450 154.050 366.900 ;
        RECT 88.950 365.400 154.050 366.450 ;
        RECT 88.950 364.950 91.050 365.400 ;
        RECT 139.950 365.250 154.050 365.400 ;
        RECT 139.950 364.800 142.050 365.250 ;
        RECT 151.950 364.800 154.050 365.250 ;
        RECT 232.950 366.600 235.050 367.050 ;
        RECT 241.950 366.600 244.050 366.900 ;
        RECT 232.950 365.400 244.050 366.600 ;
        RECT 232.950 364.950 235.050 365.400 ;
        RECT 241.950 364.800 244.050 365.400 ;
        RECT 319.950 366.600 322.050 366.900 ;
        RECT 355.950 366.600 358.050 367.050 ;
        RECT 319.950 365.400 358.050 366.600 ;
        RECT 359.400 366.600 360.600 368.400 ;
        RECT 370.950 366.600 373.050 366.900 ;
        RECT 359.400 365.400 373.050 366.600 ;
        RECT 392.400 366.600 393.600 371.100 ;
        RECT 413.400 369.600 414.600 371.100 ;
        RECT 413.400 368.400 417.600 369.600 ;
        RECT 416.400 367.050 417.600 368.400 ;
        RECT 403.950 366.600 406.050 367.050 ;
        RECT 392.400 365.400 406.050 366.600 ;
        RECT 416.400 365.400 421.050 367.050 ;
        RECT 319.950 364.800 322.050 365.400 ;
        RECT 355.950 364.950 358.050 365.400 ;
        RECT 370.950 364.800 373.050 365.400 ;
        RECT 403.950 364.950 406.050 365.400 ;
        RECT 417.000 364.950 421.050 365.400 ;
        RECT 97.950 363.600 100.050 364.050 ;
        RECT 343.950 363.600 346.050 364.050 ;
        RECT 349.950 363.600 352.050 364.050 ;
        RECT 97.950 362.400 138.600 363.600 ;
        RECT 97.950 361.950 100.050 362.400 ;
        RECT 137.400 361.050 138.600 362.400 ;
        RECT 343.950 362.400 352.050 363.600 ;
        RECT 343.950 361.950 346.050 362.400 ;
        RECT 349.950 361.950 352.050 362.400 ;
        RECT 358.950 363.600 361.050 364.050 ;
        RECT 364.950 363.600 367.050 364.050 ;
        RECT 358.950 362.400 367.050 363.600 ;
        RECT 358.950 361.950 361.050 362.400 ;
        RECT 364.950 361.950 367.050 362.400 ;
        RECT 388.950 363.600 391.050 364.050 ;
        RECT 397.950 363.600 400.050 364.050 ;
        RECT 388.950 362.400 400.050 363.600 ;
        RECT 388.950 361.950 391.050 362.400 ;
        RECT 397.950 361.950 400.050 362.400 ;
        RECT 412.950 363.600 415.050 364.050 ;
        RECT 431.400 363.600 432.600 371.100 ;
        RECT 442.950 370.950 447.600 372.600 ;
        RECT 446.400 366.600 447.600 370.950 ;
        RECT 457.950 366.600 460.050 366.900 ;
        RECT 463.950 366.600 466.050 366.900 ;
        RECT 446.400 365.400 466.050 366.600 ;
        RECT 457.950 364.800 460.050 365.400 ;
        RECT 463.950 364.800 466.050 365.400 ;
        RECT 485.400 364.050 486.600 373.950 ;
        RECT 490.950 372.600 493.050 373.200 ;
        RECT 499.950 372.600 502.050 373.200 ;
        RECT 514.950 372.600 517.050 373.050 ;
        RECT 490.950 371.400 517.050 372.600 ;
        RECT 490.950 371.100 493.050 371.400 ;
        RECT 499.950 371.100 502.050 371.400 ;
        RECT 514.950 370.950 517.050 371.400 ;
        RECT 529.950 370.950 532.050 373.050 ;
        RECT 556.950 372.750 559.050 373.200 ;
        RECT 571.950 372.750 574.050 373.200 ;
        RECT 556.950 371.550 574.050 372.750 ;
        RECT 658.950 372.600 661.050 373.200 ;
        RECT 662.400 372.600 663.600 374.400 ;
        RECT 682.950 373.950 685.050 374.400 ;
        RECT 857.400 374.400 868.050 375.600 ;
        RECT 556.950 371.100 559.050 371.550 ;
        RECT 571.950 371.100 574.050 371.550 ;
        RECT 614.400 371.400 663.600 372.600 ;
        RECT 670.950 372.600 673.050 373.050 ;
        RECT 745.950 372.600 748.050 373.050 ;
        RECT 670.950 371.400 748.050 372.600 ;
        RECT 511.950 366.600 514.050 367.050 ;
        RECT 530.400 366.600 531.600 370.950 ;
        RECT 541.950 369.600 544.050 370.050 ;
        RECT 562.950 369.600 565.050 370.050 ;
        RECT 614.400 369.600 615.600 371.400 ;
        RECT 658.950 371.100 661.050 371.400 ;
        RECT 670.950 370.950 673.050 371.400 ;
        RECT 745.950 370.950 748.050 371.400 ;
        RECT 751.950 371.100 754.050 373.200 ;
        RECT 802.950 372.750 805.050 373.200 ;
        RECT 817.950 372.750 820.050 373.200 ;
        RECT 802.950 371.550 820.050 372.750 ;
        RECT 802.950 371.100 805.050 371.550 ;
        RECT 817.950 371.100 820.050 371.550 ;
        RECT 850.950 371.100 853.050 373.200 ;
        RECT 752.400 369.600 753.600 371.100 ;
        RECT 541.950 368.400 565.050 369.600 ;
        RECT 541.950 367.950 544.050 368.400 ;
        RECT 562.950 367.950 565.050 368.400 ;
        RECT 611.400 368.400 615.600 369.600 ;
        RECT 722.400 369.000 762.600 369.600 ;
        RECT 721.950 368.400 763.050 369.000 ;
        RECT 511.950 365.400 531.600 366.600 ;
        RECT 595.950 366.600 598.050 367.050 ;
        RECT 611.400 366.900 612.600 368.400 ;
        RECT 610.950 366.600 613.050 366.900 ;
        RECT 595.950 365.400 613.050 366.600 ;
        RECT 511.950 364.950 514.050 365.400 ;
        RECT 595.950 364.950 598.050 365.400 ;
        RECT 610.950 364.800 613.050 365.400 ;
        RECT 619.950 366.450 622.050 366.900 ;
        RECT 628.950 366.450 631.050 366.900 ;
        RECT 619.950 365.250 631.050 366.450 ;
        RECT 619.950 364.800 622.050 365.250 ;
        RECT 628.950 364.800 631.050 365.250 ;
        RECT 706.950 366.450 709.050 366.900 ;
        RECT 715.950 366.450 718.050 366.900 ;
        RECT 706.950 365.250 718.050 366.450 ;
        RECT 706.950 364.800 709.050 365.250 ;
        RECT 715.950 364.800 718.050 365.250 ;
        RECT 721.950 364.950 724.050 368.400 ;
        RECT 760.950 364.950 763.050 368.400 ;
        RECT 766.950 366.450 769.050 366.900 ;
        RECT 790.950 366.450 793.050 367.050 ;
        RECT 799.950 366.450 802.050 366.900 ;
        RECT 766.950 365.250 802.050 366.450 ;
        RECT 766.950 364.800 769.050 365.250 ;
        RECT 790.950 364.950 793.050 365.250 ;
        RECT 799.950 364.800 802.050 365.250 ;
        RECT 814.950 366.450 817.050 366.900 ;
        RECT 823.950 366.450 826.050 366.900 ;
        RECT 814.950 365.250 826.050 366.450 ;
        RECT 814.950 364.800 817.050 365.250 ;
        RECT 823.950 364.800 826.050 365.250 ;
        RECT 841.950 366.600 844.050 367.050 ;
        RECT 851.400 366.600 852.600 371.100 ;
        RECT 841.950 365.400 852.600 366.600 ;
        RECT 853.950 366.600 856.050 366.900 ;
        RECT 857.400 366.600 858.600 374.400 ;
        RECT 865.950 373.950 868.050 374.400 ;
        RECT 871.950 375.600 874.050 376.050 ;
        RECT 895.950 375.600 898.050 376.050 ;
        RECT 871.950 374.400 894.600 375.600 ;
        RECT 871.950 373.950 874.050 374.400 ;
        RECT 859.950 370.950 862.050 373.050 ;
        RECT 893.400 372.600 894.600 374.400 ;
        RECT 895.950 374.400 903.600 375.600 ;
        RECT 895.950 373.950 898.050 374.400 ;
        RECT 898.950 372.600 901.050 373.200 ;
        RECT 893.400 371.400 901.050 372.600 ;
        RECT 898.950 371.100 901.050 371.400 ;
        RECT 853.950 365.400 858.600 366.600 ;
        RECT 841.950 364.950 844.050 365.400 ;
        RECT 853.950 364.800 856.050 365.400 ;
        RECT 412.950 362.400 432.600 363.600 ;
        RECT 481.950 362.400 486.600 364.050 ;
        RECT 550.950 363.600 553.050 364.050 ;
        RECT 568.950 363.600 571.050 364.050 ;
        RECT 550.950 362.400 571.050 363.600 ;
        RECT 412.950 361.950 415.050 362.400 ;
        RECT 481.950 361.950 486.000 362.400 ;
        RECT 550.950 361.950 553.050 362.400 ;
        RECT 568.950 361.950 571.050 362.400 ;
        RECT 580.950 363.600 583.050 364.050 ;
        RECT 592.950 363.600 595.050 364.050 ;
        RECT 607.950 363.600 610.050 364.050 ;
        RECT 580.950 362.400 610.050 363.600 ;
        RECT 580.950 361.950 583.050 362.400 ;
        RECT 592.950 361.950 595.050 362.400 ;
        RECT 607.950 361.950 610.050 362.400 ;
        RECT 670.950 363.600 673.050 364.050 ;
        RECT 682.950 363.600 685.050 364.050 ;
        RECT 670.950 362.400 685.050 363.600 ;
        RECT 670.950 361.950 673.050 362.400 ;
        RECT 682.950 361.950 685.050 362.400 ;
        RECT 742.950 363.600 745.050 364.050 ;
        RECT 829.950 363.600 832.050 364.050 ;
        RECT 860.400 363.600 861.600 370.950 ;
        RECT 902.400 366.900 903.600 374.400 ;
        RECT 994.950 373.950 997.050 376.050 ;
        RECT 1001.400 375.600 1002.600 382.950 ;
        RECT 1001.400 374.400 1008.600 375.600 ;
        RECT 943.950 372.600 946.050 373.200 ;
        RECT 929.400 371.400 946.050 372.600 ;
        RECT 929.400 367.050 930.600 371.400 ;
        RECT 943.950 371.100 946.050 371.400 ;
        RECT 970.950 371.100 973.050 373.200 ;
        RECT 971.400 369.600 972.600 371.100 ;
        RECT 995.400 369.600 996.600 373.950 ;
        RECT 1000.950 370.950 1003.050 373.050 ;
        RECT 965.400 369.000 972.600 369.600 ;
        RECT 980.400 369.000 996.600 369.600 ;
        RECT 964.950 368.400 972.600 369.000 ;
        RECT 979.950 368.400 996.600 369.000 ;
        RECT 901.950 366.600 904.050 366.900 ;
        RECT 916.950 366.600 919.050 366.900 ;
        RECT 901.950 365.400 919.050 366.600 ;
        RECT 901.950 364.800 904.050 365.400 ;
        RECT 916.950 364.800 919.050 365.400 ;
        RECT 928.950 364.950 931.050 367.050 ;
        RECT 964.950 364.950 967.050 368.400 ;
        RECT 979.950 364.950 982.050 368.400 ;
        RECT 1001.400 367.050 1002.600 370.950 ;
        RECT 1000.950 364.950 1003.050 367.050 ;
        RECT 742.950 363.000 750.600 363.600 ;
        RECT 742.950 362.400 751.050 363.000 ;
        RECT 742.950 361.950 745.050 362.400 ;
        RECT 103.950 360.600 106.050 361.050 ;
        RECT 115.950 360.600 118.050 361.050 ;
        RECT 103.950 359.400 118.050 360.600 ;
        RECT 103.950 358.950 106.050 359.400 ;
        RECT 115.950 358.950 118.050 359.400 ;
        RECT 136.950 360.600 139.050 361.050 ;
        RECT 145.950 360.600 148.050 361.050 ;
        RECT 136.950 359.400 148.050 360.600 ;
        RECT 136.950 358.950 139.050 359.400 ;
        RECT 145.950 358.950 148.050 359.400 ;
        RECT 454.950 360.600 457.050 361.050 ;
        RECT 472.950 360.600 475.050 361.050 ;
        RECT 454.950 359.400 475.050 360.600 ;
        RECT 454.950 358.950 457.050 359.400 ;
        RECT 472.950 358.950 475.050 359.400 ;
        RECT 517.950 360.600 520.050 361.050 ;
        RECT 551.400 360.600 552.600 361.950 ;
        RECT 517.950 359.400 552.600 360.600 ;
        RECT 583.950 360.600 586.050 361.050 ;
        RECT 592.950 360.600 595.050 360.900 ;
        RECT 583.950 359.400 595.050 360.600 ;
        RECT 517.950 358.950 520.050 359.400 ;
        RECT 583.950 358.950 586.050 359.400 ;
        RECT 592.950 358.800 595.050 359.400 ;
        RECT 652.950 360.600 655.050 361.050 ;
        RECT 658.950 360.600 661.050 361.050 ;
        RECT 721.950 360.600 724.050 361.050 ;
        RECT 652.950 359.400 661.050 360.600 ;
        RECT 652.950 358.950 655.050 359.400 ;
        RECT 658.950 358.950 661.050 359.400 ;
        RECT 695.400 359.400 724.050 360.600 ;
        RECT 334.950 357.600 337.050 358.050 ;
        RECT 403.950 357.600 406.050 358.050 ;
        RECT 415.950 357.600 418.050 358.050 ;
        RECT 553.950 357.600 556.050 358.050 ;
        RECT 601.950 357.600 604.050 358.050 ;
        RECT 613.950 357.600 616.050 358.050 ;
        RECT 676.950 357.600 679.050 358.050 ;
        RECT 695.400 357.600 696.600 359.400 ;
        RECT 721.950 358.950 724.050 359.400 ;
        RECT 748.950 358.950 751.050 362.400 ;
        RECT 829.950 362.400 861.600 363.600 ;
        RECT 865.950 363.600 868.050 364.050 ;
        RECT 886.950 363.600 889.050 364.050 ;
        RECT 865.950 362.400 889.050 363.600 ;
        RECT 829.950 361.950 832.050 362.400 ;
        RECT 865.950 361.950 868.050 362.400 ;
        RECT 886.950 361.950 889.050 362.400 ;
        RECT 931.950 363.600 934.050 364.050 ;
        RECT 946.950 363.600 949.050 364.050 ;
        RECT 931.950 362.400 949.050 363.600 ;
        RECT 931.950 361.950 934.050 362.400 ;
        RECT 946.950 361.950 949.050 362.400 ;
        RECT 961.950 363.600 964.050 364.050 ;
        RECT 973.950 363.600 976.050 364.050 ;
        RECT 961.950 362.400 976.050 363.600 ;
        RECT 961.950 361.950 964.050 362.400 ;
        RECT 973.950 361.950 976.050 362.400 ;
        RECT 994.950 363.600 997.050 364.050 ;
        RECT 1003.950 363.600 1006.050 364.050 ;
        RECT 994.950 362.400 1006.050 363.600 ;
        RECT 994.950 361.950 997.050 362.400 ;
        RECT 1003.950 361.950 1006.050 362.400 ;
        RECT 1007.400 361.050 1008.600 374.400 ;
        RECT 754.950 360.600 757.050 361.050 ;
        RECT 862.950 360.600 865.050 361.050 ;
        RECT 754.950 359.400 865.050 360.600 ;
        RECT 754.950 358.950 757.050 359.400 ;
        RECT 862.950 358.950 865.050 359.400 ;
        RECT 910.950 360.600 913.050 361.050 ;
        RECT 922.950 360.600 925.050 361.050 ;
        RECT 1005.000 360.900 1008.600 361.050 ;
        RECT 910.950 359.400 925.050 360.600 ;
        RECT 910.950 358.950 913.050 359.400 ;
        RECT 922.950 358.950 925.050 359.400 ;
        RECT 1003.950 359.400 1008.600 360.900 ;
        RECT 1003.950 358.950 1008.000 359.400 ;
        RECT 1003.950 358.800 1006.050 358.950 ;
        RECT 334.950 356.400 402.600 357.600 ;
        RECT 334.950 355.950 337.050 356.400 ;
        RECT 73.950 354.600 76.050 355.050 ;
        RECT 109.950 354.600 112.050 355.050 ;
        RECT 73.950 353.400 112.050 354.600 ;
        RECT 73.950 352.950 76.050 353.400 ;
        RECT 109.950 352.950 112.050 353.400 ;
        RECT 175.950 354.600 178.050 355.050 ;
        RECT 214.950 354.600 217.050 355.050 ;
        RECT 175.950 353.400 217.050 354.600 ;
        RECT 175.950 352.950 178.050 353.400 ;
        RECT 214.950 352.950 217.050 353.400 ;
        RECT 319.950 354.600 322.050 355.050 ;
        RECT 388.950 354.600 391.050 355.050 ;
        RECT 319.950 353.400 391.050 354.600 ;
        RECT 401.400 354.600 402.600 356.400 ;
        RECT 403.950 356.400 679.050 357.600 ;
        RECT 403.950 355.950 406.050 356.400 ;
        RECT 415.950 355.950 418.050 356.400 ;
        RECT 553.950 355.950 556.050 356.400 ;
        RECT 601.950 355.950 604.050 356.400 ;
        RECT 613.950 355.950 616.050 356.400 ;
        RECT 676.950 355.950 679.050 356.400 ;
        RECT 686.400 356.400 696.600 357.600 ;
        RECT 703.950 357.600 706.050 358.050 ;
        RECT 712.950 357.600 715.050 358.050 ;
        RECT 703.950 356.400 715.050 357.600 ;
        RECT 409.950 354.600 412.050 355.050 ;
        RECT 401.400 353.400 412.050 354.600 ;
        RECT 319.950 352.950 322.050 353.400 ;
        RECT 388.950 352.950 391.050 353.400 ;
        RECT 409.950 352.950 412.050 353.400 ;
        RECT 433.950 354.600 436.050 355.050 ;
        RECT 472.950 354.600 475.050 355.050 ;
        RECT 433.950 353.400 475.050 354.600 ;
        RECT 433.950 352.950 436.050 353.400 ;
        RECT 472.950 352.950 475.050 353.400 ;
        RECT 526.950 354.600 529.050 355.050 ;
        RECT 538.950 354.600 541.050 355.050 ;
        RECT 526.950 353.400 541.050 354.600 ;
        RECT 526.950 352.950 529.050 353.400 ;
        RECT 538.950 352.950 541.050 353.400 ;
        RECT 607.950 354.600 610.050 355.050 ;
        RECT 652.950 354.600 655.050 355.050 ;
        RECT 607.950 353.400 655.050 354.600 ;
        RECT 607.950 352.950 610.050 353.400 ;
        RECT 652.950 352.950 655.050 353.400 ;
        RECT 661.950 354.600 664.050 355.050 ;
        RECT 686.400 354.600 687.600 356.400 ;
        RECT 703.950 355.950 706.050 356.400 ;
        RECT 712.950 355.950 715.050 356.400 ;
        RECT 730.950 357.600 733.050 358.050 ;
        RECT 766.950 357.600 769.050 358.050 ;
        RECT 730.950 356.400 769.050 357.600 ;
        RECT 730.950 355.950 733.050 356.400 ;
        RECT 766.950 355.950 769.050 356.400 ;
        RECT 781.950 357.600 784.050 358.050 ;
        RECT 841.950 357.600 844.050 358.050 ;
        RECT 880.950 357.600 883.050 358.050 ;
        RECT 781.950 356.400 883.050 357.600 ;
        RECT 781.950 355.950 784.050 356.400 ;
        RECT 841.950 355.950 844.050 356.400 ;
        RECT 880.950 355.950 883.050 356.400 ;
        RECT 898.950 357.600 901.050 358.050 ;
        RECT 907.950 357.600 910.050 358.050 ;
        RECT 898.950 356.400 910.050 357.600 ;
        RECT 898.950 355.950 901.050 356.400 ;
        RECT 907.950 355.950 910.050 356.400 ;
        RECT 661.950 353.400 687.600 354.600 ;
        RECT 715.950 354.600 718.050 355.050 ;
        RECT 769.950 354.600 772.050 355.050 ;
        RECT 715.950 353.400 772.050 354.600 ;
        RECT 661.950 352.950 664.050 353.400 ;
        RECT 715.950 352.950 718.050 353.400 ;
        RECT 769.950 352.950 772.050 353.400 ;
        RECT 778.950 354.600 781.050 355.050 ;
        RECT 805.950 354.600 808.050 355.050 ;
        RECT 847.950 354.600 850.050 355.050 ;
        RECT 871.950 354.600 874.050 355.050 ;
        RECT 778.950 353.400 801.600 354.600 ;
        RECT 778.950 352.950 781.050 353.400 ;
        RECT 4.950 351.600 7.050 352.050 ;
        RECT 25.950 351.600 28.050 352.050 ;
        RECT 4.950 350.400 28.050 351.600 ;
        RECT 4.950 349.950 7.050 350.400 ;
        RECT 25.950 349.950 28.050 350.400 ;
        RECT 328.950 351.600 331.050 352.050 ;
        RECT 355.950 351.600 358.050 352.050 ;
        RECT 328.950 350.400 358.050 351.600 ;
        RECT 328.950 349.950 331.050 350.400 ;
        RECT 355.950 349.950 358.050 350.400 ;
        RECT 475.950 351.600 478.050 352.050 ;
        RECT 493.950 351.600 496.050 352.050 ;
        RECT 475.950 350.400 496.050 351.600 ;
        RECT 475.950 349.950 478.050 350.400 ;
        RECT 493.950 349.950 496.050 350.400 ;
        RECT 502.950 351.600 505.050 352.050 ;
        RECT 511.950 351.600 514.050 352.050 ;
        RECT 502.950 350.400 514.050 351.600 ;
        RECT 502.950 349.950 505.050 350.400 ;
        RECT 511.950 349.950 514.050 350.400 ;
        RECT 553.950 351.600 556.050 352.050 ;
        RECT 700.950 351.600 703.050 352.050 ;
        RECT 553.950 350.400 703.050 351.600 ;
        RECT 800.400 351.600 801.600 353.400 ;
        RECT 805.950 353.400 874.050 354.600 ;
        RECT 805.950 352.950 808.050 353.400 ;
        RECT 847.950 352.950 850.050 353.400 ;
        RECT 871.950 352.950 874.050 353.400 ;
        RECT 946.950 354.600 949.050 355.050 ;
        RECT 958.950 354.600 961.050 355.050 ;
        RECT 946.950 353.400 961.050 354.600 ;
        RECT 946.950 352.950 949.050 353.400 ;
        RECT 958.950 352.950 961.050 353.400 ;
        RECT 871.950 351.600 874.050 351.900 ;
        RECT 800.400 350.400 874.050 351.600 ;
        RECT 553.950 349.950 556.050 350.400 ;
        RECT 700.950 349.950 703.050 350.400 ;
        RECT 871.950 349.800 874.050 350.400 ;
        RECT 883.950 351.600 886.050 352.050 ;
        RECT 916.950 351.600 919.050 352.050 ;
        RECT 883.950 350.400 919.050 351.600 ;
        RECT 883.950 349.950 886.050 350.400 ;
        RECT 916.950 349.950 919.050 350.400 ;
        RECT 943.950 351.600 946.050 352.050 ;
        RECT 955.950 351.600 958.050 352.050 ;
        RECT 985.950 351.600 988.050 352.050 ;
        RECT 943.950 350.400 988.050 351.600 ;
        RECT 943.950 349.950 946.050 350.400 ;
        RECT 955.950 349.950 958.050 350.400 ;
        RECT 985.950 349.950 988.050 350.400 ;
        RECT 115.950 348.600 118.050 349.050 ;
        RECT 541.950 348.600 544.050 349.050 ;
        RECT 53.400 347.400 118.050 348.600 ;
        RECT 53.400 346.050 54.600 347.400 ;
        RECT 115.950 346.950 118.050 347.400 ;
        RECT 515.400 347.400 544.050 348.600 ;
        RECT 40.950 345.600 43.050 346.050 ;
        RECT 52.950 345.600 55.050 346.050 ;
        RECT 40.950 344.400 55.050 345.600 ;
        RECT 40.950 343.950 43.050 344.400 ;
        RECT 52.950 343.950 55.050 344.400 ;
        RECT 61.950 345.600 64.050 346.050 ;
        RECT 85.950 345.600 88.050 346.050 ;
        RECT 61.950 344.400 88.050 345.600 ;
        RECT 61.950 343.950 64.050 344.400 ;
        RECT 85.950 343.950 88.050 344.400 ;
        RECT 187.950 345.600 190.050 346.050 ;
        RECT 199.950 345.600 202.050 346.050 ;
        RECT 187.950 344.400 202.050 345.600 ;
        RECT 187.950 343.950 190.050 344.400 ;
        RECT 199.950 343.950 202.050 344.400 ;
        RECT 286.950 345.600 289.050 346.050 ;
        RECT 295.950 345.600 298.050 346.050 ;
        RECT 286.950 344.400 298.050 345.600 ;
        RECT 286.950 343.950 289.050 344.400 ;
        RECT 295.950 343.950 298.050 344.400 ;
        RECT 325.950 345.600 328.050 346.050 ;
        RECT 358.950 345.600 361.050 346.050 ;
        RECT 379.950 345.600 382.050 346.050 ;
        RECT 325.950 344.400 382.050 345.600 ;
        RECT 325.950 343.950 328.050 344.400 ;
        RECT 358.950 343.950 361.050 344.400 ;
        RECT 379.950 343.950 382.050 344.400 ;
        RECT 460.950 345.600 463.050 346.050 ;
        RECT 515.400 345.600 516.600 347.400 ;
        RECT 541.950 346.950 544.050 347.400 ;
        RECT 619.950 348.600 622.050 349.050 ;
        RECT 736.950 348.600 739.050 349.050 ;
        RECT 754.950 348.600 757.050 349.050 ;
        RECT 784.950 348.600 787.050 349.050 ;
        RECT 619.950 347.400 645.600 348.600 ;
        RECT 619.950 346.950 622.050 347.400 ;
        RECT 460.950 344.400 516.600 345.600 ;
        RECT 644.400 345.600 645.600 347.400 ;
        RECT 736.950 347.400 787.050 348.600 ;
        RECT 736.950 346.950 739.050 347.400 ;
        RECT 754.950 346.950 757.050 347.400 ;
        RECT 784.950 346.950 787.050 347.400 ;
        RECT 835.950 348.600 838.050 349.050 ;
        RECT 859.950 348.600 862.050 349.050 ;
        RECT 835.950 347.400 862.050 348.600 ;
        RECT 835.950 346.950 838.050 347.400 ;
        RECT 859.950 346.950 862.050 347.400 ;
        RECT 952.950 348.600 955.050 349.050 ;
        RECT 991.950 348.600 994.050 349.050 ;
        RECT 952.950 347.400 994.050 348.600 ;
        RECT 952.950 346.950 955.050 347.400 ;
        RECT 991.950 346.950 994.050 347.400 ;
        RECT 655.950 345.600 658.050 346.050 ;
        RECT 679.950 345.600 682.050 346.050 ;
        RECT 644.400 344.400 682.050 345.600 ;
        RECT 460.950 343.950 463.050 344.400 ;
        RECT 655.950 343.950 658.050 344.400 ;
        RECT 679.950 343.950 682.050 344.400 ;
        RECT 691.950 345.600 694.050 346.050 ;
        RECT 727.950 345.600 730.050 346.050 ;
        RECT 691.950 344.400 730.050 345.600 ;
        RECT 691.950 343.950 694.050 344.400 ;
        RECT 727.950 343.950 730.050 344.400 ;
        RECT 811.950 345.600 814.050 346.050 ;
        RECT 865.950 345.600 868.050 346.050 ;
        RECT 811.950 344.400 868.050 345.600 ;
        RECT 811.950 343.950 814.050 344.400 ;
        RECT 865.950 343.950 868.050 344.400 ;
        RECT 874.950 345.600 877.050 346.050 ;
        RECT 901.950 345.600 904.050 346.050 ;
        RECT 874.950 344.400 904.050 345.600 ;
        RECT 874.950 343.950 877.050 344.400 ;
        RECT 901.950 343.950 904.050 344.400 ;
        RECT 913.950 345.600 916.050 346.050 ;
        RECT 946.950 345.600 949.050 346.050 ;
        RECT 913.950 344.400 949.050 345.600 ;
        RECT 913.950 343.950 916.050 344.400 ;
        RECT 946.950 343.950 949.050 344.400 ;
        RECT 964.950 345.600 967.050 346.050 ;
        RECT 997.950 345.600 1000.050 346.050 ;
        RECT 964.950 344.400 1000.050 345.600 ;
        RECT 964.950 343.950 967.050 344.400 ;
        RECT 997.950 343.950 1000.050 344.400 ;
        RECT 43.950 342.600 46.050 343.050 ;
        RECT 55.950 342.600 58.050 343.050 ;
        RECT 43.950 341.400 58.050 342.600 ;
        RECT 43.950 340.950 46.050 341.400 ;
        RECT 55.950 340.950 58.050 341.400 ;
        RECT 112.950 342.600 115.050 343.050 ;
        RECT 163.950 342.600 166.050 343.050 ;
        RECT 475.950 342.600 478.050 343.050 ;
        RECT 112.950 341.400 166.050 342.600 ;
        RECT 112.950 340.950 115.050 341.400 ;
        RECT 163.950 340.950 166.050 341.400 ;
        RECT 449.400 341.400 478.050 342.600 ;
        RECT 449.400 340.200 450.600 341.400 ;
        RECT 475.950 340.950 478.050 341.400 ;
        RECT 523.950 342.600 526.050 343.050 ;
        RECT 529.950 342.600 532.050 343.050 ;
        RECT 595.950 342.600 598.050 343.050 ;
        RECT 523.950 341.400 532.050 342.600 ;
        RECT 523.950 340.950 526.050 341.400 ;
        RECT 529.950 340.950 532.050 341.400 ;
        RECT 566.400 341.400 598.050 342.600 ;
        RECT 16.950 339.600 19.050 340.200 ;
        RECT 70.950 339.600 73.050 340.050 ;
        RECT 16.950 338.400 73.050 339.600 ;
        RECT 16.950 338.100 19.050 338.400 ;
        RECT 70.950 337.950 73.050 338.400 ;
        RECT 85.950 339.600 88.050 340.200 ;
        RECT 124.950 339.600 127.050 340.200 ;
        RECT 142.950 339.750 145.050 340.200 ;
        RECT 151.950 339.750 154.050 340.200 ;
        RECT 142.950 339.600 154.050 339.750 ;
        RECT 85.950 338.400 108.600 339.600 ;
        RECT 85.950 338.100 88.050 338.400 ;
        RECT 107.400 333.900 108.600 338.400 ;
        RECT 124.950 338.550 154.050 339.600 ;
        RECT 124.950 338.400 145.050 338.550 ;
        RECT 124.950 338.100 127.050 338.400 ;
        RECT 142.950 338.100 145.050 338.400 ;
        RECT 151.950 338.100 154.050 338.550 ;
        RECT 169.950 339.600 172.050 340.200 ;
        RECT 235.950 339.600 238.050 340.200 ;
        RECT 244.950 339.600 247.050 340.050 ;
        RECT 169.950 338.400 247.050 339.600 ;
        RECT 169.950 338.100 172.050 338.400 ;
        RECT 235.950 338.100 238.050 338.400 ;
        RECT 244.950 337.950 247.050 338.400 ;
        RECT 280.950 338.100 283.050 340.200 ;
        RECT 286.950 339.750 289.050 340.200 ;
        RECT 292.950 339.750 295.050 340.200 ;
        RECT 286.950 338.550 295.050 339.750 ;
        RECT 286.950 338.100 289.050 338.550 ;
        RECT 292.950 338.100 295.050 338.550 ;
        RECT 304.950 339.600 307.050 340.200 ;
        RECT 313.950 339.600 316.050 340.050 ;
        RECT 304.950 338.400 316.050 339.600 ;
        RECT 304.950 338.100 307.050 338.400 ;
        RECT 281.400 336.600 282.600 338.100 ;
        RECT 313.950 337.950 316.050 338.400 ;
        RECT 331.950 339.600 334.050 340.200 ;
        RECT 331.950 338.400 351.600 339.600 ;
        RECT 331.950 338.100 334.050 338.400 ;
        RECT 281.400 335.400 291.600 336.600 ;
        RECT 19.950 333.600 22.050 333.900 ;
        RECT 34.950 333.600 37.050 333.900 ;
        RECT 19.950 332.400 48.600 333.600 ;
        RECT 19.950 331.800 22.050 332.400 ;
        RECT 34.950 331.800 37.050 332.400 ;
        RECT 47.400 330.600 48.600 332.400 ;
        RECT 70.950 333.450 73.050 333.900 ;
        RECT 82.950 333.450 85.050 333.900 ;
        RECT 70.950 332.250 85.050 333.450 ;
        RECT 70.950 331.800 73.050 332.250 ;
        RECT 82.950 331.800 85.050 332.250 ;
        RECT 106.950 331.800 109.050 333.900 ;
        RECT 151.950 333.600 154.050 334.050 ;
        RECT 166.950 333.600 169.050 333.900 ;
        RECT 151.950 332.400 169.050 333.600 ;
        RECT 151.950 331.950 154.050 332.400 ;
        RECT 166.950 331.800 169.050 332.400 ;
        RECT 175.950 333.450 178.050 333.900 ;
        RECT 190.950 333.450 193.050 333.900 ;
        RECT 175.950 332.250 193.050 333.450 ;
        RECT 175.950 331.800 178.050 332.250 ;
        RECT 190.950 331.800 193.050 332.250 ;
        RECT 199.950 333.450 202.050 333.900 ;
        RECT 205.950 333.450 208.050 333.900 ;
        RECT 199.950 332.250 208.050 333.450 ;
        RECT 199.950 331.800 202.050 332.250 ;
        RECT 205.950 331.800 208.050 332.250 ;
        RECT 238.950 333.450 241.050 333.900 ;
        RECT 250.950 333.450 253.050 333.900 ;
        RECT 238.950 332.250 253.050 333.450 ;
        RECT 290.400 333.600 291.600 335.400 ;
        RECT 350.400 333.900 351.600 338.400 ;
        RECT 352.950 337.950 355.050 340.050 ;
        RECT 367.950 338.100 370.050 340.200 ;
        RECT 430.950 339.750 433.050 340.200 ;
        RECT 448.950 339.750 451.050 340.200 ;
        RECT 430.950 338.550 451.050 339.750 ;
        RECT 430.950 338.100 433.050 338.550 ;
        RECT 448.950 338.100 451.050 338.550 ;
        RECT 353.400 334.050 354.600 337.950 ;
        RECT 307.950 333.600 310.050 333.900 ;
        RECT 290.400 332.400 310.050 333.600 ;
        RECT 238.950 331.800 241.050 332.250 ;
        RECT 250.950 331.800 253.050 332.250 ;
        RECT 307.950 331.800 310.050 332.400 ;
        RECT 313.950 333.450 316.050 333.900 ;
        RECT 328.950 333.450 331.050 333.900 ;
        RECT 313.950 332.250 331.050 333.450 ;
        RECT 313.950 331.800 316.050 332.250 ;
        RECT 328.950 331.800 331.050 332.250 ;
        RECT 349.800 331.800 351.900 333.900 ;
        RECT 352.950 331.950 355.050 334.050 ;
        RECT 368.400 333.600 369.600 338.100 ;
        RECT 566.400 336.600 567.600 341.400 ;
        RECT 595.950 340.950 598.050 341.400 ;
        RECT 604.950 342.600 607.050 343.050 ;
        RECT 625.950 342.600 628.050 343.050 ;
        RECT 604.950 341.400 628.050 342.600 ;
        RECT 604.950 340.950 607.050 341.400 ;
        RECT 625.950 340.950 628.050 341.400 ;
        RECT 679.950 342.600 682.050 342.900 ;
        RECT 685.950 342.600 688.050 343.050 ;
        RECT 679.950 341.400 688.050 342.600 ;
        RECT 679.950 340.800 682.050 341.400 ;
        RECT 685.950 340.950 688.050 341.400 ;
        RECT 739.950 342.600 742.050 343.050 ;
        RECT 745.950 342.600 748.050 343.050 ;
        RECT 739.950 341.400 748.050 342.600 ;
        RECT 739.950 340.950 742.050 341.400 ;
        RECT 745.950 340.950 748.050 341.400 ;
        RECT 790.950 342.600 793.050 343.050 ;
        RECT 802.950 342.600 805.050 343.050 ;
        RECT 790.950 341.400 805.050 342.600 ;
        RECT 790.950 340.950 793.050 341.400 ;
        RECT 802.950 340.950 805.050 341.400 ;
        RECT 871.950 342.600 874.050 343.050 ;
        RECT 922.950 342.600 925.050 343.050 ;
        RECT 871.950 341.400 925.050 342.600 ;
        RECT 871.950 340.950 874.050 341.400 ;
        RECT 922.950 340.950 925.050 341.400 ;
        RECT 568.950 339.600 571.050 340.200 ;
        RECT 637.950 339.600 640.050 340.050 ;
        RECT 652.950 339.600 655.050 340.200 ;
        RECT 568.950 338.400 636.600 339.600 ;
        RECT 568.950 338.100 571.050 338.400 ;
        RECT 635.400 336.600 636.600 338.400 ;
        RECT 637.950 338.400 655.050 339.600 ;
        RECT 637.950 337.950 640.050 338.400 ;
        RECT 652.950 338.100 655.050 338.400 ;
        RECT 661.950 339.600 664.050 340.050 ;
        RECT 667.950 339.600 670.050 340.200 ;
        RECT 661.950 338.400 670.050 339.600 ;
        RECT 661.950 337.950 664.050 338.400 ;
        RECT 667.950 338.100 670.050 338.400 ;
        RECT 751.950 337.950 754.050 340.050 ;
        RECT 766.950 339.600 769.050 340.050 ;
        RECT 772.950 339.600 775.050 340.050 ;
        RECT 766.950 338.400 775.050 339.600 ;
        RECT 766.950 337.950 769.050 338.400 ;
        RECT 772.950 337.950 775.050 338.400 ;
        RECT 784.950 339.600 787.050 340.200 ;
        RECT 808.950 339.600 811.050 340.200 ;
        RECT 820.950 339.600 823.050 340.050 ;
        RECT 784.950 338.400 807.600 339.600 ;
        RECT 784.950 338.100 787.050 338.400 ;
        RECT 566.400 335.400 573.600 336.600 ;
        RECT 635.400 335.400 645.600 336.600 ;
        RECT 385.950 333.600 388.050 333.900 ;
        RECT 368.400 332.400 388.050 333.600 ;
        RECT 385.950 331.800 388.050 332.400 ;
        RECT 415.950 333.600 418.050 333.900 ;
        RECT 436.950 333.600 439.050 333.900 ;
        RECT 415.950 332.400 441.600 333.600 ;
        RECT 445.950 333.450 448.050 333.900 ;
        RECT 457.950 333.450 460.050 333.900 ;
        RECT 415.950 331.800 418.050 332.400 ;
        RECT 436.950 331.800 439.050 332.400 ;
        RECT 445.950 332.250 460.050 333.450 ;
        RECT 445.950 331.800 448.050 332.250 ;
        RECT 457.950 331.800 460.050 332.250 ;
        RECT 481.950 333.600 484.050 333.900 ;
        RECT 499.950 333.600 502.050 333.900 ;
        RECT 481.950 332.400 502.050 333.600 ;
        RECT 481.950 331.800 484.050 332.400 ;
        RECT 499.950 331.800 502.050 332.400 ;
        RECT 529.950 333.600 532.050 334.050 ;
        RECT 572.400 333.900 573.600 335.400 ;
        RECT 544.950 333.600 547.050 333.900 ;
        RECT 529.950 332.400 547.050 333.600 ;
        RECT 529.950 331.950 532.050 332.400 ;
        RECT 544.950 331.800 547.050 332.400 ;
        RECT 571.950 331.800 574.050 333.900 ;
        RECT 586.950 333.450 589.050 333.900 ;
        RECT 607.950 333.450 610.050 333.900 ;
        RECT 586.950 332.250 610.050 333.450 ;
        RECT 586.950 331.800 589.050 332.250 ;
        RECT 607.950 331.800 610.050 332.250 ;
        RECT 616.950 333.600 619.050 334.050 ;
        RECT 644.400 333.900 645.600 335.400 ;
        RECT 752.400 334.050 753.600 337.950 ;
        RECT 806.400 336.600 807.600 338.400 ;
        RECT 808.950 338.400 823.050 339.600 ;
        RECT 808.950 338.100 811.050 338.400 ;
        RECT 820.950 337.950 823.050 338.400 ;
        RECT 829.950 339.600 832.050 340.200 ;
        RECT 841.950 339.750 844.050 340.200 ;
        RECT 853.950 339.750 856.050 340.200 ;
        RECT 829.950 338.400 840.600 339.600 ;
        RECT 829.950 338.100 832.050 338.400 ;
        RECT 806.400 335.400 828.600 336.600 ;
        RECT 628.950 333.600 631.050 333.900 ;
        RECT 616.950 332.400 631.050 333.600 ;
        RECT 616.950 331.950 619.050 332.400 ;
        RECT 628.950 331.800 631.050 332.400 ;
        RECT 643.950 331.800 646.050 333.900 ;
        RECT 706.950 333.450 709.050 333.900 ;
        RECT 718.950 333.450 721.050 333.900 ;
        RECT 706.950 332.250 721.050 333.450 ;
        RECT 706.950 331.800 709.050 332.250 ;
        RECT 718.950 331.800 721.050 332.250 ;
        RECT 751.950 331.950 754.050 334.050 ;
        RECT 827.400 333.900 828.600 335.400 ;
        RECT 839.400 334.050 840.600 338.400 ;
        RECT 841.950 338.550 856.050 339.750 ;
        RECT 841.950 338.100 844.050 338.550 ;
        RECT 853.950 338.100 856.050 338.550 ;
        RECT 886.950 339.600 889.050 340.200 ;
        RECT 895.950 339.600 898.050 340.050 ;
        RECT 886.950 338.400 898.050 339.600 ;
        RECT 886.950 338.100 889.050 338.400 ;
        RECT 895.950 337.950 898.050 338.400 ;
        RECT 907.950 339.600 910.050 340.200 ;
        RECT 928.950 339.600 931.050 340.050 ;
        RECT 948.000 339.600 952.050 340.050 ;
        RECT 907.950 338.400 931.050 339.600 ;
        RECT 907.950 338.100 910.050 338.400 ;
        RECT 769.950 333.450 772.050 333.900 ;
        RECT 775.950 333.600 778.050 333.900 ;
        RECT 805.950 333.600 808.050 333.900 ;
        RECT 775.950 333.450 808.050 333.600 ;
        RECT 769.950 332.400 808.050 333.450 ;
        RECT 769.950 332.250 778.050 332.400 ;
        RECT 769.950 331.800 772.050 332.250 ;
        RECT 775.950 331.800 778.050 332.250 ;
        RECT 805.950 331.800 808.050 332.400 ;
        RECT 826.950 331.800 829.050 333.900 ;
        RECT 838.950 331.950 841.050 334.050 ;
        RECT 871.950 333.450 874.050 333.900 ;
        RECT 877.950 333.450 880.050 333.900 ;
        RECT 871.950 332.250 880.050 333.450 ;
        RECT 908.400 333.600 909.600 338.100 ;
        RECT 928.950 337.950 931.050 338.400 ;
        RECT 947.400 337.950 952.050 339.600 ;
        RECT 955.950 339.600 958.050 340.050 ;
        RECT 961.950 339.600 964.050 340.200 ;
        RECT 955.950 338.400 964.050 339.600 ;
        RECT 955.950 337.950 958.050 338.400 ;
        RECT 961.950 338.100 964.050 338.400 ;
        RECT 967.950 339.600 970.050 340.050 ;
        RECT 973.950 339.600 976.050 340.050 ;
        RECT 967.950 338.400 976.050 339.600 ;
        RECT 967.950 337.950 970.050 338.400 ;
        RECT 973.950 337.950 976.050 338.400 ;
        RECT 925.950 333.600 928.050 333.900 ;
        RECT 908.400 332.400 928.050 333.600 ;
        RECT 871.950 331.800 874.050 332.250 ;
        RECT 877.950 331.800 880.050 332.250 ;
        RECT 925.950 331.800 928.050 332.400 ;
        RECT 931.950 333.600 934.050 334.050 ;
        RECT 937.950 333.600 940.050 334.050 ;
        RECT 947.400 333.900 948.600 337.950 ;
        RECT 931.950 332.400 940.050 333.600 ;
        RECT 931.950 331.950 934.050 332.400 ;
        RECT 937.950 331.950 940.050 332.400 ;
        RECT 946.950 331.800 949.050 333.900 ;
        RECT 952.950 333.450 955.050 333.900 ;
        RECT 964.950 333.450 967.050 333.900 ;
        RECT 952.950 332.250 967.050 333.450 ;
        RECT 952.950 331.800 955.050 332.250 ;
        RECT 964.950 331.800 967.050 332.250 ;
        RECT 976.950 333.600 979.050 334.050 ;
        RECT 994.950 333.600 997.050 333.900 ;
        RECT 976.950 332.400 997.050 333.600 ;
        RECT 976.950 331.950 979.050 332.400 ;
        RECT 994.950 331.800 997.050 332.400 ;
        RECT 64.950 330.600 67.050 331.050 ;
        RECT 47.400 329.400 67.050 330.600 ;
        RECT 64.950 328.950 67.050 329.400 ;
        RECT 160.950 330.600 163.050 331.050 ;
        RECT 220.950 330.600 223.050 331.050 ;
        RECT 301.950 330.600 304.050 331.050 ;
        RECT 160.950 329.400 223.050 330.600 ;
        RECT 160.950 328.950 163.050 329.400 ;
        RECT 220.950 328.950 223.050 329.400 ;
        RECT 260.400 329.400 304.050 330.600 ;
        RECT 260.400 328.050 261.600 329.400 ;
        RECT 301.950 328.950 304.050 329.400 ;
        RECT 391.950 330.600 394.050 331.050 ;
        RECT 403.950 330.600 406.050 331.050 ;
        RECT 391.950 329.400 406.050 330.600 ;
        RECT 391.950 328.950 394.050 329.400 ;
        RECT 403.950 328.950 406.050 329.400 ;
        RECT 694.950 330.600 697.050 331.050 ;
        RECT 703.950 330.600 706.050 331.050 ;
        RECT 712.950 330.600 715.050 331.050 ;
        RECT 694.950 329.400 715.050 330.600 ;
        RECT 694.950 328.950 697.050 329.400 ;
        RECT 703.950 328.950 706.050 329.400 ;
        RECT 712.950 328.950 715.050 329.400 ;
        RECT 844.950 330.600 847.050 331.050 ;
        RECT 853.950 330.600 856.050 331.050 ;
        RECT 844.950 329.400 856.050 330.600 ;
        RECT 844.950 328.950 847.050 329.400 ;
        RECT 853.950 328.950 856.050 329.400 ;
        RECT 883.950 330.600 886.050 331.050 ;
        RECT 892.950 330.600 895.050 331.050 ;
        RECT 883.950 329.400 895.050 330.600 ;
        RECT 883.950 328.950 886.050 329.400 ;
        RECT 892.950 328.950 895.050 329.400 ;
        RECT 49.950 327.600 52.050 328.050 ;
        RECT 58.950 327.600 61.050 327.900 ;
        RECT 49.950 326.400 61.050 327.600 ;
        RECT 49.950 325.950 52.050 326.400 ;
        RECT 58.950 325.800 61.050 326.400 ;
        RECT 73.950 327.600 76.050 328.050 ;
        RECT 85.800 327.600 87.900 328.050 ;
        RECT 73.950 326.400 87.900 327.600 ;
        RECT 73.950 325.950 76.050 326.400 ;
        RECT 85.800 325.950 87.900 326.400 ;
        RECT 88.950 327.600 91.050 328.050 ;
        RECT 145.950 327.600 148.050 328.050 ;
        RECT 88.950 326.400 148.050 327.600 ;
        RECT 88.950 325.950 91.050 326.400 ;
        RECT 145.950 325.950 148.050 326.400 ;
        RECT 244.950 327.600 247.050 328.050 ;
        RECT 259.950 327.600 262.050 328.050 ;
        RECT 244.950 326.400 262.050 327.600 ;
        RECT 244.950 325.950 247.050 326.400 ;
        RECT 259.950 325.950 262.050 326.400 ;
        RECT 274.950 327.600 277.050 328.050 ;
        RECT 295.950 327.600 298.050 328.050 ;
        RECT 307.950 327.600 310.050 328.050 ;
        RECT 340.950 327.600 343.050 328.050 ;
        RECT 382.800 327.600 384.900 328.050 ;
        RECT 274.950 326.400 384.900 327.600 ;
        RECT 274.950 325.950 277.050 326.400 ;
        RECT 295.950 325.950 298.050 326.400 ;
        RECT 307.950 325.950 310.050 326.400 ;
        RECT 340.950 325.950 343.050 326.400 ;
        RECT 382.800 325.950 384.900 326.400 ;
        RECT 385.950 327.600 388.050 328.050 ;
        RECT 409.950 327.600 412.050 328.050 ;
        RECT 385.950 326.400 412.050 327.600 ;
        RECT 385.950 325.950 388.050 326.400 ;
        RECT 409.950 325.950 412.050 326.400 ;
        RECT 496.950 327.600 499.050 328.050 ;
        RECT 514.950 327.600 517.050 328.050 ;
        RECT 538.950 327.600 541.050 328.050 ;
        RECT 577.950 327.600 580.050 328.050 ;
        RECT 496.950 326.400 580.050 327.600 ;
        RECT 496.950 325.950 499.050 326.400 ;
        RECT 514.950 325.950 517.050 326.400 ;
        RECT 538.950 325.950 541.050 326.400 ;
        RECT 577.950 325.950 580.050 326.400 ;
        RECT 628.950 327.600 631.050 328.050 ;
        RECT 643.950 327.600 646.050 328.050 ;
        RECT 628.950 326.400 646.050 327.600 ;
        RECT 628.950 325.950 631.050 326.400 ;
        RECT 643.950 325.950 646.050 326.400 ;
        RECT 670.950 327.600 673.050 328.050 ;
        RECT 682.950 327.600 685.050 328.050 ;
        RECT 718.950 327.600 721.050 328.050 ;
        RECT 670.950 326.400 721.050 327.600 ;
        RECT 670.950 325.950 673.050 326.400 ;
        RECT 682.950 325.950 685.050 326.400 ;
        RECT 718.950 325.950 721.050 326.400 ;
        RECT 724.950 327.600 727.050 328.050 ;
        RECT 733.950 327.600 736.050 327.900 ;
        RECT 724.950 326.400 736.050 327.600 ;
        RECT 724.950 325.950 727.050 326.400 ;
        RECT 733.950 325.800 736.050 326.400 ;
        RECT 781.950 327.600 784.050 328.050 ;
        RECT 826.950 327.600 829.050 328.050 ;
        RECT 781.950 326.400 829.050 327.600 ;
        RECT 781.950 325.950 784.050 326.400 ;
        RECT 826.950 325.950 829.050 326.400 ;
        RECT 904.950 327.600 907.050 328.050 ;
        RECT 943.950 327.600 946.050 328.050 ;
        RECT 904.950 326.400 946.050 327.600 ;
        RECT 904.950 325.950 907.050 326.400 ;
        RECT 943.950 325.950 946.050 326.400 ;
        RECT 211.950 324.600 214.050 325.050 ;
        RECT 292.950 324.600 295.050 325.050 ;
        RECT 211.950 323.400 295.050 324.600 ;
        RECT 211.950 322.950 214.050 323.400 ;
        RECT 292.950 322.950 295.050 323.400 ;
        RECT 319.950 324.600 322.050 325.050 ;
        RECT 334.950 324.600 337.050 325.050 ;
        RECT 319.950 323.400 337.050 324.600 ;
        RECT 319.950 322.950 322.050 323.400 ;
        RECT 334.950 322.950 337.050 323.400 ;
        RECT 373.950 324.600 376.050 325.050 ;
        RECT 406.950 324.600 409.050 325.050 ;
        RECT 415.950 324.600 418.050 325.050 ;
        RECT 373.950 323.400 418.050 324.600 ;
        RECT 373.950 322.950 376.050 323.400 ;
        RECT 406.950 322.950 409.050 323.400 ;
        RECT 415.950 322.950 418.050 323.400 ;
        RECT 421.950 324.600 424.050 325.050 ;
        RECT 562.950 324.600 565.050 325.050 ;
        RECT 421.950 323.400 565.050 324.600 ;
        RECT 421.950 322.950 424.050 323.400 ;
        RECT 562.950 322.950 565.050 323.400 ;
        RECT 592.950 324.600 595.050 325.050 ;
        RECT 604.950 324.600 607.050 325.050 ;
        RECT 592.950 323.400 607.050 324.600 ;
        RECT 592.950 322.950 595.050 323.400 ;
        RECT 604.950 322.950 607.050 323.400 ;
        RECT 682.950 324.600 685.050 324.900 ;
        RECT 697.950 324.600 700.050 325.050 ;
        RECT 682.950 323.400 700.050 324.600 ;
        RECT 682.950 322.800 685.050 323.400 ;
        RECT 697.950 322.950 700.050 323.400 ;
        RECT 736.950 324.600 739.050 325.050 ;
        RECT 766.950 324.600 769.050 325.050 ;
        RECT 736.950 323.400 769.050 324.600 ;
        RECT 736.950 322.950 739.050 323.400 ;
        RECT 766.950 322.950 769.050 323.400 ;
        RECT 934.950 324.600 937.050 325.050 ;
        RECT 940.950 324.600 943.050 325.050 ;
        RECT 934.950 323.400 943.050 324.600 ;
        RECT 934.950 322.950 937.050 323.400 ;
        RECT 940.950 322.950 943.050 323.400 ;
        RECT 85.950 321.600 88.050 322.050 ;
        RECT 367.950 321.600 370.050 322.050 ;
        RECT 85.950 320.400 318.600 321.600 ;
        RECT 85.950 319.950 88.050 320.400 ;
        RECT 145.950 318.600 148.050 319.050 ;
        RECT 277.950 318.600 280.050 319.050 ;
        RECT 145.950 317.400 280.050 318.600 ;
        RECT 317.400 318.600 318.600 320.400 ;
        RECT 335.400 320.400 370.050 321.600 ;
        RECT 335.400 318.600 336.600 320.400 ;
        RECT 367.950 319.950 370.050 320.400 ;
        RECT 448.950 321.600 451.050 322.050 ;
        RECT 553.950 321.600 556.050 322.050 ;
        RECT 448.950 320.400 556.050 321.600 ;
        RECT 448.950 319.950 451.050 320.400 ;
        RECT 553.950 319.950 556.050 320.400 ;
        RECT 658.950 321.600 661.050 322.050 ;
        RECT 697.950 321.600 700.050 321.900 ;
        RECT 658.950 320.400 700.050 321.600 ;
        RECT 658.950 319.950 661.050 320.400 ;
        RECT 697.950 319.800 700.050 320.400 ;
        RECT 757.950 321.600 760.050 322.050 ;
        RECT 790.950 321.600 793.050 322.050 ;
        RECT 757.950 320.400 793.050 321.600 ;
        RECT 757.950 319.950 760.050 320.400 ;
        RECT 790.950 319.950 793.050 320.400 ;
        RECT 826.950 321.600 829.050 322.050 ;
        RECT 832.950 321.600 835.050 322.050 ;
        RECT 826.950 320.400 835.050 321.600 ;
        RECT 826.950 319.950 829.050 320.400 ;
        RECT 832.950 319.950 835.050 320.400 ;
        RECT 895.950 321.600 898.050 322.050 ;
        RECT 931.950 321.600 934.050 322.050 ;
        RECT 985.950 321.600 988.050 322.050 ;
        RECT 895.950 320.400 988.050 321.600 ;
        RECT 895.950 319.950 898.050 320.400 ;
        RECT 931.950 319.950 934.050 320.400 ;
        RECT 985.950 319.950 988.050 320.400 ;
        RECT 373.950 318.600 376.050 319.050 ;
        RECT 317.400 317.400 336.600 318.600 ;
        RECT 338.400 317.400 376.050 318.600 ;
        RECT 145.950 316.950 148.050 317.400 ;
        RECT 277.950 316.950 280.050 317.400 ;
        RECT 25.950 315.600 28.050 316.050 ;
        RECT 64.950 315.600 67.050 316.050 ;
        RECT 97.950 315.600 100.050 316.050 ;
        RECT 25.950 314.400 100.050 315.600 ;
        RECT 25.950 313.950 28.050 314.400 ;
        RECT 64.950 313.950 67.050 314.400 ;
        RECT 97.950 313.950 100.050 314.400 ;
        RECT 289.950 315.600 292.050 316.050 ;
        RECT 338.400 315.600 339.600 317.400 ;
        RECT 373.950 316.950 376.050 317.400 ;
        RECT 466.950 318.600 469.050 319.050 ;
        RECT 508.950 318.600 511.050 319.050 ;
        RECT 466.950 317.400 511.050 318.600 ;
        RECT 466.950 316.950 469.050 317.400 ;
        RECT 508.950 316.950 511.050 317.400 ;
        RECT 601.950 318.600 604.050 319.050 ;
        RECT 619.950 318.600 622.050 319.050 ;
        RECT 601.950 317.400 622.050 318.600 ;
        RECT 601.950 316.950 604.050 317.400 ;
        RECT 619.950 316.950 622.050 317.400 ;
        RECT 685.950 318.600 688.050 319.050 ;
        RECT 727.950 318.600 730.050 319.050 ;
        RECT 685.950 317.400 730.050 318.600 ;
        RECT 685.950 316.950 688.050 317.400 ;
        RECT 727.950 316.950 730.050 317.400 ;
        RECT 289.950 314.400 339.600 315.600 ;
        RECT 346.950 315.600 349.050 316.050 ;
        RECT 448.950 315.600 451.050 316.050 ;
        RECT 346.950 314.400 451.050 315.600 ;
        RECT 289.950 313.950 292.050 314.400 ;
        RECT 346.950 313.950 349.050 314.400 ;
        RECT 448.950 313.950 451.050 314.400 ;
        RECT 469.950 315.600 472.050 316.050 ;
        RECT 526.950 315.600 529.050 316.050 ;
        RECT 469.950 314.400 529.050 315.600 ;
        RECT 469.950 313.950 472.050 314.400 ;
        RECT 526.950 313.950 529.050 314.400 ;
        RECT 535.950 315.600 538.050 316.050 ;
        RECT 550.950 315.600 553.050 316.050 ;
        RECT 535.950 314.400 553.050 315.600 ;
        RECT 535.950 313.950 538.050 314.400 ;
        RECT 550.950 313.950 553.050 314.400 ;
        RECT 562.950 315.600 565.050 316.050 ;
        RECT 616.950 315.600 619.050 316.050 ;
        RECT 562.950 314.400 619.050 315.600 ;
        RECT 562.950 313.950 565.050 314.400 ;
        RECT 616.950 313.950 619.050 314.400 ;
        RECT 724.950 315.600 727.050 316.050 ;
        RECT 751.950 315.600 754.050 316.050 ;
        RECT 724.950 314.400 754.050 315.600 ;
        RECT 724.950 313.950 727.050 314.400 ;
        RECT 751.950 313.950 754.050 314.400 ;
        RECT 790.950 315.600 793.050 316.050 ;
        RECT 835.950 315.600 838.050 316.050 ;
        RECT 790.950 314.400 838.050 315.600 ;
        RECT 790.950 313.950 793.050 314.400 ;
        RECT 835.950 313.950 838.050 314.400 ;
        RECT 283.950 312.600 286.050 313.050 ;
        RECT 367.950 312.600 370.050 313.050 ;
        RECT 466.950 312.600 469.050 313.050 ;
        RECT 283.950 311.400 363.600 312.600 ;
        RECT 283.950 310.950 286.050 311.400 ;
        RECT 334.950 309.600 337.050 310.050 ;
        RECT 343.950 309.600 346.050 310.050 ;
        RECT 358.950 309.600 361.050 310.050 ;
        RECT 334.950 308.400 361.050 309.600 ;
        RECT 362.400 309.600 363.600 311.400 ;
        RECT 367.950 311.400 469.050 312.600 ;
        RECT 367.950 310.950 370.050 311.400 ;
        RECT 466.950 310.950 469.050 311.400 ;
        RECT 520.950 312.600 523.050 313.050 ;
        RECT 565.950 312.600 568.050 313.050 ;
        RECT 580.950 312.600 583.050 313.050 ;
        RECT 520.950 311.400 583.050 312.600 ;
        RECT 520.950 310.950 523.050 311.400 ;
        RECT 565.950 310.950 568.050 311.400 ;
        RECT 580.950 310.950 583.050 311.400 ;
        RECT 646.950 312.600 649.050 313.050 ;
        RECT 670.950 312.600 673.050 313.050 ;
        RECT 646.950 311.400 673.050 312.600 ;
        RECT 646.950 310.950 649.050 311.400 ;
        RECT 670.950 310.950 673.050 311.400 ;
        RECT 679.950 312.600 682.050 313.050 ;
        RECT 754.950 312.600 757.050 313.050 ;
        RECT 763.950 312.600 766.050 313.050 ;
        RECT 844.950 312.600 847.050 313.050 ;
        RECT 679.950 311.400 847.050 312.600 ;
        RECT 679.950 310.950 682.050 311.400 ;
        RECT 754.950 310.950 757.050 311.400 ;
        RECT 763.950 310.950 766.050 311.400 ;
        RECT 844.950 310.950 847.050 311.400 ;
        RECT 970.950 312.600 973.050 313.050 ;
        RECT 997.950 312.600 1000.050 313.050 ;
        RECT 970.950 311.400 1000.050 312.600 ;
        RECT 970.950 310.950 973.050 311.400 ;
        RECT 997.950 310.950 1000.050 311.400 ;
        RECT 521.400 309.600 522.600 310.950 ;
        RECT 362.400 308.400 522.600 309.600 ;
        RECT 544.950 309.600 547.050 310.050 ;
        RECT 556.950 309.600 559.050 310.050 ;
        RECT 544.950 308.400 559.050 309.600 ;
        RECT 334.950 307.950 337.050 308.400 ;
        RECT 343.950 307.950 346.050 308.400 ;
        RECT 358.950 307.950 361.050 308.400 ;
        RECT 544.950 307.950 547.050 308.400 ;
        RECT 556.950 307.950 559.050 308.400 ;
        RECT 607.950 309.600 610.050 310.050 ;
        RECT 628.950 309.600 631.050 310.050 ;
        RECT 607.950 308.400 631.050 309.600 ;
        RECT 607.950 307.950 610.050 308.400 ;
        RECT 628.950 307.950 631.050 308.400 ;
        RECT 634.950 309.600 637.050 310.050 ;
        RECT 724.950 309.600 727.050 310.050 ;
        RECT 634.950 308.400 727.050 309.600 ;
        RECT 634.950 307.950 637.050 308.400 ;
        RECT 724.950 307.950 727.050 308.400 ;
        RECT 736.950 309.600 739.050 310.050 ;
        RECT 745.950 309.600 748.050 310.050 ;
        RECT 736.950 308.400 748.050 309.600 ;
        RECT 736.950 307.950 739.050 308.400 ;
        RECT 745.950 307.950 748.050 308.400 ;
        RECT 799.950 309.600 802.050 310.050 ;
        RECT 817.950 309.600 820.050 310.050 ;
        RECT 841.950 309.600 844.050 310.050 ;
        RECT 799.950 308.400 844.050 309.600 ;
        RECT 799.950 307.950 802.050 308.400 ;
        RECT 817.950 307.950 820.050 308.400 ;
        RECT 841.950 307.950 844.050 308.400 ;
        RECT 88.950 306.600 91.050 307.050 ;
        RECT 283.950 306.600 286.050 307.050 ;
        RECT 88.950 305.400 286.050 306.600 ;
        RECT 88.950 304.950 91.050 305.400 ;
        RECT 283.950 304.950 286.050 305.400 ;
        RECT 451.950 306.600 454.050 307.050 ;
        RECT 472.950 306.600 475.050 307.050 ;
        RECT 451.950 305.400 475.050 306.600 ;
        RECT 451.950 304.950 454.050 305.400 ;
        RECT 472.950 304.950 475.050 305.400 ;
        RECT 520.950 306.600 523.050 306.900 ;
        RECT 529.950 306.600 532.050 307.050 ;
        RECT 520.950 305.400 532.050 306.600 ;
        RECT 520.950 304.800 523.050 305.400 ;
        RECT 529.950 304.950 532.050 305.400 ;
        RECT 598.950 306.600 601.050 307.050 ;
        RECT 607.950 306.600 610.050 306.900 ;
        RECT 598.950 305.400 610.050 306.600 ;
        RECT 598.950 304.950 601.050 305.400 ;
        RECT 607.950 304.800 610.050 305.400 ;
        RECT 691.950 306.600 694.050 307.050 ;
        RECT 760.950 306.600 763.050 307.050 ;
        RECT 691.950 305.400 763.050 306.600 ;
        RECT 691.950 304.950 694.050 305.400 ;
        RECT 760.950 304.950 763.050 305.400 ;
        RECT 820.950 306.600 823.050 307.050 ;
        RECT 874.950 306.600 877.050 307.050 ;
        RECT 820.950 305.400 877.050 306.600 ;
        RECT 820.950 304.950 823.050 305.400 ;
        RECT 874.950 304.950 877.050 305.400 ;
        RECT 916.950 306.600 919.050 307.050 ;
        RECT 964.950 306.600 967.050 307.050 ;
        RECT 916.950 305.400 967.050 306.600 ;
        RECT 916.950 304.950 919.050 305.400 ;
        RECT 964.950 304.950 967.050 305.400 ;
        RECT 115.950 303.600 118.050 304.050 ;
        RECT 157.950 303.600 160.050 304.050 ;
        RECT 115.950 302.400 160.050 303.600 ;
        RECT 115.950 301.950 118.050 302.400 ;
        RECT 157.950 301.950 160.050 302.400 ;
        RECT 175.950 303.600 178.050 304.050 ;
        RECT 268.950 303.600 271.050 304.050 ;
        RECT 175.950 302.400 271.050 303.600 ;
        RECT 175.950 301.950 178.050 302.400 ;
        RECT 268.950 301.950 271.050 302.400 ;
        RECT 484.950 303.600 487.050 304.050 ;
        RECT 502.950 303.600 505.050 304.050 ;
        RECT 484.950 302.400 505.050 303.600 ;
        RECT 484.950 301.950 487.050 302.400 ;
        RECT 502.950 301.950 505.050 302.400 ;
        RECT 577.950 303.600 580.050 304.050 ;
        RECT 595.950 303.600 598.050 304.050 ;
        RECT 577.950 302.400 598.050 303.600 ;
        RECT 577.950 301.950 580.050 302.400 ;
        RECT 595.950 301.950 598.050 302.400 ;
        RECT 610.950 303.600 613.050 304.050 ;
        RECT 646.950 303.600 649.050 304.050 ;
        RECT 610.950 302.400 649.050 303.600 ;
        RECT 610.950 301.950 613.050 302.400 ;
        RECT 646.950 301.950 649.050 302.400 ;
        RECT 919.950 303.600 922.050 304.050 ;
        RECT 961.950 303.600 964.050 304.050 ;
        RECT 919.950 302.400 964.050 303.600 ;
        RECT 919.950 301.950 922.050 302.400 ;
        RECT 961.950 301.950 964.050 302.400 ;
        RECT 991.950 303.600 994.050 304.050 ;
        RECT 1000.950 303.600 1003.050 304.050 ;
        RECT 991.950 302.400 1003.050 303.600 ;
        RECT 991.950 301.950 994.050 302.400 ;
        RECT 1000.950 301.950 1003.050 302.400 ;
        RECT 439.950 300.600 442.050 301.050 ;
        RECT 451.950 300.600 454.050 301.050 ;
        RECT 439.950 299.400 454.050 300.600 ;
        RECT 439.950 298.950 442.050 299.400 ;
        RECT 451.950 298.950 454.050 299.400 ;
        RECT 508.950 300.600 511.050 301.050 ;
        RECT 598.950 300.600 601.050 301.050 ;
        RECT 508.950 299.400 543.600 300.600 ;
        RECT 508.950 298.950 511.050 299.400 ;
        RECT 292.950 297.600 295.050 298.050 ;
        RECT 346.950 297.600 349.050 298.050 ;
        RECT 292.950 296.400 349.050 297.600 ;
        RECT 292.950 295.950 295.050 296.400 ;
        RECT 346.950 295.950 349.050 296.400 ;
        RECT 355.950 295.950 358.050 298.050 ;
        RECT 505.950 297.600 508.050 298.050 ;
        RECT 523.950 297.600 526.050 298.050 ;
        RECT 505.950 296.400 526.050 297.600 ;
        RECT 542.400 297.600 543.600 299.400 ;
        RECT 584.400 299.400 601.050 300.600 ;
        RECT 584.400 297.600 585.600 299.400 ;
        RECT 598.950 298.950 601.050 299.400 ;
        RECT 631.950 300.600 634.050 301.050 ;
        RECT 688.950 300.600 691.050 301.050 ;
        RECT 631.950 299.400 691.050 300.600 ;
        RECT 631.950 298.950 634.050 299.400 ;
        RECT 688.950 298.950 691.050 299.400 ;
        RECT 697.950 300.600 700.050 301.050 ;
        RECT 703.950 300.600 706.050 301.050 ;
        RECT 805.950 300.600 808.050 301.050 ;
        RECT 697.950 299.400 808.050 300.600 ;
        RECT 697.950 298.950 700.050 299.400 ;
        RECT 703.950 298.950 706.050 299.400 ;
        RECT 805.950 298.950 808.050 299.400 ;
        RECT 838.950 300.600 841.050 301.050 ;
        RECT 880.950 300.600 883.050 301.050 ;
        RECT 895.950 300.600 898.050 301.050 ;
        RECT 838.950 299.400 898.050 300.600 ;
        RECT 838.950 298.950 841.050 299.400 ;
        RECT 880.950 298.950 883.050 299.400 ;
        RECT 895.950 298.950 898.050 299.400 ;
        RECT 904.950 300.600 907.050 301.050 ;
        RECT 949.950 300.600 952.050 301.050 ;
        RECT 904.950 299.400 952.050 300.600 ;
        RECT 904.950 298.950 907.050 299.400 ;
        RECT 949.950 298.950 952.050 299.400 ;
        RECT 955.950 300.600 958.050 301.050 ;
        RECT 964.950 300.600 967.050 301.050 ;
        RECT 955.950 299.400 967.050 300.600 ;
        RECT 955.950 298.950 958.050 299.400 ;
        RECT 964.950 298.950 967.050 299.400 ;
        RECT 542.400 296.400 585.600 297.600 ;
        RECT 670.950 297.600 673.050 298.050 ;
        RECT 697.950 297.600 700.050 297.900 ;
        RECT 670.950 296.400 700.050 297.600 ;
        RECT 505.950 295.950 508.050 296.400 ;
        RECT 523.950 295.950 526.050 296.400 ;
        RECT 670.950 295.950 673.050 296.400 ;
        RECT 34.950 294.750 37.050 295.200 ;
        RECT 43.950 294.750 46.050 295.200 ;
        RECT 34.950 293.550 46.050 294.750 ;
        RECT 34.950 293.100 37.050 293.550 ;
        RECT 43.950 293.100 46.050 293.550 ;
        RECT 127.950 294.600 130.050 295.200 ;
        RECT 142.950 294.600 145.050 295.200 ;
        RECT 163.950 294.600 166.050 295.050 ;
        RECT 127.950 293.400 166.050 294.600 ;
        RECT 127.950 293.100 130.050 293.400 ;
        RECT 142.950 293.100 145.050 293.400 ;
        RECT 163.950 292.950 166.050 293.400 ;
        RECT 229.950 294.750 232.050 295.200 ;
        RECT 244.950 294.750 247.050 295.200 ;
        RECT 229.950 293.550 247.050 294.750 ;
        RECT 229.950 293.100 232.050 293.550 ;
        RECT 244.950 293.100 247.050 293.550 ;
        RECT 253.950 294.750 256.050 295.200 ;
        RECT 259.950 294.750 262.050 295.200 ;
        RECT 253.950 293.550 262.050 294.750 ;
        RECT 283.950 294.600 286.050 295.200 ;
        RECT 253.950 293.100 256.050 293.550 ;
        RECT 259.950 293.100 262.050 293.550 ;
        RECT 266.400 293.400 286.050 294.600 ;
        RECT 61.950 288.600 64.050 289.050 ;
        RECT 67.950 288.600 70.050 288.900 ;
        RECT 61.950 288.450 70.050 288.600 ;
        RECT 73.950 288.450 76.050 288.900 ;
        RECT 61.950 287.400 76.050 288.450 ;
        RECT 61.950 286.950 64.050 287.400 ;
        RECT 67.950 287.250 76.050 287.400 ;
        RECT 67.950 286.800 70.050 287.250 ;
        RECT 73.950 286.800 76.050 287.250 ;
        RECT 106.950 288.450 109.050 288.900 ;
        RECT 112.950 288.450 115.050 289.050 ;
        RECT 124.950 288.450 127.050 288.900 ;
        RECT 106.950 287.250 127.050 288.450 ;
        RECT 106.950 286.800 109.050 287.250 ;
        RECT 112.950 286.950 115.050 287.250 ;
        RECT 124.950 286.800 127.050 287.250 ;
        RECT 214.950 288.450 217.050 288.900 ;
        RECT 223.950 288.450 226.050 288.900 ;
        RECT 214.950 287.250 226.050 288.450 ;
        RECT 214.950 286.800 217.050 287.250 ;
        RECT 223.950 286.800 226.050 287.250 ;
        RECT 241.950 288.600 244.050 288.900 ;
        RECT 250.950 288.600 253.050 289.050 ;
        RECT 241.950 287.400 253.050 288.600 ;
        RECT 241.950 286.800 244.050 287.400 ;
        RECT 250.950 286.950 253.050 287.400 ;
        RECT 262.950 288.600 265.050 288.900 ;
        RECT 266.400 288.600 267.600 293.400 ;
        RECT 283.950 293.100 286.050 293.400 ;
        RECT 313.950 294.750 316.050 295.200 ;
        RECT 322.950 294.750 325.050 295.200 ;
        RECT 313.950 293.550 325.050 294.750 ;
        RECT 313.950 293.100 316.050 293.550 ;
        RECT 322.950 293.100 325.050 293.550 ;
        RECT 349.950 294.600 352.050 295.200 ;
        RECT 349.950 293.400 354.600 294.600 ;
        RECT 349.950 293.100 352.050 293.400 ;
        RECT 334.950 291.600 337.050 292.050 ;
        RECT 320.400 290.400 337.050 291.600 ;
        RECT 320.400 288.900 321.600 290.400 ;
        RECT 334.950 289.950 337.050 290.400 ;
        RECT 262.950 287.400 267.600 288.600 ;
        RECT 262.950 286.800 265.050 287.400 ;
        RECT 319.950 286.800 322.050 288.900 ;
        RECT 337.950 288.600 340.050 289.050 ;
        RECT 346.950 288.600 349.050 288.900 ;
        RECT 337.950 287.400 349.050 288.600 ;
        RECT 353.400 288.600 354.600 293.400 ;
        RECT 356.400 291.600 357.600 295.950 ;
        RECT 697.950 295.800 700.050 296.400 ;
        RECT 712.950 297.600 715.050 298.050 ;
        RECT 727.950 297.600 730.050 297.900 ;
        RECT 712.950 296.400 730.050 297.600 ;
        RECT 712.950 295.950 715.050 296.400 ;
        RECT 727.950 295.800 730.050 296.400 ;
        RECT 736.950 297.600 739.050 298.050 ;
        RECT 787.950 297.600 790.050 298.050 ;
        RECT 736.950 296.400 790.050 297.600 ;
        RECT 736.950 295.950 739.050 296.400 ;
        RECT 787.950 295.950 790.050 296.400 ;
        RECT 961.950 297.600 964.050 298.050 ;
        RECT 982.950 297.600 985.050 297.900 ;
        RECT 961.950 296.400 985.050 297.600 ;
        RECT 961.950 295.950 964.050 296.400 ;
        RECT 982.950 295.800 985.050 296.400 ;
        RECT 994.950 295.950 997.050 298.050 ;
        RECT 364.950 294.750 367.050 295.200 ;
        RECT 373.950 294.750 376.050 295.200 ;
        RECT 364.950 293.550 376.050 294.750 ;
        RECT 364.950 293.100 367.050 293.550 ;
        RECT 373.950 293.100 376.050 293.550 ;
        RECT 382.950 294.600 385.050 295.200 ;
        RECT 391.950 294.600 394.050 295.200 ;
        RECT 382.950 293.400 394.050 294.600 ;
        RECT 382.950 293.100 385.050 293.400 ;
        RECT 391.950 293.100 394.050 293.400 ;
        RECT 400.950 294.600 403.050 295.200 ;
        RECT 430.950 294.750 433.050 295.200 ;
        RECT 436.950 294.750 439.050 295.200 ;
        RECT 400.950 293.400 429.600 294.600 ;
        RECT 400.950 293.100 403.050 293.400 ;
        RECT 428.400 291.600 429.600 293.400 ;
        RECT 430.950 293.550 439.050 294.750 ;
        RECT 430.950 293.100 433.050 293.550 ;
        RECT 436.950 293.100 439.050 293.550 ;
        RECT 442.950 294.600 445.050 295.200 ;
        RECT 460.950 294.600 463.050 295.200 ;
        RECT 499.950 294.600 502.050 295.050 ;
        RECT 442.950 293.400 463.050 294.600 ;
        RECT 442.950 293.100 445.050 293.400 ;
        RECT 460.950 293.100 463.050 293.400 ;
        RECT 488.400 293.400 502.050 294.600 ;
        RECT 356.400 290.400 360.600 291.600 ;
        RECT 428.400 290.400 435.600 291.600 ;
        RECT 355.950 288.600 358.050 288.900 ;
        RECT 353.400 287.400 358.050 288.600 ;
        RECT 359.400 288.600 360.600 290.400 ;
        RECT 370.950 288.600 373.050 289.050 ;
        RECT 359.400 287.400 373.050 288.600 ;
        RECT 434.400 288.600 435.600 290.400 ;
        RECT 488.400 288.900 489.600 293.400 ;
        RECT 499.950 292.950 502.050 293.400 ;
        RECT 586.950 293.100 589.050 295.200 ;
        RECT 619.950 294.600 622.050 295.200 ;
        RECT 605.400 293.400 622.050 294.600 ;
        RECT 550.950 291.600 553.050 292.050 ;
        RECT 577.950 291.600 580.050 292.050 ;
        RECT 497.400 290.400 507.600 291.600 ;
        RECT 497.400 289.050 498.600 290.400 ;
        RECT 439.950 288.600 442.050 288.900 ;
        RECT 434.400 287.400 442.050 288.600 ;
        RECT 337.950 286.950 340.050 287.400 ;
        RECT 346.950 286.800 349.050 287.400 ;
        RECT 355.950 286.800 358.050 287.400 ;
        RECT 370.950 286.950 373.050 287.400 ;
        RECT 439.950 286.800 442.050 287.400 ;
        RECT 469.950 288.450 472.050 288.900 ;
        RECT 481.950 288.450 484.050 288.900 ;
        RECT 469.950 287.250 484.050 288.450 ;
        RECT 469.950 286.800 472.050 287.250 ;
        RECT 481.950 286.800 484.050 287.250 ;
        RECT 487.950 286.800 490.050 288.900 ;
        RECT 493.950 287.400 498.600 289.050 ;
        RECT 506.400 288.900 507.600 290.400 ;
        RECT 550.950 290.400 580.050 291.600 ;
        RECT 587.400 291.600 588.600 293.100 ;
        RECT 605.400 291.600 606.600 293.400 ;
        RECT 619.950 293.100 622.050 293.400 ;
        RECT 628.950 292.950 631.050 295.050 ;
        RECT 637.950 294.600 640.050 295.050 ;
        RECT 661.950 294.600 664.050 295.050 ;
        RECT 691.950 294.600 694.050 295.050 ;
        RECT 637.950 293.400 664.050 294.600 ;
        RECT 637.950 292.950 640.050 293.400 ;
        RECT 661.950 292.950 664.050 293.400 ;
        RECT 674.400 293.400 694.050 294.600 ;
        RECT 587.400 290.400 606.600 291.600 ;
        RECT 550.950 289.950 553.050 290.400 ;
        RECT 577.950 289.950 580.050 290.400 ;
        RECT 505.950 288.600 508.050 288.900 ;
        RECT 511.950 288.600 514.050 288.900 ;
        RECT 505.950 287.400 514.050 288.600 ;
        RECT 493.950 286.950 498.000 287.400 ;
        RECT 505.950 286.800 508.050 287.400 ;
        RECT 511.950 286.800 514.050 287.400 ;
        RECT 559.950 288.600 562.050 288.900 ;
        RECT 568.950 288.600 571.050 288.900 ;
        RECT 559.950 287.400 571.050 288.600 ;
        RECT 629.400 288.600 630.600 292.950 ;
        RECT 674.400 288.900 675.600 293.400 ;
        RECT 691.950 292.950 694.050 293.400 ;
        RECT 709.950 294.750 712.050 295.200 ;
        RECT 721.950 294.750 724.050 295.200 ;
        RECT 709.950 293.550 724.050 294.750 ;
        RECT 709.950 293.100 712.050 293.550 ;
        RECT 721.950 293.100 724.050 293.550 ;
        RECT 739.950 292.950 742.050 295.050 ;
        RECT 751.950 294.600 754.050 295.050 ;
        RECT 775.950 294.600 778.050 295.050 ;
        RECT 751.950 293.400 778.050 294.600 ;
        RECT 751.950 292.950 754.050 293.400 ;
        RECT 775.950 292.950 778.050 293.400 ;
        RECT 811.950 294.600 814.050 295.200 ;
        RECT 835.950 294.600 838.050 295.200 ;
        RECT 811.950 293.400 838.050 294.600 ;
        RECT 811.950 293.100 814.050 293.400 ;
        RECT 835.950 293.100 838.050 293.400 ;
        RECT 874.950 294.600 877.050 295.200 ;
        RECT 892.950 294.600 895.050 295.050 ;
        RECT 874.950 293.400 895.050 294.600 ;
        RECT 874.950 293.100 877.050 293.400 ;
        RECT 892.950 292.950 895.050 293.400 ;
        RECT 916.950 294.750 919.050 295.200 ;
        RECT 925.950 294.750 928.050 295.200 ;
        RECT 916.950 293.550 928.050 294.750 ;
        RECT 916.950 293.100 919.050 293.550 ;
        RECT 925.950 293.100 928.050 293.550 ;
        RECT 931.950 293.100 934.050 295.200 ;
        RECT 955.950 294.600 958.050 295.200 ;
        RECT 973.950 294.600 976.050 295.200 ;
        RECT 955.950 293.400 976.050 294.600 ;
        RECT 955.950 293.100 958.050 293.400 ;
        RECT 973.950 293.100 976.050 293.400 ;
        RECT 646.950 288.600 649.050 288.900 ;
        RECT 629.400 287.400 649.050 288.600 ;
        RECT 559.950 286.800 562.050 287.400 ;
        RECT 568.950 286.800 571.050 287.400 ;
        RECT 646.950 286.800 649.050 287.400 ;
        RECT 673.950 286.800 676.050 288.900 ;
        RECT 682.950 288.600 685.050 289.050 ;
        RECT 688.950 288.600 691.050 289.050 ;
        RECT 682.950 287.400 691.050 288.600 ;
        RECT 682.950 286.950 685.050 287.400 ;
        RECT 688.950 286.950 691.050 287.400 ;
        RECT 700.950 288.600 703.050 288.900 ;
        RECT 718.950 288.600 721.050 288.900 ;
        RECT 700.950 287.400 721.050 288.600 ;
        RECT 740.400 288.600 741.600 292.950 ;
        RECT 932.400 291.600 933.600 293.100 ;
        RECT 800.400 290.400 810.600 291.600 ;
        RECT 932.400 290.400 945.600 291.600 ;
        RECT 742.950 288.600 745.050 288.900 ;
        RECT 740.400 287.400 745.050 288.600 ;
        RECT 700.950 286.800 703.050 287.400 ;
        RECT 718.950 286.800 721.050 287.400 ;
        RECT 742.950 286.800 745.050 287.400 ;
        RECT 784.950 288.600 787.050 288.900 ;
        RECT 800.400 288.600 801.600 290.400 ;
        RECT 784.950 287.400 801.600 288.600 ;
        RECT 809.400 288.600 810.600 290.400 ;
        RECT 829.950 288.600 832.050 288.900 ;
        RECT 856.950 288.600 859.050 288.900 ;
        RECT 809.400 287.400 859.050 288.600 ;
        RECT 784.950 286.800 787.050 287.400 ;
        RECT 829.950 286.800 832.050 287.400 ;
        RECT 856.950 286.800 859.050 287.400 ;
        RECT 892.950 288.450 895.050 288.900 ;
        RECT 901.950 288.450 904.050 288.900 ;
        RECT 892.950 287.250 904.050 288.450 ;
        RECT 892.950 286.800 895.050 287.250 ;
        RECT 901.950 286.800 904.050 287.250 ;
        RECT 928.950 288.600 931.050 288.900 ;
        RECT 940.950 288.600 943.050 289.050 ;
        RECT 928.950 287.400 943.050 288.600 ;
        RECT 944.400 288.600 945.600 290.400 ;
        RECT 995.400 288.900 996.600 295.950 ;
        RECT 946.950 288.600 949.050 288.900 ;
        RECT 944.400 288.450 949.050 288.600 ;
        RECT 976.950 288.450 979.050 288.900 ;
        RECT 944.400 287.400 979.050 288.450 ;
        RECT 928.950 286.800 931.050 287.400 ;
        RECT 940.950 286.950 943.050 287.400 ;
        RECT 946.950 287.250 979.050 287.400 ;
        RECT 946.950 286.800 949.050 287.250 ;
        RECT 976.950 286.800 979.050 287.250 ;
        RECT 994.950 286.800 997.050 288.900 ;
        RECT 220.950 285.600 223.050 286.050 ;
        RECT 232.950 285.600 235.050 286.050 ;
        RECT 220.950 284.400 235.050 285.600 ;
        RECT 220.950 283.950 223.050 284.400 ;
        RECT 232.950 283.950 235.050 284.400 ;
        RECT 418.950 285.600 421.050 286.050 ;
        RECT 424.950 285.600 427.050 286.050 ;
        RECT 463.950 285.600 466.050 286.050 ;
        RECT 418.950 284.400 466.050 285.600 ;
        RECT 418.950 283.950 421.050 284.400 ;
        RECT 424.950 283.950 427.050 284.400 ;
        RECT 463.950 283.950 466.050 284.400 ;
        RECT 508.950 285.600 511.050 286.050 ;
        RECT 544.950 285.600 547.050 286.050 ;
        RECT 508.950 284.400 547.050 285.600 ;
        RECT 508.950 283.950 511.050 284.400 ;
        RECT 544.950 283.950 547.050 284.400 ;
        RECT 808.950 285.600 811.050 286.050 ;
        RECT 817.950 285.600 820.050 286.050 ;
        RECT 808.950 284.400 820.050 285.600 ;
        RECT 808.950 283.950 811.050 284.400 ;
        RECT 817.950 283.950 820.050 284.400 ;
        RECT 982.950 285.600 985.050 286.050 ;
        RECT 997.950 285.600 1000.050 286.050 ;
        RECT 982.950 284.400 1000.050 285.600 ;
        RECT 982.950 283.950 985.050 284.400 ;
        RECT 997.950 283.950 1000.050 284.400 ;
        RECT 124.950 282.600 127.050 283.050 ;
        RECT 136.950 282.600 139.050 283.050 ;
        RECT 145.950 282.600 148.050 283.050 ;
        RECT 124.950 281.400 148.050 282.600 ;
        RECT 124.950 280.950 127.050 281.400 ;
        RECT 136.950 280.950 139.050 281.400 ;
        RECT 145.950 280.950 148.050 281.400 ;
        RECT 172.950 282.600 175.050 283.050 ;
        RECT 253.950 282.600 256.050 283.050 ;
        RECT 172.950 281.400 256.050 282.600 ;
        RECT 172.950 280.950 175.050 281.400 ;
        RECT 253.950 280.950 256.050 281.400 ;
        RECT 325.950 282.600 328.050 283.050 ;
        RECT 364.950 282.600 367.050 283.050 ;
        RECT 325.950 281.400 367.050 282.600 ;
        RECT 325.950 280.950 328.050 281.400 ;
        RECT 364.950 280.950 367.050 281.400 ;
        RECT 382.950 282.600 385.050 283.050 ;
        RECT 430.950 282.600 433.050 283.050 ;
        RECT 382.950 281.400 433.050 282.600 ;
        RECT 382.950 280.950 385.050 281.400 ;
        RECT 430.950 280.950 433.050 281.400 ;
        RECT 445.950 282.600 448.050 283.050 ;
        RECT 451.950 282.600 454.050 283.050 ;
        RECT 445.950 281.400 454.050 282.600 ;
        RECT 445.950 280.950 448.050 281.400 ;
        RECT 451.950 280.950 454.050 281.400 ;
        RECT 622.950 282.600 625.050 283.050 ;
        RECT 670.950 282.600 673.050 283.050 ;
        RECT 685.950 282.600 688.050 283.050 ;
        RECT 622.950 281.400 630.600 282.600 ;
        RECT 622.950 280.950 625.050 281.400 ;
        RECT 52.950 279.600 55.050 280.050 ;
        RECT 79.950 279.600 82.050 280.050 ;
        RECT 91.950 279.600 94.050 280.050 ;
        RECT 52.950 278.400 94.050 279.600 ;
        RECT 52.950 277.950 55.050 278.400 ;
        RECT 79.950 277.950 82.050 278.400 ;
        RECT 91.950 277.950 94.050 278.400 ;
        RECT 157.950 279.600 160.050 280.050 ;
        RECT 172.950 279.600 175.050 279.900 ;
        RECT 157.950 278.400 175.050 279.600 ;
        RECT 157.950 277.950 160.050 278.400 ;
        RECT 172.950 277.800 175.050 278.400 ;
        RECT 214.950 279.600 217.050 280.050 ;
        RECT 229.950 279.600 232.050 280.050 ;
        RECT 214.950 278.400 232.050 279.600 ;
        RECT 214.950 277.950 217.050 278.400 ;
        RECT 229.950 277.950 232.050 278.400 ;
        RECT 262.950 279.600 265.050 280.050 ;
        RECT 289.950 279.600 292.050 280.050 ;
        RECT 262.950 278.400 292.050 279.600 ;
        RECT 262.950 277.950 265.050 278.400 ;
        RECT 289.950 277.950 292.050 278.400 ;
        RECT 334.950 279.600 337.050 280.050 ;
        RECT 346.950 279.600 349.050 280.050 ;
        RECT 334.950 278.400 349.050 279.600 ;
        RECT 334.950 277.950 337.050 278.400 ;
        RECT 346.950 277.950 349.050 278.400 ;
        RECT 391.950 279.600 394.050 280.050 ;
        RECT 421.950 279.600 424.050 280.050 ;
        RECT 391.950 278.400 424.050 279.600 ;
        RECT 391.950 277.950 394.050 278.400 ;
        RECT 421.950 277.950 424.050 278.400 ;
        RECT 433.950 279.600 436.050 280.050 ;
        RECT 508.950 279.600 511.050 280.050 ;
        RECT 433.950 278.400 511.050 279.600 ;
        RECT 433.950 277.950 436.050 278.400 ;
        RECT 508.950 277.950 511.050 278.400 ;
        RECT 541.950 279.600 544.050 280.050 ;
        RECT 553.950 279.600 556.050 280.050 ;
        RECT 541.950 278.400 556.050 279.600 ;
        RECT 541.950 277.950 544.050 278.400 ;
        RECT 553.950 277.950 556.050 278.400 ;
        RECT 565.950 279.600 568.050 280.050 ;
        RECT 601.950 279.600 604.050 280.050 ;
        RECT 613.950 279.600 616.050 280.050 ;
        RECT 565.950 278.400 616.050 279.600 ;
        RECT 629.400 279.600 630.600 281.400 ;
        RECT 670.950 281.400 688.050 282.600 ;
        RECT 670.950 280.950 673.050 281.400 ;
        RECT 685.950 280.950 688.050 281.400 ;
        RECT 694.950 282.600 697.050 283.050 ;
        RECT 709.950 282.600 712.050 283.050 ;
        RECT 694.950 281.400 712.050 282.600 ;
        RECT 694.950 280.950 697.050 281.400 ;
        RECT 709.950 280.950 712.050 281.400 ;
        RECT 769.950 282.600 772.050 283.050 ;
        RECT 802.950 282.600 805.050 283.050 ;
        RECT 769.950 281.400 805.050 282.600 ;
        RECT 769.950 280.950 772.050 281.400 ;
        RECT 802.950 280.950 805.050 281.400 ;
        RECT 889.950 282.600 892.050 283.050 ;
        RECT 901.950 282.600 904.050 283.050 ;
        RECT 889.950 281.400 904.050 282.600 ;
        RECT 889.950 280.950 892.050 281.400 ;
        RECT 901.950 280.950 904.050 281.400 ;
        RECT 982.950 282.600 985.050 282.900 ;
        RECT 1000.950 282.600 1003.050 283.050 ;
        RECT 982.950 281.400 1003.050 282.600 ;
        RECT 982.950 280.800 985.050 281.400 ;
        RECT 1000.950 280.950 1003.050 281.400 ;
        RECT 658.950 279.600 661.050 280.050 ;
        RECT 629.400 278.400 661.050 279.600 ;
        RECT 565.950 277.950 568.050 278.400 ;
        RECT 601.950 277.950 604.050 278.400 ;
        RECT 613.950 277.950 616.050 278.400 ;
        RECT 658.950 277.950 661.050 278.400 ;
        RECT 712.950 279.600 715.050 280.050 ;
        RECT 766.950 279.600 769.050 280.050 ;
        RECT 712.950 278.400 769.050 279.600 ;
        RECT 712.950 277.950 715.050 278.400 ;
        RECT 766.950 277.950 769.050 278.400 ;
        RECT 772.950 279.600 775.050 280.050 ;
        RECT 799.950 279.600 802.050 280.050 ;
        RECT 772.950 278.400 802.050 279.600 ;
        RECT 772.950 277.950 775.050 278.400 ;
        RECT 799.950 277.950 802.050 278.400 ;
        RECT 967.950 279.600 970.050 280.050 ;
        RECT 976.950 279.600 979.050 280.050 ;
        RECT 967.950 278.400 979.050 279.600 ;
        RECT 967.950 277.950 970.050 278.400 ;
        RECT 976.950 277.950 979.050 278.400 ;
        RECT 280.950 276.600 283.050 277.050 ;
        RECT 301.950 276.600 304.050 277.050 ;
        RECT 280.950 275.400 304.050 276.600 ;
        RECT 280.950 274.950 283.050 275.400 ;
        RECT 301.950 274.950 304.050 275.400 ;
        RECT 322.950 276.600 325.050 277.050 ;
        RECT 358.950 276.600 361.050 277.050 ;
        RECT 322.950 275.400 361.050 276.600 ;
        RECT 322.950 274.950 325.050 275.400 ;
        RECT 358.950 274.950 361.050 275.400 ;
        RECT 370.950 276.600 373.050 277.050 ;
        RECT 526.950 276.600 529.050 277.050 ;
        RECT 370.950 275.400 529.050 276.600 ;
        RECT 370.950 274.950 373.050 275.400 ;
        RECT 526.950 274.950 529.050 275.400 ;
        RECT 538.950 276.600 541.050 277.050 ;
        RECT 559.950 276.600 562.050 277.050 ;
        RECT 574.800 276.600 576.900 277.050 ;
        RECT 538.950 275.400 555.600 276.600 ;
        RECT 538.950 274.950 541.050 275.400 ;
        RECT 554.400 274.050 555.600 275.400 ;
        RECT 559.950 275.400 576.900 276.600 ;
        RECT 559.950 274.950 562.050 275.400 ;
        RECT 574.800 274.950 576.900 275.400 ;
        RECT 577.950 276.600 580.050 277.050 ;
        RECT 616.950 276.600 619.050 277.050 ;
        RECT 577.950 275.400 619.050 276.600 ;
        RECT 577.950 274.950 580.050 275.400 ;
        RECT 616.950 274.950 619.050 275.400 ;
        RECT 685.950 276.600 688.050 277.050 ;
        RECT 769.950 276.600 772.050 277.050 ;
        RECT 685.950 275.400 772.050 276.600 ;
        RECT 685.950 274.950 688.050 275.400 ;
        RECT 769.950 274.950 772.050 275.400 ;
        RECT 877.950 276.600 880.050 277.050 ;
        RECT 922.950 276.600 925.050 277.050 ;
        RECT 946.950 276.600 949.050 277.050 ;
        RECT 877.950 275.400 925.050 276.600 ;
        RECT 877.950 274.950 880.050 275.400 ;
        RECT 922.950 274.950 925.050 275.400 ;
        RECT 941.400 275.400 949.050 276.600 ;
        RECT 40.950 273.600 43.050 274.050 ;
        RECT 67.950 273.600 70.050 274.050 ;
        RECT 40.950 272.400 70.050 273.600 ;
        RECT 40.950 271.950 43.050 272.400 ;
        RECT 67.950 271.950 70.050 272.400 ;
        RECT 157.950 273.600 160.050 274.050 ;
        RECT 268.950 273.600 271.050 274.050 ;
        RECT 343.950 273.600 346.050 274.050 ;
        RECT 157.950 272.400 346.050 273.600 ;
        RECT 157.950 271.950 160.050 272.400 ;
        RECT 268.950 271.950 271.050 272.400 ;
        RECT 343.950 271.950 346.050 272.400 ;
        RECT 394.950 273.600 397.050 274.050 ;
        RECT 427.950 273.600 430.050 274.050 ;
        RECT 466.950 273.600 469.050 274.050 ;
        RECT 394.950 272.400 430.050 273.600 ;
        RECT 394.950 271.950 397.050 272.400 ;
        RECT 427.950 271.950 430.050 272.400 ;
        RECT 446.400 272.400 469.050 273.600 ;
        RECT 446.400 271.050 447.600 272.400 ;
        RECT 466.950 271.950 469.050 272.400 ;
        RECT 502.950 273.600 505.050 274.050 ;
        RECT 523.950 273.600 526.050 274.050 ;
        RECT 502.950 272.400 526.050 273.600 ;
        RECT 554.400 272.400 559.050 274.050 ;
        RECT 502.950 271.950 505.050 272.400 ;
        RECT 523.950 271.950 526.050 272.400 ;
        RECT 555.000 271.950 559.050 272.400 ;
        RECT 646.950 273.600 649.050 274.050 ;
        RECT 679.950 273.600 682.050 274.050 ;
        RECT 646.950 272.400 682.050 273.600 ;
        RECT 646.950 271.950 649.050 272.400 ;
        RECT 679.950 271.950 682.050 272.400 ;
        RECT 688.950 273.600 691.050 274.050 ;
        RECT 703.950 273.600 706.050 274.050 ;
        RECT 688.950 272.400 706.050 273.600 ;
        RECT 688.950 271.950 691.050 272.400 ;
        RECT 703.950 271.950 706.050 272.400 ;
        RECT 895.950 273.600 898.050 274.050 ;
        RECT 941.400 273.600 942.600 275.400 ;
        RECT 946.950 274.950 949.050 275.400 ;
        RECT 955.950 276.600 958.050 277.050 ;
        RECT 964.950 276.600 967.050 277.050 ;
        RECT 955.950 275.400 967.050 276.600 ;
        RECT 955.950 274.950 958.050 275.400 ;
        RECT 964.950 274.950 967.050 275.400 ;
        RECT 994.950 276.600 997.050 277.050 ;
        RECT 1009.950 276.600 1012.050 277.050 ;
        RECT 994.950 275.400 1012.050 276.600 ;
        RECT 994.950 274.950 997.050 275.400 ;
        RECT 1009.950 274.950 1012.050 275.400 ;
        RECT 895.950 272.400 942.600 273.600 ;
        RECT 895.950 271.950 898.050 272.400 ;
        RECT 61.950 270.600 64.050 271.050 ;
        RECT 97.950 270.600 100.050 271.050 ;
        RECT 61.950 269.400 100.050 270.600 ;
        RECT 61.950 268.950 64.050 269.400 ;
        RECT 97.950 268.950 100.050 269.400 ;
        RECT 118.950 270.600 121.050 271.050 ;
        RECT 193.950 270.600 196.050 271.050 ;
        RECT 202.950 270.600 205.050 271.050 ;
        RECT 208.950 270.600 211.050 271.050 ;
        RECT 118.950 269.400 211.050 270.600 ;
        RECT 118.950 268.950 121.050 269.400 ;
        RECT 193.950 268.950 196.050 269.400 ;
        RECT 202.950 268.950 205.050 269.400 ;
        RECT 208.950 268.950 211.050 269.400 ;
        RECT 286.950 270.600 289.050 271.050 ;
        RECT 292.950 270.600 295.050 271.050 ;
        RECT 286.950 269.400 295.050 270.600 ;
        RECT 286.950 268.950 289.050 269.400 ;
        RECT 292.950 268.950 295.050 269.400 ;
        RECT 316.950 270.600 319.050 271.050 ;
        RECT 340.950 270.600 343.050 271.050 ;
        RECT 316.950 269.400 343.050 270.600 ;
        RECT 316.950 268.950 319.050 269.400 ;
        RECT 340.950 268.950 343.050 269.400 ;
        RECT 367.950 270.600 370.050 271.050 ;
        RECT 391.950 270.600 394.050 271.050 ;
        RECT 367.950 269.400 394.050 270.600 ;
        RECT 367.950 268.950 370.050 269.400 ;
        RECT 391.950 268.950 394.050 269.400 ;
        RECT 442.950 269.400 447.600 271.050 ;
        RECT 478.950 270.600 481.050 271.050 ;
        RECT 487.950 270.600 490.050 271.050 ;
        RECT 478.950 269.400 490.050 270.600 ;
        RECT 442.950 268.950 447.000 269.400 ;
        RECT 478.950 268.950 481.050 269.400 ;
        RECT 487.950 268.950 490.050 269.400 ;
        RECT 511.950 270.600 514.050 271.050 ;
        RECT 520.950 270.600 523.050 271.050 ;
        RECT 538.950 270.600 541.050 271.050 ;
        RECT 511.950 269.400 541.050 270.600 ;
        RECT 511.950 268.950 514.050 269.400 ;
        RECT 520.950 268.950 523.050 269.400 ;
        RECT 538.950 268.950 541.050 269.400 ;
        RECT 622.950 270.600 625.050 271.050 ;
        RECT 652.950 270.600 655.050 271.050 ;
        RECT 622.950 269.400 655.050 270.600 ;
        RECT 622.950 268.950 625.050 269.400 ;
        RECT 652.950 268.950 655.050 269.400 ;
        RECT 658.950 270.600 661.050 271.050 ;
        RECT 724.950 270.600 727.050 271.050 ;
        RECT 658.950 269.400 727.050 270.600 ;
        RECT 658.950 268.950 661.050 269.400 ;
        RECT 724.950 268.950 727.050 269.400 ;
        RECT 913.950 270.600 916.050 271.050 ;
        RECT 928.950 270.600 931.050 271.050 ;
        RECT 913.950 269.400 931.050 270.600 ;
        RECT 913.950 268.950 916.050 269.400 ;
        RECT 928.950 268.950 931.050 269.400 ;
        RECT 964.950 270.600 967.050 271.050 ;
        RECT 988.950 270.600 991.050 271.050 ;
        RECT 1000.950 270.600 1003.050 271.050 ;
        RECT 964.950 269.400 1003.050 270.600 ;
        RECT 964.950 268.950 967.050 269.400 ;
        RECT 988.950 268.950 991.050 269.400 ;
        RECT 1000.950 268.950 1003.050 269.400 ;
        RECT 121.950 267.600 124.050 268.050 ;
        RECT 148.800 267.600 150.900 268.050 ;
        RECT 121.950 266.400 150.900 267.600 ;
        RECT 121.950 265.950 124.050 266.400 ;
        RECT 148.800 265.950 150.900 266.400 ;
        RECT 151.950 267.600 154.050 268.050 ;
        RECT 190.950 267.600 193.050 268.050 ;
        RECT 151.950 266.400 193.050 267.600 ;
        RECT 151.950 265.950 154.050 266.400 ;
        RECT 190.950 265.950 193.050 266.400 ;
        RECT 427.950 267.600 430.050 268.050 ;
        RECT 439.950 267.600 442.050 268.050 ;
        RECT 427.950 266.400 442.050 267.600 ;
        RECT 427.950 265.950 430.050 266.400 ;
        RECT 439.950 265.950 442.050 266.400 ;
        RECT 499.950 267.600 502.050 268.050 ;
        RECT 541.950 267.600 544.050 268.050 ;
        RECT 499.950 266.400 544.050 267.600 ;
        RECT 499.950 265.950 502.050 266.400 ;
        RECT 541.950 265.950 544.050 266.400 ;
        RECT 556.950 267.600 559.050 268.050 ;
        RECT 565.950 267.600 568.050 268.050 ;
        RECT 556.950 266.400 568.050 267.600 ;
        RECT 556.950 265.950 559.050 266.400 ;
        RECT 565.950 265.950 568.050 266.400 ;
        RECT 583.950 267.600 586.050 268.050 ;
        RECT 589.950 267.600 592.050 268.050 ;
        RECT 583.950 266.400 592.050 267.600 ;
        RECT 583.950 265.950 586.050 266.400 ;
        RECT 589.950 265.950 592.050 266.400 ;
        RECT 775.950 267.600 778.050 268.050 ;
        RECT 787.950 267.600 790.050 268.050 ;
        RECT 817.950 267.600 820.050 268.050 ;
        RECT 775.950 266.400 820.050 267.600 ;
        RECT 775.950 265.950 778.050 266.400 ;
        RECT 787.950 265.950 790.050 266.400 ;
        RECT 817.950 265.950 820.050 266.400 ;
        RECT 877.950 267.600 880.050 268.050 ;
        RECT 895.950 267.600 898.050 268.050 ;
        RECT 877.950 266.400 898.050 267.600 ;
        RECT 877.950 265.950 880.050 266.400 ;
        RECT 895.950 265.950 898.050 266.400 ;
        RECT 16.950 264.600 19.050 265.050 ;
        RECT 31.950 264.600 34.050 265.050 ;
        RECT 16.950 263.400 34.050 264.600 ;
        RECT 16.950 262.950 19.050 263.400 ;
        RECT 31.950 262.950 34.050 263.400 ;
        RECT 46.950 264.600 49.050 265.050 ;
        RECT 61.950 264.600 64.050 265.050 ;
        RECT 46.950 263.400 64.050 264.600 ;
        RECT 46.950 262.950 49.050 263.400 ;
        RECT 61.950 262.950 64.050 263.400 ;
        RECT 226.950 264.600 229.050 265.050 ;
        RECT 250.950 264.600 253.050 265.050 ;
        RECT 226.950 263.400 253.050 264.600 ;
        RECT 226.950 262.950 229.050 263.400 ;
        RECT 250.950 262.950 253.050 263.400 ;
        RECT 307.950 264.600 310.050 265.050 ;
        RECT 325.950 264.600 328.050 265.050 ;
        RECT 307.950 263.400 328.050 264.600 ;
        RECT 307.950 262.950 310.050 263.400 ;
        RECT 325.950 262.950 328.050 263.400 ;
        RECT 391.950 264.600 394.050 265.050 ;
        RECT 406.950 264.600 409.050 265.050 ;
        RECT 391.950 263.400 409.050 264.600 ;
        RECT 391.950 262.950 394.050 263.400 ;
        RECT 406.950 262.950 409.050 263.400 ;
        RECT 454.950 264.600 457.050 265.050 ;
        RECT 475.950 264.600 478.050 265.050 ;
        RECT 454.950 263.400 478.050 264.600 ;
        RECT 454.950 262.950 457.050 263.400 ;
        RECT 475.950 262.950 478.050 263.400 ;
        RECT 526.950 264.600 529.050 265.050 ;
        RECT 535.950 264.600 538.050 265.050 ;
        RECT 526.950 263.400 538.050 264.600 ;
        RECT 526.950 262.950 529.050 263.400 ;
        RECT 535.950 262.950 538.050 263.400 ;
        RECT 571.950 264.600 574.050 265.050 ;
        RECT 580.950 264.600 583.050 265.050 ;
        RECT 571.950 263.400 583.050 264.600 ;
        RECT 571.950 262.950 574.050 263.400 ;
        RECT 580.950 262.950 583.050 263.400 ;
        RECT 595.950 264.600 598.050 265.050 ;
        RECT 604.950 264.600 607.050 265.050 ;
        RECT 595.950 263.400 607.050 264.600 ;
        RECT 595.950 262.950 598.050 263.400 ;
        RECT 604.950 262.950 607.050 263.400 ;
        RECT 736.950 264.600 739.050 265.050 ;
        RECT 763.950 264.600 766.050 265.050 ;
        RECT 736.950 263.400 766.050 264.600 ;
        RECT 736.950 262.950 739.050 263.400 ;
        RECT 763.950 262.950 766.050 263.400 ;
        RECT 943.950 264.600 946.050 265.050 ;
        RECT 949.950 264.600 952.050 265.050 ;
        RECT 943.950 263.400 952.050 264.600 ;
        RECT 943.950 262.950 946.050 263.400 ;
        RECT 949.950 262.950 952.050 263.400 ;
        RECT 64.950 261.600 67.050 262.050 ;
        RECT 53.400 260.400 67.050 261.600 ;
        RECT 53.400 255.900 54.600 260.400 ;
        RECT 64.950 259.950 67.050 260.400 ;
        RECT 79.950 260.100 82.050 262.200 ;
        RECT 103.950 261.750 106.050 262.200 ;
        RECT 112.950 261.750 115.050 262.200 ;
        RECT 103.950 260.550 115.050 261.750 ;
        RECT 103.950 260.100 106.050 260.550 ;
        RECT 112.950 260.100 115.050 260.550 ;
        RECT 121.950 260.100 124.050 262.200 ;
        RECT 133.950 261.600 136.050 262.050 ;
        RECT 128.400 260.400 136.050 261.600 ;
        RECT 80.400 256.050 81.600 260.100 ;
        RECT 52.950 253.800 55.050 255.900 ;
        RECT 80.400 254.400 85.050 256.050 ;
        RECT 81.000 253.950 85.050 254.400 ;
        RECT 106.950 255.450 109.050 255.900 ;
        RECT 115.950 255.450 118.050 255.900 ;
        RECT 106.950 254.250 118.050 255.450 ;
        RECT 106.950 253.800 109.050 254.250 ;
        RECT 115.950 253.800 118.050 254.250 ;
        RECT 122.400 253.050 123.600 260.100 ;
        RECT 124.950 255.600 127.050 255.900 ;
        RECT 128.400 255.600 129.600 260.400 ;
        RECT 133.950 259.950 136.050 260.400 ;
        RECT 190.950 261.600 193.050 262.200 ;
        RECT 199.950 261.600 202.050 262.050 ;
        RECT 190.950 260.400 202.050 261.600 ;
        RECT 190.950 260.100 193.050 260.400 ;
        RECT 199.950 259.950 202.050 260.400 ;
        RECT 235.950 261.750 238.050 262.200 ;
        RECT 241.950 261.750 244.050 262.200 ;
        RECT 235.950 260.550 244.050 261.750 ;
        RECT 235.950 260.100 238.050 260.550 ;
        RECT 241.950 260.100 244.050 260.550 ;
        RECT 271.950 261.600 274.050 262.200 ;
        RECT 283.950 261.750 286.050 262.200 ;
        RECT 292.950 261.750 295.050 262.200 ;
        RECT 271.950 260.400 282.600 261.600 ;
        RECT 271.950 260.100 274.050 260.400 ;
        RECT 281.400 258.600 282.600 260.400 ;
        RECT 283.950 260.550 295.050 261.750 ;
        RECT 283.950 260.100 286.050 260.550 ;
        RECT 292.950 260.100 295.050 260.550 ;
        RECT 298.950 261.600 301.050 262.200 ;
        RECT 334.950 261.750 337.050 262.200 ;
        RECT 349.950 261.750 352.050 262.200 ;
        RECT 334.950 261.600 352.050 261.750 ;
        RECT 373.950 261.600 376.050 262.050 ;
        RECT 298.950 260.400 318.600 261.600 ;
        RECT 298.950 260.100 301.050 260.400 ;
        RECT 281.400 257.400 297.600 258.600 ;
        RECT 124.950 254.400 129.600 255.600 ;
        RECT 130.950 255.450 133.050 255.900 ;
        RECT 139.950 255.450 142.050 255.900 ;
        RECT 124.950 253.800 127.050 254.400 ;
        RECT 130.950 254.250 142.050 255.450 ;
        RECT 130.950 253.800 133.050 254.250 ;
        RECT 139.950 253.800 142.050 254.250 ;
        RECT 145.950 255.450 148.050 255.900 ;
        RECT 160.950 255.450 163.050 255.900 ;
        RECT 145.950 254.250 163.050 255.450 ;
        RECT 145.950 253.800 148.050 254.250 ;
        RECT 160.950 253.800 163.050 254.250 ;
        RECT 193.950 255.600 196.050 255.900 ;
        RECT 211.950 255.600 214.050 255.900 ;
        RECT 193.950 254.400 214.050 255.600 ;
        RECT 193.950 253.800 196.050 254.400 ;
        RECT 211.950 253.800 214.050 254.400 ;
        RECT 223.950 255.600 226.050 256.050 ;
        RECT 296.400 255.900 297.600 257.400 ;
        RECT 317.400 255.900 318.600 260.400 ;
        RECT 334.950 260.550 376.050 261.600 ;
        RECT 334.950 260.100 337.050 260.550 ;
        RECT 349.950 260.400 376.050 260.550 ;
        RECT 349.950 260.100 352.050 260.400 ;
        RECT 373.950 259.950 376.050 260.400 ;
        RECT 403.950 261.600 406.050 262.200 ;
        RECT 418.950 261.600 421.050 262.050 ;
        RECT 433.950 261.600 436.050 262.200 ;
        RECT 403.950 260.400 421.050 261.600 ;
        RECT 403.950 260.100 406.050 260.400 ;
        RECT 418.950 259.950 421.050 260.400 ;
        RECT 422.400 260.400 436.050 261.600 ;
        RECT 415.950 258.600 418.050 259.050 ;
        RECT 422.400 258.600 423.600 260.400 ;
        RECT 433.950 260.100 436.050 260.400 ;
        RECT 451.950 261.600 454.050 262.200 ;
        RECT 472.950 261.600 475.050 262.050 ;
        RECT 451.950 260.400 475.050 261.600 ;
        RECT 451.950 260.100 454.050 260.400 ;
        RECT 472.950 259.950 475.050 260.400 ;
        RECT 487.950 261.750 490.050 262.200 ;
        RECT 499.950 261.750 502.050 262.200 ;
        RECT 487.950 260.550 502.050 261.750 ;
        RECT 487.950 260.100 490.050 260.550 ;
        RECT 499.950 260.100 502.050 260.550 ;
        RECT 517.950 261.600 520.050 262.200 ;
        RECT 523.950 261.600 526.050 262.050 ;
        RECT 517.950 260.400 526.050 261.600 ;
        RECT 517.950 260.100 520.050 260.400 ;
        RECT 523.950 259.950 526.050 260.400 ;
        RECT 544.950 261.600 547.050 262.050 ;
        RECT 562.950 261.600 565.050 262.200 ;
        RECT 544.950 260.400 565.050 261.600 ;
        RECT 544.950 259.950 547.050 260.400 ;
        RECT 562.950 260.100 565.050 260.400 ;
        RECT 592.950 261.600 595.050 262.050 ;
        RECT 601.950 261.600 604.050 262.200 ;
        RECT 592.950 260.400 604.050 261.600 ;
        RECT 592.950 259.950 595.050 260.400 ;
        RECT 601.950 260.100 604.050 260.400 ;
        RECT 607.950 261.600 610.050 262.050 ;
        RECT 613.950 261.600 616.050 262.050 ;
        RECT 607.950 260.400 616.050 261.600 ;
        RECT 607.950 259.950 610.050 260.400 ;
        RECT 613.950 259.950 616.050 260.400 ;
        RECT 661.950 261.600 664.050 262.050 ;
        RECT 667.950 261.600 670.050 262.050 ;
        RECT 661.950 260.400 670.050 261.600 ;
        RECT 661.950 259.950 664.050 260.400 ;
        RECT 667.950 259.950 670.050 260.400 ;
        RECT 697.950 260.100 700.050 262.200 ;
        RECT 415.950 257.400 423.600 258.600 ;
        RECT 568.950 258.600 571.050 259.050 ;
        RECT 619.950 258.600 622.050 259.050 ;
        RECT 698.400 258.600 699.600 260.100 ;
        RECT 709.950 259.950 712.050 262.050 ;
        RECT 715.950 261.750 718.050 262.200 ;
        RECT 724.950 261.750 727.050 262.200 ;
        RECT 715.950 260.550 727.050 261.750 ;
        RECT 715.950 260.100 718.050 260.550 ;
        RECT 724.950 260.100 727.050 260.550 ;
        RECT 778.950 261.600 781.050 262.200 ;
        RECT 808.950 261.600 811.050 262.050 ;
        RECT 778.950 260.400 811.050 261.600 ;
        RECT 778.950 260.100 781.050 260.400 ;
        RECT 808.950 259.950 811.050 260.400 ;
        RECT 832.950 261.600 835.050 262.050 ;
        RECT 838.950 261.600 841.050 262.200 ;
        RECT 832.950 260.400 841.050 261.600 ;
        RECT 832.950 259.950 835.050 260.400 ;
        RECT 838.950 260.100 841.050 260.400 ;
        RECT 844.950 261.600 847.050 262.200 ;
        RECT 865.950 261.600 868.050 262.200 ;
        RECT 844.950 260.400 868.050 261.600 ;
        RECT 844.950 260.100 847.050 260.400 ;
        RECT 865.950 260.100 868.050 260.400 ;
        RECT 871.950 261.600 874.050 262.200 ;
        RECT 889.950 261.600 892.050 262.200 ;
        RECT 913.950 261.600 916.050 262.200 ;
        RECT 871.950 260.400 916.050 261.600 ;
        RECT 871.950 260.100 874.050 260.400 ;
        RECT 568.950 257.400 585.600 258.600 ;
        RECT 415.950 256.950 418.050 257.400 ;
        RECT 568.950 256.950 571.050 257.400 ;
        RECT 232.950 255.600 235.050 255.900 ;
        RECT 223.950 254.400 235.050 255.600 ;
        RECT 223.950 253.950 226.050 254.400 ;
        RECT 232.950 253.800 235.050 254.400 ;
        RECT 262.950 255.450 265.050 255.900 ;
        RECT 274.950 255.450 277.050 255.900 ;
        RECT 262.950 254.250 277.050 255.450 ;
        RECT 262.950 253.800 265.050 254.250 ;
        RECT 274.950 253.800 277.050 254.250 ;
        RECT 295.950 253.800 298.050 255.900 ;
        RECT 316.950 253.800 319.050 255.900 ;
        RECT 346.950 255.450 349.050 255.900 ;
        RECT 361.950 255.450 364.050 255.900 ;
        RECT 346.950 254.250 364.050 255.450 ;
        RECT 346.950 253.800 349.050 254.250 ;
        RECT 361.950 253.800 364.050 254.250 ;
        RECT 373.950 255.450 376.050 255.900 ;
        RECT 379.950 255.450 382.050 255.900 ;
        RECT 373.950 254.250 382.050 255.450 ;
        RECT 373.950 253.800 376.050 254.250 ;
        RECT 379.950 253.800 382.050 254.250 ;
        RECT 385.950 255.450 388.050 255.900 ;
        RECT 391.950 255.450 394.050 255.900 ;
        RECT 385.950 254.250 394.050 255.450 ;
        RECT 385.950 253.800 388.050 254.250 ;
        RECT 391.950 253.800 394.050 254.250 ;
        RECT 418.950 255.450 421.050 255.900 ;
        RECT 424.950 255.450 427.050 255.900 ;
        RECT 418.950 254.250 427.050 255.450 ;
        RECT 418.950 253.800 421.050 254.250 ;
        RECT 424.950 253.800 427.050 254.250 ;
        RECT 460.950 255.450 463.050 255.900 ;
        RECT 490.950 255.450 493.050 256.050 ;
        RECT 496.950 255.450 499.050 255.900 ;
        RECT 460.950 254.250 499.050 255.450 ;
        RECT 460.950 253.800 463.050 254.250 ;
        RECT 490.950 253.950 493.050 254.250 ;
        RECT 496.950 253.800 499.050 254.250 ;
        RECT 514.950 255.600 517.050 255.900 ;
        RECT 526.950 255.600 529.050 256.050 ;
        RECT 514.950 254.400 529.050 255.600 ;
        RECT 514.950 253.800 517.050 254.400 ;
        RECT 526.950 253.950 529.050 254.400 ;
        RECT 538.950 255.600 541.050 255.900 ;
        RECT 559.950 255.600 562.050 255.900 ;
        RECT 538.950 254.400 562.050 255.600 ;
        RECT 538.950 253.800 541.050 254.400 ;
        RECT 559.950 253.800 562.050 254.400 ;
        RECT 571.950 255.450 574.050 256.050 ;
        RECT 580.950 255.450 583.050 255.900 ;
        RECT 571.950 254.250 583.050 255.450 ;
        RECT 584.400 255.600 585.600 257.400 ;
        RECT 619.950 258.000 702.600 258.600 ;
        RECT 619.950 257.400 703.050 258.000 ;
        RECT 619.950 256.950 622.050 257.400 ;
        RECT 586.950 255.600 589.050 255.900 ;
        RECT 604.950 255.600 607.050 255.900 ;
        RECT 584.400 254.400 607.050 255.600 ;
        RECT 571.950 253.950 574.050 254.250 ;
        RECT 580.950 253.800 583.050 254.250 ;
        RECT 586.950 253.800 589.050 254.400 ;
        RECT 604.950 253.800 607.050 254.400 ;
        RECT 616.950 255.600 619.050 256.050 ;
        RECT 661.950 255.600 664.050 256.050 ;
        RECT 616.950 254.400 664.050 255.600 ;
        RECT 616.950 253.950 619.050 254.400 ;
        RECT 661.950 253.950 664.050 254.400 ;
        RECT 676.950 255.450 679.050 255.900 ;
        RECT 685.950 255.450 688.050 255.900 ;
        RECT 676.950 254.250 688.050 255.450 ;
        RECT 676.950 253.800 679.050 254.250 ;
        RECT 685.950 253.800 688.050 254.250 ;
        RECT 700.950 253.950 703.050 257.400 ;
        RECT 710.400 255.600 711.600 259.950 ;
        RECT 829.950 258.600 832.050 259.050 ;
        RECT 818.400 257.400 832.050 258.600 ;
        RECT 712.950 255.600 715.050 255.900 ;
        RECT 710.400 254.400 715.050 255.600 ;
        RECT 712.950 253.800 715.050 254.400 ;
        RECT 739.950 255.450 742.050 255.900 ;
        RECT 745.950 255.450 748.050 255.900 ;
        RECT 739.950 254.250 748.050 255.450 ;
        RECT 739.950 253.800 742.050 254.250 ;
        RECT 745.950 253.800 748.050 254.250 ;
        RECT 754.950 255.600 757.050 255.900 ;
        RECT 775.950 255.600 778.050 255.900 ;
        RECT 754.950 254.400 778.050 255.600 ;
        RECT 754.950 253.800 757.050 254.400 ;
        RECT 775.950 253.800 778.050 254.400 ;
        RECT 781.950 255.450 784.050 255.900 ;
        RECT 787.950 255.450 790.050 255.900 ;
        RECT 781.950 254.250 790.050 255.450 ;
        RECT 781.950 253.800 784.050 254.250 ;
        RECT 787.950 253.800 790.050 254.250 ;
        RECT 802.950 255.600 805.050 255.900 ;
        RECT 818.400 255.600 819.600 257.400 ;
        RECT 829.950 256.950 832.050 257.400 ;
        RECT 875.400 256.050 876.600 260.400 ;
        RECT 889.950 260.100 892.050 260.400 ;
        RECT 913.950 260.100 916.050 260.400 ;
        RECT 925.950 261.600 928.050 262.050 ;
        RECT 937.950 261.600 940.050 262.200 ;
        RECT 925.950 260.400 940.050 261.600 ;
        RECT 958.950 261.600 961.050 265.050 ;
        RECT 979.950 264.600 982.050 265.050 ;
        RECT 985.950 264.600 988.050 265.050 ;
        RECT 979.950 263.400 988.050 264.600 ;
        RECT 991.950 264.600 994.050 268.050 ;
        RECT 1015.950 264.600 1018.050 265.050 ;
        RECT 991.950 264.000 1018.050 264.600 ;
        RECT 992.400 263.400 1018.050 264.000 ;
        RECT 979.950 262.950 982.050 263.400 ;
        RECT 985.950 262.950 988.050 263.400 ;
        RECT 1015.950 262.950 1018.050 263.400 ;
        RECT 970.950 261.600 973.050 262.200 ;
        RECT 958.950 261.000 973.050 261.600 ;
        RECT 959.400 260.400 973.050 261.000 ;
        RECT 925.950 259.950 928.050 260.400 ;
        RECT 937.950 260.100 940.050 260.400 ;
        RECT 970.950 260.100 973.050 260.400 ;
        RECT 982.950 259.950 985.050 262.050 ;
        RECT 1006.950 261.600 1009.050 262.050 ;
        RECT 992.400 260.400 1009.050 261.600 ;
        RECT 983.400 256.050 984.600 259.950 ;
        RECT 802.950 254.400 819.600 255.600 ;
        RECT 802.950 253.800 805.050 254.400 ;
        RECT 874.950 253.950 877.050 256.050 ;
        RECT 940.950 255.600 943.050 255.900 ;
        RECT 955.950 255.600 958.050 255.900 ;
        RECT 940.950 255.450 958.050 255.600 ;
        RECT 967.950 255.450 970.050 255.900 ;
        RECT 940.950 254.400 970.050 255.450 ;
        RECT 940.950 253.800 943.050 254.400 ;
        RECT 955.950 254.250 970.050 254.400 ;
        RECT 955.950 253.800 958.050 254.250 ;
        RECT 967.950 253.800 970.050 254.250 ;
        RECT 982.950 253.950 985.050 256.050 ;
        RECT 992.400 255.900 993.600 260.400 ;
        RECT 1006.950 259.950 1009.050 260.400 ;
        RECT 991.950 253.800 994.050 255.900 ;
        RECT 31.950 252.600 34.050 253.050 ;
        RECT 37.950 252.600 40.050 253.050 ;
        RECT 31.950 251.400 40.050 252.600 ;
        RECT 31.950 250.950 34.050 251.400 ;
        RECT 37.950 250.950 40.050 251.400 ;
        RECT 61.950 252.600 64.050 253.050 ;
        RECT 67.950 252.600 70.050 253.050 ;
        RECT 61.950 251.400 70.050 252.600 ;
        RECT 61.950 250.950 64.050 251.400 ;
        RECT 67.950 250.950 70.050 251.400 ;
        RECT 85.950 252.600 88.050 253.050 ;
        RECT 97.950 252.600 100.050 253.050 ;
        RECT 85.950 251.400 100.050 252.600 ;
        RECT 85.950 250.950 88.050 251.400 ;
        RECT 97.950 250.950 100.050 251.400 ;
        RECT 121.950 250.950 124.050 253.050 ;
        RECT 151.950 252.600 154.050 253.050 ;
        RECT 166.950 252.600 169.050 253.050 ;
        RECT 151.950 251.400 169.050 252.600 ;
        RECT 151.950 250.950 154.050 251.400 ;
        RECT 166.950 250.950 169.050 251.400 ;
        RECT 217.950 252.600 220.050 253.050 ;
        RECT 241.950 252.600 244.050 253.050 ;
        RECT 217.950 251.400 244.050 252.600 ;
        RECT 217.950 250.950 220.050 251.400 ;
        RECT 241.950 250.950 244.050 251.400 ;
        RECT 307.950 252.600 310.050 253.050 ;
        RECT 325.950 252.600 328.050 253.050 ;
        RECT 307.950 251.400 328.050 252.600 ;
        RECT 307.950 250.950 310.050 251.400 ;
        RECT 325.950 250.950 328.050 251.400 ;
        RECT 349.950 252.600 352.050 253.050 ;
        RECT 355.950 252.600 358.050 253.050 ;
        RECT 349.950 251.400 358.050 252.600 ;
        RECT 349.950 250.950 352.050 251.400 ;
        RECT 355.950 250.950 358.050 251.400 ;
        RECT 433.950 252.600 436.050 253.050 ;
        RECT 442.950 252.600 445.050 253.050 ;
        RECT 469.800 252.600 471.900 253.050 ;
        RECT 433.950 251.400 445.050 252.600 ;
        RECT 433.950 250.950 436.050 251.400 ;
        RECT 442.950 250.950 445.050 251.400 ;
        RECT 464.400 251.400 471.900 252.600 ;
        RECT 301.950 249.600 304.050 250.050 ;
        RECT 322.950 249.600 325.050 250.050 ;
        RECT 301.950 248.400 325.050 249.600 ;
        RECT 301.950 247.950 304.050 248.400 ;
        RECT 322.950 247.950 325.050 248.400 ;
        RECT 376.950 249.600 379.050 250.050 ;
        RECT 394.950 249.600 397.050 250.050 ;
        RECT 418.800 249.600 420.900 250.050 ;
        RECT 376.950 248.400 397.050 249.600 ;
        RECT 376.950 247.950 379.050 248.400 ;
        RECT 394.950 247.950 397.050 248.400 ;
        RECT 398.400 248.400 420.900 249.600 ;
        RECT 175.950 246.600 178.050 247.050 ;
        RECT 262.950 246.600 265.050 247.050 ;
        RECT 175.950 245.400 265.050 246.600 ;
        RECT 175.950 244.950 178.050 245.400 ;
        RECT 262.950 244.950 265.050 245.400 ;
        RECT 343.950 246.600 346.050 247.050 ;
        RECT 398.400 246.600 399.600 248.400 ;
        RECT 418.800 247.950 420.900 248.400 ;
        RECT 421.950 249.600 424.050 250.050 ;
        RECT 427.950 249.600 430.050 250.050 ;
        RECT 421.950 248.400 430.050 249.600 ;
        RECT 421.950 247.950 424.050 248.400 ;
        RECT 427.950 247.950 430.050 248.400 ;
        RECT 439.950 249.600 442.050 250.050 ;
        RECT 464.400 249.600 465.600 251.400 ;
        RECT 469.800 250.950 471.900 251.400 ;
        RECT 472.950 252.600 475.050 253.050 ;
        RECT 478.950 252.600 481.050 253.050 ;
        RECT 472.950 251.400 481.050 252.600 ;
        RECT 472.950 250.950 475.050 251.400 ;
        RECT 478.950 250.950 481.050 251.400 ;
        RECT 541.950 252.600 544.050 253.050 ;
        RECT 571.950 252.600 574.050 252.900 ;
        RECT 541.950 251.400 574.050 252.600 ;
        RECT 541.950 250.950 544.050 251.400 ;
        RECT 571.950 250.800 574.050 251.400 ;
        RECT 664.950 252.600 667.050 253.050 ;
        RECT 676.950 252.600 679.050 252.750 ;
        RECT 664.950 251.400 679.050 252.600 ;
        RECT 664.950 250.950 667.050 251.400 ;
        RECT 676.950 250.650 679.050 251.400 ;
        RECT 706.950 252.600 709.050 253.050 ;
        RECT 730.950 252.600 733.050 253.050 ;
        RECT 706.950 251.400 733.050 252.600 ;
        RECT 706.950 250.950 709.050 251.400 ;
        RECT 730.950 250.950 733.050 251.400 ;
        RECT 820.950 252.600 823.050 253.050 ;
        RECT 841.950 252.600 844.050 253.050 ;
        RECT 862.950 252.600 865.050 253.050 ;
        RECT 820.950 251.400 865.050 252.600 ;
        RECT 820.950 250.950 823.050 251.400 ;
        RECT 841.950 250.950 844.050 251.400 ;
        RECT 862.950 250.950 865.050 251.400 ;
        RECT 886.950 252.600 889.050 253.050 ;
        RECT 916.950 252.600 919.050 253.050 ;
        RECT 886.950 251.400 919.050 252.600 ;
        RECT 886.950 250.950 889.050 251.400 ;
        RECT 916.950 250.950 919.050 251.400 ;
        RECT 439.950 248.400 465.600 249.600 ;
        RECT 502.950 249.600 505.050 250.050 ;
        RECT 508.950 249.600 511.050 249.900 ;
        RECT 502.950 248.400 511.050 249.600 ;
        RECT 439.950 247.950 442.050 248.400 ;
        RECT 502.950 247.950 505.050 248.400 ;
        RECT 508.950 247.800 511.050 248.400 ;
        RECT 526.950 249.600 529.050 250.050 ;
        RECT 568.950 249.600 571.050 250.050 ;
        RECT 526.950 248.400 571.050 249.600 ;
        RECT 526.950 247.950 529.050 248.400 ;
        RECT 568.950 247.950 571.050 248.400 ;
        RECT 607.950 249.600 610.050 250.050 ;
        RECT 640.950 249.600 643.050 250.050 ;
        RECT 652.950 249.600 655.050 250.050 ;
        RECT 607.950 248.400 655.050 249.600 ;
        RECT 607.950 247.950 610.050 248.400 ;
        RECT 640.950 247.950 643.050 248.400 ;
        RECT 652.950 247.950 655.050 248.400 ;
        RECT 667.950 249.600 670.050 250.050 ;
        RECT 697.950 249.600 700.050 250.050 ;
        RECT 667.950 248.400 700.050 249.600 ;
        RECT 667.950 247.950 670.050 248.400 ;
        RECT 697.950 247.950 700.050 248.400 ;
        RECT 709.950 249.600 712.050 250.050 ;
        RECT 760.950 249.600 763.050 250.050 ;
        RECT 709.950 248.400 763.050 249.600 ;
        RECT 709.950 247.950 712.050 248.400 ;
        RECT 760.950 247.950 763.050 248.400 ;
        RECT 829.950 249.600 832.050 250.050 ;
        RECT 847.950 249.600 850.050 250.050 ;
        RECT 829.950 248.400 850.050 249.600 ;
        RECT 829.950 247.950 832.050 248.400 ;
        RECT 847.950 247.950 850.050 248.400 ;
        RECT 343.950 245.400 399.600 246.600 ;
        RECT 406.950 246.600 409.050 247.050 ;
        RECT 430.950 246.600 433.050 247.050 ;
        RECT 448.950 246.600 451.050 247.050 ;
        RECT 475.800 246.600 477.900 247.050 ;
        RECT 406.950 245.400 477.900 246.600 ;
        RECT 343.950 244.950 346.050 245.400 ;
        RECT 406.950 244.950 409.050 245.400 ;
        RECT 430.950 244.950 433.050 245.400 ;
        RECT 448.950 244.950 451.050 245.400 ;
        RECT 475.800 244.950 477.900 245.400 ;
        RECT 478.950 246.600 481.050 247.050 ;
        RECT 511.950 246.600 514.050 247.050 ;
        RECT 478.950 245.400 514.050 246.600 ;
        RECT 478.950 244.950 481.050 245.400 ;
        RECT 511.950 244.950 514.050 245.400 ;
        RECT 661.950 246.600 664.050 247.050 ;
        RECT 769.950 246.600 772.050 247.050 ;
        RECT 661.950 245.400 772.050 246.600 ;
        RECT 661.950 244.950 664.050 245.400 ;
        RECT 769.950 244.950 772.050 245.400 ;
        RECT 22.950 243.600 25.050 244.050 ;
        RECT 112.950 243.600 115.050 244.050 ;
        RECT 22.950 242.400 115.050 243.600 ;
        RECT 22.950 241.950 25.050 242.400 ;
        RECT 112.950 241.950 115.050 242.400 ;
        RECT 280.950 243.600 283.050 244.050 ;
        RECT 445.950 243.600 448.050 244.050 ;
        RECT 472.950 243.600 475.050 244.050 ;
        RECT 280.950 242.400 441.600 243.600 ;
        RECT 280.950 241.950 283.050 242.400 ;
        RECT 139.950 240.600 142.050 241.050 ;
        RECT 328.950 240.600 331.050 241.050 ;
        RECT 340.950 240.600 343.050 241.050 ;
        RECT 139.950 239.400 207.600 240.600 ;
        RECT 139.950 238.950 142.050 239.400 ;
        RECT 100.950 237.600 103.050 238.050 ;
        RECT 157.950 237.600 160.050 238.050 ;
        RECT 100.950 236.400 160.050 237.600 ;
        RECT 206.400 237.600 207.600 239.400 ;
        RECT 328.950 239.400 343.050 240.600 ;
        RECT 328.950 238.950 331.050 239.400 ;
        RECT 340.950 238.950 343.050 239.400 ;
        RECT 415.950 240.600 418.050 241.050 ;
        RECT 424.950 240.600 427.050 241.050 ;
        RECT 415.950 239.400 427.050 240.600 ;
        RECT 440.400 240.600 441.600 242.400 ;
        RECT 445.950 242.400 475.050 243.600 ;
        RECT 445.950 241.950 448.050 242.400 ;
        RECT 472.950 241.950 475.050 242.400 ;
        RECT 532.950 243.600 535.050 244.050 ;
        RECT 580.800 243.600 582.900 244.050 ;
        RECT 532.950 242.400 582.900 243.600 ;
        RECT 532.950 241.950 535.050 242.400 ;
        RECT 580.800 241.950 582.900 242.400 ;
        RECT 583.950 243.600 586.050 244.050 ;
        RECT 604.950 243.600 607.050 244.050 ;
        RECT 583.950 242.400 607.050 243.600 ;
        RECT 583.950 241.950 586.050 242.400 ;
        RECT 604.950 241.950 607.050 242.400 ;
        RECT 610.950 243.600 613.050 244.050 ;
        RECT 670.950 243.600 673.050 244.050 ;
        RECT 742.950 243.600 745.050 244.050 ;
        RECT 610.950 242.400 673.050 243.600 ;
        RECT 610.950 241.950 613.050 242.400 ;
        RECT 670.950 241.950 673.050 242.400 ;
        RECT 677.400 242.400 745.050 243.600 ;
        RECT 448.950 240.600 451.050 241.050 ;
        RECT 440.400 239.400 451.050 240.600 ;
        RECT 473.400 240.600 474.600 241.950 ;
        RECT 677.400 241.050 678.600 242.400 ;
        RECT 742.950 241.950 745.050 242.400 ;
        RECT 760.950 243.600 763.050 244.050 ;
        RECT 793.950 243.600 796.050 244.050 ;
        RECT 760.950 242.400 796.050 243.600 ;
        RECT 760.950 241.950 763.050 242.400 ;
        RECT 793.950 241.950 796.050 242.400 ;
        RECT 808.950 243.600 811.050 244.050 ;
        RECT 883.950 243.600 886.050 244.050 ;
        RECT 892.950 243.600 895.050 244.050 ;
        RECT 910.950 243.600 913.050 244.050 ;
        RECT 808.950 242.400 913.050 243.600 ;
        RECT 808.950 241.950 811.050 242.400 ;
        RECT 883.950 241.950 886.050 242.400 ;
        RECT 892.950 241.950 895.050 242.400 ;
        RECT 910.950 241.950 913.050 242.400 ;
        RECT 988.950 243.600 991.050 244.050 ;
        RECT 1000.950 243.600 1003.050 244.050 ;
        RECT 988.950 242.400 1003.050 243.600 ;
        RECT 988.950 241.950 991.050 242.400 ;
        RECT 1000.950 241.950 1003.050 242.400 ;
        RECT 505.950 240.600 508.050 241.050 ;
        RECT 473.400 239.400 508.050 240.600 ;
        RECT 415.950 238.950 418.050 239.400 ;
        RECT 424.950 238.950 427.050 239.400 ;
        RECT 448.950 238.950 451.050 239.400 ;
        RECT 505.950 238.950 508.050 239.400 ;
        RECT 511.950 240.600 514.050 241.050 ;
        RECT 565.950 240.600 568.050 241.050 ;
        RECT 511.950 239.400 568.050 240.600 ;
        RECT 511.950 238.950 514.050 239.400 ;
        RECT 565.950 238.950 568.050 239.400 ;
        RECT 571.950 240.600 574.050 241.050 ;
        RECT 607.950 240.600 610.050 241.050 ;
        RECT 571.950 239.400 610.050 240.600 ;
        RECT 571.950 238.950 574.050 239.400 ;
        RECT 607.950 238.950 610.050 239.400 ;
        RECT 652.950 240.600 655.050 241.050 ;
        RECT 658.950 240.600 661.050 241.050 ;
        RECT 652.950 239.400 661.050 240.600 ;
        RECT 652.950 238.950 655.050 239.400 ;
        RECT 658.950 238.950 661.050 239.400 ;
        RECT 673.950 239.400 678.600 241.050 ;
        RECT 697.950 240.600 700.050 241.050 ;
        RECT 802.950 240.600 805.050 241.050 ;
        RECT 697.950 239.400 805.050 240.600 ;
        RECT 673.950 238.950 678.000 239.400 ;
        RECT 697.950 238.950 700.050 239.400 ;
        RECT 802.950 238.950 805.050 239.400 ;
        RECT 901.950 240.600 904.050 241.050 ;
        RECT 940.950 240.600 943.050 241.050 ;
        RECT 901.950 239.400 943.050 240.600 ;
        RECT 901.950 238.950 904.050 239.400 ;
        RECT 940.950 238.950 943.050 239.400 ;
        RECT 955.950 240.600 958.050 241.050 ;
        RECT 979.950 240.600 982.050 241.050 ;
        RECT 955.950 239.400 982.050 240.600 ;
        RECT 955.950 238.950 958.050 239.400 ;
        RECT 979.950 238.950 982.050 239.400 ;
        RECT 985.950 240.600 988.050 241.050 ;
        RECT 991.950 240.600 994.050 241.050 ;
        RECT 985.950 239.400 994.050 240.600 ;
        RECT 985.950 238.950 988.050 239.400 ;
        RECT 991.950 238.950 994.050 239.400 ;
        RECT 280.950 237.600 283.050 238.050 ;
        RECT 206.400 236.400 283.050 237.600 ;
        RECT 100.950 235.950 103.050 236.400 ;
        RECT 157.950 235.950 160.050 236.400 ;
        RECT 280.950 235.950 283.050 236.400 ;
        RECT 349.950 237.600 352.050 238.050 ;
        RECT 496.950 237.600 499.050 238.050 ;
        RECT 349.950 236.400 499.050 237.600 ;
        RECT 506.400 237.600 507.600 238.950 ;
        RECT 541.950 237.600 544.050 238.050 ;
        RECT 506.400 236.400 544.050 237.600 ;
        RECT 349.950 235.950 352.050 236.400 ;
        RECT 496.950 235.950 499.050 236.400 ;
        RECT 541.950 235.950 544.050 236.400 ;
        RECT 553.950 237.600 556.050 238.050 ;
        RECT 568.950 237.600 571.050 237.900 ;
        RECT 553.950 236.400 571.050 237.600 ;
        RECT 553.950 235.950 556.050 236.400 ;
        RECT 568.950 235.800 571.050 236.400 ;
        RECT 574.950 237.600 577.050 238.050 ;
        RECT 703.950 237.600 706.050 238.050 ;
        RECT 712.950 237.600 715.050 238.050 ;
        RECT 574.950 236.400 639.600 237.600 ;
        RECT 574.950 235.950 577.050 236.400 ;
        RECT 76.950 234.600 79.050 235.050 ;
        RECT 91.950 234.600 94.050 235.050 ;
        RECT 112.950 234.600 115.050 235.050 ;
        RECT 76.950 233.400 115.050 234.600 ;
        RECT 76.950 232.950 79.050 233.400 ;
        RECT 91.950 232.950 94.050 233.400 ;
        RECT 112.950 232.950 115.050 233.400 ;
        RECT 259.950 234.600 262.050 235.050 ;
        RECT 268.950 234.600 271.050 235.050 ;
        RECT 259.950 233.400 271.050 234.600 ;
        RECT 259.950 232.950 262.050 233.400 ;
        RECT 268.950 232.950 271.050 233.400 ;
        RECT 301.950 234.600 304.050 235.050 ;
        RECT 460.950 234.600 463.050 235.050 ;
        RECT 301.950 233.400 463.050 234.600 ;
        RECT 638.400 234.600 639.600 236.400 ;
        RECT 703.950 236.400 715.050 237.600 ;
        RECT 703.950 235.950 706.050 236.400 ;
        RECT 712.950 235.950 715.050 236.400 ;
        RECT 976.950 237.600 979.050 238.050 ;
        RECT 1015.950 237.600 1018.050 238.050 ;
        RECT 976.950 236.400 1018.050 237.600 ;
        RECT 976.950 235.950 979.050 236.400 ;
        RECT 1015.950 235.950 1018.050 236.400 ;
        RECT 685.950 234.600 688.050 235.050 ;
        RECT 727.950 234.600 730.050 235.050 ;
        RECT 638.400 233.400 688.050 234.600 ;
        RECT 301.950 232.950 304.050 233.400 ;
        RECT 460.950 232.950 463.050 233.400 ;
        RECT 685.950 232.950 688.050 233.400 ;
        RECT 695.400 233.400 730.050 234.600 ;
        RECT 695.400 232.050 696.600 233.400 ;
        RECT 727.950 232.950 730.050 233.400 ;
        RECT 745.950 234.600 748.050 235.050 ;
        RECT 814.950 234.600 817.050 235.050 ;
        RECT 745.950 233.400 817.050 234.600 ;
        RECT 745.950 232.950 748.050 233.400 ;
        RECT 814.950 232.950 817.050 233.400 ;
        RECT 856.950 234.600 859.050 235.050 ;
        RECT 877.950 234.600 880.050 235.050 ;
        RECT 856.950 233.400 880.050 234.600 ;
        RECT 856.950 232.950 859.050 233.400 ;
        RECT 877.950 232.950 880.050 233.400 ;
        RECT 910.950 234.600 913.050 235.050 ;
        RECT 952.950 234.600 955.050 235.050 ;
        RECT 910.950 233.400 955.050 234.600 ;
        RECT 910.950 232.950 913.050 233.400 ;
        RECT 952.950 232.950 955.050 233.400 ;
        RECT 964.950 234.600 967.050 235.050 ;
        RECT 1003.950 234.600 1006.050 235.050 ;
        RECT 964.950 233.400 1006.050 234.600 ;
        RECT 964.950 232.950 967.050 233.400 ;
        RECT 1003.950 232.950 1006.050 233.400 ;
        RECT 514.950 231.600 517.050 232.050 ;
        RECT 532.950 231.600 535.050 232.050 ;
        RECT 514.950 230.400 535.050 231.600 ;
        RECT 514.950 229.950 517.050 230.400 ;
        RECT 532.950 229.950 535.050 230.400 ;
        RECT 556.950 231.600 559.050 232.050 ;
        RECT 589.950 231.600 592.050 232.050 ;
        RECT 595.950 231.600 598.050 232.050 ;
        RECT 619.950 231.600 622.050 232.050 ;
        RECT 556.950 230.400 598.050 231.600 ;
        RECT 556.950 229.950 559.050 230.400 ;
        RECT 589.950 229.950 592.050 230.400 ;
        RECT 595.950 229.950 598.050 230.400 ;
        RECT 599.400 230.400 622.050 231.600 ;
        RECT 160.950 228.600 163.050 229.050 ;
        RECT 229.950 228.600 232.050 229.050 ;
        RECT 343.800 228.600 345.900 229.050 ;
        RECT 160.950 227.400 345.900 228.600 ;
        RECT 160.950 226.950 163.050 227.400 ;
        RECT 229.950 226.950 232.050 227.400 ;
        RECT 343.800 226.950 345.900 227.400 ;
        RECT 346.950 228.600 349.050 229.050 ;
        RECT 406.950 228.600 409.050 229.050 ;
        RECT 346.950 227.400 409.050 228.600 ;
        RECT 346.950 226.950 349.050 227.400 ;
        RECT 406.950 226.950 409.050 227.400 ;
        RECT 418.950 228.600 421.050 229.050 ;
        RECT 478.950 228.600 481.050 229.050 ;
        RECT 418.950 227.400 481.050 228.600 ;
        RECT 418.950 226.950 421.050 227.400 ;
        RECT 478.950 226.950 481.050 227.400 ;
        RECT 541.950 228.600 544.050 229.050 ;
        RECT 599.400 228.600 600.600 230.400 ;
        RECT 619.950 229.950 622.050 230.400 ;
        RECT 628.950 231.600 631.050 232.050 ;
        RECT 694.950 231.600 697.050 232.050 ;
        RECT 628.950 230.400 697.050 231.600 ;
        RECT 628.950 229.950 631.050 230.400 ;
        RECT 694.950 229.950 697.050 230.400 ;
        RECT 841.950 231.600 844.050 232.050 ;
        RECT 904.950 231.600 907.050 232.050 ;
        RECT 841.950 230.400 907.050 231.600 ;
        RECT 841.950 229.950 844.050 230.400 ;
        RECT 904.950 229.950 907.050 230.400 ;
        RECT 541.950 227.400 600.600 228.600 ;
        RECT 649.950 228.600 652.050 229.050 ;
        RECT 667.950 228.600 670.050 229.050 ;
        RECT 679.950 228.600 682.050 229.050 ;
        RECT 649.950 227.400 682.050 228.600 ;
        RECT 541.950 226.950 544.050 227.400 ;
        RECT 649.950 226.950 652.050 227.400 ;
        RECT 667.950 226.950 670.050 227.400 ;
        RECT 679.950 226.950 682.050 227.400 ;
        RECT 817.950 228.600 820.050 229.050 ;
        RECT 832.950 228.600 835.050 229.050 ;
        RECT 817.950 227.400 835.050 228.600 ;
        RECT 817.950 226.950 820.050 227.400 ;
        RECT 832.950 226.950 835.050 227.400 ;
        RECT 934.950 228.600 937.050 229.050 ;
        RECT 973.950 228.600 976.050 229.050 ;
        RECT 1000.950 228.600 1003.050 229.050 ;
        RECT 934.950 227.400 1003.050 228.600 ;
        RECT 934.950 226.950 937.050 227.400 ;
        RECT 973.950 226.950 976.050 227.400 ;
        RECT 1000.950 226.950 1003.050 227.400 ;
        RECT 4.950 225.600 7.050 226.050 ;
        RECT 25.950 225.600 28.050 226.050 ;
        RECT 55.950 225.600 58.050 226.050 ;
        RECT 4.950 224.400 58.050 225.600 ;
        RECT 4.950 223.950 7.050 224.400 ;
        RECT 25.950 223.950 28.050 224.400 ;
        RECT 55.950 223.950 58.050 224.400 ;
        RECT 289.950 225.600 292.050 226.050 ;
        RECT 344.400 225.600 345.600 226.950 ;
        RECT 493.950 225.600 496.050 226.050 ;
        RECT 289.950 224.400 300.600 225.600 ;
        RECT 344.400 224.400 496.050 225.600 ;
        RECT 289.950 223.950 292.050 224.400 ;
        RECT 265.950 222.600 268.050 223.050 ;
        RECT 295.950 222.600 298.050 223.050 ;
        RECT 265.950 221.400 298.050 222.600 ;
        RECT 299.400 222.600 300.600 224.400 ;
        RECT 493.950 223.950 496.050 224.400 ;
        RECT 544.950 225.600 547.050 226.050 ;
        RECT 553.950 225.600 556.050 226.050 ;
        RECT 544.950 224.400 556.050 225.600 ;
        RECT 544.950 223.950 547.050 224.400 ;
        RECT 553.950 223.950 556.050 224.400 ;
        RECT 568.950 225.600 571.050 226.050 ;
        RECT 583.950 225.600 586.050 226.050 ;
        RECT 568.950 224.400 586.050 225.600 ;
        RECT 568.950 223.950 571.050 224.400 ;
        RECT 583.950 223.950 586.050 224.400 ;
        RECT 598.950 225.600 601.050 226.050 ;
        RECT 634.950 225.600 637.050 226.050 ;
        RECT 598.950 224.400 637.050 225.600 ;
        RECT 598.950 223.950 601.050 224.400 ;
        RECT 634.950 223.950 637.050 224.400 ;
        RECT 640.950 225.600 643.050 226.050 ;
        RECT 697.800 225.600 699.900 226.050 ;
        RECT 796.950 225.600 799.050 226.050 ;
        RECT 838.950 225.600 841.050 226.050 ;
        RECT 886.950 225.600 889.050 226.050 ;
        RECT 640.950 224.400 699.900 225.600 ;
        RECT 640.950 223.950 643.050 224.400 ;
        RECT 697.800 223.950 699.900 224.400 ;
        RECT 758.400 224.400 889.050 225.600 ;
        RECT 361.950 222.600 364.050 223.050 ;
        RECT 299.400 221.400 364.050 222.600 ;
        RECT 265.950 220.950 268.050 221.400 ;
        RECT 295.950 220.950 298.050 221.400 ;
        RECT 361.950 220.950 364.050 221.400 ;
        RECT 448.950 222.600 451.050 223.050 ;
        RECT 487.950 222.600 490.050 223.050 ;
        RECT 448.950 221.400 490.050 222.600 ;
        RECT 448.950 220.950 451.050 221.400 ;
        RECT 487.950 220.950 490.050 221.400 ;
        RECT 496.950 222.600 499.050 223.050 ;
        RECT 514.950 222.600 517.050 223.050 ;
        RECT 556.950 222.600 559.050 223.050 ;
        RECT 496.950 221.400 517.050 222.600 ;
        RECT 496.950 220.950 499.050 221.400 ;
        RECT 514.950 220.950 517.050 221.400 ;
        RECT 539.400 221.400 559.050 222.600 ;
        RECT 124.950 219.600 127.050 220.050 ;
        RECT 136.950 219.600 139.050 220.050 ;
        RECT 124.950 218.400 139.050 219.600 ;
        RECT 124.950 217.950 127.050 218.400 ;
        RECT 136.950 217.950 139.050 218.400 ;
        RECT 244.950 219.600 247.050 220.050 ;
        RECT 253.950 219.600 256.050 220.050 ;
        RECT 274.950 219.600 277.050 220.050 ;
        RECT 244.950 218.400 277.050 219.600 ;
        RECT 244.950 217.950 247.050 218.400 ;
        RECT 253.950 217.950 256.050 218.400 ;
        RECT 274.950 217.950 277.050 218.400 ;
        RECT 310.950 219.600 313.050 220.050 ;
        RECT 391.950 219.600 394.050 220.050 ;
        RECT 310.950 218.400 394.050 219.600 ;
        RECT 310.950 217.950 313.050 218.400 ;
        RECT 391.950 217.950 394.050 218.400 ;
        RECT 493.950 219.600 496.050 220.050 ;
        RECT 539.400 219.600 540.600 221.400 ;
        RECT 556.950 220.950 559.050 221.400 ;
        RECT 565.950 222.600 568.050 223.050 ;
        RECT 592.950 222.600 595.050 223.050 ;
        RECT 565.950 221.400 595.050 222.600 ;
        RECT 565.950 220.950 568.050 221.400 ;
        RECT 592.950 220.950 595.050 221.400 ;
        RECT 619.950 222.600 622.050 223.050 ;
        RECT 758.400 222.600 759.600 224.400 ;
        RECT 796.950 223.950 799.050 224.400 ;
        RECT 838.950 223.950 841.050 224.400 ;
        RECT 886.950 223.950 889.050 224.400 ;
        RECT 895.950 225.600 898.050 226.050 ;
        RECT 928.950 225.600 931.050 226.050 ;
        RECT 895.950 224.400 931.050 225.600 ;
        RECT 895.950 223.950 898.050 224.400 ;
        RECT 928.950 223.950 931.050 224.400 ;
        RECT 979.950 225.600 982.050 226.050 ;
        RECT 997.950 225.600 1000.050 226.050 ;
        RECT 979.950 224.400 1000.050 225.600 ;
        RECT 979.950 223.950 982.050 224.400 ;
        RECT 997.950 223.950 1000.050 224.400 ;
        RECT 619.950 221.400 759.600 222.600 ;
        RECT 811.950 222.600 814.050 223.050 ;
        RECT 853.950 222.600 856.050 223.050 ;
        RECT 811.950 221.400 856.050 222.600 ;
        RECT 619.950 220.950 622.050 221.400 ;
        RECT 811.950 220.950 814.050 221.400 ;
        RECT 853.950 220.950 856.050 221.400 ;
        RECT 907.950 222.600 910.050 223.050 ;
        RECT 913.950 222.600 916.050 223.050 ;
        RECT 925.950 222.600 928.050 223.050 ;
        RECT 907.950 221.400 928.050 222.600 ;
        RECT 907.950 220.950 910.050 221.400 ;
        RECT 913.950 220.950 916.050 221.400 ;
        RECT 925.950 220.950 928.050 221.400 ;
        RECT 934.950 222.600 937.050 223.050 ;
        RECT 949.950 222.600 952.050 223.050 ;
        RECT 934.950 221.400 952.050 222.600 ;
        RECT 934.950 220.950 937.050 221.400 ;
        RECT 949.950 220.950 952.050 221.400 ;
        RECT 586.950 219.600 589.050 220.050 ;
        RECT 493.950 218.400 540.600 219.600 ;
        RECT 569.400 218.400 589.050 219.600 ;
        RECT 493.950 217.950 496.050 218.400 ;
        RECT 40.950 216.600 43.050 217.200 ;
        RECT 43.950 216.600 46.050 217.050 ;
        RECT 61.950 216.600 64.050 217.200 ;
        RECT 40.950 215.400 64.050 216.600 ;
        RECT 40.950 215.100 43.050 215.400 ;
        RECT 43.950 214.950 46.050 215.400 ;
        RECT 61.950 215.100 64.050 215.400 ;
        RECT 73.950 216.750 76.050 217.200 ;
        RECT 82.950 216.750 85.050 217.200 ;
        RECT 73.950 215.550 85.050 216.750 ;
        RECT 73.950 215.100 76.050 215.550 ;
        RECT 82.950 215.100 85.050 215.550 ;
        RECT 97.950 216.600 100.050 217.050 ;
        RECT 106.950 216.600 109.050 217.200 ;
        RECT 97.950 215.400 109.050 216.600 ;
        RECT 97.950 214.950 100.050 215.400 ;
        RECT 106.950 215.100 109.050 215.400 ;
        RECT 145.950 216.600 148.050 217.050 ;
        RECT 157.950 216.600 160.050 217.200 ;
        RECT 145.950 215.400 160.050 216.600 ;
        RECT 145.950 214.950 148.050 215.400 ;
        RECT 157.950 215.100 160.050 215.400 ;
        RECT 163.950 216.750 166.050 217.200 ;
        RECT 175.950 216.750 178.050 217.200 ;
        RECT 163.950 215.550 178.050 216.750 ;
        RECT 163.950 215.100 166.050 215.550 ;
        RECT 175.950 215.100 178.050 215.550 ;
        RECT 250.950 216.600 253.050 217.200 ;
        RECT 280.950 216.600 283.050 217.200 ;
        RECT 319.950 216.600 322.050 217.200 ;
        RECT 250.950 215.400 283.050 216.600 ;
        RECT 250.950 215.100 253.050 215.400 ;
        RECT 280.950 215.100 283.050 215.400 ;
        RECT 317.400 215.400 322.050 216.600 ;
        RECT 281.400 213.600 282.600 215.100 ;
        RECT 281.400 212.400 294.600 213.600 ;
        RECT 154.950 210.600 157.050 210.900 ;
        RECT 163.950 210.600 166.050 211.050 ;
        RECT 178.950 210.600 181.050 210.900 ;
        RECT 154.950 209.400 181.050 210.600 ;
        RECT 154.950 208.800 157.050 209.400 ;
        RECT 163.950 208.950 166.050 209.400 ;
        RECT 178.950 208.800 181.050 209.400 ;
        RECT 208.950 210.600 211.050 210.900 ;
        RECT 217.950 210.600 220.050 211.050 ;
        RECT 226.950 210.600 229.050 210.900 ;
        RECT 208.950 209.400 229.050 210.600 ;
        RECT 208.950 208.800 211.050 209.400 ;
        RECT 217.950 208.950 220.050 209.400 ;
        RECT 226.950 208.800 229.050 209.400 ;
        RECT 238.950 210.450 241.050 210.900 ;
        RECT 247.950 210.450 250.050 210.900 ;
        RECT 238.950 209.250 250.050 210.450 ;
        RECT 238.950 208.800 241.050 209.250 ;
        RECT 247.950 208.800 250.050 209.250 ;
        RECT 271.950 210.600 274.050 210.900 ;
        RECT 286.950 210.600 289.050 211.050 ;
        RECT 271.950 209.400 289.050 210.600 ;
        RECT 293.400 210.600 294.600 212.400 ;
        RECT 298.950 210.600 301.050 210.900 ;
        RECT 293.400 209.400 301.050 210.600 ;
        RECT 271.950 208.800 274.050 209.400 ;
        RECT 286.950 208.950 289.050 209.400 ;
        RECT 298.950 208.800 301.050 209.400 ;
        RECT 37.950 207.600 40.050 208.050 ;
        RECT 52.950 207.600 55.050 208.050 ;
        RECT 73.950 207.600 76.050 208.050 ;
        RECT 37.950 206.400 76.050 207.600 ;
        RECT 37.950 205.950 40.050 206.400 ;
        RECT 52.950 205.950 55.050 206.400 ;
        RECT 73.950 205.950 76.050 206.400 ;
        RECT 109.950 207.600 112.050 208.050 ;
        RECT 124.950 207.600 127.050 208.050 ;
        RECT 109.950 206.400 127.050 207.600 ;
        RECT 109.950 205.950 112.050 206.400 ;
        RECT 124.950 205.950 127.050 206.400 ;
        RECT 289.950 207.600 292.050 208.050 ;
        RECT 304.950 207.600 307.050 208.050 ;
        RECT 289.950 206.400 307.050 207.600 ;
        RECT 289.950 205.950 292.050 206.400 ;
        RECT 304.950 205.950 307.050 206.400 ;
        RECT 310.950 207.600 313.050 208.050 ;
        RECT 317.400 207.600 318.600 215.400 ;
        RECT 319.950 215.100 322.050 215.400 ;
        RECT 400.950 215.100 403.050 217.200 ;
        RECT 430.950 216.750 433.050 217.200 ;
        RECT 439.950 216.750 442.050 217.200 ;
        RECT 430.950 215.550 442.050 216.750 ;
        RECT 430.950 215.100 433.050 215.550 ;
        RECT 439.950 215.100 442.050 215.550 ;
        RECT 469.950 215.100 472.050 217.200 ;
        RECT 478.950 216.750 481.050 217.200 ;
        RECT 490.950 216.750 493.050 217.200 ;
        RECT 478.950 215.550 493.050 216.750 ;
        RECT 478.950 215.100 481.050 215.550 ;
        RECT 490.950 215.100 493.050 215.550 ;
        RECT 517.950 216.600 520.050 217.200 ;
        RECT 541.950 216.600 544.050 217.050 ;
        RECT 517.950 215.400 544.050 216.600 ;
        RECT 517.950 215.100 520.050 215.400 ;
        RECT 401.400 211.050 402.600 215.100 ;
        RECT 470.400 211.050 471.600 215.100 ;
        RECT 541.950 214.950 544.050 215.400 ;
        RECT 547.950 215.100 550.050 217.200 ;
        RECT 559.950 216.600 562.050 217.050 ;
        RECT 569.400 216.600 570.600 218.400 ;
        RECT 586.950 217.950 589.050 218.400 ;
        RECT 709.950 219.600 712.050 220.050 ;
        RECT 742.950 219.600 745.050 220.050 ;
        RECT 760.950 219.600 763.050 220.050 ;
        RECT 709.950 218.400 723.600 219.600 ;
        RECT 709.950 217.950 712.050 218.400 ;
        RECT 559.950 215.400 570.600 216.600 ;
        RECT 604.950 216.750 607.050 217.200 ;
        RECT 616.950 216.750 619.050 217.200 ;
        RECT 604.950 215.550 619.050 216.750 ;
        RECT 322.950 210.600 325.050 211.050 ;
        RECT 328.950 210.600 331.050 211.050 ;
        RECT 322.950 209.400 331.050 210.600 ;
        RECT 322.950 208.950 325.050 209.400 ;
        RECT 328.950 208.950 331.050 209.400 ;
        RECT 343.950 210.450 346.050 210.900 ;
        RECT 358.950 210.450 361.050 210.900 ;
        RECT 343.950 209.250 361.050 210.450 ;
        RECT 343.950 208.800 346.050 209.250 ;
        RECT 358.950 208.800 361.050 209.250 ;
        RECT 376.950 210.600 379.050 211.050 ;
        RECT 385.950 210.600 388.050 210.900 ;
        RECT 376.950 209.400 388.050 210.600 ;
        RECT 401.400 209.400 406.050 211.050 ;
        RECT 376.950 208.950 379.050 209.400 ;
        RECT 385.950 208.800 388.050 209.400 ;
        RECT 402.000 208.950 406.050 209.400 ;
        RECT 433.950 210.600 436.050 211.050 ;
        RECT 442.950 210.600 445.050 210.900 ;
        RECT 433.950 209.400 445.050 210.600 ;
        RECT 433.950 208.950 436.050 209.400 ;
        RECT 442.950 208.800 445.050 209.400 ;
        RECT 466.950 209.400 471.600 211.050 ;
        RECT 505.950 210.600 508.050 211.050 ;
        RECT 511.950 210.600 514.050 211.050 ;
        RECT 505.950 209.400 514.050 210.600 ;
        RECT 466.950 208.950 471.000 209.400 ;
        RECT 505.950 208.950 508.050 209.400 ;
        RECT 511.950 208.950 514.050 209.400 ;
        RECT 310.950 206.400 318.600 207.600 ;
        RECT 373.950 207.600 376.050 208.050 ;
        RECT 418.950 207.600 421.050 208.050 ;
        RECT 430.950 207.600 433.050 208.050 ;
        RECT 373.950 206.400 433.050 207.600 ;
        RECT 310.950 205.950 313.050 206.400 ;
        RECT 373.950 205.950 376.050 206.400 ;
        RECT 418.950 205.950 421.050 206.400 ;
        RECT 430.950 205.950 433.050 206.400 ;
        RECT 499.950 207.600 502.050 208.050 ;
        RECT 548.400 207.600 549.600 215.100 ;
        RECT 559.950 214.950 562.050 215.400 ;
        RECT 604.950 215.100 607.050 215.550 ;
        RECT 616.950 215.100 619.050 215.550 ;
        RECT 553.950 213.600 556.050 214.050 ;
        RECT 580.950 213.600 583.050 214.050 ;
        RECT 628.950 213.600 631.050 217.050 ;
        RECT 661.950 216.600 664.050 217.200 ;
        RECT 553.950 212.400 567.600 213.600 ;
        RECT 553.950 211.950 556.050 212.400 ;
        RECT 566.400 210.600 567.600 212.400 ;
        RECT 580.950 213.000 631.050 213.600 ;
        RECT 641.400 215.400 664.050 216.600 ;
        RECT 580.950 212.400 630.600 213.000 ;
        RECT 580.950 211.950 583.050 212.400 ;
        RECT 568.950 210.600 571.050 210.900 ;
        RECT 566.400 209.400 571.050 210.600 ;
        RECT 568.950 208.800 571.050 209.400 ;
        RECT 607.950 208.950 610.050 212.400 ;
        RECT 637.950 210.600 640.050 210.900 ;
        RECT 641.400 210.600 642.600 215.400 ;
        RECT 661.950 215.100 664.050 215.400 ;
        RECT 688.950 216.600 691.050 217.200 ;
        RECT 703.950 216.600 706.050 217.050 ;
        RECT 688.950 215.400 706.050 216.600 ;
        RECT 722.400 216.600 723.600 218.400 ;
        RECT 742.950 218.400 763.050 219.600 ;
        RECT 742.950 217.950 745.050 218.400 ;
        RECT 760.950 217.950 763.050 218.400 ;
        RECT 997.950 219.600 1000.050 220.050 ;
        RECT 1006.950 219.600 1009.050 220.050 ;
        RECT 997.950 218.400 1009.050 219.600 ;
        RECT 997.950 217.950 1000.050 218.400 ;
        RECT 1006.950 217.950 1009.050 218.400 ;
        RECT 736.950 216.600 739.050 217.200 ;
        RECT 751.950 216.600 754.050 217.200 ;
        RECT 722.400 215.400 754.050 216.600 ;
        RECT 688.950 215.100 691.050 215.400 ;
        RECT 703.950 214.950 706.050 215.400 ;
        RECT 736.950 215.100 739.050 215.400 ;
        RECT 751.950 215.100 754.050 215.400 ;
        RECT 763.950 216.600 766.050 217.050 ;
        RECT 778.950 216.600 781.050 217.200 ;
        RECT 763.950 215.400 781.050 216.600 ;
        RECT 763.950 214.950 766.050 215.400 ;
        RECT 778.950 215.100 781.050 215.400 ;
        RECT 832.950 216.600 835.050 217.200 ;
        RECT 850.950 216.600 853.050 217.200 ;
        RECT 868.950 216.600 871.050 217.200 ;
        RECT 832.950 215.400 871.050 216.600 ;
        RECT 832.950 215.100 835.050 215.400 ;
        RECT 850.950 215.100 853.050 215.400 ;
        RECT 868.950 215.100 871.050 215.400 ;
        RECT 901.950 216.600 904.050 217.200 ;
        RECT 922.950 216.600 925.050 217.200 ;
        RECT 901.950 215.400 925.050 216.600 ;
        RECT 901.950 215.100 904.050 215.400 ;
        RECT 922.950 215.100 925.050 215.400 ;
        RECT 928.950 216.750 931.050 217.200 ;
        RECT 937.950 216.750 940.050 217.200 ;
        RECT 928.950 215.550 940.050 216.750 ;
        RECT 928.950 215.100 931.050 215.550 ;
        RECT 937.950 215.100 940.050 215.550 ;
        RECT 955.950 216.600 958.050 217.200 ;
        RECT 964.950 216.750 967.050 216.900 ;
        RECT 973.950 216.750 976.050 217.200 ;
        RECT 955.950 215.400 960.600 216.600 ;
        RECT 955.950 215.100 958.050 215.400 ;
        RECT 883.950 213.600 886.050 214.050 ;
        RECT 872.400 212.400 886.050 213.600 ;
        RECT 872.400 210.900 873.600 212.400 ;
        RECT 883.950 211.950 886.050 212.400 ;
        RECT 637.950 209.400 642.600 210.600 ;
        RECT 664.950 210.600 667.050 210.900 ;
        RECT 691.950 210.600 694.050 210.900 ;
        RECT 664.950 209.400 694.050 210.600 ;
        RECT 637.950 208.800 640.050 209.400 ;
        RECT 664.950 208.800 667.050 209.400 ;
        RECT 691.950 208.800 694.050 209.400 ;
        RECT 871.950 208.800 874.050 210.900 ;
        RECT 898.950 210.450 901.050 210.900 ;
        RECT 907.950 210.450 910.050 210.900 ;
        RECT 898.950 209.250 910.050 210.450 ;
        RECT 923.400 210.600 924.600 215.100 ;
        RECT 959.400 213.600 960.600 215.400 ;
        RECT 964.950 215.550 976.050 216.750 ;
        RECT 964.950 214.800 967.050 215.550 ;
        RECT 973.950 215.100 976.050 215.550 ;
        RECT 959.400 212.400 963.600 213.600 ;
        RECT 946.950 210.600 949.050 210.900 ;
        RECT 923.400 209.400 949.050 210.600 ;
        RECT 962.400 210.600 963.600 212.400 ;
        RECT 976.950 210.600 979.050 210.900 ;
        RECT 962.400 209.400 979.050 210.600 ;
        RECT 898.950 208.800 901.050 209.250 ;
        RECT 907.950 208.800 910.050 209.250 ;
        RECT 946.950 208.800 949.050 209.400 ;
        RECT 976.950 208.800 979.050 209.400 ;
        RECT 997.950 210.600 1000.050 210.900 ;
        RECT 1012.950 210.600 1015.050 211.050 ;
        RECT 997.950 209.400 1015.050 210.600 ;
        RECT 997.950 208.800 1000.050 209.400 ;
        RECT 1012.950 208.950 1015.050 209.400 ;
        RECT 499.950 206.400 549.600 207.600 ;
        RECT 613.950 207.600 616.050 208.050 ;
        RECT 649.950 207.600 652.050 208.050 ;
        RECT 673.950 207.600 676.050 208.050 ;
        RECT 613.950 206.400 652.050 207.600 ;
        RECT 499.950 205.950 502.050 206.400 ;
        RECT 613.950 205.950 616.050 206.400 ;
        RECT 649.950 205.950 652.050 206.400 ;
        RECT 662.400 206.400 676.050 207.600 ;
        RECT 22.950 204.600 25.050 205.050 ;
        RECT 58.950 204.600 61.050 205.050 ;
        RECT 22.950 203.400 61.050 204.600 ;
        RECT 22.950 202.950 25.050 203.400 ;
        RECT 58.950 202.950 61.050 203.400 ;
        RECT 253.950 204.600 256.050 205.050 ;
        RECT 259.950 204.600 262.050 205.050 ;
        RECT 253.950 203.400 262.050 204.600 ;
        RECT 253.950 202.950 256.050 203.400 ;
        RECT 259.950 202.950 262.050 203.400 ;
        RECT 484.950 204.600 487.050 205.050 ;
        RECT 547.950 204.600 550.050 205.050 ;
        RECT 484.950 203.400 550.050 204.600 ;
        RECT 484.950 202.950 487.050 203.400 ;
        RECT 547.950 202.950 550.050 203.400 ;
        RECT 568.950 204.600 571.050 205.050 ;
        RECT 646.950 204.600 649.050 205.050 ;
        RECT 568.950 203.400 649.050 204.600 ;
        RECT 568.950 202.950 571.050 203.400 ;
        RECT 646.950 202.950 649.050 203.400 ;
        RECT 655.950 204.600 658.050 205.050 ;
        RECT 662.400 204.600 663.600 206.400 ;
        RECT 673.950 205.950 676.050 206.400 ;
        RECT 715.950 207.600 718.050 208.050 ;
        RECT 772.950 207.600 775.050 208.050 ;
        RECT 715.950 206.400 775.050 207.600 ;
        RECT 715.950 205.950 718.050 206.400 ;
        RECT 772.950 205.950 775.050 206.400 ;
        RECT 805.950 207.600 808.050 208.050 ;
        RECT 913.950 207.600 916.050 208.050 ;
        RECT 925.950 207.600 928.050 208.050 ;
        RECT 805.950 206.400 819.600 207.600 ;
        RECT 805.950 205.950 808.050 206.400 ;
        RECT 818.400 205.050 819.600 206.400 ;
        RECT 913.950 206.400 928.050 207.600 ;
        RECT 913.950 205.950 916.050 206.400 ;
        RECT 925.950 205.950 928.050 206.400 ;
        RECT 985.950 207.600 988.050 208.050 ;
        RECT 1003.950 207.600 1006.050 208.050 ;
        RECT 985.950 206.400 1006.050 207.600 ;
        RECT 985.950 205.950 988.050 206.400 ;
        RECT 1003.950 205.950 1006.050 206.400 ;
        RECT 655.950 203.400 663.600 204.600 ;
        RECT 724.950 204.600 727.050 205.050 ;
        RECT 745.950 204.600 748.050 205.050 ;
        RECT 724.950 203.400 748.050 204.600 ;
        RECT 655.950 202.950 658.050 203.400 ;
        RECT 724.950 202.950 727.050 203.400 ;
        RECT 745.950 202.950 748.050 203.400 ;
        RECT 757.950 204.600 760.050 205.050 ;
        RECT 769.950 204.600 772.050 205.050 ;
        RECT 757.950 203.400 772.050 204.600 ;
        RECT 757.950 202.950 760.050 203.400 ;
        RECT 769.950 202.950 772.050 203.400 ;
        RECT 817.950 204.600 820.050 205.050 ;
        RECT 823.950 204.600 826.050 205.050 ;
        RECT 817.950 203.400 826.050 204.600 ;
        RECT 817.950 202.950 820.050 203.400 ;
        RECT 823.950 202.950 826.050 203.400 ;
        RECT 865.950 204.600 868.050 205.050 ;
        RECT 886.950 204.600 889.050 205.050 ;
        RECT 865.950 203.400 889.050 204.600 ;
        RECT 865.950 202.950 868.050 203.400 ;
        RECT 886.950 202.950 889.050 203.400 ;
        RECT 262.950 201.600 265.050 202.050 ;
        RECT 337.950 201.600 340.050 202.050 ;
        RECT 262.950 200.400 340.050 201.600 ;
        RECT 262.950 199.950 265.050 200.400 ;
        RECT 337.950 199.950 340.050 200.400 ;
        RECT 517.950 201.600 520.050 202.050 ;
        RECT 526.950 201.600 529.050 202.050 ;
        RECT 517.950 200.400 529.050 201.600 ;
        RECT 517.950 199.950 520.050 200.400 ;
        RECT 526.950 199.950 529.050 200.400 ;
        RECT 652.950 201.600 655.050 202.050 ;
        RECT 725.400 201.600 726.600 202.950 ;
        RECT 652.950 200.400 726.600 201.600 ;
        RECT 751.950 201.600 754.050 202.050 ;
        RECT 766.950 201.600 769.050 202.050 ;
        RECT 805.950 201.600 808.050 202.050 ;
        RECT 751.950 200.400 808.050 201.600 ;
        RECT 652.950 199.950 655.050 200.400 ;
        RECT 751.950 199.950 754.050 200.400 ;
        RECT 766.950 199.950 769.050 200.400 ;
        RECT 805.950 199.950 808.050 200.400 ;
        RECT 850.950 201.600 853.050 202.050 ;
        RECT 910.950 201.600 913.050 202.050 ;
        RECT 850.950 200.400 913.050 201.600 ;
        RECT 850.950 199.950 853.050 200.400 ;
        RECT 910.950 199.950 913.050 200.400 ;
        RECT 922.950 201.600 925.050 202.050 ;
        RECT 940.950 201.600 943.050 202.050 ;
        RECT 922.950 200.400 943.050 201.600 ;
        RECT 922.950 199.950 925.050 200.400 ;
        RECT 940.950 199.950 943.050 200.400 ;
        RECT 952.950 201.600 955.050 202.050 ;
        RECT 985.950 201.600 988.050 202.050 ;
        RECT 952.950 200.400 988.050 201.600 ;
        RECT 952.950 199.950 955.050 200.400 ;
        RECT 985.950 199.950 988.050 200.400 ;
        RECT 73.950 198.600 76.050 199.050 ;
        RECT 85.950 198.600 88.050 199.050 ;
        RECT 73.950 197.400 88.050 198.600 ;
        RECT 73.950 196.950 76.050 197.400 ;
        RECT 85.950 196.950 88.050 197.400 ;
        RECT 115.950 198.600 118.050 199.050 ;
        RECT 142.950 198.600 145.050 199.050 ;
        RECT 115.950 197.400 145.050 198.600 ;
        RECT 115.950 196.950 118.050 197.400 ;
        RECT 142.950 196.950 145.050 197.400 ;
        RECT 226.950 198.600 229.050 199.050 ;
        RECT 253.950 198.600 256.050 199.050 ;
        RECT 226.950 197.400 256.050 198.600 ;
        RECT 226.950 196.950 229.050 197.400 ;
        RECT 253.950 196.950 256.050 197.400 ;
        RECT 409.950 198.600 412.050 199.050 ;
        RECT 415.950 198.600 418.050 199.050 ;
        RECT 409.950 197.400 418.050 198.600 ;
        RECT 409.950 196.950 412.050 197.400 ;
        RECT 415.950 196.950 418.050 197.400 ;
        RECT 427.950 198.600 430.050 199.050 ;
        RECT 451.950 198.600 454.050 199.050 ;
        RECT 427.950 197.400 454.050 198.600 ;
        RECT 427.950 196.950 430.050 197.400 ;
        RECT 451.950 196.950 454.050 197.400 ;
        RECT 460.950 198.600 463.050 199.050 ;
        RECT 550.950 198.600 553.050 199.050 ;
        RECT 460.950 197.400 553.050 198.600 ;
        RECT 460.950 196.950 463.050 197.400 ;
        RECT 550.950 196.950 553.050 197.400 ;
        RECT 598.950 198.600 601.050 199.050 ;
        RECT 604.950 198.600 607.050 199.050 ;
        RECT 598.950 197.400 607.050 198.600 ;
        RECT 598.950 196.950 601.050 197.400 ;
        RECT 604.950 196.950 607.050 197.400 ;
        RECT 658.950 198.600 661.050 199.050 ;
        RECT 694.950 198.600 697.050 199.050 ;
        RECT 658.950 197.400 697.050 198.600 ;
        RECT 658.950 196.950 661.050 197.400 ;
        RECT 694.950 196.950 697.050 197.400 ;
        RECT 781.950 198.600 784.050 199.050 ;
        RECT 790.950 198.600 793.050 199.050 ;
        RECT 781.950 197.400 793.050 198.600 ;
        RECT 781.950 196.950 784.050 197.400 ;
        RECT 790.950 196.950 793.050 197.400 ;
        RECT 964.950 198.600 967.050 199.050 ;
        RECT 979.950 198.600 982.050 199.050 ;
        RECT 964.950 197.400 982.050 198.600 ;
        RECT 964.950 196.950 967.050 197.400 ;
        RECT 979.950 196.950 982.050 197.400 ;
        RECT 70.950 195.600 73.050 196.050 ;
        RECT 91.950 195.600 94.050 196.050 ;
        RECT 274.950 195.600 277.050 196.050 ;
        RECT 70.950 194.400 277.050 195.600 ;
        RECT 70.950 193.950 73.050 194.400 ;
        RECT 91.950 193.950 94.050 194.400 ;
        RECT 274.950 193.950 277.050 194.400 ;
        RECT 301.950 195.600 304.050 196.050 ;
        RECT 310.950 195.600 313.050 196.050 ;
        RECT 301.950 194.400 313.050 195.600 ;
        RECT 301.950 193.950 304.050 194.400 ;
        RECT 310.950 193.950 313.050 194.400 ;
        RECT 466.950 195.600 469.050 196.050 ;
        RECT 475.950 195.600 478.050 196.050 ;
        RECT 466.950 194.400 478.050 195.600 ;
        RECT 466.950 193.950 469.050 194.400 ;
        RECT 475.950 193.950 478.050 194.400 ;
        RECT 547.950 195.600 550.050 196.050 ;
        RECT 568.950 195.600 571.050 196.050 ;
        RECT 547.950 194.400 571.050 195.600 ;
        RECT 547.950 193.950 550.050 194.400 ;
        RECT 568.950 193.950 571.050 194.400 ;
        RECT 574.950 195.600 577.050 196.050 ;
        RECT 619.950 195.600 622.050 196.050 ;
        RECT 574.950 194.400 622.050 195.600 ;
        RECT 574.950 193.950 577.050 194.400 ;
        RECT 619.950 193.950 622.050 194.400 ;
        RECT 697.950 195.600 700.050 196.050 ;
        RECT 703.950 195.600 706.050 196.050 ;
        RECT 697.950 194.400 706.050 195.600 ;
        RECT 697.950 193.950 700.050 194.400 ;
        RECT 703.950 193.950 706.050 194.400 ;
        RECT 838.950 195.600 841.050 196.050 ;
        RECT 874.950 195.600 877.050 196.050 ;
        RECT 838.950 194.400 877.050 195.600 ;
        RECT 838.950 193.950 841.050 194.400 ;
        RECT 874.950 193.950 877.050 194.400 ;
        RECT 880.950 195.600 883.050 196.050 ;
        RECT 889.950 195.600 892.050 196.050 ;
        RECT 880.950 194.400 892.050 195.600 ;
        RECT 880.950 193.950 883.050 194.400 ;
        RECT 889.950 193.950 892.050 194.400 ;
        RECT 940.950 195.600 943.050 196.050 ;
        RECT 964.950 195.600 967.050 195.900 ;
        RECT 940.950 194.400 967.050 195.600 ;
        RECT 940.950 193.950 943.050 194.400 ;
        RECT 100.950 192.600 103.050 193.050 ;
        RECT 130.950 192.600 133.050 193.050 ;
        RECT 100.950 191.400 133.050 192.600 ;
        RECT 100.950 190.950 103.050 191.400 ;
        RECT 130.950 190.950 133.050 191.400 ;
        RECT 172.950 192.600 175.050 193.050 ;
        RECT 187.950 192.600 190.050 193.050 ;
        RECT 202.950 192.600 205.050 193.050 ;
        RECT 172.950 191.400 205.050 192.600 ;
        RECT 172.950 190.950 175.050 191.400 ;
        RECT 187.950 190.950 190.050 191.400 ;
        RECT 202.950 190.950 205.050 191.400 ;
        RECT 253.950 192.600 256.050 193.050 ;
        RECT 302.400 192.600 303.600 193.950 ;
        RECT 964.950 193.800 967.050 194.400 ;
        RECT 253.950 191.400 303.600 192.600 ;
        RECT 334.950 192.600 337.050 193.050 ;
        RECT 343.950 192.600 346.050 193.050 ;
        RECT 460.950 192.600 463.050 193.050 ;
        RECT 481.950 192.600 484.050 193.050 ;
        RECT 334.950 191.400 346.050 192.600 ;
        RECT 253.950 190.950 256.050 191.400 ;
        RECT 334.950 190.950 337.050 191.400 ;
        RECT 343.950 190.950 346.050 191.400 ;
        RECT 362.400 191.400 484.050 192.600 ;
        RECT 362.400 190.050 363.600 191.400 ;
        RECT 460.950 190.950 463.050 191.400 ;
        RECT 481.950 190.950 484.050 191.400 ;
        RECT 658.950 192.600 661.050 193.050 ;
        RECT 742.950 192.600 745.050 193.050 ;
        RECT 658.950 191.400 745.050 192.600 ;
        RECT 658.950 190.950 661.050 191.400 ;
        RECT 742.950 190.950 745.050 191.400 ;
        RECT 910.950 192.600 913.050 193.050 ;
        RECT 919.950 192.600 922.050 193.050 ;
        RECT 910.950 191.400 922.050 192.600 ;
        RECT 910.950 190.950 913.050 191.400 ;
        RECT 919.950 190.950 922.050 191.400 ;
        RECT 937.950 192.600 940.050 193.050 ;
        RECT 937.950 191.400 987.600 192.600 ;
        RECT 937.950 190.950 940.050 191.400 ;
        RECT 986.400 190.050 987.600 191.400 ;
        RECT 118.950 189.600 121.050 190.050 ;
        RECT 136.950 189.600 139.050 190.050 ;
        RECT 86.400 188.400 139.050 189.600 ;
        RECT 86.400 187.050 87.600 188.400 ;
        RECT 118.950 187.950 121.050 188.400 ;
        RECT 136.950 187.950 139.050 188.400 ;
        RECT 148.950 189.600 151.050 190.050 ;
        RECT 160.950 189.600 163.050 190.050 ;
        RECT 148.950 188.400 163.050 189.600 ;
        RECT 148.950 187.950 151.050 188.400 ;
        RECT 160.950 187.950 163.050 188.400 ;
        RECT 166.950 189.600 169.050 190.050 ;
        RECT 280.950 189.600 283.050 190.050 ;
        RECT 307.950 189.600 310.050 190.050 ;
        RECT 361.950 189.600 364.050 190.050 ;
        RECT 166.950 188.400 364.050 189.600 ;
        RECT 166.950 187.950 169.050 188.400 ;
        RECT 280.950 187.950 283.050 188.400 ;
        RECT 307.950 187.950 310.050 188.400 ;
        RECT 361.950 187.950 364.050 188.400 ;
        RECT 367.950 189.600 370.050 190.050 ;
        RECT 424.950 189.600 427.050 190.050 ;
        RECT 367.950 188.400 427.050 189.600 ;
        RECT 367.950 187.950 370.050 188.400 ;
        RECT 424.950 187.950 427.050 188.400 ;
        RECT 532.950 189.600 535.050 190.050 ;
        RECT 538.950 189.600 541.050 190.050 ;
        RECT 559.950 189.600 562.050 190.050 ;
        RECT 586.950 189.600 589.050 190.050 ;
        RECT 532.950 188.400 562.050 189.600 ;
        RECT 532.950 187.950 535.050 188.400 ;
        RECT 538.950 187.950 541.050 188.400 ;
        RECT 559.950 187.950 562.050 188.400 ;
        RECT 578.400 188.400 589.050 189.600 ;
        RECT 58.950 186.600 61.050 187.050 ;
        RECT 85.950 186.600 88.050 187.050 ;
        RECT 58.950 185.400 88.050 186.600 ;
        RECT 58.950 184.950 61.050 185.400 ;
        RECT 85.950 184.950 88.050 185.400 ;
        RECT 238.950 186.600 241.050 187.050 ;
        RECT 277.950 186.600 280.050 187.050 ;
        RECT 238.950 185.400 280.050 186.600 ;
        RECT 238.950 184.950 241.050 185.400 ;
        RECT 277.950 184.950 280.050 185.400 ;
        RECT 310.950 186.600 313.050 187.050 ;
        RECT 349.950 186.600 352.050 187.050 ;
        RECT 310.950 185.400 352.050 186.600 ;
        RECT 310.950 184.950 313.050 185.400 ;
        RECT 349.950 184.950 352.050 185.400 ;
        RECT 562.950 186.600 565.050 187.050 ;
        RECT 578.400 186.600 579.600 188.400 ;
        RECT 586.950 187.950 589.050 188.400 ;
        RECT 640.950 189.600 643.050 190.050 ;
        RECT 652.950 189.600 655.050 190.050 ;
        RECT 640.950 188.400 655.050 189.600 ;
        RECT 640.950 187.950 643.050 188.400 ;
        RECT 652.950 187.950 655.050 188.400 ;
        RECT 676.950 189.600 679.050 190.050 ;
        RECT 703.950 189.600 706.050 190.050 ;
        RECT 676.950 188.400 706.050 189.600 ;
        RECT 676.950 187.950 679.050 188.400 ;
        RECT 703.950 187.950 706.050 188.400 ;
        RECT 832.950 189.600 835.050 190.050 ;
        RECT 865.950 189.600 868.050 190.050 ;
        RECT 832.950 188.400 868.050 189.600 ;
        RECT 832.950 187.950 835.050 188.400 ;
        RECT 865.950 187.950 868.050 188.400 ;
        RECT 901.950 189.600 904.050 190.050 ;
        RECT 928.950 189.600 931.050 190.050 ;
        RECT 901.950 188.400 931.050 189.600 ;
        RECT 901.950 187.950 904.050 188.400 ;
        RECT 928.950 187.950 931.050 188.400 ;
        RECT 943.950 189.600 946.050 190.050 ;
        RECT 955.950 189.600 958.050 190.050 ;
        RECT 943.950 188.400 958.050 189.600 ;
        RECT 986.400 188.400 991.050 190.050 ;
        RECT 943.950 187.950 946.050 188.400 ;
        RECT 955.950 187.950 958.050 188.400 ;
        RECT 987.000 187.950 991.050 188.400 ;
        RECT 562.950 185.400 579.600 186.600 ;
        RECT 562.950 184.950 565.050 185.400 ;
        RECT 16.950 183.600 19.050 184.200 ;
        RECT 28.950 183.600 31.050 184.050 ;
        RECT 16.950 182.400 31.050 183.600 ;
        RECT 16.950 182.100 19.050 182.400 ;
        RECT 28.950 181.950 31.050 182.400 ;
        RECT 40.950 183.600 43.050 184.200 ;
        RECT 91.950 183.600 94.050 184.200 ;
        RECT 40.950 182.400 57.600 183.600 ;
        RECT 40.950 182.100 43.050 182.400 ;
        RECT 56.400 177.600 57.600 182.400 ;
        RECT 91.950 182.400 96.600 183.600 ;
        RECT 91.950 182.100 94.050 182.400 ;
        RECT 95.400 178.050 96.600 182.400 ;
        RECT 106.950 182.100 109.050 184.200 ;
        RECT 115.950 183.750 118.050 184.200 ;
        RECT 127.950 183.750 130.050 184.200 ;
        RECT 115.950 182.550 130.050 183.750 ;
        RECT 115.950 182.100 118.050 182.550 ;
        RECT 127.950 182.100 130.050 182.550 ;
        RECT 133.950 183.600 136.050 184.200 ;
        RECT 148.950 183.600 151.050 184.050 ;
        RECT 133.950 182.400 151.050 183.600 ;
        RECT 133.950 182.100 136.050 182.400 ;
        RECT 61.950 177.600 64.050 177.900 ;
        RECT 56.400 176.400 64.050 177.600 ;
        RECT 61.950 175.800 64.050 176.400 ;
        RECT 67.950 177.450 70.050 177.900 ;
        RECT 73.950 177.450 76.050 177.900 ;
        RECT 67.950 176.250 76.050 177.450 ;
        RECT 67.950 175.800 70.050 176.250 ;
        RECT 73.950 175.800 76.050 176.250 ;
        RECT 94.950 175.950 97.050 178.050 ;
        RECT 107.400 174.600 108.600 182.100 ;
        RECT 148.950 181.950 151.050 182.400 ;
        RECT 154.950 183.600 157.050 184.200 ;
        RECT 169.950 183.750 172.050 184.200 ;
        RECT 196.950 183.750 199.050 184.200 ;
        RECT 154.950 182.400 165.600 183.600 ;
        RECT 154.950 182.100 157.050 182.400 ;
        RECT 164.400 180.600 165.600 182.400 ;
        RECT 169.950 182.550 199.050 183.750 ;
        RECT 169.950 182.100 172.050 182.550 ;
        RECT 196.950 182.100 199.050 182.550 ;
        RECT 208.950 183.600 211.050 184.050 ;
        RECT 220.950 183.600 223.050 184.200 ;
        RECT 208.950 182.400 223.050 183.600 ;
        RECT 208.950 181.950 211.050 182.400 ;
        RECT 220.950 182.100 223.050 182.400 ;
        RECT 289.950 183.600 292.050 184.200 ;
        RECT 298.950 183.600 301.050 184.050 ;
        RECT 289.950 182.400 301.050 183.600 ;
        RECT 289.950 182.100 292.050 182.400 ;
        RECT 298.950 181.950 301.050 182.400 ;
        RECT 307.950 183.600 310.050 184.200 ;
        RECT 307.950 182.400 333.600 183.600 ;
        RECT 307.950 182.100 310.050 182.400 ;
        RECT 184.950 180.600 187.050 181.050 ;
        RECT 164.400 179.400 187.050 180.600 ;
        RECT 184.950 178.950 187.050 179.400 ;
        RECT 332.400 177.900 333.600 182.400 ;
        RECT 340.950 181.950 343.050 184.050 ;
        RECT 355.950 182.100 358.050 184.200 ;
        RECT 382.950 183.600 385.050 184.200 ;
        RECT 391.950 183.600 394.050 184.050 ;
        RECT 382.950 182.400 394.050 183.600 ;
        RECT 382.950 182.100 385.050 182.400 ;
        RECT 136.950 177.450 139.050 177.900 ;
        RECT 145.950 177.600 148.050 177.900 ;
        RECT 157.950 177.600 160.050 177.900 ;
        RECT 145.950 177.450 160.050 177.600 ;
        RECT 136.950 176.400 160.050 177.450 ;
        RECT 136.950 176.250 148.050 176.400 ;
        RECT 136.950 175.800 139.050 176.250 ;
        RECT 145.950 175.800 148.050 176.250 ;
        RECT 157.950 175.800 160.050 176.400 ;
        RECT 175.950 177.600 178.050 177.900 ;
        RECT 193.950 177.600 196.050 177.900 ;
        RECT 175.950 176.400 196.050 177.600 ;
        RECT 175.950 175.800 178.050 176.400 ;
        RECT 193.950 175.800 196.050 176.400 ;
        RECT 223.950 177.600 226.050 177.900 ;
        RECT 244.950 177.600 247.050 177.900 ;
        RECT 223.950 176.400 247.050 177.600 ;
        RECT 223.950 175.800 226.050 176.400 ;
        RECT 244.950 175.800 247.050 176.400 ;
        RECT 280.950 177.450 283.050 177.900 ;
        RECT 286.950 177.450 289.050 177.900 ;
        RECT 280.950 176.250 289.050 177.450 ;
        RECT 280.950 175.800 283.050 176.250 ;
        RECT 286.950 175.800 289.050 176.250 ;
        RECT 301.950 177.450 304.050 177.900 ;
        RECT 310.950 177.450 313.050 177.900 ;
        RECT 301.950 176.250 313.050 177.450 ;
        RECT 301.950 175.800 304.050 176.250 ;
        RECT 310.950 175.800 313.050 176.250 ;
        RECT 331.950 175.800 334.050 177.900 ;
        RECT 337.950 177.600 340.050 177.900 ;
        RECT 341.400 177.600 342.600 181.950 ;
        RECT 337.950 176.400 342.600 177.600 ;
        RECT 349.950 177.600 352.050 178.050 ;
        RECT 356.400 177.600 357.600 182.100 ;
        RECT 391.950 181.950 394.050 182.400 ;
        RECT 409.950 183.600 412.050 184.200 ;
        RECT 418.800 183.600 420.900 184.050 ;
        RECT 409.950 182.400 420.900 183.600 ;
        RECT 409.950 182.100 412.050 182.400 ;
        RECT 418.800 181.950 420.900 182.400 ;
        RECT 421.950 183.600 424.050 184.050 ;
        RECT 430.950 183.600 433.050 184.200 ;
        RECT 421.950 182.400 433.050 183.600 ;
        RECT 421.950 181.950 424.050 182.400 ;
        RECT 430.950 182.100 433.050 182.400 ;
        RECT 451.950 183.600 454.050 184.200 ;
        RECT 466.950 183.600 469.050 184.050 ;
        RECT 451.950 182.400 469.050 183.600 ;
        RECT 451.950 182.100 454.050 182.400 ;
        RECT 466.950 181.950 469.050 182.400 ;
        RECT 496.950 183.600 499.050 184.200 ;
        RECT 523.950 183.600 526.050 184.200 ;
        RECT 496.950 182.400 526.050 183.600 ;
        RECT 496.950 182.100 499.050 182.400 ;
        RECT 523.950 182.100 526.050 182.400 ;
        RECT 556.950 182.100 559.050 184.200 ;
        RECT 574.950 183.600 577.050 184.050 ;
        RECT 580.950 183.600 583.050 184.200 ;
        RECT 574.950 182.400 583.050 183.600 ;
        RECT 604.950 183.600 607.050 187.050 ;
        RECT 733.950 184.950 736.050 187.050 ;
        RECT 829.950 186.600 832.050 187.050 ;
        RECT 850.950 186.600 853.050 187.050 ;
        RECT 829.950 185.400 853.050 186.600 ;
        RECT 829.950 184.950 832.050 185.400 ;
        RECT 850.950 184.950 853.050 185.400 ;
        RECT 880.950 186.600 883.050 187.050 ;
        RECT 895.800 186.600 897.900 187.050 ;
        RECT 880.950 185.400 897.900 186.600 ;
        RECT 880.950 184.950 883.050 185.400 ;
        RECT 895.800 184.950 897.900 185.400 ;
        RECT 898.950 186.600 901.050 187.050 ;
        RECT 937.950 186.600 940.050 187.050 ;
        RECT 898.950 185.400 940.050 186.600 ;
        RECT 898.950 184.950 901.050 185.400 ;
        RECT 937.950 184.950 940.050 185.400 ;
        RECT 613.950 183.600 616.050 184.200 ;
        RECT 604.950 183.000 616.050 183.600 ;
        RECT 605.400 182.400 616.050 183.000 ;
        RECT 557.400 180.600 558.600 182.100 ;
        RECT 574.950 181.950 577.050 182.400 ;
        RECT 580.950 182.100 583.050 182.400 ;
        RECT 613.950 182.100 616.050 182.400 ;
        RECT 634.950 182.100 637.050 184.200 ;
        RECT 646.950 183.750 649.050 184.200 ;
        RECT 655.950 183.750 658.050 184.200 ;
        RECT 646.950 182.550 658.050 183.750 ;
        RECT 646.950 182.100 649.050 182.550 ;
        RECT 655.950 182.100 658.050 182.550 ;
        RECT 679.950 183.750 682.050 184.200 ;
        RECT 685.950 183.750 688.050 184.200 ;
        RECT 679.950 182.550 688.050 183.750 ;
        RECT 679.950 182.100 682.050 182.550 ;
        RECT 685.950 182.100 688.050 182.550 ;
        RECT 709.950 183.600 712.050 184.200 ;
        RECT 721.950 183.750 724.050 184.200 ;
        RECT 730.950 183.750 733.050 184.200 ;
        RECT 709.950 182.400 714.600 183.600 ;
        RECT 709.950 182.100 712.050 182.400 ;
        RECT 635.400 180.600 636.600 182.100 ;
        RECT 673.950 180.600 676.050 181.050 ;
        RECT 479.400 179.400 676.050 180.600 ;
        RECT 349.950 176.400 357.600 177.600 ;
        RECT 358.950 177.450 361.050 177.900 ;
        RECT 367.950 177.450 370.050 177.900 ;
        RECT 337.950 175.800 340.050 176.400 ;
        RECT 349.950 175.950 352.050 176.400 ;
        RECT 358.950 176.250 370.050 177.450 ;
        RECT 358.950 175.800 361.050 176.250 ;
        RECT 367.950 175.800 370.050 176.250 ;
        RECT 373.950 177.600 376.050 178.050 ;
        RECT 479.400 177.900 480.600 179.400 ;
        RECT 673.950 178.950 676.050 179.400 ;
        RECT 379.950 177.600 382.050 177.900 ;
        RECT 373.950 176.400 382.050 177.600 ;
        RECT 373.950 175.950 376.050 176.400 ;
        RECT 379.950 175.800 382.050 176.400 ;
        RECT 385.950 177.600 388.050 177.900 ;
        RECT 385.950 176.400 420.600 177.600 ;
        RECT 385.950 175.800 388.050 176.400 ;
        RECT 419.400 175.050 420.600 176.400 ;
        RECT 466.950 177.450 469.050 177.900 ;
        RECT 472.950 177.450 475.050 177.900 ;
        RECT 466.950 176.250 475.050 177.450 ;
        RECT 466.950 175.800 469.050 176.250 ;
        RECT 472.950 175.800 475.050 176.250 ;
        RECT 478.950 175.800 481.050 177.900 ;
        RECT 514.950 177.450 517.050 177.900 ;
        RECT 529.950 177.450 532.050 177.900 ;
        RECT 514.950 176.250 532.050 177.450 ;
        RECT 514.950 175.800 517.050 176.250 ;
        RECT 529.950 175.800 532.050 176.250 ;
        RECT 589.950 177.450 592.050 177.900 ;
        RECT 595.950 177.450 598.050 177.900 ;
        RECT 589.950 176.250 598.050 177.450 ;
        RECT 589.950 175.800 592.050 176.250 ;
        RECT 595.950 175.800 598.050 176.250 ;
        RECT 655.950 177.600 658.050 177.900 ;
        RECT 697.950 177.600 700.050 177.900 ;
        RECT 655.950 177.450 700.050 177.600 ;
        RECT 706.950 177.450 709.050 177.900 ;
        RECT 655.950 176.400 709.050 177.450 ;
        RECT 655.950 175.800 658.050 176.400 ;
        RECT 697.950 176.250 709.050 176.400 ;
        RECT 697.950 175.800 700.050 176.250 ;
        RECT 706.950 175.800 709.050 176.250 ;
        RECT 130.950 174.600 133.050 175.050 ;
        RECT 107.400 173.400 133.050 174.600 ;
        RECT 130.950 172.950 133.050 173.400 ;
        RECT 199.950 174.600 202.050 175.050 ;
        RECT 208.950 174.600 211.050 175.050 ;
        RECT 199.950 173.400 211.050 174.600 ;
        RECT 199.950 172.950 202.050 173.400 ;
        RECT 208.950 172.950 211.050 173.400 ;
        RECT 403.950 174.600 406.050 175.050 ;
        RECT 415.800 174.600 417.900 175.050 ;
        RECT 403.950 173.400 417.900 174.600 ;
        RECT 403.950 172.950 406.050 173.400 ;
        RECT 415.800 172.950 417.900 173.400 ;
        RECT 418.950 174.600 421.050 175.050 ;
        RECT 427.950 174.600 430.050 175.050 ;
        RECT 418.950 173.400 430.050 174.600 ;
        RECT 418.950 172.950 421.050 173.400 ;
        RECT 427.950 172.950 430.050 173.400 ;
        RECT 601.950 174.600 604.050 175.050 ;
        RECT 610.950 174.600 613.050 175.050 ;
        RECT 637.950 174.600 640.050 175.050 ;
        RECT 601.950 173.400 640.050 174.600 ;
        RECT 601.950 172.950 604.050 173.400 ;
        RECT 610.950 172.950 613.050 173.400 ;
        RECT 637.950 172.950 640.050 173.400 ;
        RECT 43.950 171.600 46.050 172.050 ;
        RECT 82.950 171.600 85.050 172.050 ;
        RECT 97.950 171.600 100.050 172.050 ;
        RECT 43.950 170.400 100.050 171.600 ;
        RECT 43.950 169.950 46.050 170.400 ;
        RECT 82.950 169.950 85.050 170.400 ;
        RECT 97.950 169.950 100.050 170.400 ;
        RECT 622.950 171.600 625.050 172.050 ;
        RECT 713.400 171.900 714.600 182.400 ;
        RECT 721.950 182.550 733.050 183.750 ;
        RECT 721.950 182.100 724.050 182.550 ;
        RECT 730.950 182.100 733.050 182.550 ;
        RECT 734.400 177.900 735.600 184.950 ;
        RECT 736.950 183.600 739.050 184.200 ;
        RECT 742.950 183.600 745.050 184.050 ;
        RECT 748.950 183.600 751.050 184.050 ;
        RECT 736.950 182.400 741.600 183.600 ;
        RECT 736.950 182.100 739.050 182.400 ;
        RECT 733.950 175.800 736.050 177.900 ;
        RECT 740.400 174.600 741.600 182.400 ;
        RECT 742.950 182.400 751.050 183.600 ;
        RECT 742.950 181.950 745.050 182.400 ;
        RECT 748.950 181.950 751.050 182.400 ;
        RECT 772.950 183.600 775.050 184.050 ;
        RECT 781.950 183.750 784.050 184.200 ;
        RECT 793.950 183.750 796.050 184.200 ;
        RECT 781.950 183.600 796.050 183.750 ;
        RECT 772.950 182.550 796.050 183.600 ;
        RECT 772.950 182.400 784.050 182.550 ;
        RECT 772.950 181.950 775.050 182.400 ;
        RECT 781.950 182.100 784.050 182.400 ;
        RECT 793.950 182.100 796.050 182.550 ;
        RECT 856.950 183.600 859.050 184.200 ;
        RECT 907.950 183.600 910.050 184.050 ;
        RECT 916.950 183.600 919.050 184.200 ;
        RECT 856.950 182.400 897.600 183.600 ;
        RECT 856.950 182.100 859.050 182.400 ;
        RECT 896.400 180.600 897.600 182.400 ;
        RECT 907.950 182.400 919.050 183.600 ;
        RECT 907.950 181.950 910.050 182.400 ;
        RECT 916.950 182.100 919.050 182.400 ;
        RECT 946.950 183.600 949.050 184.200 ;
        RECT 970.950 183.600 973.050 184.200 ;
        RECT 985.950 183.600 988.050 184.050 ;
        RECT 946.950 182.400 973.050 183.600 ;
        RECT 946.950 182.100 949.050 182.400 ;
        RECT 970.950 182.100 973.050 182.400 ;
        RECT 974.400 182.400 988.050 183.600 ;
        RECT 974.400 180.600 975.600 182.400 ;
        RECT 985.950 181.950 988.050 182.400 ;
        RECT 896.400 180.000 906.600 180.600 ;
        RECT 896.400 179.400 907.050 180.000 ;
        RECT 760.950 177.600 763.050 177.900 ;
        RECT 778.950 177.600 781.050 177.900 ;
        RECT 760.950 176.400 781.050 177.600 ;
        RECT 760.950 175.800 763.050 176.400 ;
        RECT 778.950 175.800 781.050 176.400 ;
        RECT 787.950 177.600 790.050 177.900 ;
        RECT 802.950 177.600 805.050 177.900 ;
        RECT 787.950 176.400 805.050 177.600 ;
        RECT 787.950 175.800 790.050 176.400 ;
        RECT 802.950 175.800 805.050 176.400 ;
        RECT 841.950 177.450 844.050 177.900 ;
        RECT 853.950 177.450 856.050 177.900 ;
        RECT 841.950 176.250 856.050 177.450 ;
        RECT 841.950 175.800 844.050 176.250 ;
        RECT 853.950 175.800 856.050 176.250 ;
        RECT 868.950 177.450 871.050 177.900 ;
        RECT 895.950 177.450 898.050 177.900 ;
        RECT 868.950 176.250 898.050 177.450 ;
        RECT 868.950 175.800 871.050 176.250 ;
        RECT 895.950 175.800 898.050 176.250 ;
        RECT 904.950 175.950 907.050 179.400 ;
        RECT 968.400 179.400 975.600 180.600 ;
        RECT 968.400 177.900 969.600 179.400 ;
        RECT 910.950 177.450 913.050 177.900 ;
        RECT 919.950 177.450 922.050 177.900 ;
        RECT 910.950 176.250 922.050 177.450 ;
        RECT 910.950 175.800 913.050 176.250 ;
        RECT 919.950 175.800 922.050 176.250 ;
        RECT 949.950 177.600 952.050 177.900 ;
        RECT 967.950 177.600 970.050 177.900 ;
        RECT 949.950 176.400 970.050 177.600 ;
        RECT 949.950 175.800 952.050 176.400 ;
        RECT 967.950 175.800 970.050 176.400 ;
        RECT 757.950 174.600 760.050 175.050 ;
        RECT 740.400 173.400 760.050 174.600 ;
        RECT 757.950 172.950 760.050 173.400 ;
        RECT 829.950 174.600 832.050 175.050 ;
        RECT 842.400 174.600 843.600 175.800 ;
        RECT 829.950 173.400 843.600 174.600 ;
        RECT 901.950 174.600 904.050 175.050 ;
        RECT 934.950 174.600 937.050 175.050 ;
        RECT 946.950 174.600 949.050 175.050 ;
        RECT 901.950 173.400 949.050 174.600 ;
        RECT 829.950 172.950 832.050 173.400 ;
        RECT 901.950 172.950 904.050 173.400 ;
        RECT 934.950 172.950 937.050 173.400 ;
        RECT 946.950 172.950 949.050 173.400 ;
        RECT 976.950 174.600 979.050 175.050 ;
        RECT 982.950 174.600 985.050 175.050 ;
        RECT 991.950 174.600 994.050 175.050 ;
        RECT 976.950 173.400 994.050 174.600 ;
        RECT 976.950 172.950 979.050 173.400 ;
        RECT 982.950 172.950 985.050 173.400 ;
        RECT 991.950 172.950 994.050 173.400 ;
        RECT 655.950 171.600 658.050 171.900 ;
        RECT 622.950 170.400 658.050 171.600 ;
        RECT 622.950 169.950 625.050 170.400 ;
        RECT 655.950 169.800 658.050 170.400 ;
        RECT 712.950 169.800 715.050 171.900 ;
        RECT 823.950 171.600 826.050 172.050 ;
        RECT 847.950 171.600 850.050 172.050 ;
        RECT 862.950 171.600 865.050 172.050 ;
        RECT 823.950 170.400 865.050 171.600 ;
        RECT 823.950 169.950 826.050 170.400 ;
        RECT 847.950 169.950 850.050 170.400 ;
        RECT 862.950 169.950 865.050 170.400 ;
        RECT 109.950 168.600 112.050 169.050 ;
        RECT 151.950 168.600 154.050 169.050 ;
        RECT 217.950 168.600 220.050 169.050 ;
        RECT 589.950 168.600 592.050 169.050 ;
        RECT 109.950 167.400 220.050 168.600 ;
        RECT 109.950 166.950 112.050 167.400 ;
        RECT 151.950 166.950 154.050 167.400 ;
        RECT 217.950 166.950 220.050 167.400 ;
        RECT 335.400 167.400 592.050 168.600 ;
        RECT 211.950 165.600 214.050 166.050 ;
        RECT 247.950 165.600 250.050 166.050 ;
        RECT 262.950 165.600 265.050 166.050 ;
        RECT 211.950 164.400 265.050 165.600 ;
        RECT 211.950 163.950 214.050 164.400 ;
        RECT 247.950 163.950 250.050 164.400 ;
        RECT 262.950 163.950 265.050 164.400 ;
        RECT 274.950 165.600 277.050 166.050 ;
        RECT 335.400 165.600 336.600 167.400 ;
        RECT 589.950 166.950 592.050 167.400 ;
        RECT 595.950 168.600 598.050 169.050 ;
        RECT 733.950 168.600 736.050 169.050 ;
        RECT 595.950 167.400 736.050 168.600 ;
        RECT 595.950 166.950 598.050 167.400 ;
        RECT 733.950 166.950 736.050 167.400 ;
        RECT 790.950 168.600 793.050 169.050 ;
        RECT 808.950 168.600 811.050 169.050 ;
        RECT 838.950 168.600 841.050 169.050 ;
        RECT 790.950 167.400 841.050 168.600 ;
        RECT 790.950 166.950 793.050 167.400 ;
        RECT 808.950 166.950 811.050 167.400 ;
        RECT 838.950 166.950 841.050 167.400 ;
        RECT 958.950 168.600 961.050 169.050 ;
        RECT 982.950 168.600 985.050 169.050 ;
        RECT 958.950 167.400 985.050 168.600 ;
        RECT 958.950 166.950 961.050 167.400 ;
        RECT 982.950 166.950 985.050 167.400 ;
        RECT 274.950 164.400 336.600 165.600 ;
        RECT 541.950 165.600 544.050 166.050 ;
        RECT 571.950 165.600 574.050 166.050 ;
        RECT 541.950 164.400 574.050 165.600 ;
        RECT 274.950 163.950 277.050 164.400 ;
        RECT 541.950 163.950 544.050 164.400 ;
        RECT 571.950 163.950 574.050 164.400 ;
        RECT 601.950 165.600 604.050 166.050 ;
        RECT 649.950 165.600 652.050 166.050 ;
        RECT 601.950 164.400 652.050 165.600 ;
        RECT 601.950 163.950 604.050 164.400 ;
        RECT 649.950 163.950 652.050 164.400 ;
        RECT 688.950 165.600 691.050 166.050 ;
        RECT 727.950 165.600 730.050 166.050 ;
        RECT 688.950 164.400 730.050 165.600 ;
        RECT 688.950 163.950 691.050 164.400 ;
        RECT 727.950 163.950 730.050 164.400 ;
        RECT 745.950 165.600 748.050 166.050 ;
        RECT 754.950 165.600 757.050 166.050 ;
        RECT 799.950 165.600 802.050 166.050 ;
        RECT 745.950 164.400 802.050 165.600 ;
        RECT 745.950 163.950 748.050 164.400 ;
        RECT 754.950 163.950 757.050 164.400 ;
        RECT 799.950 163.950 802.050 164.400 ;
        RECT 859.950 165.600 862.050 166.050 ;
        RECT 892.950 165.600 895.050 166.050 ;
        RECT 859.950 164.400 895.050 165.600 ;
        RECT 859.950 163.950 862.050 164.400 ;
        RECT 892.950 163.950 895.050 164.400 ;
        RECT 28.950 162.600 31.050 163.050 ;
        RECT 73.950 162.600 76.050 163.050 ;
        RECT 28.950 161.400 76.050 162.600 ;
        RECT 28.950 160.950 31.050 161.400 ;
        RECT 73.950 160.950 76.050 161.400 ;
        RECT 382.950 162.600 385.050 163.050 ;
        RECT 544.950 162.600 547.050 163.050 ;
        RECT 598.950 162.600 601.050 163.050 ;
        RECT 661.950 162.600 664.050 163.050 ;
        RECT 382.950 161.400 664.050 162.600 ;
        RECT 382.950 160.950 385.050 161.400 ;
        RECT 544.950 160.950 547.050 161.400 ;
        RECT 598.950 160.950 601.050 161.400 ;
        RECT 661.950 160.950 664.050 161.400 ;
        RECT 802.950 162.600 805.050 163.050 ;
        RECT 907.950 162.600 910.050 163.050 ;
        RECT 802.950 161.400 910.050 162.600 ;
        RECT 802.950 160.950 805.050 161.400 ;
        RECT 907.950 160.950 910.050 161.400 ;
        RECT 943.950 162.600 946.050 163.050 ;
        RECT 973.950 162.600 976.050 163.050 ;
        RECT 943.950 161.400 976.050 162.600 ;
        RECT 943.950 160.950 946.050 161.400 ;
        RECT 973.950 160.950 976.050 161.400 ;
        RECT 454.950 159.600 457.050 160.050 ;
        RECT 484.950 159.600 487.050 160.050 ;
        RECT 508.950 159.600 511.050 160.050 ;
        RECT 454.950 158.400 511.050 159.600 ;
        RECT 454.950 157.950 457.050 158.400 ;
        RECT 484.950 157.950 487.050 158.400 ;
        RECT 508.950 157.950 511.050 158.400 ;
        RECT 550.950 159.600 553.050 160.050 ;
        RECT 559.950 159.600 562.050 160.050 ;
        RECT 643.950 159.600 646.050 160.050 ;
        RECT 550.950 158.400 646.050 159.600 ;
        RECT 550.950 157.950 553.050 158.400 ;
        RECT 559.950 157.950 562.050 158.400 ;
        RECT 643.950 157.950 646.050 158.400 ;
        RECT 652.950 159.600 655.050 160.050 ;
        RECT 721.950 159.600 724.050 160.050 ;
        RECT 652.950 158.400 724.050 159.600 ;
        RECT 652.950 157.950 655.050 158.400 ;
        RECT 721.950 157.950 724.050 158.400 ;
        RECT 763.950 159.600 766.050 160.050 ;
        RECT 790.950 159.600 793.050 160.050 ;
        RECT 763.950 158.400 793.050 159.600 ;
        RECT 763.950 157.950 766.050 158.400 ;
        RECT 790.950 157.950 793.050 158.400 ;
        RECT 796.950 159.600 799.050 160.050 ;
        RECT 910.950 159.600 913.050 160.050 ;
        RECT 796.950 158.400 913.050 159.600 ;
        RECT 796.950 157.950 799.050 158.400 ;
        RECT 910.950 157.950 913.050 158.400 ;
        RECT 19.950 156.600 22.050 157.050 ;
        RECT 25.950 156.600 28.050 157.050 ;
        RECT 67.950 156.600 70.050 157.050 ;
        RECT 19.950 155.400 70.050 156.600 ;
        RECT 19.950 154.950 22.050 155.400 ;
        RECT 25.950 154.950 28.050 155.400 ;
        RECT 67.950 154.950 70.050 155.400 ;
        RECT 655.950 156.600 658.050 157.050 ;
        RECT 655.950 155.400 768.600 156.600 ;
        RECT 655.950 154.950 658.050 155.400 ;
        RECT 337.950 153.600 340.050 154.050 ;
        RECT 382.950 153.600 385.050 154.050 ;
        RECT 337.950 152.400 385.050 153.600 ;
        RECT 337.950 151.950 340.050 152.400 ;
        RECT 382.950 151.950 385.050 152.400 ;
        RECT 433.950 153.600 436.050 154.050 ;
        RECT 505.950 153.600 508.050 154.050 ;
        RECT 511.950 153.600 514.050 154.050 ;
        RECT 433.950 152.400 514.050 153.600 ;
        RECT 433.950 151.950 436.050 152.400 ;
        RECT 505.950 151.950 508.050 152.400 ;
        RECT 511.950 151.950 514.050 152.400 ;
        RECT 571.950 153.600 574.050 154.050 ;
        RECT 589.950 153.600 592.050 154.050 ;
        RECT 571.950 152.400 592.050 153.600 ;
        RECT 571.950 151.950 574.050 152.400 ;
        RECT 589.950 151.950 592.050 152.400 ;
        RECT 616.950 153.600 619.050 154.050 ;
        RECT 670.950 153.600 673.050 154.050 ;
        RECT 616.950 152.400 673.050 153.600 ;
        RECT 616.950 151.950 619.050 152.400 ;
        RECT 670.950 151.950 673.050 152.400 ;
        RECT 694.950 153.600 697.050 154.050 ;
        RECT 763.950 153.600 766.050 154.050 ;
        RECT 694.950 152.400 766.050 153.600 ;
        RECT 767.400 153.600 768.600 155.400 ;
        RECT 796.950 153.600 799.050 154.050 ;
        RECT 859.950 153.600 862.050 154.050 ;
        RECT 767.400 152.400 799.050 153.600 ;
        RECT 694.950 151.950 697.050 152.400 ;
        RECT 763.950 151.950 766.050 152.400 ;
        RECT 796.950 151.950 799.050 152.400 ;
        RECT 830.400 152.400 862.050 153.600 ;
        RECT 49.950 150.600 52.050 151.050 ;
        RECT 85.950 150.600 88.050 151.050 ;
        RECT 49.950 149.400 88.050 150.600 ;
        RECT 49.950 148.950 52.050 149.400 ;
        RECT 85.950 148.950 88.050 149.400 ;
        RECT 130.950 150.600 133.050 151.050 ;
        RECT 172.950 150.600 175.050 151.050 ;
        RECT 130.950 149.400 175.050 150.600 ;
        RECT 130.950 148.950 133.050 149.400 ;
        RECT 172.950 148.950 175.050 149.400 ;
        RECT 499.950 150.600 502.050 151.050 ;
        RECT 562.950 150.600 565.050 151.050 ;
        RECT 595.950 150.600 598.050 151.050 ;
        RECT 499.950 149.400 598.050 150.600 ;
        RECT 499.950 148.950 502.050 149.400 ;
        RECT 562.950 148.950 565.050 149.400 ;
        RECT 595.950 148.950 598.050 149.400 ;
        RECT 757.950 150.600 760.050 151.050 ;
        RECT 830.400 150.600 831.600 152.400 ;
        RECT 859.950 151.950 862.050 152.400 ;
        RECT 955.950 153.600 958.050 154.050 ;
        RECT 970.950 153.600 973.050 154.050 ;
        RECT 955.950 152.400 973.050 153.600 ;
        RECT 955.950 151.950 958.050 152.400 ;
        RECT 970.950 151.950 973.050 152.400 ;
        RECT 757.950 149.400 831.600 150.600 ;
        RECT 886.950 150.600 889.050 151.050 ;
        RECT 895.950 150.600 898.050 151.050 ;
        RECT 886.950 149.400 898.050 150.600 ;
        RECT 757.950 148.950 760.050 149.400 ;
        RECT 886.950 148.950 889.050 149.400 ;
        RECT 895.950 148.950 898.050 149.400 ;
        RECT 19.950 147.600 22.050 148.050 ;
        RECT 46.950 147.600 49.050 148.050 ;
        RECT 19.950 146.400 49.050 147.600 ;
        RECT 19.950 145.950 22.050 146.400 ;
        RECT 46.950 145.950 49.050 146.400 ;
        RECT 193.950 147.600 196.050 148.050 ;
        RECT 226.950 147.600 229.050 148.050 ;
        RECT 193.950 146.400 229.050 147.600 ;
        RECT 193.950 145.950 196.050 146.400 ;
        RECT 226.950 145.950 229.050 146.400 ;
        RECT 565.950 147.600 568.050 148.050 ;
        RECT 649.950 147.600 652.050 148.050 ;
        RECT 841.950 147.600 844.050 148.050 ;
        RECT 565.950 146.400 652.050 147.600 ;
        RECT 565.950 145.950 568.050 146.400 ;
        RECT 649.950 145.950 652.050 146.400 ;
        RECT 695.400 146.400 844.050 147.600 ;
        RECT 695.400 145.050 696.600 146.400 ;
        RECT 841.950 145.950 844.050 146.400 ;
        RECT 898.950 147.600 901.050 148.050 ;
        RECT 904.950 147.600 907.050 148.050 ;
        RECT 928.950 147.600 931.050 148.050 ;
        RECT 898.950 146.400 931.050 147.600 ;
        RECT 898.950 145.950 901.050 146.400 ;
        RECT 904.950 145.950 907.050 146.400 ;
        RECT 928.950 145.950 931.050 146.400 ;
        RECT 49.950 144.600 52.050 145.050 ;
        RECT 61.950 144.600 64.050 145.050 ;
        RECT 49.950 143.400 64.050 144.600 ;
        RECT 49.950 142.950 52.050 143.400 ;
        RECT 61.950 142.950 64.050 143.400 ;
        RECT 94.950 144.600 97.050 145.050 ;
        RECT 136.950 144.600 139.050 145.050 ;
        RECT 145.950 144.600 148.050 145.050 ;
        RECT 94.950 143.400 148.050 144.600 ;
        RECT 94.950 142.950 97.050 143.400 ;
        RECT 136.950 142.950 139.050 143.400 ;
        RECT 145.950 142.950 148.050 143.400 ;
        RECT 253.950 144.600 256.050 145.050 ;
        RECT 295.950 144.600 298.050 145.050 ;
        RECT 253.950 143.400 298.050 144.600 ;
        RECT 253.950 142.950 256.050 143.400 ;
        RECT 295.950 142.950 298.050 143.400 ;
        RECT 421.950 144.600 424.050 145.050 ;
        RECT 469.950 144.600 472.050 145.050 ;
        RECT 421.950 143.400 472.050 144.600 ;
        RECT 421.950 142.950 424.050 143.400 ;
        RECT 469.950 142.950 472.050 143.400 ;
        RECT 490.950 144.600 493.050 145.050 ;
        RECT 496.950 144.600 499.050 145.050 ;
        RECT 490.950 143.400 499.050 144.600 ;
        RECT 490.950 142.950 493.050 143.400 ;
        RECT 496.950 142.950 499.050 143.400 ;
        RECT 547.950 144.600 550.050 145.050 ;
        RECT 559.950 144.600 562.050 145.050 ;
        RECT 547.950 143.400 562.050 144.600 ;
        RECT 547.950 142.950 550.050 143.400 ;
        RECT 559.950 142.950 562.050 143.400 ;
        RECT 574.950 144.600 577.050 145.050 ;
        RECT 580.950 144.600 583.050 145.050 ;
        RECT 574.950 143.400 583.050 144.600 ;
        RECT 574.950 142.950 577.050 143.400 ;
        RECT 580.950 142.950 583.050 143.400 ;
        RECT 670.950 144.600 673.050 145.050 ;
        RECT 694.950 144.600 697.050 145.050 ;
        RECT 670.950 143.400 697.050 144.600 ;
        RECT 670.950 142.950 673.050 143.400 ;
        RECT 694.950 142.950 697.050 143.400 ;
        RECT 868.950 144.600 871.050 145.050 ;
        RECT 949.950 144.600 952.050 145.050 ;
        RECT 868.950 143.400 952.050 144.600 ;
        RECT 868.950 142.950 871.050 143.400 ;
        RECT 949.950 142.950 952.050 143.400 ;
        RECT 223.950 141.600 226.050 142.050 ;
        RECT 250.950 141.600 253.050 142.050 ;
        RECT 394.950 141.600 397.050 142.050 ;
        RECT 223.950 140.400 253.050 141.600 ;
        RECT 223.950 139.950 226.050 140.400 ;
        RECT 250.950 139.950 253.050 140.400 ;
        RECT 368.400 140.400 397.050 141.600 ;
        RECT 34.950 138.600 37.050 139.050 ;
        RECT 40.950 138.600 43.050 139.200 ;
        RECT 34.950 137.400 43.050 138.600 ;
        RECT 34.950 136.950 37.050 137.400 ;
        RECT 40.950 137.100 43.050 137.400 ;
        RECT 46.950 138.600 49.050 139.050 ;
        RECT 52.950 138.600 55.050 139.050 ;
        RECT 61.950 138.600 64.050 139.200 ;
        RECT 46.950 137.400 64.050 138.600 ;
        RECT 46.950 136.950 49.050 137.400 ;
        RECT 52.950 136.950 55.050 137.400 ;
        RECT 61.950 137.100 64.050 137.400 ;
        RECT 91.950 138.600 94.050 139.200 ;
        RECT 109.950 138.600 112.050 139.200 ;
        RECT 91.950 137.400 112.050 138.600 ;
        RECT 91.950 137.100 94.050 137.400 ;
        RECT 109.950 137.100 112.050 137.400 ;
        RECT 142.950 138.750 145.050 139.200 ;
        RECT 151.950 138.750 154.050 139.200 ;
        RECT 142.950 137.550 154.050 138.750 ;
        RECT 142.950 137.100 145.050 137.550 ;
        RECT 151.950 137.100 154.050 137.550 ;
        RECT 163.950 138.750 166.050 139.200 ;
        RECT 178.950 138.750 181.050 139.200 ;
        RECT 163.950 137.550 181.050 138.750 ;
        RECT 163.950 137.100 166.050 137.550 ;
        RECT 178.950 137.100 181.050 137.550 ;
        RECT 187.950 138.750 190.050 139.200 ;
        RECT 199.950 138.750 202.050 139.200 ;
        RECT 187.950 138.600 202.050 138.750 ;
        RECT 220.950 138.600 223.050 139.050 ;
        RECT 187.950 137.550 223.050 138.600 ;
        RECT 187.950 137.100 190.050 137.550 ;
        RECT 199.950 137.400 223.050 137.550 ;
        RECT 199.950 137.100 202.050 137.400 ;
        RECT 220.950 136.950 223.050 137.400 ;
        RECT 262.950 138.750 265.050 139.200 ;
        RECT 268.950 138.750 271.050 139.050 ;
        RECT 271.950 138.750 274.050 139.200 ;
        RECT 262.950 137.550 274.050 138.750 ;
        RECT 262.950 137.100 265.050 137.550 ;
        RECT 268.950 136.950 271.050 137.550 ;
        RECT 271.950 137.100 274.050 137.550 ;
        RECT 307.950 138.750 310.050 139.200 ;
        RECT 313.950 138.750 316.050 139.200 ;
        RECT 307.950 137.550 316.050 138.750 ;
        RECT 307.950 137.100 310.050 137.550 ;
        RECT 313.950 137.100 316.050 137.550 ;
        RECT 319.950 138.600 322.050 139.200 ;
        RECT 337.950 138.600 340.050 139.200 ;
        RECT 319.950 137.400 340.050 138.600 ;
        RECT 319.950 137.100 322.050 137.400 ;
        RECT 337.950 137.100 340.050 137.400 ;
        RECT 346.950 138.750 349.050 139.200 ;
        RECT 358.950 138.750 361.050 139.200 ;
        RECT 346.950 138.600 361.050 138.750 ;
        RECT 368.400 138.600 369.600 140.400 ;
        RECT 394.950 139.950 397.050 140.400 ;
        RECT 346.950 137.550 369.600 138.600 ;
        RECT 346.950 137.100 349.050 137.550 ;
        RECT 358.950 137.400 369.600 137.550 ;
        RECT 370.950 138.600 373.050 139.050 ;
        RECT 388.950 138.600 391.050 139.200 ;
        RECT 370.950 137.400 391.050 138.600 ;
        RECT 358.950 137.100 361.050 137.400 ;
        RECT 370.950 136.950 373.050 137.400 ;
        RECT 388.950 137.100 391.050 137.400 ;
        RECT 412.950 137.100 415.050 139.200 ;
        RECT 418.950 138.600 421.050 139.200 ;
        RECT 427.950 138.750 430.050 139.200 ;
        RECT 436.950 138.750 439.050 139.200 ;
        RECT 427.950 138.600 439.050 138.750 ;
        RECT 418.950 137.550 439.050 138.600 ;
        RECT 418.950 137.400 430.050 137.550 ;
        RECT 418.950 137.100 421.050 137.400 ;
        RECT 427.950 137.100 430.050 137.400 ;
        RECT 436.950 137.100 439.050 137.550 ;
        RECT 442.950 137.100 445.050 139.200 ;
        RECT 463.950 138.750 466.050 139.200 ;
        RECT 475.800 138.750 477.900 139.200 ;
        RECT 463.950 137.550 477.900 138.750 ;
        RECT 463.950 137.100 466.050 137.550 ;
        RECT 475.800 137.100 477.900 137.550 ;
        RECT 478.950 138.750 481.050 139.200 ;
        RECT 490.950 138.750 493.050 139.200 ;
        RECT 478.950 137.550 493.050 138.750 ;
        RECT 478.950 137.100 481.050 137.550 ;
        RECT 490.950 137.100 493.050 137.550 ;
        RECT 505.950 138.750 508.050 139.200 ;
        RECT 514.950 138.750 517.050 139.200 ;
        RECT 505.950 137.550 517.050 138.750 ;
        RECT 505.950 137.100 508.050 137.550 ;
        RECT 514.950 137.100 517.050 137.550 ;
        RECT 631.950 138.750 634.050 139.200 ;
        RECT 646.800 138.750 648.900 139.200 ;
        RECT 631.950 137.550 648.900 138.750 ;
        RECT 631.950 137.100 634.050 137.550 ;
        RECT 646.800 137.100 648.900 137.550 ;
        RECT 649.950 138.600 652.050 139.050 ;
        RECT 670.950 138.600 673.050 139.200 ;
        RECT 688.950 138.600 691.050 139.200 ;
        RECT 649.950 137.400 691.050 138.600 ;
        RECT 136.950 135.600 139.050 136.050 ;
        RECT 128.400 134.400 139.050 135.600 ;
        RECT 413.400 135.600 414.600 137.100 ;
        RECT 413.400 134.400 432.600 135.600 ;
        RECT 128.400 132.900 129.600 134.400 ;
        RECT 136.950 133.950 139.050 134.400 ;
        RECT 43.950 132.450 46.050 132.900 ;
        RECT 49.950 132.450 52.050 132.900 ;
        RECT 43.950 131.250 52.050 132.450 ;
        RECT 43.950 130.800 46.050 131.250 ;
        RECT 49.950 130.800 52.050 131.250 ;
        RECT 127.950 130.800 130.050 132.900 ;
        RECT 154.950 132.450 157.050 132.900 ;
        RECT 163.950 132.450 166.050 132.900 ;
        RECT 154.950 131.250 166.050 132.450 ;
        RECT 154.950 130.800 157.050 131.250 ;
        RECT 163.950 130.800 166.050 131.250 ;
        RECT 175.950 132.600 178.050 132.900 ;
        RECT 196.950 132.600 199.050 132.900 ;
        RECT 175.950 131.400 199.050 132.600 ;
        RECT 175.950 130.800 178.050 131.400 ;
        RECT 196.950 130.800 199.050 131.400 ;
        RECT 202.950 132.600 205.050 132.900 ;
        RECT 214.950 132.600 217.050 133.050 ;
        RECT 202.950 131.400 217.050 132.600 ;
        RECT 202.950 130.800 205.050 131.400 ;
        RECT 214.950 130.950 217.050 131.400 ;
        RECT 238.950 132.600 241.050 133.050 ;
        RECT 244.950 132.600 247.050 132.900 ;
        RECT 238.950 131.400 247.050 132.600 ;
        RECT 238.950 130.950 241.050 131.400 ;
        RECT 244.950 130.800 247.050 131.400 ;
        RECT 280.950 132.600 283.050 132.900 ;
        RECT 298.950 132.600 301.050 132.900 ;
        RECT 280.950 131.400 301.050 132.600 ;
        RECT 280.950 130.800 283.050 131.400 ;
        RECT 298.950 130.800 301.050 131.400 ;
        RECT 316.950 132.600 319.050 132.900 ;
        RECT 328.950 132.600 331.050 133.050 ;
        RECT 316.950 131.400 331.050 132.600 ;
        RECT 316.950 130.800 319.050 131.400 ;
        RECT 328.950 130.950 331.050 131.400 ;
        RECT 397.950 132.600 400.050 133.050 ;
        RECT 403.950 132.600 406.050 133.050 ;
        RECT 431.400 132.900 432.600 134.400 ;
        RECT 397.950 131.400 406.050 132.600 ;
        RECT 397.950 130.950 400.050 131.400 ;
        RECT 403.950 130.950 406.050 131.400 ;
        RECT 430.950 132.450 433.050 132.900 ;
        RECT 439.950 132.450 442.050 132.900 ;
        RECT 430.950 131.250 442.050 132.450 ;
        RECT 430.950 130.800 433.050 131.250 ;
        RECT 439.950 130.800 442.050 131.250 ;
        RECT 22.950 129.600 25.050 130.050 ;
        RECT 64.950 129.600 67.050 130.050 ;
        RECT 118.950 129.600 121.050 130.050 ;
        RECT 22.950 128.400 121.050 129.600 ;
        RECT 22.950 127.950 25.050 128.400 ;
        RECT 64.950 127.950 67.050 128.400 ;
        RECT 118.950 127.950 121.050 128.400 ;
        RECT 160.950 129.600 163.050 130.050 ;
        RECT 169.950 129.600 172.050 130.050 ;
        RECT 160.950 128.400 172.050 129.600 ;
        RECT 160.950 127.950 163.050 128.400 ;
        RECT 169.950 127.950 172.050 128.400 ;
        RECT 196.950 129.600 199.050 130.050 ;
        RECT 223.950 129.600 226.050 130.050 ;
        RECT 196.950 128.400 226.050 129.600 ;
        RECT 196.950 127.950 199.050 128.400 ;
        RECT 223.950 127.950 226.050 128.400 ;
        RECT 229.950 129.600 232.050 130.050 ;
        RECT 250.950 129.600 253.050 130.050 ;
        RECT 262.950 129.600 265.050 130.050 ;
        RECT 229.950 128.400 265.050 129.600 ;
        RECT 229.950 127.950 232.050 128.400 ;
        RECT 250.950 127.950 253.050 128.400 ;
        RECT 262.950 127.950 265.050 128.400 ;
        RECT 415.950 129.600 418.050 130.050 ;
        RECT 443.400 129.600 444.600 137.100 ;
        RECT 649.950 136.950 652.050 137.400 ;
        RECT 670.950 137.100 673.050 137.400 ;
        RECT 688.950 137.100 691.050 137.400 ;
        RECT 706.950 138.750 709.050 139.200 ;
        RECT 718.950 138.750 721.050 139.200 ;
        RECT 706.950 137.550 721.050 138.750 ;
        RECT 706.950 137.100 709.050 137.550 ;
        RECT 718.950 137.100 721.050 137.550 ;
        RECT 727.950 138.600 730.050 139.050 ;
        RECT 739.950 138.600 742.050 139.200 ;
        RECT 727.950 137.400 742.050 138.600 ;
        RECT 727.950 136.950 730.050 137.400 ;
        RECT 739.950 137.100 742.050 137.400 ;
        RECT 751.950 138.600 754.050 139.050 ;
        RECT 757.950 138.600 760.050 139.200 ;
        RECT 751.950 137.400 760.050 138.600 ;
        RECT 751.950 136.950 754.050 137.400 ;
        RECT 757.950 137.100 760.050 137.400 ;
        RECT 817.950 138.600 820.050 139.050 ;
        RECT 823.950 138.750 826.050 139.200 ;
        RECT 853.950 138.750 856.050 139.200 ;
        RECT 823.950 138.600 856.050 138.750 ;
        RECT 817.950 137.550 856.050 138.600 ;
        RECT 817.950 137.400 826.050 137.550 ;
        RECT 817.950 136.950 820.050 137.400 ;
        RECT 823.950 137.100 826.050 137.400 ;
        RECT 853.950 137.100 856.050 137.550 ;
        RECT 880.950 138.750 883.050 139.200 ;
        RECT 889.950 138.750 892.050 139.200 ;
        RECT 880.950 138.600 892.050 138.750 ;
        RECT 904.950 138.600 907.050 139.200 ;
        RECT 880.950 137.550 907.050 138.600 ;
        RECT 880.950 137.100 883.050 137.550 ;
        RECT 889.950 137.400 907.050 137.550 ;
        RECT 889.950 137.100 892.050 137.400 ;
        RECT 904.950 137.100 907.050 137.400 ;
        RECT 919.950 138.750 922.050 139.200 ;
        RECT 934.950 138.750 937.050 139.200 ;
        RECT 919.950 137.550 937.050 138.750 ;
        RECT 919.950 137.100 922.050 137.550 ;
        RECT 934.950 137.100 937.050 137.550 ;
        RECT 946.950 138.750 949.050 139.200 ;
        RECT 967.950 138.750 970.050 139.200 ;
        RECT 946.950 138.600 970.050 138.750 ;
        RECT 1000.950 138.600 1003.050 139.200 ;
        RECT 946.950 137.550 1003.050 138.600 ;
        RECT 946.950 137.100 949.050 137.550 ;
        RECT 967.950 137.400 1003.050 137.550 ;
        RECT 967.950 137.100 970.050 137.400 ;
        RECT 1000.950 137.100 1003.050 137.400 ;
        RECT 475.950 132.600 478.050 133.050 ;
        RECT 487.950 132.600 490.050 132.900 ;
        RECT 475.950 131.400 490.050 132.600 ;
        RECT 475.950 130.950 478.050 131.400 ;
        RECT 487.950 130.800 490.050 131.400 ;
        RECT 568.950 132.600 571.050 132.900 ;
        RECT 592.950 132.600 595.050 132.900 ;
        RECT 568.950 131.400 595.050 132.600 ;
        RECT 568.950 130.800 571.050 131.400 ;
        RECT 592.950 130.800 595.050 131.400 ;
        RECT 691.950 132.600 694.050 132.900 ;
        RECT 706.950 132.600 709.050 133.050 ;
        RECT 691.950 131.400 709.050 132.600 ;
        RECT 691.950 130.800 694.050 131.400 ;
        RECT 706.950 130.950 709.050 131.400 ;
        RECT 715.950 132.450 718.050 132.900 ;
        RECT 727.950 132.450 730.050 132.900 ;
        RECT 715.950 131.250 730.050 132.450 ;
        RECT 715.950 130.800 718.050 131.250 ;
        RECT 727.950 130.800 730.050 131.250 ;
        RECT 733.950 132.450 736.050 132.900 ;
        RECT 742.950 132.450 745.050 132.900 ;
        RECT 733.950 131.250 745.050 132.450 ;
        RECT 733.950 130.800 736.050 131.250 ;
        RECT 742.950 130.800 745.050 131.250 ;
        RECT 751.950 132.450 754.050 132.900 ;
        RECT 784.950 132.450 787.050 132.900 ;
        RECT 751.950 131.250 787.050 132.450 ;
        RECT 751.950 130.800 754.050 131.250 ;
        RECT 784.950 130.800 787.050 131.250 ;
        RECT 811.950 132.600 814.050 132.900 ;
        RECT 823.950 132.600 826.050 133.050 ;
        RECT 811.950 131.400 826.050 132.600 ;
        RECT 811.950 130.800 814.050 131.400 ;
        RECT 823.950 130.950 826.050 131.400 ;
        RECT 835.950 132.450 838.050 132.900 ;
        RECT 841.950 132.450 844.050 132.900 ;
        RECT 835.950 131.250 844.050 132.450 ;
        RECT 835.950 130.800 838.050 131.250 ;
        RECT 841.950 130.800 844.050 131.250 ;
        RECT 856.950 132.600 859.050 132.900 ;
        RECT 868.950 132.600 871.050 133.050 ;
        RECT 856.950 131.400 871.050 132.600 ;
        RECT 856.950 130.800 859.050 131.400 ;
        RECT 868.950 130.950 871.050 131.400 ;
        RECT 883.950 132.600 886.050 132.900 ;
        RECT 895.950 132.600 898.050 132.900 ;
        RECT 883.950 132.450 898.050 132.600 ;
        RECT 907.950 132.450 910.050 132.900 ;
        RECT 883.950 131.400 910.050 132.450 ;
        RECT 883.950 130.800 886.050 131.400 ;
        RECT 895.950 131.250 910.050 131.400 ;
        RECT 895.950 130.800 898.050 131.250 ;
        RECT 907.950 130.800 910.050 131.250 ;
        RECT 913.950 132.600 916.050 132.900 ;
        RECT 931.950 132.600 934.050 132.900 ;
        RECT 913.950 131.400 934.050 132.600 ;
        RECT 913.950 130.800 916.050 131.400 ;
        RECT 931.950 130.800 934.050 131.400 ;
        RECT 952.950 132.600 955.050 132.900 ;
        RECT 985.950 132.600 988.050 132.900 ;
        RECT 952.950 131.400 988.050 132.600 ;
        RECT 952.950 130.800 955.050 131.400 ;
        RECT 985.950 130.800 988.050 131.400 ;
        RECT 415.950 128.400 444.600 129.600 ;
        RECT 466.950 129.600 469.050 130.050 ;
        RECT 514.950 129.600 517.050 130.050 ;
        RECT 466.950 128.400 517.050 129.600 ;
        RECT 415.950 127.950 418.050 128.400 ;
        RECT 466.950 127.950 469.050 128.400 ;
        RECT 514.950 127.950 517.050 128.400 ;
        RECT 529.950 129.600 532.050 130.050 ;
        RECT 568.950 129.600 571.050 130.050 ;
        RECT 529.950 128.400 571.050 129.600 ;
        RECT 529.950 127.950 532.050 128.400 ;
        RECT 568.950 127.950 571.050 128.400 ;
        RECT 859.950 129.600 862.050 130.050 ;
        RECT 871.950 129.600 874.050 130.050 ;
        RECT 859.950 128.400 874.050 129.600 ;
        RECT 859.950 127.950 862.050 128.400 ;
        RECT 871.950 127.950 874.050 128.400 ;
        RECT 34.950 126.600 37.050 127.050 ;
        RECT 52.950 126.600 55.050 127.050 ;
        RECT 34.950 125.400 55.050 126.600 ;
        RECT 34.950 124.950 37.050 125.400 ;
        RECT 52.950 124.950 55.050 125.400 ;
        RECT 445.950 126.600 448.050 127.050 ;
        RECT 460.950 126.600 463.050 127.050 ;
        RECT 445.950 125.400 463.050 126.600 ;
        RECT 445.950 124.950 448.050 125.400 ;
        RECT 460.950 124.950 463.050 125.400 ;
        RECT 511.950 126.600 514.050 127.050 ;
        RECT 523.950 126.600 526.050 127.050 ;
        RECT 511.950 125.400 526.050 126.600 ;
        RECT 511.950 124.950 514.050 125.400 ;
        RECT 523.950 124.950 526.050 125.400 ;
        RECT 592.950 126.600 595.050 127.050 ;
        RECT 628.950 126.600 631.050 126.900 ;
        RECT 592.950 125.400 631.050 126.600 ;
        RECT 592.950 124.950 595.050 125.400 ;
        RECT 628.950 124.800 631.050 125.400 ;
        RECT 709.950 126.600 712.050 127.050 ;
        RECT 838.950 126.600 841.050 127.050 ;
        RECT 919.950 126.600 922.050 127.050 ;
        RECT 709.950 125.400 922.050 126.600 ;
        RECT 709.950 124.950 712.050 125.400 ;
        RECT 838.950 124.950 841.050 125.400 ;
        RECT 919.950 124.950 922.050 125.400 ;
        RECT 946.950 126.600 949.050 127.050 ;
        RECT 979.950 126.600 982.050 127.050 ;
        RECT 946.950 125.400 982.050 126.600 ;
        RECT 946.950 124.950 949.050 125.400 ;
        RECT 979.950 124.950 982.050 125.400 ;
        RECT 43.950 123.600 46.050 124.050 ;
        RECT 82.950 123.600 85.050 124.050 ;
        RECT 43.950 122.400 85.050 123.600 ;
        RECT 43.950 121.950 46.050 122.400 ;
        RECT 82.950 121.950 85.050 122.400 ;
        RECT 106.950 123.600 109.050 124.050 ;
        RECT 127.950 123.600 130.050 124.050 ;
        RECT 148.950 123.600 151.050 124.050 ;
        RECT 106.950 122.400 151.050 123.600 ;
        RECT 106.950 121.950 109.050 122.400 ;
        RECT 127.950 121.950 130.050 122.400 ;
        RECT 148.950 121.950 151.050 122.400 ;
        RECT 562.950 123.600 565.050 124.050 ;
        RECT 595.800 123.600 597.900 124.050 ;
        RECT 562.950 122.400 597.900 123.600 ;
        RECT 562.950 121.950 565.050 122.400 ;
        RECT 595.800 121.950 597.900 122.400 ;
        RECT 598.950 123.600 601.050 124.050 ;
        RECT 622.950 123.600 625.050 124.050 ;
        RECT 637.950 123.600 640.050 124.050 ;
        RECT 598.950 122.400 640.050 123.600 ;
        RECT 598.950 121.950 601.050 122.400 ;
        RECT 622.950 121.950 625.050 122.400 ;
        RECT 637.950 121.950 640.050 122.400 ;
        RECT 742.950 123.600 745.050 124.050 ;
        RECT 826.950 123.600 829.050 124.050 ;
        RECT 850.950 123.600 853.050 124.050 ;
        RECT 742.950 122.400 853.050 123.600 ;
        RECT 742.950 121.950 745.050 122.400 ;
        RECT 826.950 121.950 829.050 122.400 ;
        RECT 850.950 121.950 853.050 122.400 ;
        RECT 340.950 120.600 343.050 121.050 ;
        RECT 379.950 120.600 382.050 121.050 ;
        RECT 340.950 119.400 382.050 120.600 ;
        RECT 340.950 118.950 343.050 119.400 ;
        RECT 379.950 118.950 382.050 119.400 ;
        RECT 388.950 120.600 391.050 121.050 ;
        RECT 544.950 120.600 547.050 121.050 ;
        RECT 730.950 120.600 733.050 121.050 ;
        RECT 736.950 120.600 739.050 121.050 ;
        RECT 388.950 119.400 739.050 120.600 ;
        RECT 388.950 118.950 391.050 119.400 ;
        RECT 544.950 118.950 547.050 119.400 ;
        RECT 730.950 118.950 733.050 119.400 ;
        RECT 736.950 118.950 739.050 119.400 ;
        RECT 88.950 117.600 91.050 118.050 ;
        RECT 97.950 117.600 100.050 118.050 ;
        RECT 88.950 116.400 100.050 117.600 ;
        RECT 88.950 115.950 91.050 116.400 ;
        RECT 97.950 115.950 100.050 116.400 ;
        RECT 232.950 117.600 235.050 118.050 ;
        RECT 286.950 117.600 289.050 118.050 ;
        RECT 232.950 116.400 289.050 117.600 ;
        RECT 232.950 115.950 235.050 116.400 ;
        RECT 286.950 115.950 289.050 116.400 ;
        RECT 298.950 117.600 301.050 118.050 ;
        RECT 361.950 117.600 364.050 118.050 ;
        RECT 382.950 117.600 385.050 118.050 ;
        RECT 298.950 116.400 385.050 117.600 ;
        RECT 298.950 115.950 301.050 116.400 ;
        RECT 361.950 115.950 364.050 116.400 ;
        RECT 382.950 115.950 385.050 116.400 ;
        RECT 406.950 117.600 409.050 118.050 ;
        RECT 469.950 117.600 472.050 118.050 ;
        RECT 406.950 116.400 472.050 117.600 ;
        RECT 406.950 115.950 409.050 116.400 ;
        RECT 469.950 115.950 472.050 116.400 ;
        RECT 559.950 117.600 562.050 118.050 ;
        RECT 565.950 117.600 568.050 118.050 ;
        RECT 559.950 116.400 568.050 117.600 ;
        RECT 559.950 115.950 562.050 116.400 ;
        RECT 565.950 115.950 568.050 116.400 ;
        RECT 571.950 117.600 574.050 118.050 ;
        RECT 580.950 117.600 583.050 118.050 ;
        RECT 571.950 116.400 583.050 117.600 ;
        RECT 571.950 115.950 574.050 116.400 ;
        RECT 580.950 115.950 583.050 116.400 ;
        RECT 595.950 117.600 598.050 118.050 ;
        RECT 622.950 117.600 625.050 118.050 ;
        RECT 634.950 117.600 637.050 118.050 ;
        RECT 595.950 116.400 637.050 117.600 ;
        RECT 595.950 115.950 598.050 116.400 ;
        RECT 622.950 115.950 625.050 116.400 ;
        RECT 634.950 115.950 637.050 116.400 ;
        RECT 799.950 117.600 802.050 118.050 ;
        RECT 829.950 117.600 832.050 118.050 ;
        RECT 799.950 116.400 832.050 117.600 ;
        RECT 799.950 115.950 802.050 116.400 ;
        RECT 829.950 115.950 832.050 116.400 ;
        RECT 853.950 117.600 856.050 118.050 ;
        RECT 868.950 117.600 871.050 118.050 ;
        RECT 877.950 117.600 880.050 118.050 ;
        RECT 853.950 116.400 880.050 117.600 ;
        RECT 853.950 115.950 856.050 116.400 ;
        RECT 868.950 115.950 871.050 116.400 ;
        RECT 877.950 115.950 880.050 116.400 ;
        RECT 79.950 114.600 82.050 115.050 ;
        RECT 88.950 114.600 91.050 114.900 ;
        RECT 109.950 114.600 112.050 115.050 ;
        RECT 79.950 113.400 112.050 114.600 ;
        RECT 79.950 112.950 82.050 113.400 ;
        RECT 88.950 112.800 91.050 113.400 ;
        RECT 109.950 112.950 112.050 113.400 ;
        RECT 139.950 114.600 142.050 115.050 ;
        RECT 556.950 114.600 559.050 115.050 ;
        RECT 139.950 113.400 559.050 114.600 ;
        RECT 139.950 112.950 142.050 113.400 ;
        RECT 556.950 112.950 559.050 113.400 ;
        RECT 616.950 114.600 619.050 115.050 ;
        RECT 640.950 114.600 643.050 115.050 ;
        RECT 616.950 113.400 643.050 114.600 ;
        RECT 616.950 112.950 619.050 113.400 ;
        RECT 640.950 112.950 643.050 113.400 ;
        RECT 655.950 114.600 658.050 115.050 ;
        RECT 685.950 114.600 688.050 115.050 ;
        RECT 775.950 114.600 778.050 115.050 ;
        RECT 655.950 113.400 778.050 114.600 ;
        RECT 655.950 112.950 658.050 113.400 ;
        RECT 685.950 112.950 688.050 113.400 ;
        RECT 775.950 112.950 778.050 113.400 ;
        RECT 892.950 114.600 895.050 115.050 ;
        RECT 931.950 114.600 934.050 115.050 ;
        RECT 892.950 113.400 934.050 114.600 ;
        RECT 892.950 112.950 895.050 113.400 ;
        RECT 931.950 112.950 934.050 113.400 ;
        RECT 991.950 114.600 994.050 115.050 ;
        RECT 1000.950 114.600 1003.050 115.050 ;
        RECT 1015.950 114.600 1018.050 115.050 ;
        RECT 991.950 113.400 1018.050 114.600 ;
        RECT 991.950 112.950 994.050 113.400 ;
        RECT 1000.950 112.950 1003.050 113.400 ;
        RECT 1015.950 112.950 1018.050 113.400 ;
        RECT 73.950 111.600 76.050 112.050 ;
        RECT 133.950 111.600 136.050 112.050 ;
        RECT 73.950 110.400 136.050 111.600 ;
        RECT 73.950 109.950 76.050 110.400 ;
        RECT 133.950 109.950 136.050 110.400 ;
        RECT 259.950 111.600 262.050 112.050 ;
        RECT 292.950 111.600 295.050 112.050 ;
        RECT 259.950 110.400 295.050 111.600 ;
        RECT 259.950 109.950 262.050 110.400 ;
        RECT 292.950 109.950 295.050 110.400 ;
        RECT 340.950 111.600 343.050 112.050 ;
        RECT 346.950 111.600 349.050 112.050 ;
        RECT 340.950 110.400 349.050 111.600 ;
        RECT 340.950 109.950 343.050 110.400 ;
        RECT 346.950 109.950 349.050 110.400 ;
        RECT 361.950 111.600 364.050 112.050 ;
        RECT 370.950 111.600 373.050 112.050 ;
        RECT 361.950 110.400 373.050 111.600 ;
        RECT 361.950 109.950 364.050 110.400 ;
        RECT 370.950 109.950 373.050 110.400 ;
        RECT 379.950 111.600 382.050 112.050 ;
        RECT 415.950 111.600 418.050 112.050 ;
        RECT 379.950 110.400 418.050 111.600 ;
        RECT 379.950 109.950 382.050 110.400 ;
        RECT 415.950 109.950 418.050 110.400 ;
        RECT 421.950 111.600 424.050 112.050 ;
        RECT 460.950 111.600 463.050 112.050 ;
        RECT 478.950 111.600 481.050 112.050 ;
        RECT 526.950 111.600 529.050 112.050 ;
        RECT 421.950 110.400 529.050 111.600 ;
        RECT 421.950 109.950 424.050 110.400 ;
        RECT 460.950 109.950 463.050 110.400 ;
        RECT 478.950 109.950 481.050 110.400 ;
        RECT 526.950 109.950 529.050 110.400 ;
        RECT 580.950 111.600 583.050 112.050 ;
        RECT 604.950 111.600 607.050 112.050 ;
        RECT 580.950 110.400 607.050 111.600 ;
        RECT 580.950 109.950 583.050 110.400 ;
        RECT 604.950 109.950 607.050 110.400 ;
        RECT 673.950 111.600 676.050 112.050 ;
        RECT 766.950 111.600 769.050 112.050 ;
        RECT 673.950 110.400 769.050 111.600 ;
        RECT 673.950 109.950 676.050 110.400 ;
        RECT 766.950 109.950 769.050 110.400 ;
        RECT 874.950 111.600 877.050 112.050 ;
        RECT 889.950 111.600 892.050 112.050 ;
        RECT 979.950 111.600 982.050 112.050 ;
        RECT 988.950 111.600 991.050 112.050 ;
        RECT 874.950 110.400 991.050 111.600 ;
        RECT 874.950 109.950 877.050 110.400 ;
        RECT 889.950 109.950 892.050 110.400 ;
        RECT 979.950 109.950 982.050 110.400 ;
        RECT 988.950 109.950 991.050 110.400 ;
        RECT 28.950 108.600 31.050 109.050 ;
        RECT 37.950 108.600 40.050 109.050 ;
        RECT 28.950 107.400 40.050 108.600 ;
        RECT 28.950 106.950 31.050 107.400 ;
        RECT 37.950 106.950 40.050 107.400 ;
        RECT 184.950 108.600 187.050 109.050 ;
        RECT 202.950 108.600 205.050 109.050 ;
        RECT 213.000 108.600 217.050 109.050 ;
        RECT 223.950 108.600 226.050 109.050 ;
        RECT 184.950 107.400 205.050 108.600 ;
        RECT 212.400 107.400 226.050 108.600 ;
        RECT 184.950 106.950 187.050 107.400 ;
        RECT 202.950 106.950 205.050 107.400 ;
        RECT 213.000 106.950 217.050 107.400 ;
        RECT 223.950 106.950 226.050 107.400 ;
        RECT 376.950 108.600 379.050 109.050 ;
        RECT 403.950 108.600 406.050 109.050 ;
        RECT 376.950 107.400 406.050 108.600 ;
        RECT 376.950 106.950 379.050 107.400 ;
        RECT 403.950 106.950 406.050 107.400 ;
        RECT 556.950 108.600 559.050 109.050 ;
        RECT 568.950 108.600 571.050 109.050 ;
        RECT 607.950 108.600 610.050 109.050 ;
        RECT 556.950 107.400 610.050 108.600 ;
        RECT 556.950 106.950 559.050 107.400 ;
        RECT 568.950 106.950 571.050 107.400 ;
        RECT 607.950 106.950 610.050 107.400 ;
        RECT 745.950 108.600 748.050 109.050 ;
        RECT 754.950 108.600 757.050 109.050 ;
        RECT 745.950 107.400 757.050 108.600 ;
        RECT 745.950 106.950 748.050 107.400 ;
        RECT 754.950 106.950 757.050 107.400 ;
        RECT 16.950 105.600 19.050 106.200 ;
        RECT 25.950 105.600 28.050 106.050 ;
        RECT 16.950 104.400 28.050 105.600 ;
        RECT 16.950 104.100 19.050 104.400 ;
        RECT 25.950 103.950 28.050 104.400 ;
        RECT 37.950 105.600 40.050 106.200 ;
        RECT 61.950 105.600 64.050 106.200 ;
        RECT 37.950 104.400 64.050 105.600 ;
        RECT 37.950 104.100 40.050 104.400 ;
        RECT 61.950 104.100 64.050 104.400 ;
        RECT 67.950 105.600 70.050 106.200 ;
        RECT 79.800 105.600 81.900 106.050 ;
        RECT 67.950 104.400 81.900 105.600 ;
        RECT 67.950 104.100 70.050 104.400 ;
        RECT 79.800 103.950 81.900 104.400 ;
        RECT 82.950 105.600 85.050 106.200 ;
        RECT 115.950 105.600 118.050 106.200 ;
        RECT 121.950 105.600 124.050 106.050 ;
        RECT 82.950 104.400 93.600 105.600 ;
        RECT 82.950 104.100 85.050 104.400 ;
        RECT 92.400 100.050 93.600 104.400 ;
        RECT 115.950 104.400 124.050 105.600 ;
        RECT 115.950 104.100 118.050 104.400 ;
        RECT 121.950 103.950 124.050 104.400 ;
        RECT 154.950 105.750 157.050 106.200 ;
        RECT 160.950 105.750 163.050 106.200 ;
        RECT 154.950 104.550 163.050 105.750 ;
        RECT 154.950 104.100 157.050 104.550 ;
        RECT 160.950 104.100 163.050 104.550 ;
        RECT 169.950 105.750 172.050 106.200 ;
        RECT 178.950 105.750 181.050 106.200 ;
        RECT 169.950 104.550 181.050 105.750 ;
        RECT 169.950 104.100 172.050 104.550 ;
        RECT 178.950 104.100 181.050 104.550 ;
        RECT 199.950 105.750 202.050 106.200 ;
        RECT 208.950 105.750 211.050 106.200 ;
        RECT 199.950 104.550 211.050 105.750 ;
        RECT 199.950 104.100 202.050 104.550 ;
        RECT 208.950 104.100 211.050 104.550 ;
        RECT 247.950 105.750 250.050 106.200 ;
        RECT 256.950 105.750 259.050 106.200 ;
        RECT 247.950 104.550 259.050 105.750 ;
        RECT 247.950 104.100 250.050 104.550 ;
        RECT 256.950 104.100 259.050 104.550 ;
        RECT 274.950 105.750 277.050 106.200 ;
        RECT 280.950 105.750 283.050 106.200 ;
        RECT 274.950 104.550 283.050 105.750 ;
        RECT 274.950 104.100 277.050 104.550 ;
        RECT 280.950 104.100 283.050 104.550 ;
        RECT 295.950 105.750 298.050 106.200 ;
        RECT 301.950 105.750 304.050 106.200 ;
        RECT 295.950 105.600 304.050 105.750 ;
        RECT 328.950 105.600 331.050 106.200 ;
        RECT 295.950 104.550 372.600 105.600 ;
        RECT 295.950 104.100 298.050 104.550 ;
        RECT 301.950 104.400 372.600 104.550 ;
        RECT 301.950 104.100 304.050 104.400 ;
        RECT 328.950 104.100 331.050 104.400 ;
        RECT 127.950 102.600 130.050 103.050 ;
        RECT 113.400 101.400 130.050 102.600 ;
        RECT 371.400 102.600 372.600 104.400 ;
        RECT 421.950 104.100 424.050 106.200 ;
        RECT 487.950 105.750 490.050 106.200 ;
        RECT 493.950 105.750 496.050 106.200 ;
        RECT 487.950 104.550 496.050 105.750 ;
        RECT 487.950 104.100 490.050 104.550 ;
        RECT 493.950 104.100 496.050 104.550 ;
        RECT 505.950 105.750 508.050 106.200 ;
        RECT 511.950 105.750 514.050 106.200 ;
        RECT 505.950 104.550 514.050 105.750 ;
        RECT 505.950 104.100 508.050 104.550 ;
        RECT 511.950 104.100 514.050 104.550 ;
        RECT 517.950 105.750 520.050 106.200 ;
        RECT 523.950 105.750 526.050 106.200 ;
        RECT 517.950 105.600 526.050 105.750 ;
        RECT 532.950 105.600 535.050 106.200 ;
        RECT 517.950 104.550 535.050 105.600 ;
        RECT 517.950 104.100 520.050 104.550 ;
        RECT 523.950 104.400 535.050 104.550 ;
        RECT 523.950 104.100 526.050 104.400 ;
        RECT 532.950 104.100 535.050 104.400 ;
        RECT 538.950 105.600 541.050 106.200 ;
        RECT 550.950 105.600 553.050 106.050 ;
        RECT 538.950 104.400 553.050 105.600 ;
        RECT 538.950 104.100 541.050 104.400 ;
        RECT 415.950 102.600 418.050 103.050 ;
        RECT 422.400 102.600 423.600 104.100 ;
        RECT 550.950 103.950 553.050 104.400 ;
        RECT 562.950 103.950 565.050 106.050 ;
        RECT 586.950 105.600 589.050 106.200 ;
        RECT 595.950 105.600 598.050 106.050 ;
        RECT 586.950 104.400 598.050 105.600 ;
        RECT 586.950 104.100 589.050 104.400 ;
        RECT 595.950 103.950 598.050 104.400 ;
        RECT 604.950 105.600 607.050 106.200 ;
        RECT 604.950 104.400 618.600 105.600 ;
        RECT 604.950 104.100 607.050 104.400 ;
        RECT 371.400 101.400 423.600 102.600 ;
        RECT 481.950 102.600 484.050 103.050 ;
        RECT 502.950 102.600 505.050 103.050 ;
        RECT 481.950 101.400 505.050 102.600 ;
        RECT 19.950 99.600 22.050 99.900 ;
        RECT 34.950 99.600 37.050 99.900 ;
        RECT 19.950 98.400 37.050 99.600 ;
        RECT 19.950 97.800 22.050 98.400 ;
        RECT 34.950 97.800 37.050 98.400 ;
        RECT 52.950 99.450 55.050 99.900 ;
        RECT 58.950 99.450 61.050 99.900 ;
        RECT 52.950 98.250 61.050 99.450 ;
        RECT 92.400 98.400 97.050 100.050 ;
        RECT 113.400 99.900 114.600 101.400 ;
        RECT 127.950 100.950 130.050 101.400 ;
        RECT 415.950 100.950 418.050 101.400 ;
        RECT 481.950 100.950 484.050 101.400 ;
        RECT 502.950 100.950 505.050 101.400 ;
        RECT 52.950 97.800 55.050 98.250 ;
        RECT 58.950 97.800 61.050 98.250 ;
        RECT 93.000 97.950 97.050 98.400 ;
        RECT 112.950 97.800 115.050 99.900 ;
        RECT 124.950 99.450 127.050 99.900 ;
        RECT 142.950 99.450 145.050 99.900 ;
        RECT 124.950 98.250 145.050 99.450 ;
        RECT 124.950 97.800 127.050 98.250 ;
        RECT 142.950 97.800 145.050 98.250 ;
        RECT 163.950 99.600 166.050 99.900 ;
        RECT 181.950 99.600 184.050 99.900 ;
        RECT 163.950 98.400 184.050 99.600 ;
        RECT 163.950 97.800 166.050 98.400 ;
        RECT 181.950 97.800 184.050 98.400 ;
        RECT 187.950 99.600 190.050 99.900 ;
        RECT 205.950 99.600 208.050 99.900 ;
        RECT 187.950 98.400 208.050 99.600 ;
        RECT 187.950 97.800 190.050 98.400 ;
        RECT 205.950 97.800 208.050 98.400 ;
        RECT 223.950 99.450 226.050 99.900 ;
        RECT 235.950 99.600 238.050 99.900 ;
        RECT 253.950 99.600 256.050 99.900 ;
        RECT 235.950 99.450 256.050 99.600 ;
        RECT 223.950 98.400 256.050 99.450 ;
        RECT 223.950 98.250 238.050 98.400 ;
        RECT 223.950 97.800 226.050 98.250 ;
        RECT 235.950 97.800 238.050 98.250 ;
        RECT 253.950 97.800 256.050 98.400 ;
        RECT 259.950 99.600 262.050 99.900 ;
        RECT 295.950 99.600 298.050 100.050 ;
        RECT 304.950 99.600 307.050 99.900 ;
        RECT 316.950 99.600 319.050 100.050 ;
        RECT 259.950 98.400 298.050 99.600 ;
        RECT 259.950 97.800 262.050 98.400 ;
        RECT 295.950 97.950 298.050 98.400 ;
        RECT 302.400 98.400 319.050 99.600 ;
        RECT 100.950 96.600 103.050 97.050 ;
        RECT 136.950 96.600 139.050 97.050 ;
        RECT 100.950 95.400 139.050 96.600 ;
        RECT 100.950 94.950 103.050 95.400 ;
        RECT 136.950 94.950 139.050 95.400 ;
        RECT 283.950 96.600 286.050 97.050 ;
        RECT 302.400 96.600 303.600 98.400 ;
        RECT 304.950 97.800 307.050 98.400 ;
        RECT 316.950 97.950 319.050 98.400 ;
        RECT 424.950 99.600 427.050 99.900 ;
        RECT 439.950 99.600 442.050 99.900 ;
        RECT 424.950 98.400 442.050 99.600 ;
        RECT 424.950 97.800 427.050 98.400 ;
        RECT 439.950 97.800 442.050 98.400 ;
        RECT 496.950 99.600 499.050 99.900 ;
        RECT 505.950 99.600 508.050 100.050 ;
        RECT 496.950 98.400 508.050 99.600 ;
        RECT 496.950 97.800 499.050 98.400 ;
        RECT 505.950 97.950 508.050 98.400 ;
        RECT 526.950 99.450 529.050 99.900 ;
        RECT 535.950 99.450 538.050 99.900 ;
        RECT 526.950 98.250 538.050 99.450 ;
        RECT 526.950 97.800 529.050 98.250 ;
        RECT 535.950 97.800 538.050 98.250 ;
        RECT 559.950 99.600 562.050 99.900 ;
        RECT 563.400 99.600 564.600 103.950 ;
        RECT 617.400 102.600 618.600 104.400 ;
        RECT 622.950 102.600 625.050 106.050 ;
        RECT 634.950 105.600 637.050 106.200 ;
        RECT 643.950 105.600 646.050 105.900 ;
        RECT 634.950 104.400 646.050 105.600 ;
        RECT 634.950 104.100 637.050 104.400 ;
        RECT 643.950 103.800 646.050 104.400 ;
        RECT 661.950 105.600 664.050 106.200 ;
        RECT 667.800 105.600 669.900 106.050 ;
        RECT 661.950 104.400 669.900 105.600 ;
        RECT 661.950 104.100 664.050 104.400 ;
        RECT 667.800 103.950 669.900 104.400 ;
        RECT 670.950 105.600 673.050 106.050 ;
        RECT 679.950 105.600 682.050 106.200 ;
        RECT 670.950 104.400 682.050 105.600 ;
        RECT 670.950 103.950 673.050 104.400 ;
        RECT 679.950 104.100 682.050 104.400 ;
        RECT 703.950 105.750 706.050 106.200 ;
        RECT 718.950 105.750 721.050 106.200 ;
        RECT 703.950 104.550 721.050 105.750 ;
        RECT 703.950 104.100 706.050 104.550 ;
        RECT 718.950 104.100 721.050 104.550 ;
        RECT 730.950 104.100 733.050 106.200 ;
        RECT 781.950 105.600 784.050 106.200 ;
        RECT 787.950 105.600 790.050 106.050 ;
        RECT 781.950 104.400 790.050 105.600 ;
        RECT 781.950 104.100 784.050 104.400 ;
        RECT 731.400 102.600 732.600 104.100 ;
        RECT 787.950 103.950 790.050 104.400 ;
        RECT 793.950 105.600 796.050 106.050 ;
        RECT 802.950 105.750 805.050 106.200 ;
        RECT 811.950 105.750 814.050 106.200 ;
        RECT 802.950 105.600 814.050 105.750 ;
        RECT 793.950 104.550 814.050 105.600 ;
        RECT 793.950 104.400 805.050 104.550 ;
        RECT 793.950 103.950 796.050 104.400 ;
        RECT 802.950 104.100 805.050 104.400 ;
        RECT 811.950 104.100 814.050 104.550 ;
        RECT 823.950 104.100 826.050 106.200 ;
        RECT 847.950 105.600 850.050 106.200 ;
        RECT 886.950 105.600 889.050 106.050 ;
        RECT 847.950 104.400 889.050 105.600 ;
        RECT 847.950 104.100 850.050 104.400 ;
        RECT 617.400 101.400 621.600 102.600 ;
        RECT 622.950 102.000 633.600 102.600 ;
        RECT 725.400 102.000 732.600 102.600 ;
        RECT 623.400 101.400 633.600 102.000 ;
        RECT 559.950 98.400 564.600 99.600 ;
        RECT 568.950 99.450 571.050 99.900 ;
        RECT 583.950 99.600 586.050 99.900 ;
        RECT 601.950 99.600 604.050 99.900 ;
        RECT 583.950 99.450 604.050 99.600 ;
        RECT 568.950 98.400 604.050 99.450 ;
        RECT 620.400 99.600 621.600 101.400 ;
        RECT 632.400 99.900 633.600 101.400 ;
        RECT 724.950 101.400 732.600 102.000 ;
        RECT 625.950 99.600 628.050 99.900 ;
        RECT 620.400 98.400 628.050 99.600 ;
        RECT 559.950 97.800 562.050 98.400 ;
        RECT 568.950 98.250 586.050 98.400 ;
        RECT 568.950 97.800 571.050 98.250 ;
        RECT 583.950 97.800 586.050 98.250 ;
        RECT 601.950 97.800 604.050 98.400 ;
        RECT 625.950 97.800 628.050 98.400 ;
        RECT 631.950 97.800 634.050 99.900 ;
        RECT 658.950 99.600 661.050 99.900 ;
        RECT 673.950 99.600 676.050 99.900 ;
        RECT 658.950 99.450 676.050 99.600 ;
        RECT 682.950 99.450 685.050 99.900 ;
        RECT 658.950 98.400 685.050 99.450 ;
        RECT 658.950 97.800 661.050 98.400 ;
        RECT 673.950 98.250 685.050 98.400 ;
        RECT 673.950 97.800 676.050 98.250 ;
        RECT 682.950 97.800 685.050 98.250 ;
        RECT 700.950 99.450 703.050 99.900 ;
        RECT 706.950 99.450 709.050 99.900 ;
        RECT 700.950 98.250 709.050 99.450 ;
        RECT 700.950 97.800 703.050 98.250 ;
        RECT 706.950 97.800 709.050 98.250 ;
        RECT 724.950 97.950 727.050 101.400 ;
        RECT 733.950 99.450 736.050 99.900 ;
        RECT 742.950 99.450 745.050 99.900 ;
        RECT 733.950 98.250 745.050 99.450 ;
        RECT 733.950 97.800 736.050 98.250 ;
        RECT 742.950 97.800 745.050 98.250 ;
        RECT 766.950 99.450 769.050 99.900 ;
        RECT 772.950 99.450 775.050 99.900 ;
        RECT 766.950 98.250 775.050 99.450 ;
        RECT 766.950 97.800 769.050 98.250 ;
        RECT 772.950 97.800 775.050 98.250 ;
        RECT 784.950 99.450 787.050 99.900 ;
        RECT 799.950 99.600 802.050 99.900 ;
        RECT 824.400 99.600 825.600 104.100 ;
        RECT 886.950 103.950 889.050 104.400 ;
        RECT 898.950 105.600 901.050 106.200 ;
        RECT 907.950 105.600 910.050 106.050 ;
        RECT 898.950 104.400 910.050 105.600 ;
        RECT 898.950 104.100 901.050 104.400 ;
        RECT 907.950 103.950 910.050 104.400 ;
        RECT 925.950 105.600 928.050 106.200 ;
        RECT 955.950 105.600 958.050 106.050 ;
        RECT 964.950 105.600 967.050 106.200 ;
        RECT 970.950 105.600 973.050 106.050 ;
        RECT 925.950 104.400 973.050 105.600 ;
        RECT 925.950 104.100 928.050 104.400 ;
        RECT 955.950 103.950 958.050 104.400 ;
        RECT 964.950 104.100 967.050 104.400 ;
        RECT 970.950 103.950 973.050 104.400 ;
        RECT 799.950 99.450 825.600 99.600 ;
        RECT 784.950 98.400 825.600 99.450 ;
        RECT 838.950 99.450 841.050 99.900 ;
        RECT 844.950 99.450 847.050 99.900 ;
        RECT 784.950 98.250 802.050 98.400 ;
        RECT 784.950 97.800 787.050 98.250 ;
        RECT 799.950 97.800 802.050 98.250 ;
        RECT 838.950 98.250 847.050 99.450 ;
        RECT 838.950 97.800 841.050 98.250 ;
        RECT 844.950 97.800 847.050 98.250 ;
        RECT 850.950 99.600 853.050 99.900 ;
        RECT 862.950 99.600 865.050 99.900 ;
        RECT 850.950 99.450 865.050 99.600 ;
        RECT 871.950 99.450 874.050 99.900 ;
        RECT 850.950 98.400 874.050 99.450 ;
        RECT 850.950 97.800 853.050 98.400 ;
        RECT 862.950 98.250 874.050 98.400 ;
        RECT 862.950 97.800 865.050 98.250 ;
        RECT 871.950 97.800 874.050 98.250 ;
        RECT 901.950 99.600 904.050 99.900 ;
        RECT 910.950 99.600 913.050 99.900 ;
        RECT 901.950 99.450 913.050 99.600 ;
        RECT 916.950 99.450 919.050 99.900 ;
        RECT 901.950 98.400 919.050 99.450 ;
        RECT 901.950 97.800 904.050 98.400 ;
        RECT 910.950 98.250 919.050 98.400 ;
        RECT 910.950 97.800 913.050 98.250 ;
        RECT 916.950 97.800 919.050 98.250 ;
        RECT 949.950 99.450 952.050 99.900 ;
        RECT 955.950 99.450 958.050 99.900 ;
        RECT 949.950 98.250 958.050 99.450 ;
        RECT 949.950 97.800 952.050 98.250 ;
        RECT 955.950 97.800 958.050 98.250 ;
        RECT 970.950 99.450 973.050 99.900 ;
        RECT 988.950 99.450 991.050 99.900 ;
        RECT 970.950 98.250 991.050 99.450 ;
        RECT 970.950 97.800 973.050 98.250 ;
        RECT 988.950 97.800 991.050 98.250 ;
        RECT 283.950 95.400 303.600 96.600 ;
        RECT 304.950 96.600 307.050 96.750 ;
        RECT 310.950 96.600 313.050 97.050 ;
        RECT 334.950 96.600 337.050 97.050 ;
        RECT 304.950 95.400 337.050 96.600 ;
        RECT 283.950 94.950 286.050 95.400 ;
        RECT 304.950 94.650 307.050 95.400 ;
        RECT 310.950 94.950 313.050 95.400 ;
        RECT 334.950 94.950 337.050 95.400 ;
        RECT 502.950 96.600 505.050 97.050 ;
        RECT 514.950 96.600 517.050 97.050 ;
        RECT 502.950 95.400 517.050 96.600 ;
        RECT 502.950 94.950 505.050 95.400 ;
        RECT 514.950 94.950 517.050 95.400 ;
        RECT 652.950 96.600 655.050 97.050 ;
        RECT 688.950 96.600 691.050 97.050 ;
        RECT 712.950 96.600 715.050 97.050 ;
        RECT 652.950 95.400 715.050 96.600 ;
        RECT 652.950 94.950 655.050 95.400 ;
        RECT 688.950 94.950 691.050 95.400 ;
        RECT 712.950 94.950 715.050 95.400 ;
        RECT 721.950 96.600 724.050 97.050 ;
        RECT 727.950 96.600 730.050 97.050 ;
        RECT 721.950 95.400 730.050 96.600 ;
        RECT 721.950 94.950 724.050 95.400 ;
        RECT 727.950 94.950 730.050 95.400 ;
        RECT 811.950 96.600 814.050 97.050 ;
        RECT 820.950 96.600 823.050 97.050 ;
        RECT 811.950 95.400 823.050 96.600 ;
        RECT 811.950 94.950 814.050 95.400 ;
        RECT 820.950 94.950 823.050 95.400 ;
        RECT 40.950 93.600 43.050 94.050 ;
        RECT 52.950 93.600 55.050 94.050 ;
        RECT 40.950 92.400 55.050 93.600 ;
        RECT 40.950 91.950 43.050 92.400 ;
        RECT 52.950 91.950 55.050 92.400 ;
        RECT 121.950 93.600 124.050 94.050 ;
        RECT 169.950 93.600 172.050 94.050 ;
        RECT 121.950 92.400 172.050 93.600 ;
        RECT 121.950 91.950 124.050 92.400 ;
        RECT 169.950 91.950 172.050 92.400 ;
        RECT 181.950 93.600 184.050 94.050 ;
        RECT 211.950 93.600 214.050 94.050 ;
        RECT 181.950 92.400 214.050 93.600 ;
        RECT 181.950 91.950 184.050 92.400 ;
        RECT 211.950 91.950 214.050 92.400 ;
        RECT 232.950 93.600 235.050 94.050 ;
        RECT 247.950 93.600 250.050 94.050 ;
        RECT 232.950 92.400 250.050 93.600 ;
        RECT 232.950 91.950 235.050 92.400 ;
        RECT 247.950 91.950 250.050 92.400 ;
        RECT 445.950 93.600 448.050 94.050 ;
        RECT 472.950 93.600 475.050 94.050 ;
        RECT 445.950 92.400 475.050 93.600 ;
        RECT 445.950 91.950 448.050 92.400 ;
        RECT 472.950 91.950 475.050 92.400 ;
        RECT 487.950 93.600 490.050 94.050 ;
        RECT 541.950 93.600 544.050 94.050 ;
        RECT 487.950 92.400 544.050 93.600 ;
        RECT 487.950 91.950 490.050 92.400 ;
        RECT 541.950 91.950 544.050 92.400 ;
        RECT 550.950 93.600 553.050 94.050 ;
        RECT 637.950 93.600 640.050 94.050 ;
        RECT 550.950 92.400 640.050 93.600 ;
        RECT 550.950 91.950 553.050 92.400 ;
        RECT 637.950 91.950 640.050 92.400 ;
        RECT 655.950 93.600 658.050 94.050 ;
        RECT 685.950 93.600 688.050 94.050 ;
        RECT 655.950 92.400 688.050 93.600 ;
        RECT 713.400 93.600 714.600 94.950 ;
        RECT 745.950 93.600 748.050 94.050 ;
        RECT 713.400 92.400 748.050 93.600 ;
        RECT 655.950 91.950 658.050 92.400 ;
        RECT 685.950 91.950 688.050 92.400 ;
        RECT 745.950 91.950 748.050 92.400 ;
        RECT 787.950 93.600 790.050 94.050 ;
        RECT 826.950 93.600 829.050 93.900 ;
        RECT 877.950 93.600 880.050 94.050 ;
        RECT 895.950 93.600 898.050 94.050 ;
        RECT 787.950 93.000 810.600 93.600 ;
        RECT 787.950 92.400 811.050 93.000 ;
        RECT 787.950 91.950 790.050 92.400 ;
        RECT 34.950 90.600 37.050 91.050 ;
        RECT 64.950 90.600 67.050 91.050 ;
        RECT 34.950 89.400 67.050 90.600 ;
        RECT 34.950 88.950 37.050 89.400 ;
        RECT 64.950 88.950 67.050 89.400 ;
        RECT 193.950 90.600 196.050 91.050 ;
        RECT 229.950 90.600 232.050 91.050 ;
        RECT 193.950 89.400 232.050 90.600 ;
        RECT 193.950 88.950 196.050 89.400 ;
        RECT 229.950 88.950 232.050 89.400 ;
        RECT 577.950 90.600 580.050 91.050 ;
        RECT 589.950 90.600 592.050 91.050 ;
        RECT 577.950 89.400 592.050 90.600 ;
        RECT 577.950 88.950 580.050 89.400 ;
        RECT 589.950 88.950 592.050 89.400 ;
        RECT 595.950 90.600 598.050 91.050 ;
        RECT 634.950 90.600 637.050 90.900 ;
        RECT 595.950 89.400 637.050 90.600 ;
        RECT 595.950 88.950 598.050 89.400 ;
        RECT 634.950 88.800 637.050 89.400 ;
        RECT 646.950 90.600 649.050 91.050 ;
        RECT 652.950 90.600 655.050 91.050 ;
        RECT 646.950 89.400 655.050 90.600 ;
        RECT 646.950 88.950 649.050 89.400 ;
        RECT 652.950 88.950 655.050 89.400 ;
        RECT 658.950 90.600 661.050 91.050 ;
        RECT 700.950 90.600 703.050 91.050 ;
        RECT 658.950 89.400 703.050 90.600 ;
        RECT 658.950 88.950 661.050 89.400 ;
        RECT 700.950 88.950 703.050 89.400 ;
        RECT 706.950 90.600 709.050 91.050 ;
        RECT 784.950 90.600 787.050 91.050 ;
        RECT 706.950 89.400 787.050 90.600 ;
        RECT 706.950 88.950 709.050 89.400 ;
        RECT 784.950 88.950 787.050 89.400 ;
        RECT 808.950 88.950 811.050 92.400 ;
        RECT 826.950 92.400 898.050 93.600 ;
        RECT 826.950 91.800 829.050 92.400 ;
        RECT 877.950 91.950 880.050 92.400 ;
        RECT 895.950 91.950 898.050 92.400 ;
        RECT 934.950 93.600 937.050 94.050 ;
        RECT 982.950 93.600 985.050 94.050 ;
        RECT 934.950 92.400 985.050 93.600 ;
        RECT 934.950 91.950 937.050 92.400 ;
        RECT 982.950 91.950 985.050 92.400 ;
        RECT 943.950 90.600 946.050 91.050 ;
        RECT 958.950 90.600 961.050 91.050 ;
        RECT 943.950 89.400 961.050 90.600 ;
        RECT 943.950 88.950 946.050 89.400 ;
        RECT 958.950 88.950 961.050 89.400 ;
        RECT 244.950 87.600 247.050 88.050 ;
        RECT 265.950 87.600 268.050 88.050 ;
        RECT 244.950 86.400 268.050 87.600 ;
        RECT 244.950 85.950 247.050 86.400 ;
        RECT 265.950 85.950 268.050 86.400 ;
        RECT 415.950 87.600 418.050 88.050 ;
        RECT 466.950 87.600 469.050 88.050 ;
        RECT 415.950 86.400 469.050 87.600 ;
        RECT 415.950 85.950 418.050 86.400 ;
        RECT 466.950 85.950 469.050 86.400 ;
        RECT 655.950 87.600 658.050 88.050 ;
        RECT 718.950 87.600 721.050 88.050 ;
        RECT 763.950 87.600 766.050 88.050 ;
        RECT 655.950 86.400 766.050 87.600 ;
        RECT 655.950 85.950 658.050 86.400 ;
        RECT 718.950 85.950 721.050 86.400 ;
        RECT 763.950 85.950 766.050 86.400 ;
        RECT 601.950 84.600 604.050 85.050 ;
        RECT 697.950 84.600 700.050 85.050 ;
        RECT 601.950 83.400 700.050 84.600 ;
        RECT 601.950 82.950 604.050 83.400 ;
        RECT 697.950 82.950 700.050 83.400 ;
        RECT 805.950 84.600 808.050 85.050 ;
        RECT 814.950 84.600 817.050 85.050 ;
        RECT 805.950 83.400 817.050 84.600 ;
        RECT 805.950 82.950 808.050 83.400 ;
        RECT 814.950 82.950 817.050 83.400 ;
        RECT 358.950 81.600 361.050 82.050 ;
        RECT 376.950 81.600 379.050 82.050 ;
        RECT 385.950 81.600 388.050 82.050 ;
        RECT 358.950 80.400 388.050 81.600 ;
        RECT 358.950 79.950 361.050 80.400 ;
        RECT 376.950 79.950 379.050 80.400 ;
        RECT 385.950 79.950 388.050 80.400 ;
        RECT 430.950 81.600 433.050 82.050 ;
        RECT 454.950 81.600 457.050 82.050 ;
        RECT 430.950 80.400 457.050 81.600 ;
        RECT 430.950 79.950 433.050 80.400 ;
        RECT 454.950 79.950 457.050 80.400 ;
        RECT 574.950 81.600 577.050 82.050 ;
        RECT 592.950 81.600 595.050 82.050 ;
        RECT 721.950 81.600 724.050 82.050 ;
        RECT 574.950 80.400 724.050 81.600 ;
        RECT 574.950 79.950 577.050 80.400 ;
        RECT 592.950 79.950 595.050 80.400 ;
        RECT 721.950 79.950 724.050 80.400 ;
        RECT 19.950 78.600 22.050 79.050 ;
        RECT 25.950 78.600 28.050 79.050 ;
        RECT 52.950 78.600 55.050 79.050 ;
        RECT 19.950 77.400 55.050 78.600 ;
        RECT 19.950 76.950 22.050 77.400 ;
        RECT 25.950 76.950 28.050 77.400 ;
        RECT 52.950 76.950 55.050 77.400 ;
        RECT 466.950 78.600 469.050 79.050 ;
        RECT 526.950 78.600 529.050 79.050 ;
        RECT 466.950 77.400 529.050 78.600 ;
        RECT 466.950 76.950 469.050 77.400 ;
        RECT 526.950 76.950 529.050 77.400 ;
        RECT 622.950 78.600 625.050 79.050 ;
        RECT 649.950 78.600 652.050 79.050 ;
        RECT 622.950 77.400 652.050 78.600 ;
        RECT 622.950 76.950 625.050 77.400 ;
        RECT 649.950 76.950 652.050 77.400 ;
        RECT 790.950 78.600 793.050 79.050 ;
        RECT 811.950 78.600 814.050 79.050 ;
        RECT 790.950 77.400 814.050 78.600 ;
        RECT 790.950 76.950 793.050 77.400 ;
        RECT 811.950 76.950 814.050 77.400 ;
        RECT 97.950 75.600 100.050 76.050 ;
        RECT 184.950 75.600 187.050 76.050 ;
        RECT 199.950 75.600 202.050 76.050 ;
        RECT 208.950 75.600 211.050 76.050 ;
        RECT 97.950 74.400 211.050 75.600 ;
        RECT 97.950 73.950 100.050 74.400 ;
        RECT 184.950 73.950 187.050 74.400 ;
        RECT 199.950 73.950 202.050 74.400 ;
        RECT 208.950 73.950 211.050 74.400 ;
        RECT 232.950 75.600 235.050 76.050 ;
        RECT 391.950 75.600 394.050 76.050 ;
        RECT 403.950 75.600 406.050 76.050 ;
        RECT 232.950 74.400 406.050 75.600 ;
        RECT 232.950 73.950 235.050 74.400 ;
        RECT 391.950 73.950 394.050 74.400 ;
        RECT 403.950 73.950 406.050 74.400 ;
        RECT 454.950 75.600 457.050 76.050 ;
        RECT 613.950 75.600 616.050 76.050 ;
        RECT 454.950 74.400 616.050 75.600 ;
        RECT 454.950 73.950 457.050 74.400 ;
        RECT 613.950 73.950 616.050 74.400 ;
        RECT 145.950 72.600 148.050 73.050 ;
        RECT 157.950 72.600 160.050 73.050 ;
        RECT 178.950 72.600 181.050 73.050 ;
        RECT 145.950 71.400 181.050 72.600 ;
        RECT 145.950 70.950 148.050 71.400 ;
        RECT 157.950 70.950 160.050 71.400 ;
        RECT 178.950 70.950 181.050 71.400 ;
        RECT 220.950 72.600 223.050 73.050 ;
        RECT 259.950 72.600 262.050 73.050 ;
        RECT 220.950 71.400 262.050 72.600 ;
        RECT 220.950 70.950 223.050 71.400 ;
        RECT 259.950 70.950 262.050 71.400 ;
        RECT 268.950 72.600 271.050 73.050 ;
        RECT 355.950 72.600 358.050 73.050 ;
        RECT 268.950 71.400 358.050 72.600 ;
        RECT 268.950 70.950 271.050 71.400 ;
        RECT 355.950 70.950 358.050 71.400 ;
        RECT 478.950 72.600 481.050 73.050 ;
        RECT 487.950 72.600 490.050 73.050 ;
        RECT 478.950 71.400 490.050 72.600 ;
        RECT 478.950 70.950 481.050 71.400 ;
        RECT 487.950 70.950 490.050 71.400 ;
        RECT 523.950 72.600 526.050 73.050 ;
        RECT 538.950 72.600 541.050 73.050 ;
        RECT 523.950 71.400 541.050 72.600 ;
        RECT 523.950 70.950 526.050 71.400 ;
        RECT 538.950 70.950 541.050 71.400 ;
        RECT 580.950 72.600 583.050 73.050 ;
        RECT 667.950 72.600 670.050 73.050 ;
        RECT 580.950 71.400 670.050 72.600 ;
        RECT 580.950 70.950 583.050 71.400 ;
        RECT 667.950 70.950 670.050 71.400 ;
        RECT 76.950 69.600 79.050 70.050 ;
        RECT 85.950 69.600 88.050 70.050 ;
        RECT 76.950 68.400 88.050 69.600 ;
        RECT 76.950 67.950 79.050 68.400 ;
        RECT 85.950 67.950 88.050 68.400 ;
        RECT 121.950 69.600 124.050 70.050 ;
        RECT 136.950 69.600 139.050 70.050 ;
        RECT 121.950 68.400 139.050 69.600 ;
        RECT 121.950 67.950 124.050 68.400 ;
        RECT 136.950 67.950 139.050 68.400 ;
        RECT 166.950 69.600 169.050 70.050 ;
        RECT 202.950 69.600 205.050 70.050 ;
        RECT 205.950 69.600 208.050 70.050 ;
        RECT 364.950 69.600 367.050 70.050 ;
        RECT 412.950 69.600 415.050 70.050 ;
        RECT 436.950 69.600 439.050 70.050 ;
        RECT 166.950 68.400 367.050 69.600 ;
        RECT 166.950 67.950 169.050 68.400 ;
        RECT 202.950 67.950 205.050 68.400 ;
        RECT 205.950 67.950 208.050 68.400 ;
        RECT 364.950 67.950 367.050 68.400 ;
        RECT 371.400 68.400 439.050 69.600 ;
        RECT 97.950 66.600 100.050 67.050 ;
        RECT 106.950 66.600 109.050 67.050 ;
        RECT 124.950 66.600 127.050 67.050 ;
        RECT 97.950 65.400 127.050 66.600 ;
        RECT 97.950 64.950 100.050 65.400 ;
        RECT 106.950 64.950 109.050 65.400 ;
        RECT 124.950 64.950 127.050 65.400 ;
        RECT 247.950 66.600 250.050 67.050 ;
        RECT 304.950 66.600 307.050 67.050 ;
        RECT 337.950 66.600 340.050 67.050 ;
        RECT 247.950 65.400 340.050 66.600 ;
        RECT 247.950 64.950 250.050 65.400 ;
        RECT 304.950 64.950 307.050 65.400 ;
        RECT 337.950 64.950 340.050 65.400 ;
        RECT 352.950 66.600 355.050 67.050 ;
        RECT 371.400 66.600 372.600 68.400 ;
        RECT 412.950 67.950 415.050 68.400 ;
        RECT 436.950 67.950 439.050 68.400 ;
        RECT 460.950 69.600 463.050 70.050 ;
        RECT 490.950 69.600 493.050 70.050 ;
        RECT 508.950 69.600 511.050 70.050 ;
        RECT 460.950 68.400 511.050 69.600 ;
        RECT 460.950 67.950 463.050 68.400 ;
        RECT 490.950 67.950 493.050 68.400 ;
        RECT 508.950 67.950 511.050 68.400 ;
        RECT 724.950 69.600 727.050 70.050 ;
        RECT 775.950 69.600 778.050 70.050 ;
        RECT 724.950 68.400 778.050 69.600 ;
        RECT 724.950 67.950 727.050 68.400 ;
        RECT 775.950 67.950 778.050 68.400 ;
        RECT 886.950 69.600 889.050 70.050 ;
        RECT 925.950 69.600 928.050 70.050 ;
        RECT 946.950 69.600 949.050 70.050 ;
        RECT 886.950 68.400 949.050 69.600 ;
        RECT 886.950 67.950 889.050 68.400 ;
        RECT 925.950 67.950 928.050 68.400 ;
        RECT 946.950 67.950 949.050 68.400 ;
        RECT 352.950 65.400 372.600 66.600 ;
        RECT 577.950 66.600 580.050 67.050 ;
        RECT 607.950 66.600 610.050 67.050 ;
        RECT 577.950 65.400 610.050 66.600 ;
        RECT 352.950 64.950 355.050 65.400 ;
        RECT 577.950 64.950 580.050 65.400 ;
        RECT 607.950 64.950 610.050 65.400 ;
        RECT 661.950 66.600 664.050 67.050 ;
        RECT 706.950 66.600 709.050 67.050 ;
        RECT 661.950 65.400 709.050 66.600 ;
        RECT 661.950 64.950 664.050 65.400 ;
        RECT 706.950 64.950 709.050 65.400 ;
        RECT 49.950 63.600 52.050 64.050 ;
        RECT 67.950 63.600 70.050 64.050 ;
        RECT 49.950 62.400 70.050 63.600 ;
        RECT 49.950 61.950 52.050 62.400 ;
        RECT 67.950 61.950 70.050 62.400 ;
        RECT 94.950 63.600 97.050 64.050 ;
        RECT 130.950 63.600 133.050 64.050 ;
        RECT 154.950 63.600 157.050 64.050 ;
        RECT 172.950 63.600 175.050 64.050 ;
        RECT 196.950 63.600 199.050 64.050 ;
        RECT 226.950 63.600 229.050 64.050 ;
        RECT 94.950 62.400 229.050 63.600 ;
        RECT 94.950 61.950 97.050 62.400 ;
        RECT 130.950 61.950 133.050 62.400 ;
        RECT 154.950 61.950 157.050 62.400 ;
        RECT 172.950 61.950 175.050 62.400 ;
        RECT 196.950 61.950 199.050 62.400 ;
        RECT 226.950 61.950 229.050 62.400 ;
        RECT 424.950 63.600 427.050 64.050 ;
        RECT 460.950 63.600 463.050 64.050 ;
        RECT 424.950 62.400 463.050 63.600 ;
        RECT 424.950 61.950 427.050 62.400 ;
        RECT 460.950 61.950 463.050 62.400 ;
        RECT 844.950 63.600 847.050 64.050 ;
        RECT 877.950 63.600 880.050 64.050 ;
        RECT 901.950 63.600 904.050 64.050 ;
        RECT 844.950 62.400 904.050 63.600 ;
        RECT 844.950 61.950 847.050 62.400 ;
        RECT 877.950 61.950 880.050 62.400 ;
        RECT 901.950 61.950 904.050 62.400 ;
        RECT 88.950 60.600 91.050 61.200 ;
        RECT 112.950 60.600 115.050 61.200 ;
        RECT 121.950 60.600 124.050 61.050 ;
        RECT 88.950 59.400 124.050 60.600 ;
        RECT 88.950 59.100 91.050 59.400 ;
        RECT 112.950 59.100 115.050 59.400 ;
        RECT 121.950 58.950 124.050 59.400 ;
        RECT 238.950 59.100 241.050 61.200 ;
        RECT 244.950 60.750 247.050 61.200 ;
        RECT 253.950 60.750 256.050 61.200 ;
        RECT 244.950 59.550 256.050 60.750 ;
        RECT 244.950 59.100 247.050 59.550 ;
        RECT 253.950 59.100 256.050 59.550 ;
        RECT 271.950 60.750 274.050 61.200 ;
        RECT 280.950 60.750 283.050 61.200 ;
        RECT 271.950 59.550 283.050 60.750 ;
        RECT 271.950 59.100 274.050 59.550 ;
        RECT 280.950 59.100 283.050 59.550 ;
        RECT 286.950 59.100 289.050 61.200 ;
        RECT 310.950 60.600 313.050 61.200 ;
        RECT 322.950 60.750 325.050 61.200 ;
        RECT 331.950 60.750 334.050 61.200 ;
        RECT 322.950 60.600 334.050 60.750 ;
        RECT 310.950 59.550 334.050 60.600 ;
        RECT 310.950 59.400 325.050 59.550 ;
        RECT 310.950 59.100 313.050 59.400 ;
        RECT 322.950 59.100 325.050 59.400 ;
        RECT 331.950 59.100 334.050 59.550 ;
        RECT 355.950 60.750 358.050 61.200 ;
        RECT 364.950 60.750 367.050 61.200 ;
        RECT 355.950 60.600 367.050 60.750 ;
        RECT 385.950 60.600 388.050 61.200 ;
        RECT 355.950 59.550 388.050 60.600 ;
        RECT 355.950 59.100 358.050 59.550 ;
        RECT 364.950 59.400 388.050 59.550 ;
        RECT 364.950 59.100 367.050 59.400 ;
        RECT 385.950 59.100 388.050 59.400 ;
        RECT 406.950 60.750 409.050 61.200 ;
        RECT 418.950 60.750 421.050 61.200 ;
        RECT 406.950 60.600 421.050 60.750 ;
        RECT 442.950 60.750 445.050 61.200 ;
        RECT 448.950 60.750 451.050 61.200 ;
        RECT 406.950 59.550 435.600 60.600 ;
        RECT 406.950 59.100 409.050 59.550 ;
        RECT 418.950 59.400 435.600 59.550 ;
        RECT 418.950 59.100 421.050 59.400 ;
        RECT 49.950 57.600 52.050 58.050 ;
        RECT 17.400 56.400 52.050 57.600 ;
        RECT 17.400 54.900 18.600 56.400 ;
        RECT 49.950 55.950 52.050 56.400 ;
        RECT 16.950 52.800 19.050 54.900 ;
        RECT 31.950 54.450 34.050 54.900 ;
        RECT 40.950 54.450 43.050 54.900 ;
        RECT 31.950 53.250 43.050 54.450 ;
        RECT 31.950 52.800 34.050 53.250 ;
        RECT 40.950 52.800 43.050 53.250 ;
        RECT 52.950 54.450 55.050 54.900 ;
        RECT 58.950 54.450 61.050 54.900 ;
        RECT 52.950 53.250 61.050 54.450 ;
        RECT 52.950 52.800 55.050 53.250 ;
        RECT 58.950 52.800 61.050 53.250 ;
        RECT 64.950 54.600 67.050 54.900 ;
        RECT 76.800 54.600 78.900 55.050 ;
        RECT 64.950 53.400 78.900 54.600 ;
        RECT 64.950 52.800 67.050 53.400 ;
        RECT 76.800 52.950 78.900 53.400 ;
        RECT 79.950 54.600 82.050 55.050 ;
        RECT 85.950 54.600 88.050 54.900 ;
        RECT 79.950 54.450 88.050 54.600 ;
        RECT 100.950 54.450 103.050 54.900 ;
        RECT 79.950 53.400 103.050 54.450 ;
        RECT 79.950 52.950 82.050 53.400 ;
        RECT 85.950 53.250 103.050 53.400 ;
        RECT 85.950 52.800 88.050 53.250 ;
        RECT 100.950 52.800 103.050 53.250 ;
        RECT 172.950 54.450 175.050 54.900 ;
        RECT 181.950 54.450 184.050 54.900 ;
        RECT 172.950 53.250 184.050 54.450 ;
        RECT 172.950 52.800 175.050 53.250 ;
        RECT 181.950 52.800 184.050 53.250 ;
        RECT 187.950 54.600 190.050 54.900 ;
        RECT 193.800 54.600 195.900 55.050 ;
        RECT 187.950 53.400 195.900 54.600 ;
        RECT 187.950 52.800 190.050 53.400 ;
        RECT 193.800 52.950 195.900 53.400 ;
        RECT 196.950 54.450 199.050 54.900 ;
        RECT 205.950 54.450 208.050 54.900 ;
        RECT 196.950 53.250 208.050 54.450 ;
        RECT 196.950 52.800 199.050 53.250 ;
        RECT 205.950 52.800 208.050 53.250 ;
        RECT 211.950 54.600 214.050 54.900 ;
        RECT 229.950 54.600 232.050 54.900 ;
        RECT 211.950 53.400 232.050 54.600 ;
        RECT 239.400 54.600 240.600 59.100 ;
        RECT 287.400 57.600 288.600 59.100 ;
        RECT 295.950 57.600 298.050 58.050 ;
        RECT 287.400 56.400 298.050 57.600 ;
        RECT 295.950 55.950 298.050 56.400 ;
        RECT 256.950 54.600 259.050 54.900 ;
        RECT 239.400 53.400 259.050 54.600 ;
        RECT 211.950 52.800 214.050 53.400 ;
        RECT 229.950 52.800 232.050 53.400 ;
        RECT 256.950 52.800 259.050 53.400 ;
        RECT 262.950 54.600 265.050 54.900 ;
        RECT 268.950 54.600 271.050 55.050 ;
        RECT 262.950 53.400 271.050 54.600 ;
        RECT 262.950 52.800 265.050 53.400 ;
        RECT 268.950 52.950 271.050 53.400 ;
        RECT 289.950 54.600 292.050 54.900 ;
        RECT 307.950 54.600 310.050 54.900 ;
        RECT 334.950 54.600 337.050 54.900 ;
        RECT 289.950 53.400 337.050 54.600 ;
        RECT 289.950 52.800 292.050 53.400 ;
        RECT 307.950 52.800 310.050 53.400 ;
        RECT 334.950 52.800 337.050 53.400 ;
        RECT 340.950 54.600 343.050 54.900 ;
        RECT 352.950 54.600 355.050 55.050 ;
        RECT 434.400 54.900 435.600 59.400 ;
        RECT 442.950 59.550 451.050 60.750 ;
        RECT 442.950 59.100 445.050 59.550 ;
        RECT 448.950 59.100 451.050 59.550 ;
        RECT 454.950 58.950 457.050 61.050 ;
        RECT 484.950 60.750 487.050 61.200 ;
        RECT 496.950 60.750 499.050 61.200 ;
        RECT 484.950 59.550 499.050 60.750 ;
        RECT 484.950 59.100 487.050 59.550 ;
        RECT 496.950 59.100 499.050 59.550 ;
        RECT 517.950 60.600 520.050 61.200 ;
        RECT 532.950 60.600 535.050 61.200 ;
        RECT 517.950 59.400 535.050 60.600 ;
        RECT 517.950 59.100 520.050 59.400 ;
        RECT 532.950 59.100 535.050 59.400 ;
        RECT 571.950 60.750 574.050 61.200 ;
        RECT 586.950 60.750 589.050 61.200 ;
        RECT 571.950 59.550 589.050 60.750 ;
        RECT 571.950 59.100 574.050 59.550 ;
        RECT 586.950 59.100 589.050 59.550 ;
        RECT 634.950 60.600 637.050 61.200 ;
        RECT 655.950 60.600 658.050 61.200 ;
        RECT 634.950 59.400 658.050 60.600 ;
        RECT 634.950 59.100 637.050 59.400 ;
        RECT 655.950 59.100 658.050 59.400 ;
        RECT 673.950 60.750 676.050 61.200 ;
        RECT 679.950 60.750 682.050 61.200 ;
        RECT 673.950 59.550 682.050 60.750 ;
        RECT 706.950 60.600 709.050 61.200 ;
        RECT 673.950 59.100 676.050 59.550 ;
        RECT 679.950 59.100 682.050 59.550 ;
        RECT 701.400 59.400 709.050 60.600 ;
        RECT 340.950 53.400 355.050 54.600 ;
        RECT 340.950 52.800 343.050 53.400 ;
        RECT 352.950 52.950 355.050 53.400 ;
        RECT 376.950 54.450 379.050 54.900 ;
        RECT 388.950 54.450 391.050 54.900 ;
        RECT 376.950 53.250 391.050 54.450 ;
        RECT 376.950 52.800 379.050 53.250 ;
        RECT 388.950 52.800 391.050 53.250 ;
        RECT 403.950 54.450 406.050 54.900 ;
        RECT 409.950 54.450 412.050 54.900 ;
        RECT 403.950 53.250 412.050 54.450 ;
        RECT 403.950 52.800 406.050 53.250 ;
        RECT 409.950 52.800 412.050 53.250 ;
        RECT 433.950 52.800 436.050 54.900 ;
        RECT 439.950 54.600 442.050 54.900 ;
        RECT 455.400 54.600 456.600 58.950 ;
        RECT 526.950 57.600 529.050 58.050 ;
        RECT 598.950 57.600 601.050 58.050 ;
        RECT 526.950 56.400 537.600 57.600 ;
        RECT 526.950 55.950 529.050 56.400 ;
        RECT 439.950 53.400 456.600 54.600 ;
        RECT 463.950 54.600 466.050 54.900 ;
        RECT 496.950 54.600 499.050 55.050 ;
        RECT 536.400 54.900 537.600 56.400 ;
        RECT 598.950 56.400 615.600 57.600 ;
        RECT 598.950 55.950 601.050 56.400 ;
        RECT 514.950 54.600 517.050 54.900 ;
        RECT 463.950 53.400 517.050 54.600 ;
        RECT 439.950 52.800 442.050 53.400 ;
        RECT 463.950 52.800 466.050 53.400 ;
        RECT 496.950 52.950 499.050 53.400 ;
        RECT 514.950 52.800 517.050 53.400 ;
        RECT 535.950 52.800 538.050 54.900 ;
        RECT 541.950 52.800 544.050 54.900 ;
        RECT 562.950 54.450 565.050 54.900 ;
        RECT 574.950 54.450 577.050 54.900 ;
        RECT 562.950 53.250 577.050 54.450 ;
        RECT 562.950 52.800 565.050 53.250 ;
        RECT 574.950 52.800 577.050 53.250 ;
        RECT 601.950 54.450 604.050 54.900 ;
        RECT 610.950 54.450 613.050 54.900 ;
        RECT 601.950 53.250 613.050 54.450 ;
        RECT 614.400 54.600 615.600 56.400 ;
        RECT 631.950 54.600 634.050 54.900 ;
        RECT 614.400 53.400 634.050 54.600 ;
        RECT 601.950 52.800 604.050 53.250 ;
        RECT 610.950 52.800 613.050 53.250 ;
        RECT 631.950 52.800 634.050 53.400 ;
        RECT 652.950 54.450 655.050 54.900 ;
        RECT 658.950 54.450 661.050 54.900 ;
        RECT 652.950 53.250 661.050 54.450 ;
        RECT 652.950 52.800 655.050 53.250 ;
        RECT 658.950 52.800 661.050 53.250 ;
        RECT 415.950 51.600 418.050 52.050 ;
        RECT 463.950 51.600 466.050 52.050 ;
        RECT 415.950 50.400 466.050 51.600 ;
        RECT 415.950 49.950 418.050 50.400 ;
        RECT 463.950 49.950 466.050 50.400 ;
        RECT 472.950 51.600 475.050 52.050 ;
        RECT 487.950 51.600 490.050 52.050 ;
        RECT 472.950 50.400 490.050 51.600 ;
        RECT 472.950 49.950 475.050 50.400 ;
        RECT 487.950 49.950 490.050 50.400 ;
        RECT 16.950 48.600 19.050 49.050 ;
        RECT 46.950 48.600 49.050 49.050 ;
        RECT 73.950 48.600 76.050 49.050 ;
        RECT 109.950 48.600 112.050 49.050 ;
        RECT 16.950 47.400 112.050 48.600 ;
        RECT 16.950 46.950 19.050 47.400 ;
        RECT 46.950 46.950 49.050 47.400 ;
        RECT 73.950 46.950 76.050 47.400 ;
        RECT 109.950 46.950 112.050 47.400 ;
        RECT 133.950 48.600 136.050 49.050 ;
        RECT 247.950 48.600 250.050 49.050 ;
        RECT 133.950 47.400 250.050 48.600 ;
        RECT 133.950 46.950 136.050 47.400 ;
        RECT 247.950 46.950 250.050 47.400 ;
        RECT 262.950 48.600 265.050 49.050 ;
        RECT 295.950 48.600 298.050 49.050 ;
        RECT 358.950 48.600 361.050 49.050 ;
        RECT 430.950 48.600 433.050 49.050 ;
        RECT 436.950 48.600 439.050 49.050 ;
        RECT 457.950 48.600 460.050 49.050 ;
        RECT 262.950 47.400 429.600 48.600 ;
        RECT 262.950 46.950 265.050 47.400 ;
        RECT 295.950 46.950 298.050 47.400 ;
        RECT 358.950 46.950 361.050 47.400 ;
        RECT 313.950 45.600 316.050 46.050 ;
        RECT 361.950 45.600 364.050 46.050 ;
        RECT 313.950 44.400 364.050 45.600 ;
        RECT 313.950 43.950 316.050 44.400 ;
        RECT 361.950 43.950 364.050 44.400 ;
        RECT 367.950 45.600 370.050 46.050 ;
        RECT 424.950 45.600 427.050 46.050 ;
        RECT 367.950 44.400 427.050 45.600 ;
        RECT 428.400 45.600 429.600 47.400 ;
        RECT 430.950 47.400 460.050 48.600 ;
        RECT 430.950 46.950 433.050 47.400 ;
        RECT 436.950 46.950 439.050 47.400 ;
        RECT 457.950 46.950 460.050 47.400 ;
        RECT 484.950 48.600 487.050 49.050 ;
        RECT 542.400 48.600 543.600 52.800 ;
        RECT 701.400 52.050 702.600 59.400 ;
        RECT 706.950 59.100 709.050 59.400 ;
        RECT 712.950 59.100 715.050 61.200 ;
        RECT 748.950 60.750 751.050 61.200 ;
        RECT 781.950 60.750 784.050 61.200 ;
        RECT 748.950 59.550 784.050 60.750 ;
        RECT 748.950 59.100 751.050 59.550 ;
        RECT 781.950 59.100 784.050 59.550 ;
        RECT 793.950 60.750 796.050 61.200 ;
        RECT 799.950 60.750 802.050 61.200 ;
        RECT 793.950 59.550 802.050 60.750 ;
        RECT 793.950 59.100 796.050 59.550 ;
        RECT 799.950 59.100 802.050 59.550 ;
        RECT 826.950 60.600 829.050 61.200 ;
        RECT 844.950 60.600 847.050 61.200 ;
        RECT 826.950 59.400 847.050 60.600 ;
        RECT 826.950 59.100 829.050 59.400 ;
        RECT 844.950 59.100 847.050 59.400 ;
        RECT 850.950 59.100 853.050 61.200 ;
        RECT 862.950 60.750 865.050 61.200 ;
        RECT 871.950 60.750 874.050 61.200 ;
        RECT 862.950 59.550 874.050 60.750 ;
        RECT 862.950 59.100 865.050 59.550 ;
        RECT 871.950 59.100 874.050 59.550 ;
        RECT 886.950 60.750 889.050 61.200 ;
        RECT 895.950 60.750 898.050 61.200 ;
        RECT 886.950 59.550 898.050 60.750 ;
        RECT 886.950 59.100 889.050 59.550 ;
        RECT 895.950 59.100 898.050 59.550 ;
        RECT 919.950 60.600 922.050 61.200 ;
        RECT 940.950 60.600 943.050 61.200 ;
        RECT 919.950 59.400 943.050 60.600 ;
        RECT 919.950 59.100 922.050 59.400 ;
        RECT 940.950 59.100 943.050 59.400 ;
        RECT 958.950 60.750 961.050 61.200 ;
        RECT 964.950 60.750 967.050 61.200 ;
        RECT 958.950 59.550 967.050 60.750 ;
        RECT 958.950 59.100 961.050 59.550 ;
        RECT 964.950 59.100 967.050 59.550 ;
        RECT 979.950 60.750 982.050 61.200 ;
        RECT 997.950 60.750 1000.050 61.200 ;
        RECT 979.950 59.550 1000.050 60.750 ;
        RECT 979.950 59.100 982.050 59.550 ;
        RECT 997.950 59.100 1000.050 59.550 ;
        RECT 713.400 57.600 714.600 59.100 ;
        RECT 724.950 57.600 727.050 58.050 ;
        RECT 713.400 56.400 727.050 57.600 ;
        RECT 724.950 55.950 727.050 56.400 ;
        RECT 851.400 55.050 852.600 59.100 ;
        RECT 748.950 54.450 751.050 54.900 ;
        RECT 760.950 54.450 763.050 54.900 ;
        RECT 748.950 53.250 763.050 54.450 ;
        RECT 748.950 52.800 751.050 53.250 ;
        RECT 760.950 52.800 763.050 53.250 ;
        RECT 808.950 54.600 811.050 54.900 ;
        RECT 841.950 54.600 844.050 54.900 ;
        RECT 808.950 53.400 844.050 54.600 ;
        RECT 851.400 53.400 855.900 55.050 ;
        RECT 808.950 52.800 811.050 53.400 ;
        RECT 841.950 52.800 844.050 53.400 ;
        RECT 852.000 52.950 855.900 53.400 ;
        RECT 856.950 54.600 859.050 55.050 ;
        RECT 892.950 54.600 895.050 54.900 ;
        RECT 856.950 53.400 895.050 54.600 ;
        RECT 856.950 52.950 859.050 53.400 ;
        RECT 892.950 52.800 895.050 53.400 ;
        RECT 922.950 54.450 925.050 54.900 ;
        RECT 931.950 54.600 934.050 54.900 ;
        RECT 943.950 54.600 946.050 54.900 ;
        RECT 931.950 54.450 946.050 54.600 ;
        RECT 922.950 53.400 946.050 54.450 ;
        RECT 922.950 53.250 934.050 53.400 ;
        RECT 922.950 52.800 925.050 53.250 ;
        RECT 931.950 52.800 934.050 53.250 ;
        RECT 943.950 52.800 946.050 53.400 ;
        RECT 967.950 54.600 970.050 54.900 ;
        RECT 982.950 54.600 985.050 55.050 ;
        RECT 967.950 53.400 985.050 54.600 ;
        RECT 967.950 52.800 970.050 53.400 ;
        RECT 982.950 52.950 985.050 53.400 ;
        RECT 586.950 51.600 589.050 52.050 ;
        RECT 643.950 51.600 646.050 52.050 ;
        RECT 649.950 51.600 652.050 52.050 ;
        RECT 586.950 50.400 652.050 51.600 ;
        RECT 586.950 49.950 589.050 50.400 ;
        RECT 643.950 49.950 646.050 50.400 ;
        RECT 649.950 49.950 652.050 50.400 ;
        RECT 700.950 49.950 703.050 52.050 ;
        RECT 802.950 51.600 805.050 52.050 ;
        RECT 814.950 51.600 817.050 52.050 ;
        RECT 802.950 50.400 817.050 51.600 ;
        RECT 802.950 49.950 805.050 50.400 ;
        RECT 814.950 49.950 817.050 50.400 ;
        RECT 847.950 51.600 850.050 52.050 ;
        RECT 862.950 51.600 865.050 52.050 ;
        RECT 898.950 51.600 901.050 52.050 ;
        RECT 958.950 51.600 961.050 52.050 ;
        RECT 847.950 50.400 961.050 51.600 ;
        RECT 847.950 49.950 850.050 50.400 ;
        RECT 862.950 49.950 865.050 50.400 ;
        RECT 898.950 49.950 901.050 50.400 ;
        RECT 958.950 49.950 961.050 50.400 ;
        RECT 484.950 47.400 543.600 48.600 ;
        RECT 550.950 48.600 553.050 49.050 ;
        RECT 616.950 48.600 619.050 49.050 ;
        RECT 769.950 48.600 772.050 49.050 ;
        RECT 793.950 48.600 796.050 49.050 ;
        RECT 550.950 47.400 796.050 48.600 ;
        RECT 484.950 46.950 487.050 47.400 ;
        RECT 550.950 46.950 553.050 47.400 ;
        RECT 616.950 46.950 619.050 47.400 ;
        RECT 769.950 46.950 772.050 47.400 ;
        RECT 793.950 46.950 796.050 47.400 ;
        RECT 853.950 48.600 856.050 49.050 ;
        RECT 874.950 48.600 877.050 49.050 ;
        RECT 886.950 48.600 889.050 49.050 ;
        RECT 910.950 48.600 913.050 49.050 ;
        RECT 853.950 47.400 913.050 48.600 ;
        RECT 853.950 46.950 856.050 47.400 ;
        RECT 874.950 46.950 877.050 47.400 ;
        RECT 886.950 46.950 889.050 47.400 ;
        RECT 910.950 46.950 913.050 47.400 ;
        RECT 541.950 45.600 544.050 46.050 ;
        RECT 428.400 44.400 544.050 45.600 ;
        RECT 367.950 43.950 370.050 44.400 ;
        RECT 424.950 43.950 427.050 44.400 ;
        RECT 541.950 43.950 544.050 44.400 ;
        RECT 796.950 45.600 799.050 46.050 ;
        RECT 844.950 45.600 847.050 46.050 ;
        RECT 796.950 44.400 847.050 45.600 ;
        RECT 796.950 43.950 799.050 44.400 ;
        RECT 844.950 43.950 847.050 44.400 ;
        RECT 859.950 45.600 862.050 46.050 ;
        RECT 868.950 45.600 871.050 46.050 ;
        RECT 859.950 44.400 871.050 45.600 ;
        RECT 859.950 43.950 862.050 44.400 ;
        RECT 868.950 43.950 871.050 44.400 ;
        RECT 955.950 45.600 958.050 46.050 ;
        RECT 994.950 45.600 997.050 46.050 ;
        RECT 955.950 44.400 997.050 45.600 ;
        RECT 955.950 43.950 958.050 44.400 ;
        RECT 994.950 43.950 997.050 44.400 ;
        RECT 115.950 42.600 118.050 43.050 ;
        RECT 187.950 42.600 190.050 43.050 ;
        RECT 208.950 42.600 211.050 43.050 ;
        RECT 115.950 41.400 211.050 42.600 ;
        RECT 115.950 40.950 118.050 41.400 ;
        RECT 187.950 40.950 190.050 41.400 ;
        RECT 208.950 40.950 211.050 41.400 ;
        RECT 235.950 42.600 238.050 43.050 ;
        RECT 244.950 42.600 247.050 43.050 ;
        RECT 268.950 42.600 271.050 43.050 ;
        RECT 235.950 41.400 271.050 42.600 ;
        RECT 362.400 42.600 363.600 43.950 ;
        RECT 448.950 42.600 451.050 43.050 ;
        RECT 362.400 41.400 451.050 42.600 ;
        RECT 235.950 40.950 238.050 41.400 ;
        RECT 244.950 40.950 247.050 41.400 ;
        RECT 268.950 40.950 271.050 41.400 ;
        RECT 448.950 40.950 451.050 41.400 ;
        RECT 496.950 42.600 499.050 43.050 ;
        RECT 550.950 42.600 553.050 43.050 ;
        RECT 496.950 41.400 553.050 42.600 ;
        RECT 496.950 40.950 499.050 41.400 ;
        RECT 550.950 40.950 553.050 41.400 ;
        RECT 574.950 42.600 577.050 43.050 ;
        RECT 580.950 42.600 583.050 43.050 ;
        RECT 574.950 41.400 583.050 42.600 ;
        RECT 574.950 40.950 577.050 41.400 ;
        RECT 580.950 40.950 583.050 41.400 ;
        RECT 619.950 42.600 622.050 43.050 ;
        RECT 658.800 42.600 660.900 43.050 ;
        RECT 619.950 41.400 660.900 42.600 ;
        RECT 619.950 40.950 622.050 41.400 ;
        RECT 658.800 40.950 660.900 41.400 ;
        RECT 661.950 42.600 664.050 43.050 ;
        RECT 670.950 42.600 673.050 43.050 ;
        RECT 661.950 41.400 673.050 42.600 ;
        RECT 661.950 40.950 664.050 41.400 ;
        RECT 670.950 40.950 673.050 41.400 ;
        RECT 790.950 42.600 793.050 43.050 ;
        RECT 799.950 42.600 802.050 43.050 ;
        RECT 790.950 41.400 802.050 42.600 ;
        RECT 790.950 40.950 793.050 41.400 ;
        RECT 799.950 40.950 802.050 41.400 ;
        RECT 826.950 42.600 829.050 43.050 ;
        RECT 838.950 42.600 841.050 43.050 ;
        RECT 826.950 41.400 841.050 42.600 ;
        RECT 826.950 40.950 829.050 41.400 ;
        RECT 838.950 40.950 841.050 41.400 ;
        RECT 892.950 42.600 895.050 43.050 ;
        RECT 916.950 42.600 919.050 43.050 ;
        RECT 934.950 42.600 937.050 43.050 ;
        RECT 892.950 41.400 937.050 42.600 ;
        RECT 892.950 40.950 895.050 41.400 ;
        RECT 916.950 40.950 919.050 41.400 ;
        RECT 934.950 40.950 937.050 41.400 ;
        RECT 22.950 39.600 25.050 40.050 ;
        RECT 145.950 39.600 148.050 40.050 ;
        RECT 175.950 39.600 178.050 40.050 ;
        RECT 22.950 38.400 178.050 39.600 ;
        RECT 22.950 37.950 25.050 38.400 ;
        RECT 145.950 37.950 148.050 38.400 ;
        RECT 175.950 37.950 178.050 38.400 ;
        RECT 274.950 39.600 277.050 40.050 ;
        RECT 310.950 39.600 313.050 40.050 ;
        RECT 535.800 39.600 537.900 40.050 ;
        RECT 274.950 38.400 303.600 39.600 ;
        RECT 274.950 37.950 277.050 38.400 ;
        RECT 302.400 37.050 303.600 38.400 ;
        RECT 310.950 38.400 537.900 39.600 ;
        RECT 310.950 37.950 313.050 38.400 ;
        RECT 535.800 37.950 537.900 38.400 ;
        RECT 538.950 39.600 541.050 40.050 ;
        RECT 577.950 39.600 580.050 40.050 ;
        RECT 538.950 38.400 580.050 39.600 ;
        RECT 538.950 37.950 541.050 38.400 ;
        RECT 577.950 37.950 580.050 38.400 ;
        RECT 616.950 39.600 619.050 40.050 ;
        RECT 664.950 39.600 667.050 40.050 ;
        RECT 673.950 39.600 676.050 40.050 ;
        RECT 616.950 38.400 676.050 39.600 ;
        RECT 616.950 37.950 619.050 38.400 ;
        RECT 664.950 37.950 667.050 38.400 ;
        RECT 673.950 37.950 676.050 38.400 ;
        RECT 778.950 39.600 781.050 40.050 ;
        RECT 808.950 39.600 811.050 40.050 ;
        RECT 823.950 39.600 826.050 40.050 ;
        RECT 853.950 39.600 856.050 40.050 ;
        RECT 973.950 39.600 976.050 40.050 ;
        RECT 778.950 38.400 976.050 39.600 ;
        RECT 778.950 37.950 781.050 38.400 ;
        RECT 808.950 37.950 811.050 38.400 ;
        RECT 823.950 37.950 826.050 38.400 ;
        RECT 853.950 37.950 856.050 38.400 ;
        RECT 973.950 37.950 976.050 38.400 ;
        RECT 31.950 36.600 34.050 37.050 ;
        RECT 97.800 36.600 99.900 37.050 ;
        RECT 31.950 35.400 99.900 36.600 ;
        RECT 31.950 34.950 34.050 35.400 ;
        RECT 97.800 34.950 99.900 35.400 ;
        RECT 100.950 36.600 103.050 37.050 ;
        RECT 136.950 36.600 139.050 37.050 ;
        RECT 283.950 36.600 286.050 37.050 ;
        RECT 100.950 35.400 123.600 36.600 ;
        RECT 100.950 34.950 103.050 35.400 ;
        RECT 85.950 33.600 88.050 34.050 ;
        RECT 94.950 33.600 97.050 34.050 ;
        RECT 85.950 32.400 97.050 33.600 ;
        RECT 122.400 33.600 123.600 35.400 ;
        RECT 136.950 35.400 286.050 36.600 ;
        RECT 136.950 34.950 139.050 35.400 ;
        RECT 283.950 34.950 286.050 35.400 ;
        RECT 301.950 36.600 304.050 37.050 ;
        RECT 331.950 36.600 334.050 37.050 ;
        RECT 589.950 36.600 592.050 37.050 ;
        RECT 301.950 35.400 592.050 36.600 ;
        RECT 301.950 34.950 304.050 35.400 ;
        RECT 331.950 34.950 334.050 35.400 ;
        RECT 589.950 34.950 592.050 35.400 ;
        RECT 634.950 36.600 637.050 37.050 ;
        RECT 706.950 36.600 709.050 37.050 ;
        RECT 715.950 36.600 718.050 37.050 ;
        RECT 634.950 35.400 690.600 36.600 ;
        RECT 634.950 34.950 637.050 35.400 ;
        RECT 689.400 34.050 690.600 35.400 ;
        RECT 706.950 35.400 718.050 36.600 ;
        RECT 706.950 34.950 709.050 35.400 ;
        RECT 715.950 34.950 718.050 35.400 ;
        RECT 865.950 36.600 868.050 37.050 ;
        RECT 871.950 36.600 874.050 37.050 ;
        RECT 865.950 35.400 874.050 36.600 ;
        RECT 865.950 34.950 868.050 35.400 ;
        RECT 871.950 34.950 874.050 35.400 ;
        RECT 898.950 36.600 901.050 37.050 ;
        RECT 913.950 36.600 916.050 37.050 ;
        RECT 898.950 35.400 916.050 36.600 ;
        RECT 898.950 34.950 901.050 35.400 ;
        RECT 913.950 34.950 916.050 35.400 ;
        RECT 934.950 36.600 937.050 37.050 ;
        RECT 988.950 36.600 991.050 37.050 ;
        RECT 934.950 35.400 991.050 36.600 ;
        RECT 934.950 34.950 937.050 35.400 ;
        RECT 988.950 34.950 991.050 35.400 ;
        RECT 196.950 33.600 199.050 34.050 ;
        RECT 220.950 33.600 223.050 34.050 ;
        RECT 122.400 32.400 135.600 33.600 ;
        RECT 85.950 31.950 88.050 32.400 ;
        RECT 94.950 31.950 97.050 32.400 ;
        RECT 61.950 30.600 64.050 31.050 ;
        RECT 79.950 30.600 82.050 31.050 ;
        RECT 61.950 29.400 82.050 30.600 ;
        RECT 134.400 30.600 135.600 32.400 ;
        RECT 152.400 32.400 223.050 33.600 ;
        RECT 152.400 30.600 153.600 32.400 ;
        RECT 196.950 31.950 199.050 32.400 ;
        RECT 220.950 31.950 223.050 32.400 ;
        RECT 250.950 33.600 253.050 34.050 ;
        RECT 256.950 33.600 259.050 34.050 ;
        RECT 250.950 32.400 259.050 33.600 ;
        RECT 250.950 31.950 253.050 32.400 ;
        RECT 256.950 31.950 259.050 32.400 ;
        RECT 349.950 33.600 352.050 34.050 ;
        RECT 367.950 33.600 370.050 34.050 ;
        RECT 349.950 32.400 370.050 33.600 ;
        RECT 349.950 31.950 352.050 32.400 ;
        RECT 367.950 31.950 370.050 32.400 ;
        RECT 457.950 33.600 460.050 34.050 ;
        RECT 484.950 33.600 487.050 34.050 ;
        RECT 613.950 33.600 616.050 34.050 ;
        RECT 457.950 32.400 487.050 33.600 ;
        RECT 457.950 31.950 460.050 32.400 ;
        RECT 484.950 31.950 487.050 32.400 ;
        RECT 548.400 32.400 616.050 33.600 ;
        RECT 548.400 31.050 549.600 32.400 ;
        RECT 613.950 31.950 616.050 32.400 ;
        RECT 658.950 33.600 661.050 34.050 ;
        RECT 664.950 33.600 667.050 34.050 ;
        RECT 682.950 33.600 685.050 34.050 ;
        RECT 658.950 32.400 685.050 33.600 ;
        RECT 658.950 31.950 661.050 32.400 ;
        RECT 664.950 31.950 667.050 32.400 ;
        RECT 682.950 31.950 685.050 32.400 ;
        RECT 688.950 33.600 691.050 34.050 ;
        RECT 724.950 33.600 727.050 34.050 ;
        RECT 733.950 33.600 736.050 34.050 ;
        RECT 688.950 32.400 736.050 33.600 ;
        RECT 688.950 31.950 691.050 32.400 ;
        RECT 724.950 31.950 727.050 32.400 ;
        RECT 733.950 31.950 736.050 32.400 ;
        RECT 748.950 33.600 751.050 34.050 ;
        RECT 781.950 33.600 784.050 34.050 ;
        RECT 748.950 32.400 784.050 33.600 ;
        RECT 748.950 31.950 751.050 32.400 ;
        RECT 781.950 31.950 784.050 32.400 ;
        RECT 805.950 33.600 808.050 34.050 ;
        RECT 826.950 33.600 829.050 34.050 ;
        RECT 805.950 32.400 829.050 33.600 ;
        RECT 805.950 31.950 808.050 32.400 ;
        RECT 826.950 31.950 829.050 32.400 ;
        RECT 832.950 33.600 835.050 34.050 ;
        RECT 931.950 33.600 934.050 34.050 ;
        RECT 832.950 32.400 934.050 33.600 ;
        RECT 832.950 31.950 835.050 32.400 ;
        RECT 931.950 31.950 934.050 32.400 ;
        RECT 134.400 29.400 153.600 30.600 ;
        RECT 226.950 30.600 229.050 31.050 ;
        RECT 259.950 30.600 262.050 31.050 ;
        RECT 271.950 30.600 274.050 31.050 ;
        RECT 346.950 30.600 349.050 31.050 ;
        RECT 226.950 29.400 349.050 30.600 ;
        RECT 61.950 28.950 64.050 29.400 ;
        RECT 79.950 28.950 82.050 29.400 ;
        RECT 226.950 28.950 229.050 29.400 ;
        RECT 259.950 28.950 262.050 29.400 ;
        RECT 271.950 28.950 274.050 29.400 ;
        RECT 346.950 28.950 349.050 29.400 ;
        RECT 535.950 30.600 538.050 31.050 ;
        RECT 547.950 30.600 550.050 31.050 ;
        RECT 535.950 29.400 550.050 30.600 ;
        RECT 535.950 28.950 538.050 29.400 ;
        RECT 547.950 28.950 550.050 29.400 ;
        RECT 562.950 30.600 565.050 31.050 ;
        RECT 580.950 30.600 583.050 31.050 ;
        RECT 598.950 30.600 601.050 31.050 ;
        RECT 562.950 29.400 601.050 30.600 ;
        RECT 562.950 28.950 565.050 29.400 ;
        RECT 580.950 28.950 583.050 29.400 ;
        RECT 598.950 28.950 601.050 29.400 ;
        RECT 610.950 30.600 613.050 31.050 ;
        RECT 619.950 30.600 622.050 31.050 ;
        RECT 610.950 29.400 622.050 30.600 ;
        RECT 610.950 28.950 613.050 29.400 ;
        RECT 619.950 28.950 622.050 29.400 ;
        RECT 646.950 30.600 649.050 31.050 ;
        RECT 652.950 30.600 655.050 31.050 ;
        RECT 646.950 29.400 738.600 30.600 ;
        RECT 646.950 28.950 649.050 29.400 ;
        RECT 652.950 28.950 655.050 29.400 ;
        RECT 737.400 28.200 738.600 29.400 ;
        RECT 55.950 27.600 58.050 28.200 ;
        RECT 73.950 27.600 76.050 28.050 ;
        RECT 55.950 26.400 76.050 27.600 ;
        RECT 55.950 26.100 58.050 26.400 ;
        RECT 73.950 25.950 76.050 26.400 ;
        RECT 94.950 27.750 97.050 28.200 ;
        RECT 106.950 27.750 109.050 28.200 ;
        RECT 94.950 26.550 109.050 27.750 ;
        RECT 94.950 26.100 97.050 26.550 ;
        RECT 106.950 26.100 109.050 26.550 ;
        RECT 112.950 27.600 115.050 28.200 ;
        RECT 130.950 27.600 133.050 28.200 ;
        RECT 154.950 27.600 157.050 28.200 ;
        RECT 112.950 26.400 157.050 27.600 ;
        RECT 112.950 26.100 115.050 26.400 ;
        RECT 130.950 26.100 133.050 26.400 ;
        RECT 154.950 26.100 157.050 26.400 ;
        RECT 160.950 27.600 163.050 28.200 ;
        RECT 202.950 27.600 205.050 28.200 ;
        RECT 211.950 27.600 214.050 28.050 ;
        RECT 244.950 27.600 247.050 28.200 ;
        RECT 286.950 27.600 289.050 28.050 ;
        RECT 160.950 26.400 201.600 27.600 ;
        RECT 160.950 26.100 163.050 26.400 ;
        RECT 200.400 24.600 201.600 26.400 ;
        RECT 202.950 26.400 214.050 27.600 ;
        RECT 202.950 26.100 205.050 26.400 ;
        RECT 211.950 25.950 214.050 26.400 ;
        RECT 218.400 26.400 289.050 27.600 ;
        RECT 218.400 24.600 219.600 26.400 ;
        RECT 244.950 26.100 247.050 26.400 ;
        RECT 286.950 25.950 289.050 26.400 ;
        RECT 295.950 27.600 298.050 28.200 ;
        RECT 310.950 27.600 313.050 28.050 ;
        RECT 316.950 27.600 319.050 28.200 ;
        RECT 295.950 26.400 313.050 27.600 ;
        RECT 295.950 26.100 298.050 26.400 ;
        RECT 310.950 25.950 313.050 26.400 ;
        RECT 314.400 26.400 319.050 27.600 ;
        RECT 200.400 23.400 219.600 24.600 ;
        RECT 46.950 21.450 49.050 21.900 ;
        RECT 52.950 21.450 55.050 21.900 ;
        RECT 46.950 20.250 55.050 21.450 ;
        RECT 46.950 19.800 49.050 20.250 ;
        RECT 52.950 19.800 55.050 20.250 ;
        RECT 97.950 21.450 100.050 21.900 ;
        RECT 103.950 21.450 106.050 21.900 ;
        RECT 97.950 20.250 106.050 21.450 ;
        RECT 97.950 19.800 100.050 20.250 ;
        RECT 103.950 19.800 106.050 20.250 ;
        RECT 109.950 21.450 112.050 21.900 ;
        RECT 121.950 21.450 124.050 21.900 ;
        RECT 109.950 20.250 124.050 21.450 ;
        RECT 109.950 19.800 112.050 20.250 ;
        RECT 121.950 19.800 124.050 20.250 ;
        RECT 145.950 21.450 148.050 21.900 ;
        RECT 157.950 21.450 160.050 21.900 ;
        RECT 145.950 20.250 160.050 21.450 ;
        RECT 145.950 19.800 148.050 20.250 ;
        RECT 157.950 19.800 160.050 20.250 ;
        RECT 187.950 21.450 190.050 21.900 ;
        RECT 193.950 21.450 196.050 21.900 ;
        RECT 187.950 20.250 196.050 21.450 ;
        RECT 187.950 19.800 190.050 20.250 ;
        RECT 193.950 19.800 196.050 20.250 ;
        RECT 211.950 21.450 214.050 21.900 ;
        RECT 247.950 21.450 250.050 21.900 ;
        RECT 211.950 20.250 250.050 21.450 ;
        RECT 211.950 19.800 214.050 20.250 ;
        RECT 247.950 19.800 250.050 20.250 ;
        RECT 259.950 21.450 262.050 21.900 ;
        RECT 271.950 21.450 274.050 21.900 ;
        RECT 259.950 20.250 274.050 21.450 ;
        RECT 259.950 19.800 262.050 20.250 ;
        RECT 271.950 19.800 274.050 20.250 ;
        RECT 277.950 21.450 280.050 21.900 ;
        RECT 283.950 21.600 286.050 21.900 ;
        RECT 292.950 21.600 295.050 21.900 ;
        RECT 283.950 21.450 295.050 21.600 ;
        RECT 277.950 20.400 295.050 21.450 ;
        RECT 277.950 20.250 286.050 20.400 ;
        RECT 277.950 19.800 280.050 20.250 ;
        RECT 283.950 19.800 286.050 20.250 ;
        RECT 292.950 19.800 295.050 20.400 ;
        RECT 298.950 21.600 301.050 21.900 ;
        RECT 314.400 21.600 315.600 26.400 ;
        RECT 316.950 26.100 319.050 26.400 ;
        RECT 352.950 27.600 355.050 28.200 ;
        RECT 364.950 27.600 367.050 28.050 ;
        RECT 352.950 26.400 367.050 27.600 ;
        RECT 352.950 26.100 355.050 26.400 ;
        RECT 364.950 25.950 367.050 26.400 ;
        RECT 394.950 27.600 397.050 28.200 ;
        RECT 400.950 27.600 403.050 28.050 ;
        RECT 394.950 26.400 403.050 27.600 ;
        RECT 394.950 26.100 397.050 26.400 ;
        RECT 400.950 25.950 403.050 26.400 ;
        RECT 463.950 27.750 466.050 28.200 ;
        RECT 469.950 27.750 472.050 28.200 ;
        RECT 463.950 26.550 472.050 27.750 ;
        RECT 463.950 26.100 466.050 26.550 ;
        RECT 469.950 26.100 472.050 26.550 ;
        RECT 493.950 27.600 496.050 28.050 ;
        RECT 502.950 27.600 505.050 28.200 ;
        RECT 493.950 26.400 505.050 27.600 ;
        RECT 493.950 25.950 496.050 26.400 ;
        RECT 502.950 26.100 505.050 26.400 ;
        RECT 508.950 27.600 511.050 28.200 ;
        RECT 532.950 27.600 535.050 28.200 ;
        RECT 508.950 26.400 535.050 27.600 ;
        RECT 508.950 26.100 511.050 26.400 ;
        RECT 532.950 26.100 535.050 26.400 ;
        RECT 544.950 27.600 547.050 28.050 ;
        RECT 556.950 27.600 559.050 28.200 ;
        RECT 604.950 27.600 607.050 28.200 ;
        RECT 615.000 27.600 619.050 28.050 ;
        RECT 544.950 26.400 559.050 27.600 ;
        RECT 533.400 24.600 534.600 26.100 ;
        RECT 544.950 25.950 547.050 26.400 ;
        RECT 556.950 26.100 559.050 26.400 ;
        RECT 560.400 26.400 607.050 27.600 ;
        RECT 560.400 24.600 561.600 26.400 ;
        RECT 604.950 26.100 607.050 26.400 ;
        RECT 533.400 23.400 561.600 24.600 ;
        RECT 614.400 25.950 619.050 27.600 ;
        RECT 622.950 27.600 625.050 28.050 ;
        RECT 628.950 27.600 631.050 28.200 ;
        RECT 622.950 26.400 631.050 27.600 ;
        RECT 622.950 25.950 625.050 26.400 ;
        RECT 628.950 26.100 631.050 26.400 ;
        RECT 667.950 27.600 670.050 28.050 ;
        RECT 679.950 27.600 682.050 28.200 ;
        RECT 691.950 27.600 694.050 28.050 ;
        RECT 667.950 26.400 678.600 27.600 ;
        RECT 667.950 25.950 670.050 26.400 ;
        RECT 614.400 21.900 615.600 25.950 ;
        RECT 619.950 24.600 622.050 25.050 ;
        RECT 677.400 24.600 678.600 26.400 ;
        RECT 679.950 26.400 694.050 27.600 ;
        RECT 679.950 26.100 682.050 26.400 ;
        RECT 691.950 25.950 694.050 26.400 ;
        RECT 709.950 24.600 712.050 28.050 ;
        RECT 736.950 27.750 739.050 28.200 ;
        RECT 742.950 27.750 745.050 28.200 ;
        RECT 736.950 26.550 745.050 27.750 ;
        RECT 736.950 26.100 739.050 26.550 ;
        RECT 742.950 26.100 745.050 26.550 ;
        RECT 820.950 27.600 823.050 28.200 ;
        RECT 844.950 27.600 847.050 28.200 ;
        RECT 886.950 27.600 889.050 28.200 ;
        RECT 820.950 26.400 889.050 27.600 ;
        RECT 820.950 26.100 823.050 26.400 ;
        RECT 844.950 26.100 847.050 26.400 ;
        RECT 886.950 26.100 889.050 26.400 ;
        RECT 937.950 27.600 940.050 28.200 ;
        RECT 964.950 27.600 967.050 28.200 ;
        RECT 991.950 27.750 994.050 28.200 ;
        RECT 1009.950 27.750 1012.050 28.200 ;
        RECT 991.950 27.600 1012.050 27.750 ;
        RECT 937.950 26.550 1012.050 27.600 ;
        RECT 937.950 26.400 994.050 26.550 ;
        RECT 937.950 26.100 940.050 26.400 ;
        RECT 964.950 26.100 967.050 26.400 ;
        RECT 991.950 26.100 994.050 26.400 ;
        RECT 1009.950 26.100 1012.050 26.550 ;
        RECT 619.950 23.400 663.600 24.600 ;
        RECT 677.400 24.000 712.050 24.600 ;
        RECT 677.400 23.400 711.600 24.000 ;
        RECT 619.950 22.950 622.050 23.400 ;
        RECT 662.400 21.900 663.600 23.400 ;
        RECT 698.400 21.900 699.600 23.400 ;
        RECT 298.950 20.400 315.600 21.600 ;
        RECT 343.950 21.450 346.050 21.900 ;
        RECT 358.950 21.450 361.050 21.900 ;
        RECT 298.950 19.800 301.050 20.400 ;
        RECT 343.950 20.250 361.050 21.450 ;
        RECT 343.950 19.800 346.050 20.250 ;
        RECT 358.950 19.800 361.050 20.250 ;
        RECT 397.950 21.450 400.050 21.900 ;
        RECT 454.950 21.450 457.050 21.900 ;
        RECT 397.950 20.250 457.050 21.450 ;
        RECT 397.950 19.800 400.050 20.250 ;
        RECT 454.950 19.800 457.050 20.250 ;
        RECT 511.950 21.600 514.050 21.900 ;
        RECT 535.950 21.600 538.050 21.900 ;
        RECT 511.950 20.400 538.050 21.600 ;
        RECT 511.950 19.800 514.050 20.400 ;
        RECT 535.950 19.800 538.050 20.400 ;
        RECT 547.950 21.450 550.050 21.900 ;
        RECT 553.950 21.450 556.050 21.900 ;
        RECT 547.950 20.250 556.050 21.450 ;
        RECT 547.950 19.800 550.050 20.250 ;
        RECT 553.950 19.800 556.050 20.250 ;
        RECT 559.950 21.600 562.050 21.900 ;
        RECT 574.950 21.600 577.050 21.900 ;
        RECT 559.950 21.450 577.050 21.600 ;
        RECT 583.950 21.450 586.050 21.900 ;
        RECT 559.950 20.400 586.050 21.450 ;
        RECT 559.950 19.800 562.050 20.400 ;
        RECT 574.950 20.250 586.050 20.400 ;
        RECT 574.950 19.800 577.050 20.250 ;
        RECT 583.950 19.800 586.050 20.250 ;
        RECT 613.950 19.800 616.050 21.900 ;
        RECT 631.950 21.600 634.050 21.900 ;
        RECT 655.950 21.600 658.050 21.900 ;
        RECT 631.950 21.000 660.600 21.600 ;
        RECT 661.950 21.450 664.050 21.900 ;
        RECT 670.950 21.450 673.050 21.900 ;
        RECT 631.950 20.400 661.050 21.000 ;
        RECT 631.950 19.800 634.050 20.400 ;
        RECT 655.950 19.800 658.050 20.400 ;
        RECT 73.950 18.600 76.050 19.050 ;
        RECT 91.950 18.600 94.050 19.050 ;
        RECT 73.950 17.400 94.050 18.600 ;
        RECT 73.950 16.950 76.050 17.400 ;
        RECT 91.950 16.950 94.050 17.400 ;
        RECT 127.950 18.600 130.050 19.050 ;
        RECT 146.400 18.600 147.600 19.800 ;
        RECT 127.950 17.400 147.600 18.600 ;
        RECT 178.950 18.600 181.050 19.050 ;
        RECT 199.950 18.600 202.050 19.050 ;
        RECT 205.950 18.600 208.050 19.050 ;
        RECT 178.950 17.400 208.050 18.600 ;
        RECT 127.950 16.950 130.050 17.400 ;
        RECT 178.950 16.950 181.050 17.400 ;
        RECT 199.950 16.950 202.050 17.400 ;
        RECT 205.950 16.950 208.050 17.400 ;
        RECT 301.950 18.600 304.050 19.050 ;
        RECT 319.950 18.600 322.050 19.050 ;
        RECT 301.950 17.400 322.050 18.600 ;
        RECT 301.950 16.950 304.050 17.400 ;
        RECT 319.950 16.950 322.050 17.400 ;
        RECT 460.950 18.600 463.050 19.050 ;
        RECT 493.950 18.600 496.050 19.050 ;
        RECT 460.950 17.400 496.050 18.600 ;
        RECT 460.950 16.950 463.050 17.400 ;
        RECT 493.950 16.950 496.050 17.400 ;
        RECT 535.950 18.600 538.050 19.050 ;
        RECT 544.950 18.600 547.050 19.050 ;
        RECT 535.950 17.400 547.050 18.600 ;
        RECT 535.950 16.950 538.050 17.400 ;
        RECT 544.950 16.950 547.050 17.400 ;
        RECT 658.950 16.950 661.050 20.400 ;
        RECT 661.950 20.250 673.050 21.450 ;
        RECT 661.950 19.800 664.050 20.250 ;
        RECT 670.950 19.800 673.050 20.250 ;
        RECT 697.950 19.800 700.050 21.900 ;
        RECT 703.950 21.600 706.050 21.900 ;
        RECT 721.950 21.600 724.050 21.900 ;
        RECT 703.950 20.400 724.050 21.600 ;
        RECT 703.950 19.800 706.050 20.400 ;
        RECT 721.950 19.800 724.050 20.400 ;
        RECT 733.950 21.450 736.050 21.900 ;
        RECT 751.950 21.450 754.050 21.900 ;
        RECT 733.950 20.250 754.050 21.450 ;
        RECT 733.950 19.800 736.050 20.250 ;
        RECT 751.950 19.800 754.050 20.250 ;
        RECT 772.950 21.600 775.050 21.900 ;
        RECT 790.950 21.600 793.050 21.900 ;
        RECT 772.950 20.400 793.050 21.600 ;
        RECT 772.950 19.800 775.050 20.400 ;
        RECT 790.950 19.800 793.050 20.400 ;
        RECT 796.950 21.450 799.050 21.900 ;
        RECT 805.800 21.450 807.900 21.900 ;
        RECT 796.950 20.250 807.900 21.450 ;
        RECT 796.950 19.800 799.050 20.250 ;
        RECT 805.800 19.800 807.900 20.250 ;
        RECT 808.950 21.450 811.050 21.900 ;
        RECT 817.950 21.450 820.050 21.900 ;
        RECT 808.950 20.250 820.050 21.450 ;
        RECT 808.950 19.800 811.050 20.250 ;
        RECT 817.950 19.800 820.050 20.250 ;
        RECT 823.950 21.600 826.050 21.900 ;
        RECT 832.950 21.600 835.050 21.900 ;
        RECT 823.950 21.450 835.050 21.600 ;
        RECT 841.950 21.450 844.050 21.900 ;
        RECT 823.950 20.400 844.050 21.450 ;
        RECT 823.950 19.800 826.050 20.400 ;
        RECT 832.950 20.250 844.050 20.400 ;
        RECT 832.950 19.800 835.050 20.250 ;
        RECT 841.950 19.800 844.050 20.250 ;
        RECT 865.950 21.600 868.050 21.900 ;
        RECT 871.950 21.600 874.050 22.050 ;
        RECT 865.950 20.400 874.050 21.600 ;
        RECT 865.950 19.800 868.050 20.400 ;
        RECT 871.950 19.950 874.050 20.400 ;
        RECT 889.950 21.450 892.050 21.900 ;
        RECT 898.950 21.600 901.050 22.050 ;
        RECT 904.800 21.600 906.900 22.050 ;
        RECT 898.950 21.450 906.900 21.600 ;
        RECT 889.950 20.400 906.900 21.450 ;
        RECT 889.950 20.250 901.050 20.400 ;
        RECT 889.950 19.800 892.050 20.250 ;
        RECT 898.950 19.950 901.050 20.250 ;
        RECT 904.800 19.950 906.900 20.400 ;
        RECT 907.950 21.600 910.050 21.900 ;
        RECT 934.950 21.600 937.050 21.900 ;
        RECT 907.950 20.400 937.050 21.600 ;
        RECT 907.950 19.800 910.050 20.400 ;
        RECT 934.950 19.800 937.050 20.400 ;
        RECT 949.950 21.450 952.050 21.900 ;
        RECT 961.950 21.600 964.050 21.900 ;
        RECT 994.950 21.600 997.050 21.900 ;
        RECT 961.950 21.450 997.050 21.600 ;
        RECT 949.950 20.400 997.050 21.450 ;
        RECT 949.950 20.250 964.050 20.400 ;
        RECT 949.950 19.800 952.050 20.250 ;
        RECT 961.950 19.800 964.050 20.250 ;
        RECT 994.950 19.800 997.050 20.400 ;
        RECT 745.950 18.600 748.050 19.050 ;
        RECT 713.400 17.400 748.050 18.600 ;
        RECT 34.950 15.600 37.050 16.050 ;
        RECT 58.950 15.600 61.050 16.050 ;
        RECT 34.950 14.400 61.050 15.600 ;
        RECT 34.950 13.950 37.050 14.400 ;
        RECT 58.950 13.950 61.050 14.400 ;
        RECT 109.950 15.600 112.050 16.050 ;
        RECT 133.950 15.600 136.050 16.050 ;
        RECT 151.950 15.600 154.050 16.050 ;
        RECT 109.950 14.400 154.050 15.600 ;
        RECT 109.950 13.950 112.050 14.400 ;
        RECT 133.950 13.950 136.050 14.400 ;
        RECT 151.950 13.950 154.050 14.400 ;
        RECT 286.950 15.600 289.050 16.050 ;
        RECT 298.950 15.600 301.050 16.050 ;
        RECT 286.950 14.400 301.050 15.600 ;
        RECT 320.400 15.600 321.600 16.950 ;
        RECT 349.950 15.600 352.050 16.050 ;
        RECT 320.400 14.400 352.050 15.600 ;
        RECT 286.950 13.950 289.050 14.400 ;
        RECT 298.950 13.950 301.050 14.400 ;
        RECT 349.950 13.950 352.050 14.400 ;
        RECT 364.950 15.600 367.050 16.050 ;
        RECT 589.950 15.600 592.050 16.050 ;
        RECT 607.950 15.600 610.050 16.050 ;
        RECT 364.950 14.400 610.050 15.600 ;
        RECT 364.950 13.950 367.050 14.400 ;
        RECT 589.950 13.950 592.050 14.400 ;
        RECT 607.950 13.950 610.050 14.400 ;
        RECT 691.950 15.600 694.050 16.050 ;
        RECT 713.400 15.600 714.600 17.400 ;
        RECT 745.950 16.950 748.050 17.400 ;
        RECT 691.950 14.400 714.600 15.600 ;
        RECT 715.950 15.600 718.050 16.050 ;
        RECT 898.950 15.600 901.050 16.050 ;
        RECT 715.950 14.400 901.050 15.600 ;
        RECT 691.950 13.950 694.050 14.400 ;
        RECT 715.950 13.950 718.050 14.400 ;
        RECT 898.950 13.950 901.050 14.400 ;
        RECT 904.950 15.600 907.050 16.050 ;
        RECT 913.950 15.600 916.050 16.050 ;
        RECT 904.950 14.400 916.050 15.600 ;
        RECT 904.950 13.950 907.050 14.400 ;
        RECT 913.950 13.950 916.050 14.400 ;
        RECT 13.950 12.600 16.050 13.050 ;
        RECT 88.950 12.600 91.050 13.050 ;
        RECT 94.950 12.600 97.050 13.050 ;
        RECT 13.950 11.400 97.050 12.600 ;
        RECT 13.950 10.950 16.050 11.400 ;
        RECT 88.950 10.950 91.050 11.400 ;
        RECT 94.950 10.950 97.050 11.400 ;
        RECT 247.950 12.600 250.050 13.050 ;
        RECT 295.950 12.600 298.050 13.050 ;
        RECT 247.950 11.400 298.050 12.600 ;
        RECT 247.950 10.950 250.050 11.400 ;
        RECT 295.950 10.950 298.050 11.400 ;
        RECT 433.950 12.600 436.050 13.050 ;
        RECT 481.950 12.600 484.050 13.050 ;
        RECT 433.950 11.400 484.050 12.600 ;
        RECT 433.950 10.950 436.050 11.400 ;
        RECT 481.950 10.950 484.050 11.400 ;
        RECT 505.950 12.600 508.050 13.050 ;
        RECT 529.950 12.600 532.050 13.050 ;
        RECT 646.950 12.600 649.050 13.050 ;
        RECT 505.950 11.400 649.050 12.600 ;
        RECT 505.950 10.950 508.050 11.400 ;
        RECT 529.950 10.950 532.050 11.400 ;
        RECT 646.950 10.950 649.050 11.400 ;
        RECT 469.950 6.600 472.050 7.050 ;
        RECT 622.950 6.600 625.050 7.050 ;
        RECT 469.950 5.400 625.050 6.600 ;
        RECT 469.950 4.950 472.050 5.400 ;
        RECT 622.950 4.950 625.050 5.400 ;
        RECT 781.950 6.600 784.050 7.050 ;
        RECT 883.950 6.600 886.050 7.050 ;
        RECT 967.950 6.600 970.050 7.050 ;
        RECT 988.950 6.600 991.050 7.050 ;
        RECT 781.950 5.400 991.050 6.600 ;
        RECT 781.950 4.950 784.050 5.400 ;
        RECT 883.950 4.950 886.050 5.400 ;
        RECT 967.950 4.950 970.050 5.400 ;
        RECT 988.950 4.950 991.050 5.400 ;
  END
END fir_pe
END LIBRARY


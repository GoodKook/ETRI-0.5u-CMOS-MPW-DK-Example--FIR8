/* Verilog module written by vlog2Verilog (qflow) */

module fir_pe(
    input [7:0] Cin,
    input [7:0] Xin,
    output [7:0] Xout,
    input [15:0] Yin,
    output [15:0] Yout,
    input clk
);

wire vdd = 1'b1;
wire gnd = 1'b0;

wire [15:0] y ;
wire _588_ ;
wire _168_ ;
wire _60_ ;
wire _397_ ;
wire _703_ ;
wire _19_ ;
wire _512_ ;
wire _741_ ;
wire _321_ ;
wire _57_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _415_ ;
wire _95_ ;
wire _644_ ;
wire _224_ ;
wire _453_ ;
wire _509_ ;
wire _682_ ;
wire _262_ ;
wire _738_ ;
wire _318_ ;
wire _491_ ;
wire _547_ ;
wire _127_ ;
wire _356_ ;
wire _585_ ;
wire _165_ ;
wire _394_ ;
wire _679_ ;
wire _259_ ;
wire _488_ ;
wire _700_ ;
wire _297_ ;
wire _16_ ;
wire _54_ ;
wire _603_ ;
wire _412_ ;
wire _92_ ;
wire _641_ ;
wire _221_ ;
wire _450_ ;
wire _506_ ;
wire _735_ ;
wire _315_ ;
wire _544_ ;
wire _124_ ;
wire _353_ ;
wire _409_ ;
wire _89_ ;
wire _582_ ;
wire _162_ ;
wire _638_ ;
wire _218_ ;
wire _391_ ;
wire _447_ ;
wire _676_ ;
wire _256_ ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire _388_ ;
wire _600_ ;
wire _197_ ;
wire _7_ ;
wire _503_ ;
wire _732_ ;
wire _312_ ;
wire _48_ ;
wire _541_ ;
wire _121_ ;
wire _350_ ;
wire _406_ ;
wire _86_ ;
wire _635_ ;
wire _215_ ;
wire _444_ ;
wire _673_ ;
wire _253_ ;
wire _729_ ;
wire _309_ ;
wire _482_ ;
wire _538_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _347_ ;
wire _576_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire _479_ ;
wire _288_ ;
wire _4_ ;
wire _500_ ;
wire _45_ ;
wire _403_ ;
wire _83_ ;
wire _632_ ;
wire _212_ ;
wire _441_ ;
wire _670_ ;
wire _250_ ;
wire _726_ ;
wire _306_ ;
wire _535_ ;
wire _115_ ;
wire _344_ ;
wire _573_ ;
wire _153_ ;
wire _629_ ;
wire _209_ ;
wire Xin_5_bF$buf0 ;
wire Xin_5_bF$buf1 ;
wire Xin_5_bF$buf2 ;
wire Xin_5_bF$buf3 ;
wire _382_ ;
wire _438_ ;
wire _191_ ;
wire _667_ ;
wire _247_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire _285_ ;
wire _1_ ;
wire _42_ ;
wire _379_ ;
wire _188_ ;
wire _400_ ;
wire _80_ ;
wire _723_ ;
wire _303_ ;
wire _39_ ;
wire _532_ ;
wire _112_ ;
wire _341_ ;
wire clk ;
wire _77_ ;
wire _570_ ;
wire _150_ ;
wire _626_ ;
wire _206_ ;
wire _435_ ;
wire _664_ ;
wire _244_ ;
wire _473_ ;
wire _529_ ;
wire _109_ ;
wire _282_ ;
wire _338_ ;
wire _567_ ;
wire _147_ ;
wire _376_ ;
wire _185_ ;
wire _699_ ;
wire _279_ ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire _74_ ;
wire _623_ ;
wire _203_ ;
wire _432_ ;
wire _661_ ;
wire _241_ ;
wire _717_ ;
wire _470_ ;
wire _526_ ;
wire _106_ ;
wire [15:0] _755_ ;
wire _335_ ;
wire _564_ ;
wire _144_ ;
wire _373_ ;
wire _429_ ;
wire _182_ ;
wire _658_ ;
wire _238_ ;
wire _467_ ;
wire _696_ ;
wire _276_ ;
wire _33_ ;
wire _599_ ;
wire _179_ ;
wire _71_ ;
wire _620_ ;
wire _200_ ;
wire _714_ ;
wire _523_ ;
wire _103_ ;
wire [15:0] _752_ ;
wire _332_ ;
wire _68_ ;
wire _561_ ;
wire _141_ ;
wire _617_ ;
wire _370_ ;
wire _426_ ;
wire _655_ ;
wire _235_ ;
wire _464_ ;
wire _693_ ;
wire _273_ ;
wire [15:0] _749_ ;
wire _329_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _367_ ;
wire _596_ ;
wire _176_ ;
wire _499_ ;
wire _711_ ;
wire _27_ ;
wire _520_ ;
wire _100_ ;
wire _65_ ;
wire _614_ ;
wire _423_ ;
wire _652_ ;
wire _232_ ;
wire _708_ ;
wire _461_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _746_ ;
wire _326_ ;
wire _555_ ;
wire _135_ ;
wire _364_ ;
wire _593_ ;
wire _173_ ;
wire _649_ ;
wire _229_ ;
wire _458_ ;
wire _687_ ;
wire _267_ ;
wire _496_ ;
wire _24_ ;
wire _62_ ;
wire _399_ ;
wire _611_ ;
wire _420_ ;
wire _705_ ;
wire _514_ ;
wire _743_ ;
wire _323_ ;
wire _59_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _361_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _646_ ;
wire _226_ ;
wire _455_ ;
wire _684_ ;
wire _264_ ;
wire _493_ ;
wire _549_ ;
wire _129_ ;
wire _21_ ;
wire _358_ ;
wire _587_ ;
wire _167_ ;
wire _396_ ;
wire _702_ ;
wire _299_ ;
wire _18_ ;
wire _511_ ;
wire _740_ ;
wire _320_ ;
wire _56_ ;
wire _605_ ;
wire _414_ ;
wire _94_ ;
wire _643_ ;
wire _223_ ;
wire _452_ ;
wire _508_ ;
wire _681_ ;
wire _261_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _546_ ;
wire _126_ ;
wire _355_ ;
wire _584_ ;
wire _164_ ;
wire _393_ ;
wire _449_ ;
wire _678_ ;
wire _258_ ;
wire _487_ ;
wire _296_ ;
wire _15_ ;
wire _53_ ;
wire _602_ ;
wire _199_ ;
wire _411_ ;
wire _91_ ;
wire _640_ ;
wire _220_ ;
wire _9_ ;
wire _505_ ;
wire _734_ ;
wire _314_ ;
wire _543_ ;
wire _123_ ;
wire _352_ ;
wire _408_ ;
wire _88_ ;
wire _581_ ;
wire _161_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _446_ ;
wire [15:0] Yin ;
wire _675_ ;
wire _255_ ;
wire _484_ ;
wire _293_ ;
wire _12_ ;
wire _349_ ;
wire _578_ ;
wire _158_ ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire _6_ ;
wire _502_ ;
wire _731_ ;
wire _311_ ;
wire _47_ ;
wire _540_ ;
wire _120_ ;
wire _405_ ;
wire _85_ ;
wire _634_ ;
wire _214_ ;
wire _443_ ;
wire _672_ ;
wire _252_ ;
wire _728_ ;
wire _308_ ;
wire _481_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _346_ ;
wire _575_ ;
wire _155_ ;
wire _384_ ;
wire _193_ ;
wire _669_ ;
wire _249_ ;
wire _478_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _402_ ;
wire _82_ ;
wire _631_ ;
wire _211_ ;
wire _440_ ;
wire _725_ ;
wire _305_ ;
wire _534_ ;
wire _114_ ;
wire _343_ ;
wire _79_ ;
wire _572_ ;
wire _152_ ;
wire _628_ ;
wire _208_ ;
wire _381_ ;
wire _437_ ;
wire _190_ ;
wire _666_ ;
wire _246_ ;
wire _475_ ;
wire _284_ ;
wire _0_ ;
wire _569_ ;
wire _149_ ;
wire _41_ ;
wire _378_ ;
wire _187_ ;
wire [15:0] Yout ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _531_ ;
wire _111_ ;
wire _340_ ;
wire _76_ ;
wire _625_ ;
wire _205_ ;
wire _434_ ;
wire _663_ ;
wire _243_ ;
wire _719_ ;
wire _472_ ;
wire _528_ ;
wire _108_ ;
wire _281_ ;
wire _337_ ;
wire _566_ ;
wire _146_ ;
wire _375_ ;
wire _184_ ;
wire _469_ ;
wire _698_ ;
wire _278_ ;
wire _35_ ;
wire [7:0] Xout ;
wire _73_ ;
wire _622_ ;
wire _202_ ;
wire _431_ ;
wire _660_ ;
wire _240_ ;
wire _716_ ;
wire _525_ ;
wire _105_ ;
wire [7:0] _754_ ;
wire _334_ ;
wire _563_ ;
wire _143_ ;
wire _619_ ;
wire _372_ ;
wire _428_ ;
wire _181_ ;
wire _657_ ;
wire _237_ ;
wire _466_ ;
wire _695_ ;
wire _275_ ;
wire _32_ ;
wire _369_ ;
wire _598_ ;
wire _178_ ;
wire _70_ ;
wire _713_ ;
wire _29_ ;
wire _522_ ;
wire _102_ ;
wire [15:0] _751_ ;
wire _331_ ;
wire _67_ ;
wire _560_ ;
wire _140_ ;
wire _616_ ;
wire _425_ ;
wire _654_ ;
wire _234_ ;
wire _463_ ;
wire _519_ ;
wire _692_ ;
wire _272_ ;
wire [15:0] _748_ ;
wire _328_ ;
wire _557_ ;
wire _137_ ;
wire _366_ ;
wire _595_ ;
wire _175_ ;
wire _689_ ;
wire _269_ ;
wire _498_ ;
wire _710_ ;
wire _26_ ;
wire Cin_0_bF$buf0 ;
wire Cin_0_bF$buf1 ;
wire Cin_0_bF$buf2 ;
wire Cin_0_bF$buf3 ;
wire _64_ ;
wire _613_ ;
wire _422_ ;
wire _651_ ;
wire _231_ ;
wire _707_ ;
wire _460_ ;
wire _516_ ;
wire _745_ ;
wire _325_ ;
wire _554_ ;
wire _134_ ;
wire _363_ ;
wire _419_ ;
wire _99_ ;
wire _592_ ;
wire _172_ ;
wire _648_ ;
wire _228_ ;
wire _457_ ;
wire _686_ ;
wire _266_ ;
wire _495_ ;
wire _23_ ;
wire _589_ ;
wire _169_ ;
wire _61_ ;
wire _398_ ;
wire _610_ ;
wire _704_ ;
wire _513_ ;
wire _742_ ;
wire _322_ ;
wire _58_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _360_ ;
wire _416_ ;
wire _96_ ;
wire [7:0] Cin ;
wire _645_ ;
wire _225_ ;
wire _454_ ;
wire _683_ ;
wire _263_ ;
wire _739_ ;
wire _319_ ;
wire _492_ ;
wire _548_ ;
wire _128_ ;
wire _20_ ;
wire _357_ ;
wire _586_ ;
wire _166_ ;
wire _395_ ;
wire _489_ ;
wire _701_ ;
wire _298_ ;
wire _17_ ;
wire _510_ ;
wire _55_ ;
wire _604_ ;
wire _413_ ;
wire _93_ ;
wire _642_ ;
wire _222_ ;
wire _451_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _736_ ;
wire _316_ ;
wire _545_ ;
wire _125_ ;
wire _354_ ;
wire _583_ ;
wire _163_ ;
wire _639_ ;
wire _219_ ;
wire _392_ ;
wire _448_ ;
wire _677_ ;
wire _257_ ;
wire _486_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _601_ ;
wire _198_ ;
wire _410_ ;
wire _90_ ;
wire _8_ ;
wire _504_ ;
wire _733_ ;
wire _313_ ;
wire _49_ ;
wire _542_ ;
wire _122_ ;
wire _351_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _636_ ;
wire _216_ ;
wire _445_ ;
wire _674_ ;
wire _254_ ;
wire _483_ ;
wire _539_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _348_ ;
wire _577_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire _289_ ;
wire _5_ ;
wire _501_ ;
wire _730_ ;
wire _310_ ;
wire _46_ ;
wire _404_ ;
wire _84_ ;
wire _633_ ;
wire _213_ ;
wire _442_ ;
wire _671_ ;
wire _251_ ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire _536_ ;
wire _116_ ;
wire _345_ ;
wire _574_ ;
wire _154_ ;
wire _383_ ;
wire _439_ ;
wire _192_ ;
wire _668_ ;
wire _248_ ;
wire _477_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire _189_ ;
wire _401_ ;
wire _81_ ;
wire _630_ ;
wire _210_ ;
wire _724_ ;
wire _304_ ;
wire _533_ ;
wire _113_ ;
wire _342_ ;
wire _78_ ;
wire _571_ ;
wire _151_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _436_ ;
wire [7:0] Xin ;
wire _665_ ;
wire _245_ ;
wire _474_ ;
wire _283_ ;
wire _339_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire _377_ ;
wire _186_ ;
wire _721_ ;
wire _301_ ;
wire _37_ ;
wire _530_ ;
wire _110_ ;
wire _75_ ;
wire _624_ ;
wire _204_ ;
wire _433_ ;
wire _662_ ;
wire _242_ ;
wire _718_ ;
wire _471_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _336_ ;
wire _565_ ;
wire _145_ ;
wire _374_ ;
wire _183_ ;
wire _659_ ;
wire _239_ ;
wire _468_ ;
wire _697_ ;
wire _277_ ;
wire _34_ ;
wire _72_ ;
wire _621_ ;
wire _201_ ;
wire _430_ ;
wire _715_ ;
wire _524_ ;
wire _104_ ;
wire [15:0] _753_ ;
wire _333_ ;
wire _69_ ;
wire _562_ ;
wire _142_ ;
wire _618_ ;
wire _371_ ;
wire _427_ ;
wire _180_ ;
wire _656_ ;
wire _236_ ;
wire _465_ ;
wire _694_ ;
wire _274_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _368_ ;
wire _597_ ;
wire _177_ ;
wire _712_ ;
wire _28_ ;
wire _521_ ;
wire _101_ ;
wire [15:0] _750_ ;
wire _330_ ;
wire _66_ ;
wire _615_ ;
wire _424_ ;
wire _653_ ;
wire _233_ ;
wire _709_ ;
wire _462_ ;
wire _518_ ;
wire _691_ ;
wire _271_ ;
wire _747_ ;
wire _327_ ;
wire _556_ ;
wire _136_ ;
wire _365_ ;
wire _594_ ;
wire _174_ ;
wire _459_ ;
wire _688_ ;
wire _268_ ;
wire _497_ ;
wire Xin_3_bF$buf0 ;
wire Xin_3_bF$buf1 ;
wire Xin_3_bF$buf2 ;
wire Xin_3_bF$buf3 ;
wire _25_ ;
wire _63_ ;
wire _612_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire _706_ ;
wire _515_ ;
wire _744_ ;
wire _324_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _362_ ;
wire _418_ ;
wire _98_ ;
wire _591_ ;
wire _171_ ;
wire _647_ ;
wire _227_ ;
wire _456_ ;
wire _685_ ;
wire _265_ ;
wire _494_ ;
wire _22_ ;
wire _359_ ;

BUFX2 BUFX2_insert17 (
    .A(Xin[5]),
    .Y(Xin_5_bF$buf0)
);

BUFX2 BUFX2_insert16 (
    .A(Xin[5]),
    .Y(Xin_5_bF$buf1)
);

BUFX2 BUFX2_insert15 (
    .A(Xin[5]),
    .Y(Xin_5_bF$buf2)
);

BUFX2 BUFX2_insert14 (
    .A(Xin[5]),
    .Y(Xin_5_bF$buf3)
);

BUFX2 BUFX2_insert13 (
    .A(Xin[3]),
    .Y(Xin_3_bF$buf0)
);

BUFX2 BUFX2_insert12 (
    .A(Xin[3]),
    .Y(Xin_3_bF$buf1)
);

BUFX2 BUFX2_insert11 (
    .A(Xin[3]),
    .Y(Xin_3_bF$buf2)
);

BUFX2 BUFX2_insert10 (
    .A(Xin[3]),
    .Y(Xin_3_bF$buf3)
);

BUFX2 BUFX2_insert9 (
    .A(Cin[0]),
    .Y(Cin_0_bF$buf0)
);

BUFX2 BUFX2_insert8 (
    .A(Cin[0]),
    .Y(Cin_0_bF$buf1)
);

BUFX2 BUFX2_insert7 (
    .A(Cin[0]),
    .Y(Cin_0_bF$buf2)
);

BUFX2 BUFX2_insert6 (
    .A(Cin[0]),
    .Y(Cin_0_bF$buf3)
);

CLKBUF1 CLKBUF1_insert5 (
    .A(clk),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert4 (
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert3 (
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert2 (
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert1 (
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert0 (
    .A(clk),
    .Y(clk_bF$buf5)
);

AOI21X1 _1000_ (
    .A(_190_),
    .B(_189_),
    .C(_188_),
    .Y(_191_)
);

OAI21X1 _1001_ (
    .A(_191_),
    .B(_187_),
    .C(_139_),
    .Y(_192_)
);

INVX1 _1002_ (
    .A(_116_),
    .Y(_193_)
);

AOI21X1 _1003_ (
    .A(_81_),
    .B(_120_),
    .C(_193_),
    .Y(_194_)
);

NAND3X1 _1004_ (
    .A(_188_),
    .B(_189_),
    .C(_190_),
    .Y(_195_)
);

NAND3X1 _1005_ (
    .A(_144_),
    .B(_180_),
    .C(_186_),
    .Y(_196_)
);

NAND3X1 _1006_ (
    .A(_195_),
    .B(_196_),
    .C(_194_),
    .Y(_197_)
);

AOI21X1 _1007_ (
    .A(_197_),
    .B(_192_),
    .C(_137_),
    .Y(_198_)
);

INVX1 _1008_ (
    .A(_137_),
    .Y(_199_)
);

NAND3X1 _1009_ (
    .A(_195_),
    .B(_196_),
    .C(_139_),
    .Y(_200_)
);

OAI21X1 _1010_ (
    .A(_187_),
    .B(_191_),
    .C(_194_),
    .Y(_201_)
);

AOI21X1 _1011_ (
    .A(_201_),
    .B(_200_),
    .C(_199_),
    .Y(_202_)
);

OAI21X1 _1012_ (
    .A(_202_),
    .B(_198_),
    .C(_127_),
    .Y(_203_)
);

INVX1 _1013_ (
    .A(_127_),
    .Y(_204_)
);

NAND3X1 _1014_ (
    .A(_199_),
    .B(_200_),
    .C(_201_),
    .Y(_205_)
);

NAND3X1 _1015_ (
    .A(_137_),
    .B(_192_),
    .C(_197_),
    .Y(_206_)
);

NAND3X1 _1016_ (
    .A(_204_),
    .B(_205_),
    .C(_206_),
    .Y(_207_)
);

NAND3X1 _1017_ (
    .A(_136_),
    .B(_207_),
    .C(_203_),
    .Y(_208_)
);

INVX1 _1018_ (
    .A(_208_),
    .Y(_209_)
);

AOI21X1 _1019_ (
    .A(_203_),
    .B(_207_),
    .C(_136_),
    .Y(_210_)
);

NOR2X1 _1020_ (
    .A(_210_),
    .B(_209_),
    .Y(_753_[6])
);

NAND2X1 _1021_ (
    .A(_207_),
    .B(_208_),
    .Y(_211_)
);

AOI21X1 _1022_ (
    .A(_195_),
    .B(_196_),
    .C(_139_),
    .Y(_212_)
);

OAI21X1 _1023_ (
    .A(_137_),
    .B(_212_),
    .C(_200_),
    .Y(_213_)
);

NAND2X1 _1024_ (
    .A(_142_),
    .B(_143_),
    .Y(_214_)
);

INVX1 _1025_ (
    .A(_214_),
    .Y(_215_)
);

AOI21X1 _1026_ (
    .A(_184_),
    .B(_185_),
    .C(_146_),
    .Y(_216_)
);

OAI21X1 _1027_ (
    .A(_144_),
    .B(_216_),
    .C(_189_),
    .Y(_217_)
);

NAND2X1 _1028_ (
    .A(_140_),
    .B(_78_),
    .Y(_218_)
);

INVX1 _1029_ (
    .A(_218_),
    .Y(_219_)
);

NAND2X1 _1030_ (
    .A(Xin[0]),
    .B(Cin[7]),
    .Y(_220_)
);

INVX1 _1031_ (
    .A(_220_),
    .Y(_221_)
);

AND2X2 _1032_ (
    .A(Xin[2]),
    .B(Cin[5]),
    .Y(_222_)
);

NAND2X1 _1033_ (
    .A(_140_),
    .B(_222_),
    .Y(_223_)
);

NAND2X1 _1034_ (
    .A(Xin[1]),
    .B(Cin[6]),
    .Y(_224_)
);

OAI21X1 _1035_ (
    .A(_47_),
    .B(_77_),
    .C(_224_),
    .Y(_225_)
);

NAND3X1 _1036_ (
    .A(_225_),
    .B(_221_),
    .C(_223_),
    .Y(_226_)
);

NAND2X1 _1037_ (
    .A(Xin[2]),
    .B(Cin[5]),
    .Y(_227_)
);

NAND2X1 _1038_ (
    .A(_227_),
    .B(_140_),
    .Y(_228_)
);

NAND2X1 _1039_ (
    .A(_224_),
    .B(_222_),
    .Y(_229_)
);

NAND3X1 _1040_ (
    .A(_220_),
    .B(_228_),
    .C(_229_),
    .Y(_230_)
);

NAND2X1 _1041_ (
    .A(Cin[2]),
    .B(Xin[4]),
    .Y(_231_)
);

AND2X2 _1042_ (
    .A(_152_),
    .B(_231_),
    .Y(_232_)
);

OAI21X1 _1043_ (
    .A(_147_),
    .B(_232_),
    .C(_150_),
    .Y(_233_)
);

NAND3X1 _1044_ (
    .A(_226_),
    .B(_230_),
    .C(_233_),
    .Y(_234_)
);

AOI21X1 _1045_ (
    .A(_228_),
    .B(_229_),
    .C(_220_),
    .Y(_235_)
);

AOI22X1 _1046_ (
    .A(Xin[0]),
    .B(Cin[7]),
    .C(_223_),
    .D(_225_),
    .Y(_236_)
);

NOR2X1 _1047_ (
    .A(_152_),
    .B(_231_),
    .Y(_237_)
);

AOI21X1 _1048_ (
    .A(_148_),
    .B(_153_),
    .C(_237_),
    .Y(_238_)
);

OAI21X1 _1049_ (
    .A(_236_),
    .B(_235_),
    .C(_238_),
    .Y(_239_)
);

NAND3X1 _1050_ (
    .A(_219_),
    .B(_234_),
    .C(_239_),
    .Y(_240_)
);

NAND3X1 _1051_ (
    .A(_226_),
    .B(_230_),
    .C(_238_),
    .Y(_241_)
);

OAI21X1 _1052_ (
    .A(_236_),
    .B(_235_),
    .C(_233_),
    .Y(_242_)
);

NAND3X1 _1053_ (
    .A(_218_),
    .B(_241_),
    .C(_242_),
    .Y(_243_)
);

AND2X2 _1054_ (
    .A(_240_),
    .B(_243_),
    .Y(_244_)
);

AOI21X1 _1055_ (
    .A(_174_),
    .B(_173_),
    .C(_160_),
    .Y(_245_)
);

OAI21X1 _1056_ (
    .A(_245_),
    .B(_158_),
    .C(_177_),
    .Y(_246_)
);

NAND2X1 _1057_ (
    .A(Xin_3_bF$buf3),
    .B(Cin[4]),
    .Y(_247_)
);

INVX1 _1058_ (
    .A(_247_),
    .Y(_248_)
);

AND2X2 _1059_ (
    .A(Cin[3]),
    .B(Xin[4]),
    .Y(_249_)
);

AND2X2 _1060_ (
    .A(Cin[2]),
    .B(Xin_5_bF$buf3),
    .Y(_250_)
);

NAND2X1 _1061_ (
    .A(_249_),
    .B(_250_),
    .Y(_251_)
);

NAND2X1 _1062_ (
    .A(Cin[2]),
    .B(Xin_5_bF$buf2),
    .Y(_252_)
);

OAI21X1 _1063_ (
    .A(_740_),
    .B(_151_),
    .C(_252_),
    .Y(_253_)
);

NAND3X1 _1064_ (
    .A(_253_),
    .B(_248_),
    .C(_251_),
    .Y(_254_)
);

NAND2X1 _1065_ (
    .A(_252_),
    .B(_249_),
    .Y(_255_)
);

OAI21X1 _1066_ (
    .A(_740_),
    .B(_151_),
    .C(_250_),
    .Y(_256_)
);

NAND3X1 _1067_ (
    .A(_247_),
    .B(_255_),
    .C(_256_),
    .Y(_257_)
);

AND2X2 _1068_ (
    .A(_257_),
    .B(_254_),
    .Y(_258_)
);

AOI21X1 _1069_ (
    .A(Cin_0_bF$buf3),
    .B(Xin[6]),
    .C(Yin[6]),
    .Y(_259_)
);

OAI21X1 _1070_ (
    .A(_161_),
    .B(_259_),
    .C(_168_),
    .Y(_260_)
);

NAND2X1 _1071_ (
    .A(Cin[1]),
    .B(Xin[6]),
    .Y(_261_)
);

INVX1 _1072_ (
    .A(_261_),
    .Y(_262_)
);

NAND3X1 _1073_ (
    .A(Cin_0_bF$buf2),
    .B(Xin[7]),
    .C(Yin[7]),
    .Y(_263_)
);

INVX1 _1074_ (
    .A(Yin[7]),
    .Y(_264_)
);

NAND2X1 _1075_ (
    .A(Cin_0_bF$buf1),
    .B(Xin[7]),
    .Y(_265_)
);

NAND2X1 _1076_ (
    .A(_264_),
    .B(_265_),
    .Y(_266_)
);

NAND3X1 _1077_ (
    .A(_263_),
    .B(_262_),
    .C(_266_),
    .Y(_267_)
);

NAND2X1 _1078_ (
    .A(Yin[7]),
    .B(_265_),
    .Y(_268_)
);

NAND3X1 _1079_ (
    .A(Cin_0_bF$buf0),
    .B(Xin[7]),
    .C(_264_),
    .Y(_269_)
);

NAND3X1 _1080_ (
    .A(_261_),
    .B(_268_),
    .C(_269_),
    .Y(_270_)
);

NAND3X1 _1081_ (
    .A(_260_),
    .B(_267_),
    .C(_270_),
    .Y(_271_)
);

INVX1 _1082_ (
    .A(_260_),
    .Y(_272_)
);

AOI21X1 _1083_ (
    .A(_269_),
    .B(_268_),
    .C(_261_),
    .Y(_273_)
);

AOI21X1 _1084_ (
    .A(_266_),
    .B(_263_),
    .C(_262_),
    .Y(_274_)
);

OAI21X1 _1085_ (
    .A(_274_),
    .B(_273_),
    .C(_272_),
    .Y(_275_)
);

NAND3X1 _1086_ (
    .A(_271_),
    .B(_275_),
    .C(_258_),
    .Y(_276_)
);

NAND2X1 _1087_ (
    .A(_254_),
    .B(_257_),
    .Y(_277_)
);

OAI21X1 _1088_ (
    .A(_274_),
    .B(_273_),
    .C(_260_),
    .Y(_278_)
);

NAND3X1 _1089_ (
    .A(_267_),
    .B(_270_),
    .C(_272_),
    .Y(_279_)
);

NAND3X1 _1090_ (
    .A(_277_),
    .B(_279_),
    .C(_278_),
    .Y(_280_)
);

NAND3X1 _1091_ (
    .A(_280_),
    .B(_246_),
    .C(_276_),
    .Y(_281_)
);

INVX1 _1092_ (
    .A(_177_),
    .Y(_282_)
);

AOI21X1 _1093_ (
    .A(_183_),
    .B(_178_),
    .C(_282_),
    .Y(_283_)
);

AOI21X1 _1094_ (
    .A(_278_),
    .B(_279_),
    .C(_277_),
    .Y(_284_)
);

AOI22X1 _1095_ (
    .A(_254_),
    .B(_257_),
    .C(_275_),
    .D(_271_),
    .Y(_285_)
);

OAI21X1 _1096_ (
    .A(_284_),
    .B(_285_),
    .C(_283_),
    .Y(_286_)
);

NAND3X1 _1097_ (
    .A(_281_),
    .B(_286_),
    .C(_244_),
    .Y(_287_)
);

NAND2X1 _1098_ (
    .A(_240_),
    .B(_243_),
    .Y(_288_)
);

OAI21X1 _1099_ (
    .A(_285_),
    .B(_284_),
    .C(_246_),
    .Y(_289_)
);

NAND3X1 _1100_ (
    .A(_276_),
    .B(_280_),
    .C(_283_),
    .Y(_290_)
);

NAND3X1 _1101_ (
    .A(_288_),
    .B(_289_),
    .C(_290_),
    .Y(_291_)
);

NAND3X1 _1102_ (
    .A(_291_),
    .B(_287_),
    .C(_217_),
    .Y(_292_)
);

INVX1 _1103_ (
    .A(_189_),
    .Y(_293_)
);

AOI21X1 _1104_ (
    .A(_188_),
    .B(_190_),
    .C(_293_),
    .Y(_294_)
);

AOI21X1 _1105_ (
    .A(_290_),
    .B(_289_),
    .C(_288_),
    .Y(_295_)
);

AOI21X1 _1106_ (
    .A(_281_),
    .B(_286_),
    .C(_244_),
    .Y(_296_)
);

OAI21X1 _1107_ (
    .A(_295_),
    .B(_296_),
    .C(_294_),
    .Y(_297_)
);

NAND3X1 _1108_ (
    .A(_215_),
    .B(_292_),
    .C(_297_),
    .Y(_298_)
);

OAI21X1 _1109_ (
    .A(_295_),
    .B(_296_),
    .C(_217_),
    .Y(_299_)
);

NAND3X1 _1110_ (
    .A(_287_),
    .B(_291_),
    .C(_294_),
    .Y(_300_)
);

NAND3X1 _1111_ (
    .A(_214_),
    .B(_299_),
    .C(_300_),
    .Y(_301_)
);

NAND3X1 _1112_ (
    .A(_213_),
    .B(_298_),
    .C(_301_),
    .Y(_302_)
);

INVX1 _1113_ (
    .A(_200_),
    .Y(_303_)
);

AOI21X1 _1114_ (
    .A(_199_),
    .B(_201_),
    .C(_303_),
    .Y(_304_)
);

AOI21X1 _1115_ (
    .A(_300_),
    .B(_299_),
    .C(_214_),
    .Y(_305_)
);

AOI21X1 _1116_ (
    .A(_297_),
    .B(_292_),
    .C(_215_),
    .Y(_306_)
);

OAI21X1 _1117_ (
    .A(_306_),
    .B(_305_),
    .C(_304_),
    .Y(_307_)
);

NAND2X1 _1118_ (
    .A(_302_),
    .B(_307_),
    .Y(_308_)
);

XNOR2X1 _1119_ (
    .A(_211_),
    .B(_308_),
    .Y(_753_[7])
);

INVX1 _1120_ (
    .A(_307_),
    .Y(_309_)
);

AND2X2 _1121_ (
    .A(_302_),
    .B(_207_),
    .Y(_310_)
);

OAI22X1 _1122_ (
    .A(_309_),
    .B(_310_),
    .C(_308_),
    .D(_208_),
    .Y(_311_)
);

INVX1 _1123_ (
    .A(_292_),
    .Y(_312_)
);

AOI21X1 _1124_ (
    .A(_215_),
    .B(_297_),
    .C(_312_),
    .Y(_313_)
);

NAND2X1 _1125_ (
    .A(_234_),
    .B(_240_),
    .Y(_314_)
);

INVX1 _1126_ (
    .A(_314_),
    .Y(_315_)
);

AOI21X1 _1127_ (
    .A(_276_),
    .B(_280_),
    .C(_246_),
    .Y(_316_)
);

OAI21X1 _1128_ (
    .A(_288_),
    .B(_316_),
    .C(_281_),
    .Y(_317_)
);

OAI21X1 _1129_ (
    .A(_224_),
    .B(_227_),
    .C(_226_),
    .Y(_318_)
);

NAND2X1 _1130_ (
    .A(Xin[1]),
    .B(Cin[7]),
    .Y(_319_)
);

INVX1 _1131_ (
    .A(_319_),
    .Y(_320_)
);

AND2X2 _1132_ (
    .A(Xin[2]),
    .B(Cin[6]),
    .Y(_321_)
);

AND2X2 _1133_ (
    .A(Xin_3_bF$buf2),
    .B(Cin[5]),
    .Y(_322_)
);

NAND2X1 _1134_ (
    .A(_321_),
    .B(_322_),
    .Y(_323_)
);

INVX1 _1135_ (
    .A(Cin[6]),
    .Y(_324_)
);

NAND2X1 _1136_ (
    .A(Xin_3_bF$buf1),
    .B(Cin[5]),
    .Y(_325_)
);

OAI21X1 _1137_ (
    .A(_47_),
    .B(_324_),
    .C(_325_),
    .Y(_326_)
);

NAND3X1 _1138_ (
    .A(_326_),
    .B(_320_),
    .C(_323_),
    .Y(_327_)
);

OAI21X1 _1139_ (
    .A(_87_),
    .B(_77_),
    .C(_321_),
    .Y(_328_)
);

OAI21X1 _1140_ (
    .A(_47_),
    .B(_324_),
    .C(_322_),
    .Y(_329_)
);

NAND3X1 _1141_ (
    .A(_319_),
    .B(_328_),
    .C(_329_),
    .Y(_330_)
);

AOI22X1 _1142_ (
    .A(Cin[2]),
    .B(Xin_5_bF$buf1),
    .C(Cin[3]),
    .D(Xin[4]),
    .Y(_331_)
);

OAI21X1 _1143_ (
    .A(_247_),
    .B(_331_),
    .C(_251_),
    .Y(_332_)
);

NAND3X1 _1144_ (
    .A(_332_),
    .B(_327_),
    .C(_330_),
    .Y(_333_)
);

AOI21X1 _1145_ (
    .A(_328_),
    .B(_329_),
    .C(_319_),
    .Y(_334_)
);

AOI21X1 _1146_ (
    .A(_323_),
    .B(_326_),
    .C(_320_),
    .Y(_335_)
);

NAND2X1 _1147_ (
    .A(Cin[3]),
    .B(Xin_5_bF$buf0),
    .Y(_336_)
);

INVX1 _1148_ (
    .A(_336_),
    .Y(_337_)
);

AOI22X1 _1149_ (
    .A(_149_),
    .B(_337_),
    .C(_253_),
    .D(_248_),
    .Y(_338_)
);

OAI21X1 _1150_ (
    .A(_335_),
    .B(_334_),
    .C(_338_),
    .Y(_339_)
);

NAND3X1 _1151_ (
    .A(_318_),
    .B(_333_),
    .C(_339_),
    .Y(_340_)
);

AND2X2 _1152_ (
    .A(_226_),
    .B(_223_),
    .Y(_341_)
);

NAND3X1 _1153_ (
    .A(_327_),
    .B(_338_),
    .C(_330_),
    .Y(_342_)
);

OAI21X1 _1154_ (
    .A(_335_),
    .B(_334_),
    .C(_332_),
    .Y(_343_)
);

NAND3X1 _1155_ (
    .A(_341_),
    .B(_342_),
    .C(_343_),
    .Y(_344_)
);

NAND2X1 _1156_ (
    .A(_340_),
    .B(_344_),
    .Y(_345_)
);

AOI21X1 _1157_ (
    .A(_270_),
    .B(_267_),
    .C(_260_),
    .Y(_346_)
);

OAI21X1 _1158_ (
    .A(_346_),
    .B(_277_),
    .C(_271_),
    .Y(_347_)
);

NAND2X1 _1159_ (
    .A(Xin[4]),
    .B(Cin[4]),
    .Y(_348_)
);

INVX1 _1160_ (
    .A(_348_),
    .Y(_349_)
);

AND2X2 _1161_ (
    .A(Cin[3]),
    .B(Xin[6]),
    .Y(_350_)
);

NAND2X1 _1162_ (
    .A(_250_),
    .B(_350_),
    .Y(_351_)
);

INVX1 _1163_ (
    .A(Xin[6]),
    .Y(_352_)
);

OAI21X1 _1164_ (
    .A(_590_),
    .B(_352_),
    .C(_336_),
    .Y(_353_)
);

NAND3X1 _1165_ (
    .A(_353_),
    .B(_349_),
    .C(_351_),
    .Y(_354_)
);

NAND2X1 _1166_ (
    .A(Cin[2]),
    .B(Xin[6]),
    .Y(_355_)
);

NAND3X1 _1167_ (
    .A(Cin[3]),
    .B(Xin_5_bF$buf3),
    .C(_355_),
    .Y(_356_)
);

NAND3X1 _1168_ (
    .A(Cin[2]),
    .B(Xin[6]),
    .C(_336_),
    .Y(_357_)
);

NAND3X1 _1169_ (
    .A(_348_),
    .B(_356_),
    .C(_357_),
    .Y(_358_)
);

NAND2X1 _1170_ (
    .A(_358_),
    .B(_354_),
    .Y(_359_)
);

AOI21X1 _1171_ (
    .A(Cin_0_bF$buf3),
    .B(Xin[7]),
    .C(Yin[7]),
    .Y(_360_)
);

OAI21X1 _1172_ (
    .A(_261_),
    .B(_360_),
    .C(_263_),
    .Y(_361_)
);

NAND3X1 _1173_ (
    .A(Cin[1]),
    .B(Xin[7]),
    .C(Yin[8]),
    .Y(_362_)
);

INVX1 _1174_ (
    .A(_362_),
    .Y(_363_)
);

AOI21X1 _1175_ (
    .A(Cin[1]),
    .B(Xin[7]),
    .C(Yin[8]),
    .Y(_364_)
);

OAI21X1 _1176_ (
    .A(_363_),
    .B(_364_),
    .C(_361_),
    .Y(_365_)
);

NOR2X1 _1177_ (
    .A(_364_),
    .B(_363_),
    .Y(_366_)
);

NAND3X1 _1178_ (
    .A(_263_),
    .B(_267_),
    .C(_366_),
    .Y(_367_)
);

AOI21X1 _1179_ (
    .A(_367_),
    .B(_365_),
    .C(_359_),
    .Y(_368_)
);

NAND2X1 _1180_ (
    .A(_361_),
    .B(_366_),
    .Y(_369_)
);

INVX1 _1181_ (
    .A(_364_),
    .Y(_370_)
);

NAND2X1 _1182_ (
    .A(_362_),
    .B(_370_),
    .Y(_371_)
);

NAND3X1 _1183_ (
    .A(_263_),
    .B(_267_),
    .C(_371_),
    .Y(_372_)
);

AOI22X1 _1184_ (
    .A(_354_),
    .B(_358_),
    .C(_369_),
    .D(_372_),
    .Y(_373_)
);

OAI21X1 _1185_ (
    .A(_373_),
    .B(_368_),
    .C(_347_),
    .Y(_374_)
);

INVX1 _1186_ (
    .A(_271_),
    .Y(_375_)
);

AOI21X1 _1187_ (
    .A(_258_),
    .B(_275_),
    .C(_375_),
    .Y(_376_)
);

AND2X2 _1188_ (
    .A(_354_),
    .B(_358_),
    .Y(_377_)
);

NAND3X1 _1189_ (
    .A(_369_),
    .B(_372_),
    .C(_377_),
    .Y(_378_)
);

NAND3X1 _1190_ (
    .A(_365_),
    .B(_359_),
    .C(_367_),
    .Y(_379_)
);

NAND3X1 _1191_ (
    .A(_378_),
    .B(_379_),
    .C(_376_),
    .Y(_380_)
);

AOI21X1 _1192_ (
    .A(_380_),
    .B(_374_),
    .C(_345_),
    .Y(_381_)
);

AND2X2 _1193_ (
    .A(_340_),
    .B(_344_),
    .Y(_382_)
);

NAND3X1 _1194_ (
    .A(_379_),
    .B(_347_),
    .C(_378_),
    .Y(_383_)
);

OAI21X1 _1195_ (
    .A(_368_),
    .B(_373_),
    .C(_376_),
    .Y(_384_)
);

AOI21X1 _1196_ (
    .A(_383_),
    .B(_384_),
    .C(_382_),
    .Y(_385_)
);

OAI21X1 _1197_ (
    .A(_381_),
    .B(_385_),
    .C(_317_),
    .Y(_387_)
);

INVX1 _1198_ (
    .A(_281_),
    .Y(_388_)
);

AOI21X1 _1199_ (
    .A(_244_),
    .B(_286_),
    .C(_388_),
    .Y(_389_)
);

NAND3X1 _1200_ (
    .A(_383_),
    .B(_384_),
    .C(_382_),
    .Y(_390_)
);

NAND3X1 _1201_ (
    .A(_345_),
    .B(_374_),
    .C(_380_),
    .Y(_391_)
);

NAND3X1 _1202_ (
    .A(_390_),
    .B(_391_),
    .C(_389_),
    .Y(_392_)
);

AOI21X1 _1203_ (
    .A(_392_),
    .B(_387_),
    .C(_315_),
    .Y(_393_)
);

NAND3X1 _1204_ (
    .A(_391_),
    .B(_317_),
    .C(_390_),
    .Y(_394_)
);

OAI21X1 _1205_ (
    .A(_381_),
    .B(_385_),
    .C(_389_),
    .Y(_395_)
);

AOI21X1 _1206_ (
    .A(_395_),
    .B(_394_),
    .C(_314_),
    .Y(_396_)
);

OAI21X1 _1207_ (
    .A(_396_),
    .B(_393_),
    .C(_313_),
    .Y(_398_)
);

AOI21X1 _1208_ (
    .A(_287_),
    .B(_291_),
    .C(_217_),
    .Y(_399_)
);

OAI21X1 _1209_ (
    .A(_214_),
    .B(_399_),
    .C(_292_),
    .Y(_400_)
);

NAND3X1 _1210_ (
    .A(_314_),
    .B(_394_),
    .C(_395_),
    .Y(_401_)
);

NAND3X1 _1211_ (
    .A(_315_),
    .B(_387_),
    .C(_392_),
    .Y(_402_)
);

NAND3X1 _1212_ (
    .A(_400_),
    .B(_401_),
    .C(_402_),
    .Y(_403_)
);

NAND2X1 _1213_ (
    .A(_403_),
    .B(_398_),
    .Y(_404_)
);

XNOR2X1 _1214_ (
    .A(_311_),
    .B(_404_),
    .Y(_753_[8])
);

INVX1 _1215_ (
    .A(_311_),
    .Y(_405_)
);

OAI21X1 _1216_ (
    .A(_404_),
    .B(_405_),
    .C(_403_),
    .Y(_406_)
);

AOI21X1 _1217_ (
    .A(_390_),
    .B(_391_),
    .C(_317_),
    .Y(_408_)
);

OAI21X1 _1218_ (
    .A(_315_),
    .B(_408_),
    .C(_394_),
    .Y(_409_)
);

NAND2X1 _1219_ (
    .A(_333_),
    .B(_340_),
    .Y(_410_)
);

AOI21X1 _1220_ (
    .A(_378_),
    .B(_379_),
    .C(_347_),
    .Y(_411_)
);

OAI21X1 _1221_ (
    .A(_345_),
    .B(_411_),
    .C(_383_),
    .Y(_412_)
);

NAND2X1 _1222_ (
    .A(Xin_3_bF$buf0),
    .B(Cin[6]),
    .Y(_413_)
);

OAI21X1 _1223_ (
    .A(_227_),
    .B(_413_),
    .C(_327_),
    .Y(_414_)
);

NAND2X1 _1224_ (
    .A(Xin[2]),
    .B(Cin[7]),
    .Y(_415_)
);

AOI22X1 _1225_ (
    .A(Xin_3_bF$buf3),
    .B(Cin[6]),
    .C(Xin[4]),
    .D(Cin[5]),
    .Y(_416_)
);

NAND2X1 _1226_ (
    .A(Xin[4]),
    .B(Cin[6]),
    .Y(_417_)
);

NOR2X1 _1227_ (
    .A(_325_),
    .B(_417_),
    .Y(_419_)
);

OAI21X1 _1228_ (
    .A(_416_),
    .B(_419_),
    .C(_415_),
    .Y(_420_)
);

INVX1 _1229_ (
    .A(_415_),
    .Y(_421_)
);

INVX1 _1230_ (
    .A(_416_),
    .Y(_422_)
);

AND2X2 _1231_ (
    .A(Xin[4]),
    .B(Cin[6]),
    .Y(_423_)
);

NAND2X1 _1232_ (
    .A(_322_),
    .B(_423_),
    .Y(_424_)
);

NAND3X1 _1233_ (
    .A(_421_),
    .B(_422_),
    .C(_424_),
    .Y(_425_)
);

AND2X2 _1234_ (
    .A(_336_),
    .B(_355_),
    .Y(_426_)
);

OAI21X1 _1235_ (
    .A(_348_),
    .B(_426_),
    .C(_351_),
    .Y(_427_)
);

NAND3X1 _1236_ (
    .A(_425_),
    .B(_420_),
    .C(_427_),
    .Y(_428_)
);

AOI21X1 _1237_ (
    .A(_424_),
    .B(_422_),
    .C(_421_),
    .Y(_430_)
);

NOR3X1 _1238_ (
    .A(_415_),
    .B(_416_),
    .C(_419_),
    .Y(_431_)
);

AOI22X1 _1239_ (
    .A(_250_),
    .B(_350_),
    .C(_353_),
    .D(_349_),
    .Y(_432_)
);

OAI21X1 _1240_ (
    .A(_430_),
    .B(_431_),
    .C(_432_),
    .Y(_433_)
);

NAND3X1 _1241_ (
    .A(_414_),
    .B(_428_),
    .C(_433_),
    .Y(_434_)
);

AND2X2 _1242_ (
    .A(_327_),
    .B(_323_),
    .Y(_435_)
);

NAND3X1 _1243_ (
    .A(_425_),
    .B(_432_),
    .C(_420_),
    .Y(_436_)
);

OAI21X1 _1244_ (
    .A(_430_),
    .B(_431_),
    .C(_427_),
    .Y(_437_)
);

NAND3X1 _1245_ (
    .A(_435_),
    .B(_436_),
    .C(_437_),
    .Y(_438_)
);

AND2X2 _1246_ (
    .A(_434_),
    .B(_438_),
    .Y(_439_)
);

NOR2X1 _1247_ (
    .A(_361_),
    .B(_366_),
    .Y(_441_)
);

OAI21X1 _1248_ (
    .A(_359_),
    .B(_441_),
    .C(_369_),
    .Y(_442_)
);

NAND2X1 _1249_ (
    .A(Xin_5_bF$buf2),
    .B(Cin[4]),
    .Y(_443_)
);

INVX1 _1250_ (
    .A(_443_),
    .Y(_444_)
);

AND2X2 _1251_ (
    .A(Cin[2]),
    .B(Xin[7]),
    .Y(_445_)
);

NAND2X1 _1252_ (
    .A(_350_),
    .B(_445_),
    .Y(_446_)
);

INVX1 _1253_ (
    .A(Xin[7]),
    .Y(_447_)
);

OAI22X1 _1254_ (
    .A(_590_),
    .B(_447_),
    .C(_740_),
    .D(_352_),
    .Y(_448_)
);

NAND3X1 _1255_ (
    .A(_444_),
    .B(_448_),
    .C(_446_),
    .Y(_449_)
);

OAI21X1 _1256_ (
    .A(_590_),
    .B(_447_),
    .C(_350_),
    .Y(_450_)
);

OAI21X1 _1257_ (
    .A(_740_),
    .B(_352_),
    .C(_445_),
    .Y(_451_)
);

NAND3X1 _1258_ (
    .A(_443_),
    .B(_450_),
    .C(_451_),
    .Y(_452_)
);

XNOR2X1 _1259_ (
    .A(_362_),
    .B(Yin[9]),
    .Y(_453_)
);

NAND3X1 _1260_ (
    .A(_453_),
    .B(_449_),
    .C(_452_),
    .Y(_454_)
);

NAND2X1 _1261_ (
    .A(_449_),
    .B(_452_),
    .Y(_455_)
);

INVX1 _1262_ (
    .A(_453_),
    .Y(_456_)
);

NAND2X1 _1263_ (
    .A(_456_),
    .B(_455_),
    .Y(_457_)
);

NAND3X1 _1264_ (
    .A(_454_),
    .B(_457_),
    .C(_442_),
    .Y(_458_)
);

AOI21X1 _1265_ (
    .A(_263_),
    .B(_267_),
    .C(_371_),
    .Y(_459_)
);

AOI21X1 _1266_ (
    .A(_377_),
    .B(_372_),
    .C(_459_),
    .Y(_460_)
);

NAND2X1 _1267_ (
    .A(_454_),
    .B(_457_),
    .Y(_462_)
);

NAND2X1 _1268_ (
    .A(_460_),
    .B(_462_),
    .Y(_463_)
);

NAND3X1 _1269_ (
    .A(_458_),
    .B(_463_),
    .C(_439_),
    .Y(_464_)
);

NAND2X1 _1270_ (
    .A(_434_),
    .B(_438_),
    .Y(_465_)
);

NOR2X1 _1271_ (
    .A(_460_),
    .B(_462_),
    .Y(_466_)
);

AOI21X1 _1272_ (
    .A(_454_),
    .B(_457_),
    .C(_442_),
    .Y(_467_)
);

OAI21X1 _1273_ (
    .A(_467_),
    .B(_466_),
    .C(_465_),
    .Y(_468_)
);

NAND3X1 _1274_ (
    .A(_412_),
    .B(_464_),
    .C(_468_),
    .Y(_469_)
);

INVX1 _1275_ (
    .A(_383_),
    .Y(_470_)
);

AOI21X1 _1276_ (
    .A(_382_),
    .B(_384_),
    .C(_470_),
    .Y(_471_)
);

NAND2X1 _1277_ (
    .A(_442_),
    .B(_462_),
    .Y(_473_)
);

NAND3X1 _1278_ (
    .A(_454_),
    .B(_457_),
    .C(_460_),
    .Y(_474_)
);

AOI21X1 _1279_ (
    .A(_473_),
    .B(_474_),
    .C(_465_),
    .Y(_475_)
);

AOI22X1 _1280_ (
    .A(_434_),
    .B(_438_),
    .C(_463_),
    .D(_458_),
    .Y(_476_)
);

OAI21X1 _1281_ (
    .A(_475_),
    .B(_476_),
    .C(_471_),
    .Y(_477_)
);

NAND3X1 _1282_ (
    .A(_410_),
    .B(_469_),
    .C(_477_),
    .Y(_478_)
);

INVX1 _1283_ (
    .A(_410_),
    .Y(_479_)
);

OAI21X1 _1284_ (
    .A(_476_),
    .B(_475_),
    .C(_412_),
    .Y(_480_)
);

NAND3X1 _1285_ (
    .A(_464_),
    .B(_468_),
    .C(_471_),
    .Y(_481_)
);

NAND3X1 _1286_ (
    .A(_479_),
    .B(_480_),
    .C(_481_),
    .Y(_482_)
);

NAND3X1 _1287_ (
    .A(_409_),
    .B(_478_),
    .C(_482_),
    .Y(_484_)
);

INVX1 _1288_ (
    .A(_394_),
    .Y(_485_)
);

AOI21X1 _1289_ (
    .A(_314_),
    .B(_395_),
    .C(_485_),
    .Y(_486_)
);

AOI21X1 _1290_ (
    .A(_481_),
    .B(_480_),
    .C(_479_),
    .Y(_487_)
);

AOI21X1 _1291_ (
    .A(_477_),
    .B(_469_),
    .C(_410_),
    .Y(_488_)
);

OAI21X1 _1292_ (
    .A(_487_),
    .B(_488_),
    .C(_486_),
    .Y(_489_)
);

NAND2X1 _1293_ (
    .A(_484_),
    .B(_489_),
    .Y(_490_)
);

XNOR2X1 _1294_ (
    .A(_406_),
    .B(_490_),
    .Y(_753_[9])
);

INVX1 _1295_ (
    .A(_489_),
    .Y(_491_)
);

OAI21X1 _1296_ (
    .A(_403_),
    .B(_491_),
    .C(_484_),
    .Y(_492_)
);

NOR2X1 _1297_ (
    .A(_404_),
    .B(_490_),
    .Y(_494_)
);

AOI21X1 _1298_ (
    .A(_311_),
    .B(_494_),
    .C(_492_),
    .Y(_495_)
);

NOR3X1 _1299_ (
    .A(_475_),
    .B(_476_),
    .C(_471_),
    .Y(_496_)
);

AOI21X1 _1300_ (
    .A(_410_),
    .B(_477_),
    .C(_496_),
    .Y(_497_)
);

NAND2X1 _1301_ (
    .A(_428_),
    .B(_434_),
    .Y(_498_)
);

INVX1 _1302_ (
    .A(_498_),
    .Y(_499_)
);

OAI21X1 _1303_ (
    .A(_467_),
    .B(_465_),
    .C(_458_),
    .Y(_500_)
);

OAI21X1 _1304_ (
    .A(_415_),
    .B(_416_),
    .C(_424_),
    .Y(_501_)
);

NAND2X1 _1305_ (
    .A(Xin_3_bF$buf2),
    .B(Cin[7]),
    .Y(_502_)
);

NAND2X1 _1306_ (
    .A(Xin_5_bF$buf1),
    .B(Cin[5]),
    .Y(_503_)
);

NOR2X1 _1307_ (
    .A(_417_),
    .B(_503_),
    .Y(_505_)
);

AOI22X1 _1308_ (
    .A(Xin_5_bF$buf0),
    .B(Cin[5]),
    .C(Xin[4]),
    .D(Cin[6]),
    .Y(_506_)
);

OAI21X1 _1309_ (
    .A(_506_),
    .B(_505_),
    .C(_502_),
    .Y(_507_)
);

INVX1 _1310_ (
    .A(_502_),
    .Y(_508_)
);

AND2X2 _1311_ (
    .A(Xin_5_bF$buf3),
    .B(Cin[5]),
    .Y(_509_)
);

NAND2X1 _1312_ (
    .A(_423_),
    .B(_509_),
    .Y(_510_)
);

INVX1 _1313_ (
    .A(_506_),
    .Y(_511_)
);

NAND3X1 _1314_ (
    .A(_508_),
    .B(_511_),
    .C(_510_),
    .Y(_512_)
);

NOR2X1 _1315_ (
    .A(_350_),
    .B(_445_),
    .Y(_513_)
);

OAI21X1 _1316_ (
    .A(_443_),
    .B(_513_),
    .C(_446_),
    .Y(_514_)
);

NAND3X1 _1317_ (
    .A(_507_),
    .B(_512_),
    .C(_514_),
    .Y(_516_)
);

AOI21X1 _1318_ (
    .A(_510_),
    .B(_511_),
    .C(_508_),
    .Y(_517_)
);

NOR3X1 _1319_ (
    .A(_502_),
    .B(_506_),
    .C(_505_),
    .Y(_518_)
);

AND2X2 _1320_ (
    .A(_350_),
    .B(_445_),
    .Y(_519_)
);

AOI21X1 _1321_ (
    .A(_444_),
    .B(_448_),
    .C(_519_),
    .Y(_520_)
);

OAI21X1 _1322_ (
    .A(_517_),
    .B(_518_),
    .C(_520_),
    .Y(_521_)
);

NAND3X1 _1323_ (
    .A(_501_),
    .B(_516_),
    .C(_521_),
    .Y(_522_)
);

INVX1 _1324_ (
    .A(_501_),
    .Y(_523_)
);

NAND3X1 _1325_ (
    .A(_512_),
    .B(_507_),
    .C(_520_),
    .Y(_524_)
);

OAI21X1 _1326_ (
    .A(_517_),
    .B(_518_),
    .C(_514_),
    .Y(_525_)
);

NAND3X1 _1327_ (
    .A(_523_),
    .B(_524_),
    .C(_525_),
    .Y(_527_)
);

NAND2X1 _1328_ (
    .A(_522_),
    .B(_527_),
    .Y(_528_)
);

NAND2X1 _1329_ (
    .A(Yin[9]),
    .B(_363_),
    .Y(_529_)
);

NAND2X1 _1330_ (
    .A(_529_),
    .B(_454_),
    .Y(_530_)
);

AOI22X1 _1331_ (
    .A(Cin[3]),
    .B(Xin[7]),
    .C(Cin[4]),
    .D(Xin[6]),
    .Y(_531_)
);

AND2X2 _1332_ (
    .A(Cin[4]),
    .B(Xin[7]),
    .Y(_532_)
);

AOI21X1 _1333_ (
    .A(_350_),
    .B(_532_),
    .C(_531_),
    .Y(_533_)
);

NAND2X1 _1334_ (
    .A(Yin[10]),
    .B(_533_),
    .Y(_534_)
);

INVX1 _1335_ (
    .A(Yin[10]),
    .Y(_535_)
);

AND2X2 _1336_ (
    .A(_350_),
    .B(_532_),
    .Y(_536_)
);

OAI21X1 _1337_ (
    .A(_531_),
    .B(_536_),
    .C(_535_),
    .Y(_538_)
);

NAND2X1 _1338_ (
    .A(_534_),
    .B(_538_),
    .Y(_539_)
);

XOR2X1 _1339_ (
    .A(_530_),
    .B(_539_),
    .Y(_540_)
);

NOR2X1 _1340_ (
    .A(_528_),
    .B(_540_),
    .Y(_541_)
);

AND2X2 _1341_ (
    .A(_522_),
    .B(_527_),
    .Y(_542_)
);

NAND2X1 _1342_ (
    .A(_539_),
    .B(_530_),
    .Y(_543_)
);

AND2X2 _1343_ (
    .A(_538_),
    .B(_534_),
    .Y(_544_)
);

NAND3X1 _1344_ (
    .A(_529_),
    .B(_454_),
    .C(_544_),
    .Y(_545_)
);

NAND2X1 _1345_ (
    .A(_543_),
    .B(_545_),
    .Y(_546_)
);

NOR2X1 _1346_ (
    .A(_546_),
    .B(_542_),
    .Y(_547_)
);

OAI21X1 _1347_ (
    .A(_541_),
    .B(_547_),
    .C(_500_),
    .Y(_549_)
);

AOI21X1 _1348_ (
    .A(_439_),
    .B(_463_),
    .C(_466_),
    .Y(_550_)
);

NAND3X1 _1349_ (
    .A(_522_),
    .B(_527_),
    .C(_546_),
    .Y(_551_)
);

NAND2X1 _1350_ (
    .A(_528_),
    .B(_540_),
    .Y(_552_)
);

NAND3X1 _1351_ (
    .A(_551_),
    .B(_552_),
    .C(_550_),
    .Y(_553_)
);

AOI21X1 _1352_ (
    .A(_549_),
    .B(_553_),
    .C(_499_),
    .Y(_554_)
);

NAND3X1 _1353_ (
    .A(_551_),
    .B(_552_),
    .C(_500_),
    .Y(_555_)
);

OAI21X1 _1354_ (
    .A(_541_),
    .B(_547_),
    .C(_550_),
    .Y(_556_)
);

AOI21X1 _1355_ (
    .A(_556_),
    .B(_555_),
    .C(_498_),
    .Y(_557_)
);

OAI21X1 _1356_ (
    .A(_554_),
    .B(_557_),
    .C(_497_),
    .Y(_558_)
);

AOI21X1 _1357_ (
    .A(_468_),
    .B(_464_),
    .C(_412_),
    .Y(_560_)
);

OAI21X1 _1358_ (
    .A(_479_),
    .B(_560_),
    .C(_469_),
    .Y(_561_)
);

NAND3X1 _1359_ (
    .A(_555_),
    .B(_498_),
    .C(_556_),
    .Y(_562_)
);

NAND3X1 _1360_ (
    .A(_499_),
    .B(_553_),
    .C(_549_),
    .Y(_563_)
);

NAND3X1 _1361_ (
    .A(_562_),
    .B(_563_),
    .C(_561_),
    .Y(_564_)
);

NAND2X1 _1362_ (
    .A(_564_),
    .B(_558_),
    .Y(_565_)
);

XOR2X1 _1363_ (
    .A(_495_),
    .B(_565_),
    .Y(_753_[10])
);

OAI21X1 _1364_ (
    .A(_565_),
    .B(_495_),
    .C(_564_),
    .Y(_566_)
);

INVX1 _1365_ (
    .A(_555_),
    .Y(_567_)
);

AOI21X1 _1366_ (
    .A(_498_),
    .B(_556_),
    .C(_567_),
    .Y(_568_)
);

NAND2X1 _1367_ (
    .A(_516_),
    .B(_522_),
    .Y(_570_)
);

INVX1 _1368_ (
    .A(_570_),
    .Y(_571_)
);

NAND2X1 _1369_ (
    .A(_544_),
    .B(_530_),
    .Y(_572_)
);

OAI21X1 _1370_ (
    .A(_528_),
    .B(_540_),
    .C(_572_),
    .Y(_573_)
);

OAI21X1 _1371_ (
    .A(_502_),
    .B(_506_),
    .C(_510_),
    .Y(_574_)
);

INVX1 _1372_ (
    .A(Cin[7]),
    .Y(_575_)
);

NAND2X1 _1373_ (
    .A(Xin[6]),
    .B(Cin[6]),
    .Y(_576_)
);

INVX1 _1374_ (
    .A(Xin_5_bF$buf2),
    .Y(_577_)
);

NAND2X1 _1375_ (
    .A(Cin[5]),
    .B(Xin[6]),
    .Y(_578_)
);

OAI21X1 _1376_ (
    .A(_577_),
    .B(_324_),
    .C(_578_),
    .Y(_579_)
);

OAI21X1 _1377_ (
    .A(_503_),
    .B(_576_),
    .C(_579_),
    .Y(_580_)
);

OAI21X1 _1378_ (
    .A(_151_),
    .B(_575_),
    .C(_580_),
    .Y(_581_)
);

NAND2X1 _1379_ (
    .A(Xin[4]),
    .B(Cin[7]),
    .Y(_582_)
);

INVX1 _1380_ (
    .A(_582_),
    .Y(_583_)
);

NOR2X1 _1381_ (
    .A(_503_),
    .B(_576_),
    .Y(_584_)
);

INVX1 _1382_ (
    .A(_584_),
    .Y(_585_)
);

NAND3X1 _1383_ (
    .A(_583_),
    .B(_579_),
    .C(_585_),
    .Y(_586_)
);

NAND3X1 _1384_ (
    .A(_536_),
    .B(_581_),
    .C(_586_),
    .Y(_587_)
);

INVX1 _1385_ (
    .A(_536_),
    .Y(_588_)
);

AOI21X1 _1386_ (
    .A(_585_),
    .B(_579_),
    .C(_583_),
    .Y(_589_)
);

NOR2X1 _1387_ (
    .A(_582_),
    .B(_580_),
    .Y(_591_)
);

OAI21X1 _1388_ (
    .A(_591_),
    .B(_589_),
    .C(_588_),
    .Y(_592_)
);

NAND3X1 _1389_ (
    .A(_574_),
    .B(_587_),
    .C(_592_),
    .Y(_593_)
);

INVX1 _1390_ (
    .A(_574_),
    .Y(_594_)
);

NAND3X1 _1391_ (
    .A(_588_),
    .B(_581_),
    .C(_586_),
    .Y(_595_)
);

OAI21X1 _1392_ (
    .A(_591_),
    .B(_589_),
    .C(_536_),
    .Y(_596_)
);

NAND3X1 _1393_ (
    .A(_594_),
    .B(_595_),
    .C(_596_),
    .Y(_597_)
);

XNOR2X1 _1394_ (
    .A(_532_),
    .B(Yin[11]),
    .Y(_598_)
);

NAND2X1 _1395_ (
    .A(_598_),
    .B(_534_),
    .Y(_599_)
);

OR2X2 _1396_ (
    .A(_534_),
    .B(_598_),
    .Y(_600_)
);

NAND2X1 _1397_ (
    .A(_599_),
    .B(_600_),
    .Y(_602_)
);

INVX1 _1398_ (
    .A(_602_),
    .Y(_603_)
);

NAND3X1 _1399_ (
    .A(_593_),
    .B(_597_),
    .C(_603_),
    .Y(_604_)
);

AOI21X1 _1400_ (
    .A(_596_),
    .B(_595_),
    .C(_594_),
    .Y(_605_)
);

AOI21X1 _1401_ (
    .A(_592_),
    .B(_587_),
    .C(_574_),
    .Y(_606_)
);

OAI21X1 _1402_ (
    .A(_605_),
    .B(_606_),
    .C(_602_),
    .Y(_607_)
);

NAND2X1 _1403_ (
    .A(_604_),
    .B(_607_),
    .Y(_608_)
);

NAND2X1 _1404_ (
    .A(_573_),
    .B(_608_),
    .Y(_609_)
);

INVX1 _1405_ (
    .A(_572_),
    .Y(_610_)
);

AOI21X1 _1406_ (
    .A(_542_),
    .B(_546_),
    .C(_610_),
    .Y(_611_)
);

NAND3X1 _1407_ (
    .A(_604_),
    .B(_607_),
    .C(_611_),
    .Y(_613_)
);

AOI21X1 _1408_ (
    .A(_609_),
    .B(_613_),
    .C(_571_),
    .Y(_614_)
);

NAND3X1 _1409_ (
    .A(_604_),
    .B(_607_),
    .C(_573_),
    .Y(_615_)
);

NAND2X1 _1410_ (
    .A(_611_),
    .B(_608_),
    .Y(_616_)
);

AOI21X1 _1411_ (
    .A(_616_),
    .B(_615_),
    .C(_570_),
    .Y(_617_)
);

OAI21X1 _1412_ (
    .A(_614_),
    .B(_617_),
    .C(_568_),
    .Y(_618_)
);

AOI21X1 _1413_ (
    .A(_552_),
    .B(_551_),
    .C(_500_),
    .Y(_619_)
);

OAI21X1 _1414_ (
    .A(_499_),
    .B(_619_),
    .C(_555_),
    .Y(_620_)
);

NAND3X1 _1415_ (
    .A(_570_),
    .B(_615_),
    .C(_616_),
    .Y(_621_)
);

NAND3X1 _1416_ (
    .A(_571_),
    .B(_613_),
    .C(_609_),
    .Y(_622_)
);

NAND3X1 _1417_ (
    .A(_620_),
    .B(_621_),
    .C(_622_),
    .Y(_624_)
);

NAND2X1 _1418_ (
    .A(_624_),
    .B(_618_),
    .Y(_625_)
);

INVX1 _1419_ (
    .A(_625_),
    .Y(_626_)
);

XOR2X1 _1420_ (
    .A(_566_),
    .B(_626_),
    .Y(_753_[11])
);

NOR2X1 _1421_ (
    .A(_625_),
    .B(_565_),
    .Y(_627_)
);

NAND3X1 _1422_ (
    .A(_494_),
    .B(_311_),
    .C(_627_),
    .Y(_628_)
);

INVX1 _1423_ (
    .A(_565_),
    .Y(_629_)
);

NAND3X1 _1424_ (
    .A(_626_),
    .B(_629_),
    .C(_492_),
    .Y(_630_)
);

NAND2X1 _1425_ (
    .A(_624_),
    .B(_564_),
    .Y(_631_)
);

NAND2X1 _1426_ (
    .A(_618_),
    .B(_631_),
    .Y(_632_)
);

NAND3X1 _1427_ (
    .A(_630_),
    .B(_632_),
    .C(_628_),
    .Y(_634_)
);

NAND2X1 _1428_ (
    .A(_587_),
    .B(_593_),
    .Y(_635_)
);

INVX1 _1429_ (
    .A(_635_),
    .Y(_636_)
);

AND2X2 _1430_ (
    .A(_604_),
    .B(_600_),
    .Y(_637_)
);

OAI21X1 _1431_ (
    .A(_582_),
    .B(_580_),
    .C(_585_),
    .Y(_638_)
);

NAND2X1 _1432_ (
    .A(Cin[6]),
    .B(Xin[7]),
    .Y(_639_)
);

OAI21X1 _1433_ (
    .A(_77_),
    .B(_447_),
    .C(_576_),
    .Y(_640_)
);

OAI21X1 _1434_ (
    .A(_578_),
    .B(_639_),
    .C(_640_),
    .Y(_641_)
);

OAI21X1 _1435_ (
    .A(_577_),
    .B(_575_),
    .C(_641_),
    .Y(_642_)
);

NAND2X1 _1436_ (
    .A(Xin_5_bF$buf1),
    .B(Cin[7]),
    .Y(_643_)
);

OR2X2 _1437_ (
    .A(_641_),
    .B(_643_),
    .Y(_645_)
);

NAND3X1 _1438_ (
    .A(_638_),
    .B(_642_),
    .C(_645_),
    .Y(_646_)
);

INVX1 _1439_ (
    .A(_646_),
    .Y(_647_)
);

AOI21X1 _1440_ (
    .A(_645_),
    .B(_642_),
    .C(_638_),
    .Y(_648_)
);

NOR2X1 _1441_ (
    .A(_648_),
    .B(_647_),
    .Y(_649_)
);

INVX1 _1442_ (
    .A(Yin[12]),
    .Y(_650_)
);

NAND2X1 _1443_ (
    .A(Yin[11]),
    .B(_532_),
    .Y(_651_)
);

OR2X2 _1444_ (
    .A(_651_),
    .B(_650_),
    .Y(_652_)
);

NAND2X1 _1445_ (
    .A(_650_),
    .B(_651_),
    .Y(_653_)
);

NAND2X1 _1446_ (
    .A(_653_),
    .B(_652_),
    .Y(_654_)
);

INVX1 _1447_ (
    .A(_654_),
    .Y(_656_)
);

NAND2X1 _1448_ (
    .A(_656_),
    .B(_649_),
    .Y(_657_)
);

OAI21X1 _1449_ (
    .A(_648_),
    .B(_647_),
    .C(_654_),
    .Y(_658_)
);

NAND2X1 _1450_ (
    .A(_658_),
    .B(_657_),
    .Y(_659_)
);

NAND2X1 _1451_ (
    .A(_637_),
    .B(_659_),
    .Y(_660_)
);

INVX1 _1452_ (
    .A(_660_),
    .Y(_661_)
);

NOR2X1 _1453_ (
    .A(_637_),
    .B(_659_),
    .Y(_662_)
);

OAI21X1 _1454_ (
    .A(_662_),
    .B(_661_),
    .C(_636_),
    .Y(_663_)
);

OR2X2 _1455_ (
    .A(_659_),
    .B(_637_),
    .Y(_664_)
);

NAND3X1 _1456_ (
    .A(_635_),
    .B(_660_),
    .C(_664_),
    .Y(_665_)
);

NAND2X1 _1457_ (
    .A(_665_),
    .B(_663_),
    .Y(_667_)
);

NAND3X1 _1458_ (
    .A(_615_),
    .B(_621_),
    .C(_667_),
    .Y(_668_)
);

OAI21X1 _1459_ (
    .A(_611_),
    .B(_608_),
    .C(_621_),
    .Y(_669_)
);

NAND3X1 _1460_ (
    .A(_669_),
    .B(_665_),
    .C(_663_),
    .Y(_670_)
);

NAND2X1 _1461_ (
    .A(_670_),
    .B(_668_),
    .Y(_671_)
);

XNOR2X1 _1462_ (
    .A(_634_),
    .B(_671_),
    .Y(_753_[12])
);

INVX1 _1463_ (
    .A(_634_),
    .Y(_672_)
);

OAI21X1 _1464_ (
    .A(_671_),
    .B(_672_),
    .C(_670_),
    .Y(_673_)
);

AOI21X1 _1465_ (
    .A(_635_),
    .B(_660_),
    .C(_662_),
    .Y(_674_)
);

OAI22X1 _1466_ (
    .A(_578_),
    .B(_639_),
    .C(_643_),
    .D(_641_),
    .Y(_675_)
);

INVX1 _1467_ (
    .A(_576_),
    .Y(_677_)
);

NOR2X1 _1468_ (
    .A(_447_),
    .B(_575_),
    .Y(_678_)
);

NAND2X1 _1469_ (
    .A(_677_),
    .B(_678_),
    .Y(_679_)
);

OAI21X1 _1470_ (
    .A(_352_),
    .B(_575_),
    .C(_639_),
    .Y(_680_)
);

AND2X2 _1471_ (
    .A(_679_),
    .B(_680_),
    .Y(_681_)
);

XOR2X1 _1472_ (
    .A(_681_),
    .B(_675_),
    .Y(_682_)
);

XNOR2X1 _1473_ (
    .A(_682_),
    .B(Yin[13]),
    .Y(_683_)
);

NAND3X1 _1474_ (
    .A(_652_),
    .B(_657_),
    .C(_683_),
    .Y(_684_)
);

INVX1 _1475_ (
    .A(_684_),
    .Y(_685_)
);

AOI21X1 _1476_ (
    .A(_652_),
    .B(_657_),
    .C(_683_),
    .Y(_686_)
);

OAI21X1 _1477_ (
    .A(_686_),
    .B(_685_),
    .C(_646_),
    .Y(_688_)
);

OAI21X1 _1478_ (
    .A(_650_),
    .B(_651_),
    .C(_657_),
    .Y(_689_)
);

INVX1 _1479_ (
    .A(_683_),
    .Y(_690_)
);

NAND2X1 _1480_ (
    .A(_689_),
    .B(_690_),
    .Y(_691_)
);

NAND3X1 _1481_ (
    .A(_647_),
    .B(_684_),
    .C(_691_),
    .Y(_692_)
);

NAND2X1 _1482_ (
    .A(_692_),
    .B(_688_),
    .Y(_693_)
);

XOR2X1 _1483_ (
    .A(_693_),
    .B(_674_),
    .Y(_694_)
);

XOR2X1 _1484_ (
    .A(_673_),
    .B(_694_),
    .Y(_753_[13])
);

NAND2X1 _1485_ (
    .A(_674_),
    .B(_693_),
    .Y(_695_)
);

NAND3X1 _1486_ (
    .A(_668_),
    .B(_670_),
    .C(_694_),
    .Y(_696_)
);

INVX1 _1487_ (
    .A(_696_),
    .Y(_698_)
);

OAI21X1 _1488_ (
    .A(_674_),
    .B(_693_),
    .C(_670_),
    .Y(_699_)
);

AOI22X1 _1489_ (
    .A(_695_),
    .B(_699_),
    .C(_634_),
    .D(_698_),
    .Y(_700_)
);

INVX1 _1490_ (
    .A(_692_),
    .Y(_701_)
);

NOR2X1 _1491_ (
    .A(_686_),
    .B(_701_),
    .Y(_702_)
);

NAND3X1 _1492_ (
    .A(Yin[14]),
    .B(_576_),
    .C(_678_),
    .Y(_703_)
);

INVX1 _1493_ (
    .A(Yin[14]),
    .Y(_704_)
);

INVX1 _1494_ (
    .A(_678_),
    .Y(_705_)
);

OAI21X1 _1495_ (
    .A(_677_),
    .B(_705_),
    .C(_704_),
    .Y(_706_)
);

NAND2X1 _1496_ (
    .A(_703_),
    .B(_706_),
    .Y(_707_)
);

NAND2X1 _1497_ (
    .A(_675_),
    .B(_681_),
    .Y(_709_)
);

NAND2X1 _1498_ (
    .A(Yin[13]),
    .B(_682_),
    .Y(_710_)
);

NAND2X1 _1499_ (
    .A(_709_),
    .B(_710_),
    .Y(_711_)
);

XNOR2X1 _1500_ (
    .A(_711_),
    .B(_707_),
    .Y(_712_)
);

XNOR2X1 _1501_ (
    .A(_702_),
    .B(_712_),
    .Y(_713_)
);

INVX1 _1502_ (
    .A(_713_),
    .Y(_714_)
);

XOR2X1 _1503_ (
    .A(_700_),
    .B(_714_),
    .Y(_753_[14])
);

OAI21X1 _1504_ (
    .A(_686_),
    .B(_701_),
    .C(_712_),
    .Y(_715_)
);

OAI21X1 _1505_ (
    .A(_714_),
    .B(_700_),
    .C(_715_),
    .Y(_716_)
);

NAND3X1 _1506_ (
    .A(_703_),
    .B(_706_),
    .C(_711_),
    .Y(_717_)
);

OAI21X1 _1507_ (
    .A(Yin[14]),
    .B(_677_),
    .C(_678_),
    .Y(_719_)
);

XNOR2X1 _1508_ (
    .A(_719_),
    .B(Yin[15]),
    .Y(_720_)
);

XOR2X1 _1509_ (
    .A(_717_),
    .B(_720_),
    .Y(_721_)
);

NAND2X1 _1510_ (
    .A(_721_),
    .B(_716_),
    .Y(_722_)
);

AOI22X1 _1511_ (
    .A(_618_),
    .B(_631_),
    .C(_627_),
    .D(_492_),
    .Y(_723_)
);

AOI21X1 _1512_ (
    .A(_723_),
    .B(_628_),
    .C(_696_),
    .Y(_724_)
);

AND2X2 _1513_ (
    .A(_699_),
    .B(_695_),
    .Y(_725_)
);

OAI21X1 _1514_ (
    .A(_725_),
    .B(_724_),
    .C(_713_),
    .Y(_726_)
);

INVX1 _1515_ (
    .A(_721_),
    .Y(_727_)
);

NAND3X1 _1516_ (
    .A(_715_),
    .B(_727_),
    .C(_726_),
    .Y(_728_)
);

NAND2X1 _1517_ (
    .A(_728_),
    .B(_722_),
    .Y(_753_[15])
);

OAI21X1 _1518_ (
    .A(_739_),
    .B(_20_),
    .C(_24_),
    .Y(_730_)
);

XOR2X1 _1519_ (
    .A(_730_),
    .B(_72_),
    .Y(_752_[4])
);

DFFPOSX1 _1520_ (
    .CLK(clk_bF$buf5),
    .D(Xin[0]),
    .Q(_754_[0])
);

DFFPOSX1 _1521_ (
    .CLK(clk_bF$buf4),
    .D(Xin[1]),
    .Q(_754_[1])
);

DFFPOSX1 _1522_ (
    .CLK(clk_bF$buf3),
    .D(Xin[2]),
    .Q(_754_[2])
);

DFFPOSX1 _1523_ (
    .CLK(clk_bF$buf2),
    .D(Xin_3_bF$buf1),
    .Q(_754_[3])
);

DFFPOSX1 _1524_ (
    .CLK(clk_bF$buf1),
    .D(Xin[4]),
    .Q(_754_[4])
);

DFFPOSX1 _1525_ (
    .CLK(clk_bF$buf0),
    .D(Xin_5_bF$buf0),
    .Q(_754_[5])
);

DFFPOSX1 _1526_ (
    .CLK(clk_bF$buf5),
    .D(Xin[6]),
    .Q(_754_[6])
);

DFFPOSX1 _1527_ (
    .CLK(clk_bF$buf4),
    .D(Xin[7]),
    .Q(_754_[7])
);

DFFPOSX1 _1528_ (
    .CLK(clk_bF$buf3),
    .D(y[0]),
    .Q(_755_[0])
);

DFFPOSX1 _1529_ (
    .CLK(clk_bF$buf2),
    .D(y[1]),
    .Q(_755_[1])
);

DFFPOSX1 _1530_ (
    .CLK(clk_bF$buf1),
    .D(y[2]),
    .Q(_755_[2])
);

DFFPOSX1 _1531_ (
    .CLK(clk_bF$buf0),
    .D(y[3]),
    .Q(_755_[3])
);

DFFPOSX1 _1532_ (
    .CLK(clk_bF$buf5),
    .D(y[4]),
    .Q(_755_[4])
);

DFFPOSX1 _1533_ (
    .CLK(clk_bF$buf4),
    .D(y[5]),
    .Q(_755_[5])
);

DFFPOSX1 _1534_ (
    .CLK(clk_bF$buf3),
    .D(y[6]),
    .Q(_755_[6])
);

DFFPOSX1 _1535_ (
    .CLK(clk_bF$buf2),
    .D(y[7]),
    .Q(_755_[7])
);

DFFPOSX1 _1536_ (
    .CLK(clk_bF$buf1),
    .D(y[8]),
    .Q(_755_[8])
);

DFFPOSX1 _1537_ (
    .CLK(clk_bF$buf0),
    .D(y[9]),
    .Q(_755_[9])
);

DFFPOSX1 _1538_ (
    .CLK(clk_bF$buf5),
    .D(y[10]),
    .Q(_755_[10])
);

DFFPOSX1 _1539_ (
    .CLK(clk_bF$buf4),
    .D(y[11]),
    .Q(_755_[11])
);

DFFPOSX1 _1540_ (
    .CLK(clk_bF$buf3),
    .D(y[12]),
    .Q(_755_[12])
);

DFFPOSX1 _1541_ (
    .CLK(clk_bF$buf2),
    .D(y[13]),
    .Q(_755_[13])
);

DFFPOSX1 _1542_ (
    .CLK(clk_bF$buf1),
    .D(y[14]),
    .Q(_755_[14])
);

DFFPOSX1 _1543_ (
    .CLK(clk_bF$buf0),
    .D(y[15]),
    .Q(_755_[15])
);

DFFPOSX1 _1544_ (
    .CLK(clk_bF$buf5),
    .D(_748_[0]),
    .Q(y[0])
);

DFFPOSX1 _1545_ (
    .CLK(clk_bF$buf4),
    .D(_749_[1]),
    .Q(y[1])
);

DFFPOSX1 _1546_ (
    .CLK(clk_bF$buf3),
    .D(_750_[2]),
    .Q(y[2])
);

DFFPOSX1 _1547_ (
    .CLK(clk_bF$buf2),
    .D(_751_[3]),
    .Q(y[3])
);

DFFPOSX1 _1548_ (
    .CLK(clk_bF$buf1),
    .D(_752_[4]),
    .Q(y[4])
);

DFFPOSX1 _1549_ (
    .CLK(clk_bF$buf0),
    .D(_753_[5]),
    .Q(y[5])
);

DFFPOSX1 _1550_ (
    .CLK(clk_bF$buf5),
    .D(_753_[6]),
    .Q(y[6])
);

DFFPOSX1 _1551_ (
    .CLK(clk_bF$buf4),
    .D(_753_[7]),
    .Q(y[7])
);

DFFPOSX1 _1552_ (
    .CLK(clk_bF$buf3),
    .D(_753_[8]),
    .Q(y[8])
);

DFFPOSX1 _1553_ (
    .CLK(clk_bF$buf2),
    .D(_753_[9]),
    .Q(y[9])
);

DFFPOSX1 _1554_ (
    .CLK(clk_bF$buf1),
    .D(_753_[10]),
    .Q(y[10])
);

DFFPOSX1 _1555_ (
    .CLK(clk_bF$buf0),
    .D(_753_[11]),
    .Q(y[11])
);

DFFPOSX1 _1556_ (
    .CLK(clk_bF$buf5),
    .D(_753_[12]),
    .Q(y[12])
);

DFFPOSX1 _1557_ (
    .CLK(clk_bF$buf4),
    .D(_753_[13]),
    .Q(y[13])
);

DFFPOSX1 _1558_ (
    .CLK(clk_bF$buf3),
    .D(_753_[14]),
    .Q(y[14])
);

DFFPOSX1 _1559_ (
    .CLK(clk_bF$buf2),
    .D(_753_[15]),
    .Q(y[15])
);

BUFX2 _1560_ (
    .A(_754_[0]),
    .Y(Xout[0])
);

BUFX2 _1561_ (
    .A(_754_[1]),
    .Y(Xout[1])
);

BUFX2 _1562_ (
    .A(_754_[2]),
    .Y(Xout[2])
);

BUFX2 _1563_ (
    .A(_754_[3]),
    .Y(Xout[3])
);

BUFX2 _1564_ (
    .A(_754_[4]),
    .Y(Xout[4])
);

BUFX2 _1565_ (
    .A(_754_[5]),
    .Y(Xout[5])
);

BUFX2 _1566_ (
    .A(_754_[6]),
    .Y(Xout[6])
);

BUFX2 _1567_ (
    .A(_754_[7]),
    .Y(Xout[7])
);

BUFX2 _1568_ (
    .A(_755_[0]),
    .Y(Yout[0])
);

BUFX2 _1569_ (
    .A(_755_[1]),
    .Y(Yout[1])
);

BUFX2 _1570_ (
    .A(_755_[10]),
    .Y(Yout[10])
);

BUFX2 _1571_ (
    .A(_755_[11]),
    .Y(Yout[11])
);

BUFX2 _1572_ (
    .A(_755_[12]),
    .Y(Yout[12])
);

BUFX2 _1573_ (
    .A(_755_[13]),
    .Y(Yout[13])
);

BUFX2 _1574_ (
    .A(_755_[14]),
    .Y(Yout[14])
);

BUFX2 _1575_ (
    .A(_755_[15]),
    .Y(Yout[15])
);

BUFX2 _1576_ (
    .A(_755_[2]),
    .Y(Yout[2])
);

BUFX2 _1577_ (
    .A(_755_[3]),
    .Y(Yout[3])
);

BUFX2 _1578_ (
    .A(_755_[4]),
    .Y(Yout[4])
);

BUFX2 _1579_ (
    .A(_755_[5]),
    .Y(Yout[5])
);

BUFX2 _1580_ (
    .A(_755_[6]),
    .Y(Yout[6])
);

BUFX2 _1581_ (
    .A(_755_[7]),
    .Y(Yout[7])
);

BUFX2 _1582_ (
    .A(_755_[8]),
    .Y(Yout[8])
);

BUFX2 _1583_ (
    .A(_755_[9]),
    .Y(Yout[9])
);

INVX1 _756_ (
    .A(Cin_0_bF$buf2),
    .Y(_386_)
);

INVX1 _757_ (
    .A(Xin[0]),
    .Y(_397_)
);

NOR2X1 _758_ (
    .A(_386_),
    .B(_397_),
    .Y(_407_)
);

NAND2X1 _759_ (
    .A(Yin[0]),
    .B(_407_),
    .Y(_418_)
);

INVX1 _760_ (
    .A(_418_),
    .Y(_429_)
);

NOR2X1 _761_ (
    .A(Yin[0]),
    .B(_407_),
    .Y(_440_)
);

NOR2X1 _762_ (
    .A(_440_),
    .B(_429_),
    .Y(_748_[0])
);

NAND2X1 _763_ (
    .A(Xin[0]),
    .B(Cin[1]),
    .Y(_461_)
);

INVX1 _764_ (
    .A(_461_),
    .Y(_472_)
);

NAND3X1 _765_ (
    .A(Cin_0_bF$buf1),
    .B(Xin[1]),
    .C(Yin[1]),
    .Y(_483_)
);

AOI21X1 _766_ (
    .A(Cin_0_bF$buf0),
    .B(Xin[1]),
    .C(Yin[1]),
    .Y(_493_)
);

INVX1 _767_ (
    .A(_493_),
    .Y(_504_)
);

NAND3X1 _768_ (
    .A(_472_),
    .B(_483_),
    .C(_504_),
    .Y(_515_)
);

INVX1 _769_ (
    .A(_483_),
    .Y(_526_)
);

OAI21X1 _770_ (
    .A(_493_),
    .B(_526_),
    .C(_461_),
    .Y(_537_)
);

NAND3X1 _771_ (
    .A(_515_),
    .B(_537_),
    .C(_429_),
    .Y(_548_)
);

INVX1 _772_ (
    .A(_548_),
    .Y(_559_)
);

AOI21X1 _773_ (
    .A(_515_),
    .B(_537_),
    .C(_429_),
    .Y(_569_)
);

NOR2X1 _774_ (
    .A(_569_),
    .B(_559_),
    .Y(_749_[1])
);

INVX2 _775_ (
    .A(Cin[2]),
    .Y(_590_)
);

NOR2X1 _776_ (
    .A(_397_),
    .B(_590_),
    .Y(_601_)
);

OAI21X1 _777_ (
    .A(_461_),
    .B(_493_),
    .C(_483_),
    .Y(_612_)
);

NAND2X1 _778_ (
    .A(Xin[1]),
    .B(Cin[1]),
    .Y(_623_)
);

INVX1 _779_ (
    .A(_623_),
    .Y(_633_)
);

NAND3X1 _780_ (
    .A(Cin_0_bF$buf3),
    .B(Xin[2]),
    .C(Yin[2]),
    .Y(_644_)
);

AOI21X1 _781_ (
    .A(Cin_0_bF$buf2),
    .B(Xin[2]),
    .C(Yin[2]),
    .Y(_655_)
);

INVX1 _782_ (
    .A(_655_),
    .Y(_666_)
);

NAND3X1 _783_ (
    .A(_633_),
    .B(_644_),
    .C(_666_),
    .Y(_676_)
);

INVX1 _784_ (
    .A(_644_),
    .Y(_687_)
);

OAI21X1 _785_ (
    .A(_655_),
    .B(_687_),
    .C(_623_),
    .Y(_697_)
);

NAND3X1 _786_ (
    .A(_612_),
    .B(_676_),
    .C(_697_),
    .Y(_708_)
);

AOI21X1 _787_ (
    .A(_697_),
    .B(_676_),
    .C(_612_),
    .Y(_718_)
);

INVX1 _788_ (
    .A(_718_),
    .Y(_729_)
);

NAND3X1 _789_ (
    .A(_601_),
    .B(_708_),
    .C(_729_),
    .Y(_731_)
);

INVX1 _790_ (
    .A(_601_),
    .Y(_732_)
);

INVX1 _791_ (
    .A(_708_),
    .Y(_733_)
);

OAI21X1 _792_ (
    .A(_718_),
    .B(_733_),
    .C(_732_),
    .Y(_734_)
);

NAND3X1 _793_ (
    .A(_559_),
    .B(_734_),
    .C(_731_),
    .Y(_735_)
);

INVX1 _794_ (
    .A(_735_),
    .Y(_736_)
);

AOI21X1 _795_ (
    .A(_731_),
    .B(_734_),
    .C(_559_),
    .Y(_737_)
);

NOR2X1 _796_ (
    .A(_737_),
    .B(_736_),
    .Y(_750_[2])
);

OAI21X1 _797_ (
    .A(_732_),
    .B(_718_),
    .C(_708_),
    .Y(_738_)
);

INVX1 _798_ (
    .A(_738_),
    .Y(_739_)
);

INVX2 _799_ (
    .A(Cin[3]),
    .Y(_740_)
);

NAND2X1 _800_ (
    .A(Xin[1]),
    .B(Cin[2]),
    .Y(_741_)
);

OAI21X1 _801_ (
    .A(_397_),
    .B(_740_),
    .C(_741_),
    .Y(_742_)
);

AND2X2 _802_ (
    .A(Xin[1]),
    .B(Cin[3]),
    .Y(_743_)
);

NAND2X1 _803_ (
    .A(_743_),
    .B(_601_),
    .Y(_744_)
);

AND2X2 _804_ (
    .A(_744_),
    .B(_742_),
    .Y(_745_)
);

OAI21X1 _805_ (
    .A(_623_),
    .B(_655_),
    .C(_644_),
    .Y(_746_)
);

NAND2X1 _806_ (
    .A(Cin[1]),
    .B(Xin[2]),
    .Y(_747_)
);

INVX1 _807_ (
    .A(_747_),
    .Y(_0_)
);

NAND3X1 _808_ (
    .A(Cin_0_bF$buf1),
    .B(Xin_3_bF$buf0),
    .C(Yin[3]),
    .Y(_1_)
);

INVX1 _809_ (
    .A(Yin[3]),
    .Y(_2_)
);

NAND2X1 _810_ (
    .A(Cin_0_bF$buf0),
    .B(Xin_3_bF$buf3),
    .Y(_3_)
);

NAND2X1 _811_ (
    .A(_2_),
    .B(_3_),
    .Y(_4_)
);

NAND3X1 _812_ (
    .A(_1_),
    .B(_0_),
    .C(_4_),
    .Y(_5_)
);

NAND2X1 _813_ (
    .A(Yin[3]),
    .B(_3_),
    .Y(_6_)
);

NAND3X1 _814_ (
    .A(Cin_0_bF$buf3),
    .B(Xin_3_bF$buf2),
    .C(_2_),
    .Y(_7_)
);

NAND3X1 _815_ (
    .A(_747_),
    .B(_6_),
    .C(_7_),
    .Y(_8_)
);

NAND3X1 _816_ (
    .A(_746_),
    .B(_5_),
    .C(_8_),
    .Y(_9_)
);

INVX1 _817_ (
    .A(_746_),
    .Y(_10_)
);

AOI21X1 _818_ (
    .A(_7_),
    .B(_6_),
    .C(_747_),
    .Y(_11_)
);

AOI21X1 _819_ (
    .A(_4_),
    .B(_1_),
    .C(_0_),
    .Y(_12_)
);

OAI21X1 _820_ (
    .A(_12_),
    .B(_11_),
    .C(_10_),
    .Y(_13_)
);

NAND3X1 _821_ (
    .A(_9_),
    .B(_13_),
    .C(_745_),
    .Y(_14_)
);

NAND2X1 _822_ (
    .A(Xin[1]),
    .B(Cin[3]),
    .Y(_15_)
);

OAI21X1 _823_ (
    .A(_15_),
    .B(_732_),
    .C(_742_),
    .Y(_16_)
);

INVX1 _824_ (
    .A(_9_),
    .Y(_17_)
);

AOI21X1 _825_ (
    .A(_8_),
    .B(_5_),
    .C(_746_),
    .Y(_18_)
);

OAI21X1 _826_ (
    .A(_18_),
    .B(_17_),
    .C(_16_),
    .Y(_19_)
);

NAND2X1 _827_ (
    .A(_14_),
    .B(_19_),
    .Y(_20_)
);

NOR2X1 _828_ (
    .A(_739_),
    .B(_20_),
    .Y(_21_)
);

AOI21X1 _829_ (
    .A(_19_),
    .B(_14_),
    .C(_738_),
    .Y(_22_)
);

NOR3X1 _830_ (
    .A(_735_),
    .B(_22_),
    .C(_21_),
    .Y(_23_)
);

INVX1 _831_ (
    .A(_23_),
    .Y(_24_)
);

OAI21X1 _832_ (
    .A(_22_),
    .B(_21_),
    .C(_735_),
    .Y(_25_)
);

AND2X2 _833_ (
    .A(_24_),
    .B(_25_),
    .Y(_751_[3])
);

INVX1 _834_ (
    .A(_744_),
    .Y(_26_)
);

OAI21X1 _835_ (
    .A(_18_),
    .B(_16_),
    .C(_9_),
    .Y(_27_)
);

AOI21X1 _836_ (
    .A(Cin_0_bF$buf2),
    .B(Xin_3_bF$buf1),
    .C(Yin[3]),
    .Y(_28_)
);

OAI21X1 _837_ (
    .A(_747_),
    .B(_28_),
    .C(_1_),
    .Y(_29_)
);

NAND3X1 _838_ (
    .A(Cin_0_bF$buf1),
    .B(Xin[4]),
    .C(Yin[4]),
    .Y(_30_)
);

AOI21X1 _839_ (
    .A(Cin_0_bF$buf0),
    .B(Xin[4]),
    .C(Yin[4]),
    .Y(_31_)
);

INVX1 _840_ (
    .A(_31_),
    .Y(_32_)
);

NAND2X1 _841_ (
    .A(Cin[1]),
    .B(Xin_3_bF$buf0),
    .Y(_33_)
);

INVX1 _842_ (
    .A(_33_),
    .Y(_34_)
);

NAND3X1 _843_ (
    .A(_30_),
    .B(_34_),
    .C(_32_),
    .Y(_35_)
);

INVX1 _844_ (
    .A(_30_),
    .Y(_36_)
);

OAI21X1 _845_ (
    .A(_31_),
    .B(_36_),
    .C(_33_),
    .Y(_37_)
);

NAND3X1 _846_ (
    .A(_29_),
    .B(_35_),
    .C(_37_),
    .Y(_38_)
);

INVX1 _847_ (
    .A(_1_),
    .Y(_39_)
);

AOI21X1 _848_ (
    .A(_0_),
    .B(_4_),
    .C(_39_),
    .Y(_40_)
);

OAI21X1 _849_ (
    .A(_31_),
    .B(_36_),
    .C(_34_),
    .Y(_41_)
);

NAND3X1 _850_ (
    .A(_30_),
    .B(_33_),
    .C(_32_),
    .Y(_42_)
);

NAND3X1 _851_ (
    .A(_42_),
    .B(_41_),
    .C(_40_),
    .Y(_43_)
);

NAND2X1 _852_ (
    .A(Xin[0]),
    .B(Cin[4]),
    .Y(_44_)
);

AND2X2 _853_ (
    .A(Xin[2]),
    .B(Cin[2]),
    .Y(_45_)
);

NAND2X1 _854_ (
    .A(_743_),
    .B(_45_),
    .Y(_46_)
);

INVX2 _855_ (
    .A(Xin[2]),
    .Y(_47_)
);

OAI21X1 _856_ (
    .A(_47_),
    .B(_590_),
    .C(_15_),
    .Y(_48_)
);

NAND3X1 _857_ (
    .A(_44_),
    .B(_48_),
    .C(_46_),
    .Y(_49_)
);

INVX1 _858_ (
    .A(_44_),
    .Y(_50_)
);

INVX1 _859_ (
    .A(Xin[1]),
    .Y(_51_)
);

OAI21X1 _860_ (
    .A(_51_),
    .B(_740_),
    .C(_45_),
    .Y(_52_)
);

OAI21X1 _861_ (
    .A(_47_),
    .B(_590_),
    .C(_743_),
    .Y(_53_)
);

NAND3X1 _862_ (
    .A(_50_),
    .B(_52_),
    .C(_53_),
    .Y(_54_)
);

NAND2X1 _863_ (
    .A(_49_),
    .B(_54_),
    .Y(_55_)
);

NAND3X1 _864_ (
    .A(_38_),
    .B(_55_),
    .C(_43_),
    .Y(_56_)
);

AOI21X1 _865_ (
    .A(_41_),
    .B(_42_),
    .C(_40_),
    .Y(_57_)
);

AOI21X1 _866_ (
    .A(_37_),
    .B(_35_),
    .C(_29_),
    .Y(_58_)
);

NAND3X1 _867_ (
    .A(_48_),
    .B(_50_),
    .C(_46_),
    .Y(_59_)
);

NAND3X1 _868_ (
    .A(_44_),
    .B(_52_),
    .C(_53_),
    .Y(_60_)
);

NAND2X1 _869_ (
    .A(_59_),
    .B(_60_),
    .Y(_61_)
);

OAI21X1 _870_ (
    .A(_57_),
    .B(_58_),
    .C(_61_),
    .Y(_62_)
);

NAND3X1 _871_ (
    .A(_27_),
    .B(_56_),
    .C(_62_),
    .Y(_63_)
);

AOI21X1 _872_ (
    .A(_745_),
    .B(_13_),
    .C(_17_),
    .Y(_64_)
);

OAI21X1 _873_ (
    .A(_57_),
    .B(_58_),
    .C(_55_),
    .Y(_65_)
);

NAND3X1 _874_ (
    .A(_38_),
    .B(_61_),
    .C(_43_),
    .Y(_66_)
);

NAND3X1 _875_ (
    .A(_65_),
    .B(_66_),
    .C(_64_),
    .Y(_67_)
);

NAND3X1 _876_ (
    .A(_26_),
    .B(_63_),
    .C(_67_),
    .Y(_68_)
);

AOI22X1 _877_ (
    .A(_9_),
    .B(_14_),
    .C(_65_),
    .D(_66_),
    .Y(_69_)
);

AOI21X1 _878_ (
    .A(_62_),
    .B(_56_),
    .C(_27_),
    .Y(_70_)
);

OAI21X1 _879_ (
    .A(_69_),
    .B(_70_),
    .C(_744_),
    .Y(_71_)
);

AND2X2 _880_ (
    .A(_71_),
    .B(_68_),
    .Y(_72_)
);

NAND2X1 _881_ (
    .A(_72_),
    .B(_23_),
    .Y(_73_)
);

NAND3X1 _882_ (
    .A(_68_),
    .B(_21_),
    .C(_71_),
    .Y(_74_)
);

INVX1 _883_ (
    .A(_74_),
    .Y(_75_)
);

OAI21X1 _884_ (
    .A(_744_),
    .B(_70_),
    .C(_63_),
    .Y(_76_)
);

INVX1 _885_ (
    .A(Cin[5]),
    .Y(_77_)
);

NOR2X1 _886_ (
    .A(_397_),
    .B(_77_),
    .Y(_78_)
);

NAND2X1 _887_ (
    .A(Xin[2]),
    .B(Cin[3]),
    .Y(_79_)
);

OAI21X1 _888_ (
    .A(_741_),
    .B(_79_),
    .C(_59_),
    .Y(_80_)
);

XOR2X1 _889_ (
    .A(_80_),
    .B(_78_),
    .Y(_81_)
);

OAI21X1 _890_ (
    .A(_61_),
    .B(_58_),
    .C(_38_),
    .Y(_82_)
);

NAND2X1 _891_ (
    .A(Xin[1]),
    .B(Cin[4]),
    .Y(_83_)
);

INVX1 _892_ (
    .A(_83_),
    .Y(_84_)
);

AND2X2 _893_ (
    .A(Xin_3_bF$buf3),
    .B(Cin[3]),
    .Y(_85_)
);

NAND2X1 _894_ (
    .A(_45_),
    .B(_85_),
    .Y(_86_)
);

INVX1 _895_ (
    .A(Xin_3_bF$buf2),
    .Y(_87_)
);

OAI21X1 _896_ (
    .A(_590_),
    .B(_87_),
    .C(_79_),
    .Y(_88_)
);

NAND3X1 _897_ (
    .A(_84_),
    .B(_88_),
    .C(_86_),
    .Y(_89_)
);

NAND3X1 _898_ (
    .A(Cin[2]),
    .B(Xin_3_bF$buf1),
    .C(_79_),
    .Y(_90_)
);

NAND2X1 _899_ (
    .A(Cin[2]),
    .B(Xin_3_bF$buf0),
    .Y(_91_)
);

NAND3X1 _900_ (
    .A(Xin[2]),
    .B(Cin[3]),
    .C(_91_),
    .Y(_92_)
);

NAND3X1 _901_ (
    .A(_83_),
    .B(_90_),
    .C(_92_),
    .Y(_93_)
);

AND2X2 _902_ (
    .A(_89_),
    .B(_93_),
    .Y(_94_)
);

OAI21X1 _903_ (
    .A(_33_),
    .B(_31_),
    .C(_30_),
    .Y(_95_)
);

NAND2X1 _904_ (
    .A(Cin[1]),
    .B(Xin[4]),
    .Y(_96_)
);

INVX1 _905_ (
    .A(_96_),
    .Y(_97_)
);

NAND3X1 _906_ (
    .A(Cin_0_bF$buf3),
    .B(Xin_5_bF$buf3),
    .C(Yin[5]),
    .Y(_98_)
);

INVX1 _907_ (
    .A(Yin[5]),
    .Y(_99_)
);

NAND2X1 _908_ (
    .A(Cin_0_bF$buf2),
    .B(Xin_5_bF$buf2),
    .Y(_100_)
);

NAND2X1 _909_ (
    .A(_99_),
    .B(_100_),
    .Y(_101_)
);

NAND3X1 _910_ (
    .A(_98_),
    .B(_97_),
    .C(_101_),
    .Y(_102_)
);

NAND2X1 _911_ (
    .A(Yin[5]),
    .B(_100_),
    .Y(_103_)
);

NAND3X1 _912_ (
    .A(Cin_0_bF$buf1),
    .B(Xin_5_bF$buf1),
    .C(_99_),
    .Y(_104_)
);

NAND3X1 _913_ (
    .A(_96_),
    .B(_103_),
    .C(_104_),
    .Y(_105_)
);

NAND3X1 _914_ (
    .A(_95_),
    .B(_102_),
    .C(_105_),
    .Y(_106_)
);

INVX1 _915_ (
    .A(_95_),
    .Y(_107_)
);

AOI21X1 _916_ (
    .A(_104_),
    .B(_103_),
    .C(_96_),
    .Y(_108_)
);

AOI21X1 _917_ (
    .A(_101_),
    .B(_98_),
    .C(_97_),
    .Y(_109_)
);

OAI21X1 _918_ (
    .A(_109_),
    .B(_108_),
    .C(_107_),
    .Y(_110_)
);

NAND3X1 _919_ (
    .A(_106_),
    .B(_110_),
    .C(_94_),
    .Y(_111_)
);

NAND2X1 _920_ (
    .A(_93_),
    .B(_89_),
    .Y(_112_)
);

OAI21X1 _921_ (
    .A(_109_),
    .B(_108_),
    .C(_95_),
    .Y(_113_)
);

NAND3X1 _922_ (
    .A(_102_),
    .B(_105_),
    .C(_107_),
    .Y(_114_)
);

NAND3X1 _923_ (
    .A(_112_),
    .B(_114_),
    .C(_113_),
    .Y(_115_)
);

NAND3X1 _924_ (
    .A(_115_),
    .B(_111_),
    .C(_82_),
    .Y(_116_)
);

AOI21X1 _925_ (
    .A(_43_),
    .B(_55_),
    .C(_57_),
    .Y(_117_)
);

AOI21X1 _926_ (
    .A(_113_),
    .B(_114_),
    .C(_112_),
    .Y(_118_)
);

AOI22X1 _927_ (
    .A(_89_),
    .B(_93_),
    .C(_110_),
    .D(_106_),
    .Y(_119_)
);

OAI21X1 _928_ (
    .A(_119_),
    .B(_118_),
    .C(_117_),
    .Y(_120_)
);

NAND3X1 _929_ (
    .A(_81_),
    .B(_116_),
    .C(_120_),
    .Y(_121_)
);

INVX1 _930_ (
    .A(_78_),
    .Y(_122_)
);

XOR2X1 _931_ (
    .A(_80_),
    .B(_122_),
    .Y(_123_)
);

OAI21X1 _932_ (
    .A(_119_),
    .B(_118_),
    .C(_82_),
    .Y(_124_)
);

NAND3X1 _933_ (
    .A(_115_),
    .B(_111_),
    .C(_117_),
    .Y(_125_)
);

NAND3X1 _934_ (
    .A(_123_),
    .B(_125_),
    .C(_124_),
    .Y(_126_)
);

NAND3X1 _935_ (
    .A(_121_),
    .B(_126_),
    .C(_76_),
    .Y(_127_)
);

AOI21X1 _936_ (
    .A(_67_),
    .B(_26_),
    .C(_69_),
    .Y(_128_)
);

AOI21X1 _937_ (
    .A(_124_),
    .B(_125_),
    .C(_123_),
    .Y(_129_)
);

AOI21X1 _938_ (
    .A(_120_),
    .B(_116_),
    .C(_81_),
    .Y(_130_)
);

OAI21X1 _939_ (
    .A(_129_),
    .B(_130_),
    .C(_128_),
    .Y(_131_)
);

NAND3X1 _940_ (
    .A(_127_),
    .B(_131_),
    .C(_75_),
    .Y(_132_)
);

AOI22X1 _941_ (
    .A(_127_),
    .B(_131_),
    .C(_72_),
    .D(_21_),
    .Y(_133_)
);

INVX1 _942_ (
    .A(_133_),
    .Y(_134_)
);

NAND2X1 _943_ (
    .A(_132_),
    .B(_134_),
    .Y(_135_)
);

XOR2X1 _944_ (
    .A(_135_),
    .B(_73_),
    .Y(_753_[5])
);

OAI21X1 _945_ (
    .A(_73_),
    .B(_133_),
    .C(_132_),
    .Y(_136_)
);

NAND2X1 _946_ (
    .A(_78_),
    .B(_80_),
    .Y(_137_)
);

AOI21X1 _947_ (
    .A(_111_),
    .B(_115_),
    .C(_82_),
    .Y(_138_)
);

OAI21X1 _948_ (
    .A(_123_),
    .B(_138_),
    .C(_116_),
    .Y(_139_)
);

AND2X2 _949_ (
    .A(Xin[1]),
    .B(Cin[6]),
    .Y(_140_)
);

AOI22X1 _950_ (
    .A(Xin[0]),
    .B(Cin[6]),
    .C(Xin[1]),
    .D(Cin[5]),
    .Y(_141_)
);

AOI21X1 _951_ (
    .A(_78_),
    .B(_140_),
    .C(_141_),
    .Y(_142_)
);

OAI21X1 _952_ (
    .A(_79_),
    .B(_91_),
    .C(_89_),
    .Y(_143_)
);

XNOR2X1 _953_ (
    .A(_143_),
    .B(_142_),
    .Y(_144_)
);

AOI21X1 _954_ (
    .A(_105_),
    .B(_102_),
    .C(_95_),
    .Y(_145_)
);

OAI21X1 _955_ (
    .A(_112_),
    .B(_145_),
    .C(_106_),
    .Y(_146_)
);

NAND2X1 _956_ (
    .A(Xin[2]),
    .B(Cin[4]),
    .Y(_147_)
);

INVX1 _957_ (
    .A(_147_),
    .Y(_148_)
);

AND2X2 _958_ (
    .A(Cin[2]),
    .B(Xin[4]),
    .Y(_149_)
);

NAND2X1 _959_ (
    .A(_85_),
    .B(_149_),
    .Y(_150_)
);

INVX2 _960_ (
    .A(Xin[4]),
    .Y(_151_)
);

NAND2X1 _961_ (
    .A(Xin_3_bF$buf3),
    .B(Cin[3]),
    .Y(_152_)
);

OAI21X1 _962_ (
    .A(_590_),
    .B(_151_),
    .C(_152_),
    .Y(_153_)
);

NAND3X1 _963_ (
    .A(_153_),
    .B(_148_),
    .C(_150_),
    .Y(_154_)
);

OAI21X1 _964_ (
    .A(_590_),
    .B(_151_),
    .C(_85_),
    .Y(_155_)
);

OAI21X1 _965_ (
    .A(_87_),
    .B(_740_),
    .C(_149_),
    .Y(_156_)
);

NAND3X1 _966_ (
    .A(_147_),
    .B(_155_),
    .C(_156_),
    .Y(_157_)
);

NAND2X1 _967_ (
    .A(_154_),
    .B(_157_),
    .Y(_158_)
);

AOI21X1 _968_ (
    .A(Cin_0_bF$buf0),
    .B(Xin_5_bF$buf0),
    .C(Yin[5]),
    .Y(_159_)
);

OAI21X1 _969_ (
    .A(_96_),
    .B(_159_),
    .C(_98_),
    .Y(_160_)
);

NAND2X1 _970_ (
    .A(Cin[1]),
    .B(Xin_5_bF$buf3),
    .Y(_161_)
);

NAND2X1 _971_ (
    .A(Cin_0_bF$buf3),
    .B(Xin[6]),
    .Y(_162_)
);

NAND2X1 _972_ (
    .A(Yin[6]),
    .B(_162_),
    .Y(_163_)
);

INVX1 _973_ (
    .A(Yin[6]),
    .Y(_164_)
);

NAND3X1 _974_ (
    .A(Cin_0_bF$buf2),
    .B(Xin[6]),
    .C(_164_),
    .Y(_165_)
);

AOI21X1 _975_ (
    .A(_165_),
    .B(_163_),
    .C(_161_),
    .Y(_166_)
);

INVX1 _976_ (
    .A(_161_),
    .Y(_167_)
);

NAND3X1 _977_ (
    .A(Cin_0_bF$buf1),
    .B(Xin[6]),
    .C(Yin[6]),
    .Y(_168_)
);

NAND2X1 _978_ (
    .A(_164_),
    .B(_162_),
    .Y(_169_)
);

AOI21X1 _979_ (
    .A(_169_),
    .B(_168_),
    .C(_167_),
    .Y(_170_)
);

OAI21X1 _980_ (
    .A(_170_),
    .B(_166_),
    .C(_160_),
    .Y(_171_)
);

INVX1 _981_ (
    .A(_160_),
    .Y(_172_)
);

NAND3X1 _982_ (
    .A(_168_),
    .B(_167_),
    .C(_169_),
    .Y(_173_)
);

NAND3X1 _983_ (
    .A(_161_),
    .B(_163_),
    .C(_165_),
    .Y(_174_)
);

NAND3X1 _984_ (
    .A(_173_),
    .B(_174_),
    .C(_172_),
    .Y(_175_)
);

AOI21X1 _985_ (
    .A(_171_),
    .B(_175_),
    .C(_158_),
    .Y(_176_)
);

NAND3X1 _986_ (
    .A(_160_),
    .B(_173_),
    .C(_174_),
    .Y(_177_)
);

OAI21X1 _987_ (
    .A(_170_),
    .B(_166_),
    .C(_172_),
    .Y(_178_)
);

AOI22X1 _988_ (
    .A(_154_),
    .B(_157_),
    .C(_178_),
    .D(_177_),
    .Y(_179_)
);

OAI21X1 _989_ (
    .A(_179_),
    .B(_176_),
    .C(_146_),
    .Y(_180_)
);

INVX1 _990_ (
    .A(_106_),
    .Y(_181_)
);

AOI21X1 _991_ (
    .A(_94_),
    .B(_110_),
    .C(_181_),
    .Y(_182_)
);

AND2X2 _992_ (
    .A(_157_),
    .B(_154_),
    .Y(_183_)
);

NAND3X1 _993_ (
    .A(_177_),
    .B(_178_),
    .C(_183_),
    .Y(_184_)
);

NAND3X1 _994_ (
    .A(_158_),
    .B(_171_),
    .C(_175_),
    .Y(_185_)
);

NAND3X1 _995_ (
    .A(_184_),
    .B(_185_),
    .C(_182_),
    .Y(_186_)
);

AOI21X1 _996_ (
    .A(_186_),
    .B(_180_),
    .C(_144_),
    .Y(_187_)
);

XOR2X1 _997_ (
    .A(_143_),
    .B(_142_),
    .Y(_188_)
);

NAND3X1 _998_ (
    .A(_146_),
    .B(_185_),
    .C(_184_),
    .Y(_189_)
);

OAI21X1 _999_ (
    .A(_176_),
    .B(_179_),
    .C(_182_),
    .Y(_190_)
);

endmodule
